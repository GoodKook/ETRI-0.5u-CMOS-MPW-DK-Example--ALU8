magic
tech scmos
magscale 1 60
timestamp 1709419192
<< checkpaint >>
rect -1200 -1200 381200 381200
<< metal1 >>
rect 287000 199270 291700 199400
rect 287000 199090 290930 199270
rect 291110 199090 291290 199270
rect 291470 199090 291700 199270
rect 287000 198910 291700 199090
rect 287000 198730 290930 198910
rect 291110 198730 291290 198910
rect 291470 198730 291700 198910
rect 287000 198550 291700 198730
rect 287000 198370 290930 198550
rect 291110 198370 291290 198550
rect 291470 198370 291700 198550
rect 287000 198190 291700 198370
rect 287000 198010 290930 198190
rect 291110 198010 291290 198190
rect 291470 198010 291700 198190
rect 287000 197830 291700 198010
rect 287000 197650 290930 197830
rect 291110 197650 291290 197830
rect 291470 197650 291700 197830
rect 287000 197470 291700 197650
rect 287000 197290 290930 197470
rect 291110 197290 291290 197470
rect 291470 197290 291700 197470
rect 287000 197110 291700 197290
rect 287000 196930 290930 197110
rect 291110 196930 291290 197110
rect 291470 196930 291700 197110
rect 287000 196750 291700 196930
rect 88400 196520 96400 196700
rect 88400 196340 88530 196520
rect 88710 196340 88890 196520
rect 89070 196340 96400 196520
rect 88400 196160 96400 196340
rect 88400 195980 88530 196160
rect 88710 195980 88890 196160
rect 89070 195980 96400 196160
rect 88400 195800 96400 195980
rect 88400 195620 88530 195800
rect 88710 195620 88890 195800
rect 89070 195620 96400 195800
rect 88400 195440 96400 195620
rect 88400 195260 88530 195440
rect 88710 195260 88890 195440
rect 89070 195260 96400 195440
rect 88400 195080 96400 195260
rect 88400 194900 88530 195080
rect 88710 194900 88890 195080
rect 89070 194900 96400 195080
rect 88400 194720 96400 194900
rect 88400 194540 88530 194720
rect 88710 194540 88890 194720
rect 89070 194540 96400 194720
rect 88400 194360 96400 194540
rect 88400 194180 88530 194360
rect 88710 194180 88890 194360
rect 89070 194180 96400 194360
rect 88400 194000 96400 194180
rect 88400 193820 88530 194000
rect 88710 193820 88890 194000
rect 89070 193820 96400 194000
rect 88400 193640 96400 193820
rect 88400 193460 88530 193640
rect 88710 193460 88890 193640
rect 89070 193460 96400 193640
rect 88400 193280 96400 193460
rect 88400 193100 88530 193280
rect 88710 193100 88890 193280
rect 89070 193100 96400 193280
rect 88400 192920 96400 193100
rect 88400 192740 88530 192920
rect 88710 192740 88890 192920
rect 89070 192740 96400 192920
rect 88400 192560 96400 192740
rect 88400 192380 88530 192560
rect 88710 192380 88890 192560
rect 89070 192380 96400 192560
rect 88400 192200 96400 192380
rect 88400 192020 88530 192200
rect 88710 192020 88890 192200
rect 89070 192020 96400 192200
rect 88400 191840 96400 192020
rect 88400 191660 88530 191840
rect 88710 191660 88890 191840
rect 89070 191660 96400 191840
rect 88400 191480 96400 191660
rect 88400 191300 88530 191480
rect 88710 191300 88890 191480
rect 89070 191300 96400 191480
rect 88400 191120 96400 191300
rect 88400 190940 88530 191120
rect 88710 190940 88890 191120
rect 89070 190940 96400 191120
rect 88400 190760 96400 190940
rect 88400 190580 88530 190760
rect 88710 190580 88890 190760
rect 89070 190580 96400 190760
rect 88400 190400 96400 190580
rect 88400 190220 88530 190400
rect 88710 190220 88890 190400
rect 89070 190220 96400 190400
rect 88400 190040 96400 190220
rect 88400 189860 88530 190040
rect 88710 189860 88890 190040
rect 89070 189860 96400 190040
rect 88400 189680 96400 189860
rect 88400 189500 88530 189680
rect 88710 189500 88890 189680
rect 89070 189500 96400 189680
rect 88400 189320 96400 189500
rect 88400 189140 88530 189320
rect 88710 189140 88890 189320
rect 89070 189140 96400 189320
rect 88400 188960 96400 189140
rect 88400 188780 88530 188960
rect 88710 188780 88890 188960
rect 89070 188780 96400 188960
rect 88400 188600 96400 188780
rect 88400 188420 88530 188600
rect 88710 188420 88890 188600
rect 89070 188420 96400 188600
rect 88400 188240 96400 188420
rect 88400 188060 88530 188240
rect 88710 188060 88890 188240
rect 89070 188060 96400 188240
rect 88400 187880 96400 188060
rect 88400 187700 88530 187880
rect 88710 187700 88890 187880
rect 89070 187700 96400 187880
rect 88400 187520 96400 187700
rect 88400 187340 88530 187520
rect 88710 187340 88890 187520
rect 89070 187340 96400 187520
rect 88400 187160 96400 187340
rect 88400 186980 88530 187160
rect 88710 186980 88890 187160
rect 89070 186980 96400 187160
rect 88400 186800 96400 186980
rect 88400 186620 88530 186800
rect 88710 186620 88890 186800
rect 89070 186620 96400 186800
rect 88400 186440 96400 186620
rect 88400 186260 88530 186440
rect 88710 186260 88890 186440
rect 89070 186260 96400 186440
rect 88400 186080 96400 186260
rect 88400 185900 88530 186080
rect 88710 185900 88890 186080
rect 89070 185900 96400 186080
rect 88400 185720 96400 185900
rect 88400 185540 88530 185720
rect 88710 185540 88890 185720
rect 89070 185540 96400 185720
rect 88400 185360 96400 185540
rect 88400 185180 88530 185360
rect 88710 185180 88890 185360
rect 89070 185180 96400 185360
rect 88400 185000 96400 185180
rect 88400 184820 88530 185000
rect 88710 184820 88890 185000
rect 89070 184820 96400 185000
rect 88400 184640 96400 184820
rect 88400 184460 88530 184640
rect 88710 184460 88890 184640
rect 89070 184460 96400 184640
rect 88400 184280 96400 184460
rect 88400 184100 88530 184280
rect 88710 184100 88890 184280
rect 89070 184100 96400 184280
rect 88400 183920 96400 184100
rect 88400 183740 88530 183920
rect 88710 183740 88890 183920
rect 89070 183740 96400 183920
rect 88400 183560 96400 183740
rect 88400 183380 88530 183560
rect 88710 183380 88890 183560
rect 89070 183380 96400 183560
rect 88400 183200 96400 183380
rect 287000 196570 290930 196750
rect 291110 196570 291290 196750
rect 291470 196570 291700 196750
rect 287000 196390 291700 196570
rect 287000 196210 290930 196390
rect 291110 196210 291290 196390
rect 291470 196210 291700 196390
rect 287000 196030 291700 196210
rect 287000 195850 290930 196030
rect 291110 195850 291290 196030
rect 291470 195850 291700 196030
rect 287000 195670 291700 195850
rect 287000 195490 290930 195670
rect 291110 195490 291290 195670
rect 291470 195490 291700 195670
rect 287000 195310 291700 195490
rect 287000 195130 290930 195310
rect 291110 195130 291290 195310
rect 291470 195130 291700 195310
rect 287000 194950 291700 195130
rect 287000 194770 290930 194950
rect 291110 194770 291290 194950
rect 291470 194770 291700 194950
rect 287000 194590 291700 194770
rect 287000 194410 290930 194590
rect 291110 194410 291290 194590
rect 291470 194410 291700 194590
rect 287000 194230 291700 194410
rect 287000 194050 290930 194230
rect 291110 194050 291290 194230
rect 291470 194050 291700 194230
rect 287000 193870 291700 194050
rect 287000 193690 290930 193870
rect 291110 193690 291290 193870
rect 291470 193690 291700 193870
rect 287000 193510 291700 193690
rect 287000 193330 290930 193510
rect 291110 193330 291290 193510
rect 291470 193330 291700 193510
rect 287000 193150 291700 193330
rect 287000 192970 290930 193150
rect 291110 192970 291290 193150
rect 291470 192970 291700 193150
rect 287000 192790 291700 192970
rect 287000 192610 290930 192790
rect 291110 192610 291290 192790
rect 291470 192610 291700 192790
rect 287000 192430 291700 192610
rect 287000 192250 290930 192430
rect 291110 192250 291290 192430
rect 291470 192250 291700 192430
rect 287000 192070 291700 192250
rect 287000 191890 290930 192070
rect 291110 191890 291290 192070
rect 291470 191890 291700 192070
rect 287000 191710 291700 191890
rect 287000 191530 290930 191710
rect 291110 191530 291290 191710
rect 291470 191530 291700 191710
rect 287000 191350 291700 191530
rect 287000 191170 290930 191350
rect 291110 191170 291290 191350
rect 291470 191170 291700 191350
rect 287000 190990 291700 191170
rect 287000 190810 290930 190990
rect 291110 190810 291290 190990
rect 291470 190810 291700 190990
rect 287000 190630 291700 190810
rect 287000 190450 290930 190630
rect 291110 190450 291290 190630
rect 291470 190450 291700 190630
rect 287000 190270 291700 190450
rect 287000 190090 290930 190270
rect 291110 190090 291290 190270
rect 291470 190090 291700 190270
rect 287000 189910 291700 190090
rect 287000 189730 290930 189910
rect 291110 189730 291290 189910
rect 291470 189730 291700 189910
rect 287000 189550 291700 189730
rect 287000 189370 290930 189550
rect 291110 189370 291290 189550
rect 291470 189370 291700 189550
rect 287000 189190 291700 189370
rect 287000 189010 290930 189190
rect 291110 189010 291290 189190
rect 291470 189010 291700 189190
rect 287000 188830 291700 189010
rect 287000 188650 290930 188830
rect 291110 188650 291290 188830
rect 291470 188650 291700 188830
rect 287000 188470 291700 188650
rect 287000 188290 290930 188470
rect 291110 188290 291290 188470
rect 291470 188290 291700 188470
rect 287000 188110 291700 188290
rect 287000 187930 290930 188110
rect 291110 187930 291290 188110
rect 291470 187930 291700 188110
rect 287000 187750 291700 187930
rect 287000 187570 290930 187750
rect 291110 187570 291290 187750
rect 291470 187570 291700 187750
rect 287000 187390 291700 187570
rect 287000 187210 290930 187390
rect 291110 187210 291290 187390
rect 291470 187210 291700 187390
rect 287000 187030 291700 187210
rect 287000 186850 290930 187030
rect 291110 186850 291290 187030
rect 291470 186850 291700 187030
rect 287000 186670 291700 186850
rect 287000 186490 290930 186670
rect 291110 186490 291290 186670
rect 291470 186490 291700 186670
rect 287000 186310 291700 186490
rect 287000 186130 290930 186310
rect 291110 186130 291290 186310
rect 291470 186130 291700 186310
rect 287000 185950 291700 186130
rect 287000 185770 290930 185950
rect 291110 185770 291290 185950
rect 291470 185770 291700 185950
rect 287000 185590 291700 185770
rect 287000 185410 290930 185590
rect 291110 185410 291290 185590
rect 291470 185410 291700 185590
rect 287000 185230 291700 185410
rect 287000 185050 290930 185230
rect 291110 185050 291290 185230
rect 291470 185050 291700 185230
rect 287000 184870 291700 185050
rect 287000 184690 290930 184870
rect 291110 184690 291290 184870
rect 291470 184690 291700 184870
rect 287000 184510 291700 184690
rect 287000 184330 290930 184510
rect 291110 184330 291290 184510
rect 291470 184330 291700 184510
rect 287000 184150 291700 184330
rect 287000 183970 290930 184150
rect 291110 183970 291290 184150
rect 291470 183970 291700 184150
rect 287000 183790 291700 183970
rect 287000 183610 290930 183790
rect 291110 183610 291290 183790
rect 291470 183610 291700 183790
rect 287000 183430 291700 183610
rect 287000 183250 290930 183430
rect 291110 183250 291290 183430
rect 291470 183250 291700 183430
rect 287000 183070 291700 183250
rect 287000 182890 290930 183070
rect 291110 182890 291290 183070
rect 291470 182890 291700 183070
rect 287000 182710 291700 182890
rect 287000 182530 290930 182710
rect 291110 182530 291290 182710
rect 291470 182530 291700 182710
rect 287000 182350 291700 182530
rect 287000 182170 290930 182350
rect 291110 182170 291290 182350
rect 291470 182170 291700 182350
rect 287000 181990 291700 182170
rect 287000 181810 290930 181990
rect 291110 181810 291290 181990
rect 291470 181810 291700 181990
rect 287000 181630 291700 181810
rect 287000 181450 290930 181630
rect 291110 181450 291290 181630
rect 291470 181450 291700 181630
rect 287000 181270 291700 181450
rect 287000 181090 290930 181270
rect 291110 181090 291290 181270
rect 291470 181090 291700 181270
rect 287000 180910 291700 181090
rect 287000 180730 290930 180910
rect 291110 180730 291290 180910
rect 291470 180730 291700 180910
rect 287000 180600 291700 180730
<< m2contact >>
rect 290930 199090 291110 199270
rect 291290 199090 291470 199270
rect 290930 198730 291110 198910
rect 291290 198730 291470 198910
rect 290930 198370 291110 198550
rect 291290 198370 291470 198550
rect 290930 198010 291110 198190
rect 291290 198010 291470 198190
rect 290930 197650 291110 197830
rect 291290 197650 291470 197830
rect 290930 197290 291110 197470
rect 291290 197290 291470 197470
rect 290930 196930 291110 197110
rect 291290 196930 291470 197110
rect 88530 196340 88710 196520
rect 88890 196340 89070 196520
rect 88530 195980 88710 196160
rect 88890 195980 89070 196160
rect 88530 195620 88710 195800
rect 88890 195620 89070 195800
rect 88530 195260 88710 195440
rect 88890 195260 89070 195440
rect 88530 194900 88710 195080
rect 88890 194900 89070 195080
rect 88530 194540 88710 194720
rect 88890 194540 89070 194720
rect 88530 194180 88710 194360
rect 88890 194180 89070 194360
rect 88530 193820 88710 194000
rect 88890 193820 89070 194000
rect 88530 193460 88710 193640
rect 88890 193460 89070 193640
rect 88530 193100 88710 193280
rect 88890 193100 89070 193280
rect 88530 192740 88710 192920
rect 88890 192740 89070 192920
rect 88530 192380 88710 192560
rect 88890 192380 89070 192560
rect 88530 192020 88710 192200
rect 88890 192020 89070 192200
rect 88530 191660 88710 191840
rect 88890 191660 89070 191840
rect 88530 191300 88710 191480
rect 88890 191300 89070 191480
rect 88530 190940 88710 191120
rect 88890 190940 89070 191120
rect 88530 190580 88710 190760
rect 88890 190580 89070 190760
rect 88530 190220 88710 190400
rect 88890 190220 89070 190400
rect 88530 189860 88710 190040
rect 88890 189860 89070 190040
rect 88530 189500 88710 189680
rect 88890 189500 89070 189680
rect 88530 189140 88710 189320
rect 88890 189140 89070 189320
rect 88530 188780 88710 188960
rect 88890 188780 89070 188960
rect 88530 188420 88710 188600
rect 88890 188420 89070 188600
rect 88530 188060 88710 188240
rect 88890 188060 89070 188240
rect 88530 187700 88710 187880
rect 88890 187700 89070 187880
rect 88530 187340 88710 187520
rect 88890 187340 89070 187520
rect 88530 186980 88710 187160
rect 88890 186980 89070 187160
rect 88530 186620 88710 186800
rect 88890 186620 89070 186800
rect 88530 186260 88710 186440
rect 88890 186260 89070 186440
rect 88530 185900 88710 186080
rect 88890 185900 89070 186080
rect 88530 185540 88710 185720
rect 88890 185540 89070 185720
rect 88530 185180 88710 185360
rect 88890 185180 89070 185360
rect 88530 184820 88710 185000
rect 88890 184820 89070 185000
rect 88530 184460 88710 184640
rect 88890 184460 89070 184640
rect 88530 184100 88710 184280
rect 88890 184100 89070 184280
rect 88530 183740 88710 183920
rect 88890 183740 89070 183920
rect 88530 183380 88710 183560
rect 88890 183380 89070 183560
rect 290930 196570 291110 196750
rect 291290 196570 291470 196750
rect 290930 196210 291110 196390
rect 291290 196210 291470 196390
rect 290930 195850 291110 196030
rect 291290 195850 291470 196030
rect 290930 195490 291110 195670
rect 291290 195490 291470 195670
rect 290930 195130 291110 195310
rect 291290 195130 291470 195310
rect 290930 194770 291110 194950
rect 291290 194770 291470 194950
rect 290930 194410 291110 194590
rect 291290 194410 291470 194590
rect 290930 194050 291110 194230
rect 291290 194050 291470 194230
rect 290930 193690 291110 193870
rect 291290 193690 291470 193870
rect 290930 193330 291110 193510
rect 291290 193330 291470 193510
rect 290930 192970 291110 193150
rect 291290 192970 291470 193150
rect 290930 192610 291110 192790
rect 291290 192610 291470 192790
rect 290930 192250 291110 192430
rect 291290 192250 291470 192430
rect 290930 191890 291110 192070
rect 291290 191890 291470 192070
rect 290930 191530 291110 191710
rect 291290 191530 291470 191710
rect 290930 191170 291110 191350
rect 291290 191170 291470 191350
rect 290930 190810 291110 190990
rect 291290 190810 291470 190990
rect 290930 190450 291110 190630
rect 291290 190450 291470 190630
rect 290930 190090 291110 190270
rect 291290 190090 291470 190270
rect 290930 189730 291110 189910
rect 291290 189730 291470 189910
rect 290930 189370 291110 189550
rect 291290 189370 291470 189550
rect 290930 189010 291110 189190
rect 291290 189010 291470 189190
rect 290930 188650 291110 188830
rect 291290 188650 291470 188830
rect 290930 188290 291110 188470
rect 291290 188290 291470 188470
rect 290930 187930 291110 188110
rect 291290 187930 291470 188110
rect 290930 187570 291110 187750
rect 291290 187570 291470 187750
rect 290930 187210 291110 187390
rect 291290 187210 291470 187390
rect 290930 186850 291110 187030
rect 291290 186850 291470 187030
rect 290930 186490 291110 186670
rect 291290 186490 291470 186670
rect 290930 186130 291110 186310
rect 291290 186130 291470 186310
rect 290930 185770 291110 185950
rect 291290 185770 291470 185950
rect 290930 185410 291110 185590
rect 291290 185410 291470 185590
rect 290930 185050 291110 185230
rect 291290 185050 291470 185230
rect 290930 184690 291110 184870
rect 291290 184690 291470 184870
rect 290930 184330 291110 184510
rect 291290 184330 291470 184510
rect 290930 183970 291110 184150
rect 291290 183970 291470 184150
rect 290930 183610 291110 183790
rect 291290 183610 291470 183790
rect 290930 183250 291110 183430
rect 291290 183250 291470 183430
rect 290930 182890 291110 183070
rect 291290 182890 291470 183070
rect 290930 182530 291110 182710
rect 291290 182530 291470 182710
rect 290930 182170 291110 182350
rect 291290 182170 291470 182350
rect 290930 181810 291110 181990
rect 291290 181810 291470 181990
rect 290930 181450 291110 181630
rect 291290 181450 291470 181630
rect 290930 181090 291110 181270
rect 291290 181090 291470 181270
rect 290930 180730 291110 180910
rect 291290 180730 291470 180910
<< metal2 >>
rect 119600 291400 120400 291800
rect 94200 290600 120400 291400
rect 88200 259600 93600 260400
rect 88200 232600 92400 233400
rect 88200 227200 91200 228000
rect 90600 211350 91200 227200
rect 91800 217350 92400 232600
rect 93000 232950 93600 259600
rect 94200 237550 94800 290600
rect 146600 289800 147200 291800
rect 114000 289000 147200 289800
rect 114000 286000 114800 289000
rect 173600 288200 174400 291800
rect 127200 287400 174400 288200
rect 127200 286000 128000 287400
rect 200600 286600 201400 291800
rect 227600 291400 228400 291800
rect 154200 285800 201400 286600
rect 217200 290800 228400 291400
rect 217200 285800 217800 290800
rect 254600 290200 255400 291800
rect 221400 289600 255400 290200
rect 221400 286000 222000 289600
rect 281600 289000 282300 291800
rect 228600 288300 282300 289000
rect 228600 285800 229400 288300
rect 230400 286900 291200 287600
rect 230400 285800 231100 286900
rect 236500 285800 290100 286500
rect 94200 237370 94410 237550
rect 94590 237370 94800 237550
rect 94200 237190 94800 237370
rect 94200 237010 94410 237190
rect 94590 237010 94800 237190
rect 94200 236830 94800 237010
rect 94200 236650 94410 236830
rect 94590 236650 94800 236830
rect 94200 236400 94800 236650
rect 288400 259650 289000 259800
rect 288400 259470 288610 259650
rect 288790 259470 289000 259650
rect 288400 259290 289000 259470
rect 288400 259110 288610 259290
rect 288790 259110 289000 259290
rect 288400 258930 289000 259110
rect 288400 258750 288610 258930
rect 288790 258750 289000 258930
rect 93000 232770 93210 232950
rect 93390 232770 93600 232950
rect 93000 232590 93600 232770
rect 93000 232410 93210 232590
rect 93390 232410 93600 232590
rect 93000 232230 93600 232410
rect 93000 232050 93210 232230
rect 93390 232050 93600 232230
rect 93000 231800 93600 232050
rect 91800 217170 92010 217350
rect 92190 217170 92400 217350
rect 91800 216990 92400 217170
rect 91800 216810 92010 216990
rect 92190 216810 92400 216990
rect 91800 216630 92400 216810
rect 91800 216450 92010 216630
rect 92190 216450 92400 216630
rect 91800 216200 92400 216450
rect 90600 211170 90810 211350
rect 90990 211170 91200 211350
rect 90600 210990 91200 211170
rect 90600 210810 90810 210990
rect 90990 210810 91200 210990
rect 90600 210630 91200 210810
rect 90600 210450 90810 210630
rect 90990 210450 91200 210630
rect 90600 210200 91200 210450
rect 288400 206400 289000 258750
rect 289500 233400 290100 285800
rect 290600 260400 291200 286900
rect 290600 259700 291800 260400
rect 289500 232800 291800 233400
rect 288400 205700 291700 206400
rect 290700 199270 291700 199400
rect 290700 199090 290930 199270
rect 291110 199090 291290 199270
rect 291470 199090 291700 199270
rect 290700 198910 291700 199090
rect 290700 198730 290930 198910
rect 291110 198730 291290 198910
rect 291470 198730 291700 198910
rect 290700 198550 291700 198730
rect 290700 198370 290930 198550
rect 291110 198370 291290 198550
rect 291470 198370 291700 198550
rect 290700 198190 291700 198370
rect 290700 198010 290930 198190
rect 291110 198010 291290 198190
rect 291470 198010 291700 198190
rect 290700 197830 291700 198010
rect 290700 197650 290930 197830
rect 291110 197650 291290 197830
rect 291470 197650 291700 197830
rect 290700 197470 291700 197650
rect 290700 197290 290930 197470
rect 291110 197290 291290 197470
rect 291470 197290 291700 197470
rect 290700 197110 291700 197290
rect 290700 196930 290930 197110
rect 291110 196930 291290 197110
rect 291470 196930 291700 197110
rect 290700 196750 291700 196930
rect 88400 196520 89200 196700
rect 88400 196340 88530 196520
rect 88710 196340 88890 196520
rect 89070 196340 89200 196520
rect 88400 196160 89200 196340
rect 88400 195980 88530 196160
rect 88710 195980 88890 196160
rect 89070 195980 89200 196160
rect 88400 195800 89200 195980
rect 88400 195620 88530 195800
rect 88710 195620 88890 195800
rect 89070 195620 89200 195800
rect 88400 195440 89200 195620
rect 88400 195260 88530 195440
rect 88710 195260 88890 195440
rect 89070 195260 89200 195440
rect 88400 195080 89200 195260
rect 88400 194900 88530 195080
rect 88710 194900 88890 195080
rect 89070 194900 89200 195080
rect 88400 194720 89200 194900
rect 88400 194540 88530 194720
rect 88710 194540 88890 194720
rect 89070 194540 89200 194720
rect 88400 194360 89200 194540
rect 88400 194180 88530 194360
rect 88710 194180 88890 194360
rect 89070 194180 89200 194360
rect 88400 194000 89200 194180
rect 88400 193820 88530 194000
rect 88710 193820 88890 194000
rect 89070 193820 89200 194000
rect 88400 193640 89200 193820
rect 88400 193460 88530 193640
rect 88710 193460 88890 193640
rect 89070 193460 89200 193640
rect 88400 193280 89200 193460
rect 88400 193100 88530 193280
rect 88710 193100 88890 193280
rect 89070 193100 89200 193280
rect 88400 192920 89200 193100
rect 88400 192740 88530 192920
rect 88710 192740 88890 192920
rect 89070 192740 89200 192920
rect 88400 192560 89200 192740
rect 88400 192380 88530 192560
rect 88710 192380 88890 192560
rect 89070 192380 89200 192560
rect 88400 192200 89200 192380
rect 88400 192020 88530 192200
rect 88710 192020 88890 192200
rect 89070 192020 89200 192200
rect 88400 191840 89200 192020
rect 88400 191660 88530 191840
rect 88710 191660 88890 191840
rect 89070 191660 89200 191840
rect 88400 191480 89200 191660
rect 88400 191300 88530 191480
rect 88710 191300 88890 191480
rect 89070 191300 89200 191480
rect 88400 191120 89200 191300
rect 88400 190940 88530 191120
rect 88710 190940 88890 191120
rect 89070 190940 89200 191120
rect 88400 190760 89200 190940
rect 88400 190580 88530 190760
rect 88710 190580 88890 190760
rect 89070 190580 89200 190760
rect 88400 190400 89200 190580
rect 88400 190220 88530 190400
rect 88710 190220 88890 190400
rect 89070 190220 89200 190400
rect 88400 190040 89200 190220
rect 88400 189860 88530 190040
rect 88710 189860 88890 190040
rect 89070 189860 89200 190040
rect 88400 189680 89200 189860
rect 88400 189500 88530 189680
rect 88710 189500 88890 189680
rect 89070 189500 89200 189680
rect 88400 189320 89200 189500
rect 88400 189140 88530 189320
rect 88710 189140 88890 189320
rect 89070 189140 89200 189320
rect 88400 188960 89200 189140
rect 88400 188780 88530 188960
rect 88710 188780 88890 188960
rect 89070 188780 89200 188960
rect 88400 188600 89200 188780
rect 88400 188420 88530 188600
rect 88710 188420 88890 188600
rect 89070 188420 89200 188600
rect 88400 188240 89200 188420
rect 88400 188060 88530 188240
rect 88710 188060 88890 188240
rect 89070 188060 89200 188240
rect 88400 187880 89200 188060
rect 88400 187700 88530 187880
rect 88710 187700 88890 187880
rect 89070 187700 89200 187880
rect 88400 187520 89200 187700
rect 88400 187340 88530 187520
rect 88710 187340 88890 187520
rect 89070 187340 89200 187520
rect 88400 187160 89200 187340
rect 88400 186980 88530 187160
rect 88710 186980 88890 187160
rect 89070 186980 89200 187160
rect 88400 186800 89200 186980
rect 88400 186620 88530 186800
rect 88710 186620 88890 186800
rect 89070 186620 89200 186800
rect 88400 186440 89200 186620
rect 88400 186260 88530 186440
rect 88710 186260 88890 186440
rect 89070 186260 89200 186440
rect 88400 186080 89200 186260
rect 88400 185900 88530 186080
rect 88710 185900 88890 186080
rect 89070 185900 89200 186080
rect 88400 185720 89200 185900
rect 88400 185540 88530 185720
rect 88710 185540 88890 185720
rect 89070 185540 89200 185720
rect 88400 185360 89200 185540
rect 88400 185180 88530 185360
rect 88710 185180 88890 185360
rect 89070 185180 89200 185360
rect 88400 185000 89200 185180
rect 88400 184820 88530 185000
rect 88710 184820 88890 185000
rect 89070 184820 89200 185000
rect 88400 184640 89200 184820
rect 88400 184460 88530 184640
rect 88710 184460 88890 184640
rect 89070 184460 89200 184640
rect 88400 184280 89200 184460
rect 88400 184100 88530 184280
rect 88710 184100 88890 184280
rect 89070 184100 89200 184280
rect 88400 183920 89200 184100
rect 88400 183740 88530 183920
rect 88710 183740 88890 183920
rect 89070 183740 89200 183920
rect 88400 183560 89200 183740
rect 88400 183380 88530 183560
rect 88710 183380 88890 183560
rect 89070 183380 89200 183560
rect 88400 183200 89200 183380
rect 290700 196570 290930 196750
rect 291110 196570 291290 196750
rect 291470 196570 291700 196750
rect 290700 196390 291700 196570
rect 290700 196210 290930 196390
rect 291110 196210 291290 196390
rect 291470 196210 291700 196390
rect 290700 196030 291700 196210
rect 290700 195850 290930 196030
rect 291110 195850 291290 196030
rect 291470 195850 291700 196030
rect 290700 195670 291700 195850
rect 290700 195490 290930 195670
rect 291110 195490 291290 195670
rect 291470 195490 291700 195670
rect 290700 195310 291700 195490
rect 290700 195130 290930 195310
rect 291110 195130 291290 195310
rect 291470 195130 291700 195310
rect 290700 194950 291700 195130
rect 290700 194770 290930 194950
rect 291110 194770 291290 194950
rect 291470 194770 291700 194950
rect 290700 194590 291700 194770
rect 290700 194410 290930 194590
rect 291110 194410 291290 194590
rect 291470 194410 291700 194590
rect 290700 194230 291700 194410
rect 290700 194050 290930 194230
rect 291110 194050 291290 194230
rect 291470 194050 291700 194230
rect 290700 193870 291700 194050
rect 290700 193690 290930 193870
rect 291110 193690 291290 193870
rect 291470 193690 291700 193870
rect 290700 193510 291700 193690
rect 290700 193330 290930 193510
rect 291110 193330 291290 193510
rect 291470 193330 291700 193510
rect 290700 193150 291700 193330
rect 290700 192970 290930 193150
rect 291110 192970 291290 193150
rect 291470 192970 291700 193150
rect 290700 192790 291700 192970
rect 290700 192610 290930 192790
rect 291110 192610 291290 192790
rect 291470 192610 291700 192790
rect 290700 192430 291700 192610
rect 290700 192250 290930 192430
rect 291110 192250 291290 192430
rect 291470 192250 291700 192430
rect 290700 192070 291700 192250
rect 290700 191890 290930 192070
rect 291110 191890 291290 192070
rect 291470 191890 291700 192070
rect 290700 191710 291700 191890
rect 290700 191530 290930 191710
rect 291110 191530 291290 191710
rect 291470 191530 291700 191710
rect 290700 191350 291700 191530
rect 290700 191170 290930 191350
rect 291110 191170 291290 191350
rect 291470 191170 291700 191350
rect 290700 190990 291700 191170
rect 290700 190810 290930 190990
rect 291110 190810 291290 190990
rect 291470 190810 291700 190990
rect 290700 190630 291700 190810
rect 290700 190450 290930 190630
rect 291110 190450 291290 190630
rect 291470 190450 291700 190630
rect 290700 190270 291700 190450
rect 290700 190090 290930 190270
rect 291110 190090 291290 190270
rect 291470 190090 291700 190270
rect 290700 189910 291700 190090
rect 290700 189730 290930 189910
rect 291110 189730 291290 189910
rect 291470 189730 291700 189910
rect 290700 189550 291700 189730
rect 290700 189370 290930 189550
rect 291110 189370 291290 189550
rect 291470 189370 291700 189550
rect 290700 189190 291700 189370
rect 290700 189010 290930 189190
rect 291110 189010 291290 189190
rect 291470 189010 291700 189190
rect 290700 188830 291700 189010
rect 290700 188650 290930 188830
rect 291110 188650 291290 188830
rect 291470 188650 291700 188830
rect 290700 188470 291700 188650
rect 290700 188290 290930 188470
rect 291110 188290 291290 188470
rect 291470 188290 291700 188470
rect 290700 188110 291700 188290
rect 290700 187930 290930 188110
rect 291110 187930 291290 188110
rect 291470 187930 291700 188110
rect 290700 187750 291700 187930
rect 290700 187570 290930 187750
rect 291110 187570 291290 187750
rect 291470 187570 291700 187750
rect 290700 187390 291700 187570
rect 290700 187210 290930 187390
rect 291110 187210 291290 187390
rect 291470 187210 291700 187390
rect 290700 187030 291700 187210
rect 290700 186850 290930 187030
rect 291110 186850 291290 187030
rect 291470 186850 291700 187030
rect 290700 186670 291700 186850
rect 290700 186490 290930 186670
rect 291110 186490 291290 186670
rect 291470 186490 291700 186670
rect 290700 186310 291700 186490
rect 290700 186130 290930 186310
rect 291110 186130 291290 186310
rect 291470 186130 291700 186310
rect 290700 185950 291700 186130
rect 290700 185770 290930 185950
rect 291110 185770 291290 185950
rect 291470 185770 291700 185950
rect 290700 185590 291700 185770
rect 290700 185410 290930 185590
rect 291110 185410 291290 185590
rect 291470 185410 291700 185590
rect 290700 185230 291700 185410
rect 290700 185050 290930 185230
rect 291110 185050 291290 185230
rect 291470 185050 291700 185230
rect 290700 184870 291700 185050
rect 290700 184690 290930 184870
rect 291110 184690 291290 184870
rect 291470 184690 291700 184870
rect 290700 184510 291700 184690
rect 290700 184330 290930 184510
rect 291110 184330 291290 184510
rect 291470 184330 291700 184510
rect 290700 184150 291700 184330
rect 290700 183970 290930 184150
rect 291110 183970 291290 184150
rect 291470 183970 291700 184150
rect 290700 183790 291700 183970
rect 290700 183610 290930 183790
rect 291110 183610 291290 183790
rect 291470 183610 291700 183790
rect 290700 183430 291700 183610
rect 290700 183250 290930 183430
rect 291110 183250 291290 183430
rect 291470 183250 291700 183430
rect 290700 183070 291700 183250
rect 290700 182890 290930 183070
rect 291110 182890 291290 183070
rect 291470 182890 291700 183070
rect 290700 182710 291700 182890
rect 290700 182530 290930 182710
rect 291110 182530 291290 182710
rect 291470 182530 291700 182710
rect 290700 182350 291700 182530
rect 290700 182170 290930 182350
rect 291110 182170 291290 182350
rect 291470 182170 291700 182350
rect 290700 181990 291700 182170
rect 290700 181810 290930 181990
rect 291110 181810 291290 181990
rect 291470 181810 291700 181990
rect 290700 181630 291700 181810
rect 290700 181450 290930 181630
rect 291110 181450 291290 181630
rect 291470 181450 291700 181630
rect 290700 181270 291700 181450
rect 290700 181090 290930 181270
rect 291110 181090 291290 181270
rect 291470 181090 291700 181270
rect 290700 180910 291700 181090
rect 290700 180730 290930 180910
rect 291110 180730 291290 180910
rect 291470 180730 291700 180910
rect 290700 180600 291700 180730
rect 92300 179150 92900 179400
rect 92300 178970 92510 179150
rect 92690 178970 92900 179150
rect 92300 178790 92900 178970
rect 92300 178610 92510 178790
rect 92690 178610 92900 178790
rect 92300 178430 92900 178610
rect 92300 178250 92510 178430
rect 92690 178250 92900 178430
rect 90600 171480 91200 171600
rect 90600 171300 90810 171480
rect 90990 171300 91200 171480
rect 90600 171120 91200 171300
rect 90600 170940 90810 171120
rect 90990 170940 91200 171120
rect 90600 170760 91200 170940
rect 90600 170580 90810 170760
rect 90990 170580 91200 170760
rect 90600 170400 91200 170580
rect 90600 170220 90810 170400
rect 90990 170220 91200 170400
rect 90600 152400 91200 170220
rect 88200 151600 91200 152400
rect 92300 147000 92900 178250
rect 88200 146200 92900 147000
rect 93800 177450 94400 177700
rect 93800 177270 94010 177450
rect 94190 177270 94400 177450
rect 93800 177090 94400 177270
rect 93800 176910 94010 177090
rect 94190 176910 94400 177090
rect 93800 176730 94400 176910
rect 93800 176550 94010 176730
rect 94190 176550 94400 176730
rect 93800 120000 94400 176550
rect 88200 119200 94400 120000
rect 99600 89500 100200 96500
rect 102100 91903 102700 96400
rect 102098 91900 102700 91903
rect 102100 90703 102700 91900
rect 104500 91903 105100 96400
rect 108100 93103 108700 96400
rect 117000 94303 117600 96400
rect 132100 95503 132700 96400
rect 132100 95500 232900 95503
rect 132100 94900 233708 95500
rect 117000 93700 206700 94303
rect 108096 93100 179700 93103
rect 108100 92500 179700 93100
rect 104500 91300 152700 91903
rect 102100 90100 125700 90703
rect 98000 88886 100200 89500
rect 98000 88300 98700 88886
rect 125000 88300 125700 90100
rect 152000 88300 152700 91300
rect 179000 88300 179700 92500
rect 206000 88300 206700 93700
rect 233000 89002 233708 94900
rect 232994 88876 233708 89002
rect 232994 88294 233703 88876
<< m3contact >>
rect 94410 237370 94590 237550
rect 94410 237010 94590 237190
rect 94410 236650 94590 236830
rect 288610 259470 288790 259650
rect 288610 259110 288790 259290
rect 288610 258750 288790 258930
rect 93210 232770 93390 232950
rect 93210 232410 93390 232590
rect 93210 232050 93390 232230
rect 92010 217170 92190 217350
rect 92010 216810 92190 216990
rect 92010 216450 92190 216630
rect 90810 211170 90990 211350
rect 90810 210810 90990 210990
rect 90810 210450 90990 210630
rect 92510 178970 92690 179150
rect 92510 178610 92690 178790
rect 92510 178250 92690 178430
rect 90810 171300 90990 171480
rect 90810 170940 90990 171120
rect 90810 170580 90990 170760
rect 90810 170220 90990 170400
rect 94010 177270 94190 177450
rect 94010 176910 94190 177090
rect 94010 176550 94190 176730
<< metal3 >>
rect 288400 259720 289000 259800
rect 284980 259650 289000 259720
rect 284980 259480 288610 259650
rect 288400 259470 288610 259480
rect 288790 259470 289000 259650
rect 288400 259290 289000 259470
rect 288400 259110 288610 259290
rect 288790 259110 289000 259290
rect 288400 258930 289000 259110
rect 288400 258750 288610 258930
rect 288790 258750 289000 258930
rect 288400 258600 289000 258750
rect 94200 237550 94800 237800
rect 94200 237370 94410 237550
rect 94590 237370 94800 237550
rect 94200 237190 94800 237370
rect 94200 237010 94410 237190
rect 94590 237010 94800 237190
rect 94200 236830 94800 237010
rect 94200 236650 94410 236830
rect 94590 236680 94800 236830
rect 94590 236650 98520 236680
rect 94200 236440 98520 236650
rect 94200 236400 94800 236440
rect 93000 232950 93600 233200
rect 93000 232770 93210 232950
rect 93390 232770 93600 232950
rect 93000 232590 93600 232770
rect 93000 232410 93210 232590
rect 93390 232410 93600 232590
rect 93000 232230 93600 232410
rect 93000 232050 93210 232230
rect 93390 232120 93600 232230
rect 93390 232050 98320 232120
rect 93000 231880 98320 232050
rect 93000 231800 93600 231880
rect 91800 217350 92400 217600
rect 91800 217170 92010 217350
rect 92190 217170 92400 217350
rect 91800 216990 92400 217170
rect 91800 216810 92010 216990
rect 92190 216810 92400 216990
rect 91800 216630 92400 216810
rect 91800 216450 92010 216630
rect 92190 216520 92400 216630
rect 92190 216450 98520 216520
rect 91800 216280 98520 216450
rect 91800 216200 92400 216280
rect 90600 211350 91200 211600
rect 90600 211170 90810 211350
rect 90990 211170 91200 211350
rect 90600 210990 91200 211170
rect 90600 210810 90810 210990
rect 90990 210810 91200 210990
rect 90600 210630 91200 210810
rect 90600 210450 90810 210630
rect 90990 210520 91200 210630
rect 90990 210450 98320 210520
rect 90600 210280 98320 210450
rect 90600 210200 91200 210280
rect 92300 179320 92900 179400
rect 92300 179150 98720 179320
rect 92300 178970 92510 179150
rect 92690 179080 98720 179150
rect 92690 178970 92900 179080
rect 92300 178790 92900 178970
rect 92300 178610 92510 178790
rect 92690 178610 92900 178790
rect 92300 178430 92900 178610
rect 92300 178250 92510 178430
rect 92690 178250 92900 178430
rect 92300 178000 92900 178250
rect 93800 177580 94400 177700
rect 93800 177450 97320 177580
rect 93800 177270 94010 177450
rect 94190 177340 97320 177450
rect 94190 177270 94400 177340
rect 93800 177090 94400 177270
rect 93800 176910 94010 177090
rect 94190 176910 94400 177090
rect 93800 176730 94400 176910
rect 93800 176550 94010 176730
rect 94190 176550 94400 176730
rect 93800 176300 94400 176550
rect 90600 171480 97000 171600
rect 90600 171300 90810 171480
rect 90990 171300 97000 171480
rect 90600 171200 97000 171300
rect 90600 171120 91200 171200
rect 90600 170940 90810 171120
rect 90990 170940 91200 171120
rect 90600 170760 91200 170940
rect 90600 170580 90810 170760
rect 90990 170580 91200 170760
rect 90600 170400 91200 170580
rect 90600 170220 90810 170400
rect 90990 170220 91200 170400
rect 90600 170100 91200 170220
<< comment >>
rect 0 0 380000 380000
<< end >>
