magic
tech scmos
magscale 1 2
timestamp 1709017741
<< error_s >>
rect 4 6244 6236 6256
rect 4 5984 6236 5996
rect 4 5724 6236 5736
rect 4 5464 6236 5476
rect 4 5204 6236 5216
rect 4 4944 6236 4956
rect 4 4684 6236 4696
rect 4 4424 6236 4436
rect 4 4164 6236 4176
rect 4 3904 6236 3916
rect 4 3644 6236 3656
rect 4 3384 6236 3396
rect 4 3124 6236 3136
rect 4 2864 6236 2876
rect 4 2604 6236 2616
rect 4 2344 6236 2356
rect 4 2084 6236 2096
rect 4 1824 6236 1836
rect 4 1564 6236 1576
rect 4 1304 6236 1316
rect 4 1044 6236 1056
rect 4 784 6236 796
rect 4 524 6236 536
rect 4 264 6236 276
rect 4 4 6236 16
<< nwell >>
rect 5873 5676 5889 5684
<< metal1 >>
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 2827 6173 2833 6187
rect 2067 6137 2193 6143
rect 2627 6137 2673 6143
rect 2980 6123 2993 6127
rect 2977 6113 2993 6123
rect 5327 6117 5353 6123
rect 2977 6087 2983 6113
rect 1977 6080 2013 6083
rect 1973 6077 2013 6080
rect 1973 6067 1987 6077
rect 2967 6077 2983 6087
rect 2967 6073 2980 6077
rect 3747 6057 3833 6063
rect 3887 6057 3933 6063
rect 5587 6057 5653 6063
rect 3387 6017 3413 6023
rect 6243 5998 6303 6258
rect 6210 5982 6303 5998
rect 2327 5937 2373 5943
rect 1987 5917 2013 5923
rect 3497 5897 3533 5903
rect 3497 5863 3503 5897
rect 3967 5897 3993 5903
rect 5027 5903 5040 5907
rect 5027 5893 5043 5903
rect 5167 5903 5180 5907
rect 5920 5903 5933 5907
rect 5167 5893 5183 5903
rect 3477 5857 3503 5863
rect 527 5837 613 5843
rect 2167 5837 2193 5843
rect 3477 5843 3483 5857
rect 3427 5837 3483 5843
rect 4647 5837 4693 5843
rect 5037 5843 5043 5893
rect 5037 5837 5093 5843
rect 5177 5846 5183 5893
rect 5917 5893 5933 5903
rect 6047 5903 6060 5907
rect 6047 5893 6063 5903
rect 5917 5867 5923 5893
rect 5917 5857 5933 5867
rect 5920 5853 5933 5857
rect 6057 5863 6063 5893
rect 6057 5857 6083 5863
rect 6077 5843 6083 5857
rect 6027 5837 6133 5843
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 87 5617 113 5623
rect 187 5617 233 5623
rect 3227 5617 3263 5623
rect 467 5603 480 5607
rect 880 5603 893 5607
rect 467 5593 483 5603
rect 477 5547 483 5593
rect 877 5593 893 5603
rect 1317 5597 1353 5603
rect 877 5567 883 5593
rect 1317 5567 1323 5597
rect 1480 5603 1493 5607
rect 1477 5593 1493 5603
rect 2697 5597 2733 5603
rect 877 5557 893 5567
rect 880 5553 893 5557
rect 1307 5557 1323 5567
rect 1307 5553 1320 5557
rect 627 5537 673 5543
rect 1477 5543 1483 5593
rect 2697 5567 2703 5597
rect 3140 5603 3153 5607
rect 3137 5593 3153 5603
rect 3257 5603 3263 5617
rect 4080 5603 4093 5607
rect 3257 5597 3283 5603
rect 2687 5557 2703 5567
rect 3137 5567 3143 5593
rect 3137 5557 3153 5567
rect 2687 5553 2700 5557
rect 3140 5553 3153 5557
rect 3277 5563 3283 5597
rect 4077 5593 4093 5603
rect 5687 5597 5713 5603
rect 4077 5567 4083 5593
rect 3277 5560 3303 5563
rect 3277 5557 3307 5560
rect 4077 5557 4093 5567
rect 3293 5547 3307 5557
rect 4080 5553 4093 5557
rect 1427 5537 1483 5543
rect 2247 5537 2333 5543
rect 3527 5537 3553 5543
rect 6243 5478 6303 5982
rect 6210 5462 6303 5478
rect 337 5397 373 5403
rect 337 5343 343 5397
rect 733 5383 747 5393
rect 1377 5397 1413 5403
rect 1377 5383 1383 5397
rect 1627 5397 1653 5403
rect 3157 5397 3233 5403
rect 717 5380 747 5383
rect 717 5377 743 5380
rect 1357 5377 1383 5383
rect 717 5347 723 5377
rect 337 5337 363 5343
rect 357 5327 363 5337
rect 707 5337 723 5347
rect 1357 5347 1363 5377
rect 1967 5383 1980 5387
rect 2000 5383 2013 5387
rect 1967 5373 1983 5383
rect 1977 5347 1983 5373
rect 1357 5337 1373 5347
rect 707 5333 720 5337
rect 1360 5333 1373 5337
rect 1967 5337 1983 5347
rect 1997 5373 2013 5383
rect 2567 5377 2593 5383
rect 1997 5343 2003 5373
rect 3157 5347 3163 5397
rect 3487 5397 3553 5403
rect 4967 5397 5013 5403
rect 6127 5397 6193 5403
rect 3360 5383 3373 5387
rect 1997 5337 2023 5343
rect 1967 5333 1980 5337
rect 67 5317 93 5323
rect 357 5317 373 5327
rect 360 5313 373 5317
rect 1627 5317 1653 5323
rect 1827 5317 1873 5323
rect 2017 5323 2023 5337
rect 3147 5337 3163 5347
rect 3357 5373 3373 5383
rect 3497 5377 3533 5383
rect 3357 5347 3363 5373
rect 3497 5347 3503 5377
rect 3357 5337 3373 5347
rect 3147 5333 3160 5337
rect 3360 5333 3373 5337
rect 3487 5337 3503 5347
rect 4077 5347 4083 5393
rect 4187 5383 4200 5387
rect 4480 5383 4493 5387
rect 4187 5373 4203 5383
rect 4077 5337 4093 5347
rect 3487 5333 3500 5337
rect 4080 5333 4093 5337
rect 4197 5343 4203 5373
rect 4477 5373 4493 5383
rect 4477 5347 4483 5373
rect 4197 5337 4233 5343
rect 4467 5337 4483 5347
rect 4467 5333 4480 5337
rect 2017 5317 2053 5323
rect 3407 5313 3413 5327
rect 3487 5317 3553 5323
rect 3647 5317 3693 5323
rect 4207 5317 4253 5323
rect 1667 5297 1693 5303
rect 4587 5297 4633 5303
rect 3487 5257 3533 5263
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 953 5123 967 5133
rect 953 5120 993 5123
rect 957 5117 993 5120
rect 4327 5117 4353 5123
rect 4707 5117 4733 5123
rect 5507 5117 5613 5123
rect 1087 5097 1113 5103
rect 1587 5097 1713 5103
rect 1333 5083 1347 5093
rect 1813 5083 1827 5093
rect 1333 5080 1363 5083
rect 1337 5077 1363 5080
rect 1357 5047 1363 5077
rect 1797 5080 1827 5083
rect 1957 5097 1993 5103
rect 1797 5077 1823 5080
rect 1797 5047 1803 5077
rect 1357 5037 1373 5047
rect 1360 5033 1373 5037
rect 1797 5037 1813 5047
rect 1800 5033 1813 5037
rect 1920 5043 1933 5047
rect 1917 5033 1933 5043
rect 317 5007 323 5033
rect 607 5017 673 5023
rect 1917 5023 1923 5033
rect 1957 5027 1963 5097
rect 2600 5103 2613 5107
rect 2597 5093 2613 5103
rect 3147 5097 3213 5103
rect 4787 5097 4833 5103
rect 2077 5043 2083 5093
rect 2260 5083 2273 5087
rect 2257 5073 2273 5083
rect 2597 5083 2603 5093
rect 2900 5083 2913 5087
rect 2577 5077 2603 5083
rect 2077 5037 2113 5043
rect 2257 5046 2263 5073
rect 2577 5047 2583 5077
rect 2897 5073 2913 5083
rect 2897 5047 2903 5073
rect 3297 5047 3303 5093
rect 5547 5097 5613 5103
rect 6127 5097 6163 5103
rect 3700 5083 3713 5087
rect 3697 5073 3713 5083
rect 3827 5083 3840 5087
rect 3827 5073 3843 5083
rect 2577 5037 2593 5047
rect 2580 5033 2593 5037
rect 2897 5037 2913 5047
rect 2900 5033 2913 5037
rect 3287 5037 3303 5047
rect 3287 5033 3300 5037
rect 3697 5043 3703 5073
rect 3837 5047 3843 5073
rect 3957 5077 3993 5083
rect 3957 5047 3963 5077
rect 5257 5077 5293 5083
rect 4177 5047 4183 5073
rect 5257 5047 5263 5077
rect 6157 5083 6163 5097
rect 6157 5077 6183 5083
rect 6177 5047 6183 5077
rect 3667 5037 3703 5043
rect 3827 5037 3843 5047
rect 3827 5033 3840 5037
rect 3947 5037 3963 5047
rect 3947 5033 3960 5037
rect 4167 5037 4183 5047
rect 4167 5033 4180 5037
rect 5247 5037 5263 5047
rect 5247 5033 5260 5037
rect 6167 5037 6183 5047
rect 6167 5033 6180 5037
rect 1940 5026 1963 5027
rect 1867 5017 1923 5023
rect 317 4997 333 5007
rect 320 4993 333 4997
rect 773 5003 787 5013
rect 1947 5017 1963 5026
rect 1947 5013 1960 5017
rect 2227 5017 2313 5023
rect 5387 5017 5433 5023
rect 773 5000 833 5003
rect 777 4997 833 5000
rect 1927 4977 1953 4983
rect 6243 4958 6303 5462
rect 6210 4942 6303 4958
rect 5247 4917 5273 4923
rect 227 4897 313 4903
rect 5687 4877 5713 4883
rect 1627 4863 1640 4867
rect 3320 4863 3333 4867
rect 1627 4853 1643 4863
rect 1637 4827 1643 4853
rect 3317 4853 3333 4863
rect 3807 4863 3820 4867
rect 3807 4853 3823 4863
rect 4327 4863 4340 4867
rect 4600 4863 4613 4867
rect 4327 4853 4343 4863
rect 3317 4827 3323 4853
rect 3817 4827 3823 4853
rect 4237 4827 4243 4853
rect 4337 4827 4343 4853
rect 4597 4853 4613 4863
rect 5100 4863 5113 4867
rect 5097 4853 5113 4863
rect 5387 4863 5400 4867
rect 5387 4853 5403 4863
rect 5527 4863 5540 4867
rect 5527 4853 5543 4863
rect 5827 4863 5840 4867
rect 5827 4853 5843 4863
rect 4597 4827 4603 4853
rect 1627 4817 1643 4827
rect 1627 4813 1640 4817
rect 3317 4817 3333 4827
rect 3320 4813 3333 4817
rect 3807 4817 3823 4827
rect 3807 4813 3820 4817
rect 4327 4817 4343 4827
rect 4327 4813 4340 4817
rect 4587 4817 4603 4827
rect 5097 4823 5103 4853
rect 5397 4827 5403 4853
rect 5077 4817 5103 4823
rect 4587 4813 4600 4817
rect 367 4797 413 4803
rect 867 4797 933 4803
rect 767 4783 813 4789
rect 1407 4797 1493 4803
rect 2187 4797 2233 4803
rect 2407 4797 2513 4803
rect 2587 4797 2613 4803
rect 3007 4797 3033 4803
rect 3057 4787 3063 4813
rect 4093 4803 4107 4813
rect 4093 4800 4133 4803
rect 4097 4797 4133 4800
rect 4207 4797 4253 4803
rect 5077 4803 5083 4817
rect 5387 4817 5403 4827
rect 5537 4823 5543 4853
rect 5837 4827 5843 4853
rect 5537 4817 5573 4823
rect 5387 4813 5400 4817
rect 5827 4817 5843 4827
rect 5827 4813 5840 4817
rect 5027 4797 5083 4803
rect 5467 4797 5553 4803
rect 5567 4797 5633 4803
rect 5787 4797 5873 4803
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 5927 4597 5973 4603
rect 1267 4577 1293 4583
rect 2847 4577 2893 4583
rect 3807 4577 3873 4583
rect 3887 4577 3913 4583
rect 4807 4577 4833 4583
rect 5547 4577 5593 4583
rect 5607 4577 5633 4583
rect 5907 4577 5963 4583
rect 360 4563 373 4567
rect 357 4553 373 4563
rect 357 4527 363 4553
rect 357 4517 373 4527
rect 360 4513 373 4517
rect 497 4523 503 4573
rect 747 4563 760 4567
rect 4240 4563 4253 4567
rect 747 4553 763 4563
rect 467 4517 503 4523
rect 757 4506 763 4553
rect 4237 4553 4253 4563
rect 4607 4557 4653 4563
rect 5420 4563 5433 4567
rect 5417 4553 5433 4563
rect 5820 4563 5833 4567
rect 5817 4553 5833 4563
rect 4237 4527 4243 4553
rect 3407 4517 3433 4523
rect 4227 4517 4243 4527
rect 4227 4513 4240 4517
rect 2707 4497 2753 4503
rect 3767 4497 3833 4503
rect 3967 4497 4033 4503
rect 4727 4497 4813 4503
rect 4827 4497 4853 4503
rect 5417 4503 5423 4553
rect 5817 4527 5823 4553
rect 5957 4527 5963 4577
rect 5807 4517 5823 4527
rect 5807 4513 5820 4517
rect 5947 4517 5963 4527
rect 5947 4513 5960 4517
rect 5367 4497 5423 4503
rect 6243 4438 6303 4942
rect 6210 4422 6303 4438
rect 2807 4397 2833 4403
rect 6167 4397 6213 4403
rect 3787 4377 3813 4383
rect 5967 4377 6013 4383
rect 2287 4357 2313 4363
rect 3807 4357 3833 4363
rect 5967 4357 6023 4363
rect 3173 4343 3187 4353
rect 3173 4340 3203 4343
rect 3177 4337 3203 4340
rect 3047 4297 3073 4303
rect 3197 4303 3203 4337
rect 5087 4337 5113 4343
rect 5620 4343 5633 4347
rect 5617 4333 5633 4343
rect 5760 4343 5773 4347
rect 5757 4333 5773 4343
rect 3197 4300 3223 4303
rect 3197 4297 3227 4300
rect 3213 4287 3227 4297
rect 4937 4303 4943 4333
rect 4907 4297 4943 4303
rect 5617 4307 5623 4333
rect 5757 4307 5763 4333
rect 5617 4297 5633 4307
rect 5620 4293 5633 4297
rect 5747 4297 5763 4307
rect 6017 4307 6023 4357
rect 6157 4357 6193 4363
rect 6157 4307 6163 4357
rect 6017 4297 6033 4307
rect 5747 4293 5760 4297
rect 6020 4293 6033 4297
rect 6147 4297 6163 4307
rect 6147 4293 6160 4297
rect 507 4277 533 4283
rect 1267 4277 1333 4283
rect 4207 4277 4253 4283
rect 4547 4277 4613 4283
rect 4627 4277 4693 4283
rect 5727 4277 5773 4283
rect 5967 4277 6073 4283
rect 5327 4237 5353 4243
rect 3067 4217 3093 4223
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 787 4097 813 4103
rect 6117 4100 6173 4103
rect 6113 4097 6173 4100
rect 6113 4087 6127 4097
rect 4507 4077 4573 4083
rect 1167 4057 1213 4063
rect 2627 4057 2683 4063
rect 197 4037 233 4043
rect 197 4007 203 4037
rect 1187 4043 1200 4047
rect 2040 4043 2053 4047
rect 1187 4033 1203 4043
rect 187 3997 203 4007
rect 187 3993 200 3997
rect 1027 3992 1058 3998
rect 1052 3983 1058 3992
rect 1052 3977 1073 3983
rect 1197 3986 1203 4033
rect 2037 4033 2053 4043
rect 2147 4043 2160 4047
rect 2420 4043 2433 4047
rect 2147 4033 2163 4043
rect 2037 4007 2043 4033
rect 2157 4007 2163 4033
rect 2417 4033 2433 4043
rect 2677 4043 2683 4057
rect 2727 4057 2753 4063
rect 2767 4057 2773 4063
rect 5107 4057 5153 4063
rect 5767 4057 5853 4063
rect 2860 4043 2873 4047
rect 2677 4037 2703 4043
rect 2417 4007 2423 4033
rect 2557 4007 2563 4033
rect 1727 3997 1763 4003
rect 1687 3977 1733 3983
rect 1757 3967 1763 3997
rect 2027 3997 2043 4007
rect 2027 3993 2040 3997
rect 2147 3997 2163 4007
rect 2147 3993 2160 3997
rect 2407 3997 2423 4007
rect 2407 3993 2420 3997
rect 2547 3997 2563 4007
rect 2697 4003 2703 4037
rect 2857 4033 2873 4043
rect 3580 4043 3593 4047
rect 3577 4033 3593 4043
rect 3707 4043 3720 4047
rect 3707 4033 3723 4043
rect 2857 4007 2863 4033
rect 2697 3997 2733 4003
rect 2547 3993 2560 3997
rect 2857 3997 2873 4007
rect 2860 3993 2873 3997
rect 3577 4003 3583 4033
rect 3547 3997 3583 4003
rect 3717 4007 3723 4033
rect 3717 3997 3733 4007
rect 3720 3993 3733 3997
rect 4397 3987 4403 4053
rect 4853 4043 4867 4053
rect 4837 4040 4867 4043
rect 4837 4037 4863 4040
rect 4837 4007 4843 4037
rect 4967 4037 4993 4043
rect 5120 4043 5133 4047
rect 5117 4033 5133 4043
rect 5327 4043 5340 4047
rect 6140 4043 6153 4047
rect 5327 4033 5343 4043
rect 5117 4007 5123 4033
rect 4827 3997 4843 4007
rect 4827 3993 4840 3997
rect 5107 3997 5123 4007
rect 5337 4006 5343 4033
rect 6137 4033 6153 4043
rect 5107 3993 5120 3997
rect 6137 4003 6143 4033
rect 6107 3997 6143 4003
rect 2627 3977 2693 3983
rect 4397 3986 4420 3987
rect 4397 3977 4413 3986
rect 4400 3973 4413 3977
rect 747 3957 773 3963
rect 1027 3957 1053 3963
rect 6243 3918 6303 4422
rect 6210 3902 6303 3918
rect 447 3837 493 3843
rect 287 3823 300 3827
rect 700 3823 713 3827
rect 287 3813 303 3823
rect 297 3787 303 3813
rect 697 3813 713 3823
rect 697 3787 703 3813
rect 297 3777 313 3787
rect 300 3773 313 3777
rect 687 3777 703 3787
rect 837 3787 843 3853
rect 4933 3843 4947 3853
rect 4933 3840 5033 3843
rect 4937 3837 5033 3840
rect 6067 3837 6163 3843
rect 967 3823 980 3827
rect 967 3813 983 3823
rect 1427 3823 1440 3827
rect 1427 3813 1443 3823
rect 2160 3823 2173 3827
rect 2157 3813 2173 3823
rect 2297 3817 2333 3823
rect 837 3777 853 3787
rect 687 3773 700 3777
rect 840 3773 853 3777
rect 977 3783 983 3813
rect 1437 3787 1443 3813
rect 977 3777 1003 3783
rect 997 3767 1003 3777
rect 1427 3777 1443 3787
rect 1427 3773 1440 3777
rect 387 3757 493 3763
rect 997 3757 1013 3767
rect 1000 3753 1013 3757
rect 1087 3757 1153 3763
rect 1457 3763 1463 3793
rect 1977 3783 1983 3813
rect 2157 3787 2163 3813
rect 2297 3787 2303 3817
rect 2447 3823 2460 3827
rect 2600 3823 2613 3827
rect 2447 3813 2463 3823
rect 2457 3787 2463 3813
rect 1977 3777 2033 3783
rect 2157 3777 2173 3787
rect 2160 3773 2173 3777
rect 2287 3777 2303 3787
rect 2287 3773 2300 3777
rect 2447 3777 2463 3787
rect 2597 3813 2613 3823
rect 3620 3823 3633 3827
rect 3617 3813 3633 3823
rect 4960 3823 4973 3827
rect 4957 3813 4973 3823
rect 5120 3823 5133 3827
rect 5117 3813 5133 3823
rect 5293 3823 5307 3833
rect 5247 3820 5307 3823
rect 5247 3817 5303 3820
rect 5547 3823 5560 3827
rect 5547 3813 5563 3823
rect 2447 3773 2460 3777
rect 1407 3757 1463 3763
rect 2427 3757 2493 3763
rect 2597 3763 2603 3813
rect 3617 3787 3623 3813
rect 3877 3787 3883 3813
rect 3607 3777 3623 3787
rect 3607 3773 3620 3777
rect 3867 3777 3883 3787
rect 4957 3787 4963 3813
rect 5117 3787 5123 3813
rect 5557 3787 5563 3813
rect 4957 3777 4973 3787
rect 3867 3773 3880 3777
rect 4960 3773 4973 3777
rect 5117 3777 5133 3787
rect 5120 3773 5133 3777
rect 5557 3777 5573 3787
rect 5560 3773 5573 3777
rect 6157 3786 6163 3837
rect 2547 3757 2603 3763
rect 3987 3757 4013 3763
rect 4307 3757 4333 3763
rect 4507 3757 4533 3763
rect 5407 3757 5473 3763
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 3247 3577 3293 3583
rect 4587 3557 4693 3563
rect 627 3523 640 3527
rect 673 3523 687 3533
rect 820 3523 833 3527
rect 627 3513 643 3523
rect 637 3467 643 3513
rect 657 3520 687 3523
rect 657 3517 683 3520
rect 657 3487 663 3517
rect 817 3513 833 3523
rect 947 3523 960 3527
rect 1100 3523 1113 3527
rect 947 3513 963 3523
rect 817 3487 823 3513
rect 957 3487 963 3513
rect 657 3477 673 3487
rect 660 3473 673 3477
rect 817 3477 833 3487
rect 820 3473 833 3477
rect 947 3477 963 3487
rect 1097 3513 1113 3523
rect 1187 3523 1200 3527
rect 1187 3513 1203 3523
rect 1427 3523 1440 3527
rect 1427 3513 1443 3523
rect 1097 3487 1103 3513
rect 1197 3487 1203 3513
rect 1437 3487 1443 3513
rect 1097 3477 1113 3487
rect 947 3473 960 3477
rect 1100 3473 1113 3477
rect 1187 3477 1203 3487
rect 1187 3473 1200 3477
rect 1427 3477 1443 3487
rect 1457 3487 1463 3533
rect 4587 3537 4643 3543
rect 4507 3523 4520 3527
rect 4637 3523 4643 3537
rect 4787 3537 4843 3543
rect 4507 3513 4523 3523
rect 4637 3517 4663 3523
rect 4517 3487 4523 3513
rect 4657 3487 4663 3517
rect 4807 3523 4820 3527
rect 4807 3513 4823 3523
rect 1457 3477 1473 3487
rect 1427 3473 1440 3477
rect 1460 3473 1473 3477
rect 4507 3477 4523 3487
rect 4507 3473 4520 3477
rect 4647 3477 4663 3487
rect 4817 3486 4823 3513
rect 4647 3473 4660 3477
rect 1047 3457 1093 3463
rect 4837 3463 4843 3537
rect 5887 3537 5943 3543
rect 5197 3517 5233 3523
rect 4807 3457 4843 3463
rect 4927 3457 5033 3463
rect 5197 3463 5203 3517
rect 5487 3523 5500 3527
rect 5487 3513 5503 3523
rect 5497 3487 5503 3513
rect 5637 3517 5673 3523
rect 5637 3487 5643 3517
rect 5787 3523 5800 3527
rect 5787 3513 5803 3523
rect 5797 3487 5803 3513
rect 5497 3477 5513 3487
rect 5500 3473 5513 3477
rect 5627 3477 5643 3487
rect 5627 3473 5640 3477
rect 5787 3477 5803 3487
rect 5937 3487 5943 3537
rect 5937 3477 5953 3487
rect 5787 3473 5800 3477
rect 5940 3473 5953 3477
rect 6077 3483 6083 3533
rect 6077 3477 6113 3483
rect 5087 3457 5203 3463
rect 6047 3457 6073 3463
rect 6243 3398 6303 3902
rect 6210 3382 6303 3398
rect 3807 3357 3853 3363
rect 1260 3303 1273 3307
rect 1257 3300 1273 3303
rect 1253 3293 1273 3300
rect 1387 3303 1400 3307
rect 1387 3293 1403 3303
rect 1253 3286 1267 3293
rect 1397 3267 1403 3293
rect 1387 3257 1403 3267
rect 1387 3253 1400 3257
rect 1417 3243 1423 3313
rect 4420 3303 4433 3307
rect 4417 3293 4433 3303
rect 4920 3303 4933 3307
rect 4917 3293 4933 3303
rect 5047 3303 5060 3307
rect 5320 3303 5333 3307
rect 5047 3293 5063 3303
rect 4417 3267 4423 3293
rect 1367 3237 1423 3243
rect 4417 3257 4433 3267
rect 4420 3253 4433 3257
rect 3833 3243 3847 3253
rect 3833 3240 3873 3243
rect 3837 3237 3873 3240
rect 4917 3237 4923 3293
rect 5057 3267 5063 3293
rect 5317 3293 5333 3303
rect 5317 3283 5323 3293
rect 5297 3277 5323 3283
rect 5297 3267 5303 3277
rect 5057 3257 5073 3267
rect 5060 3253 5073 3257
rect 5287 3257 5303 3267
rect 5287 3253 5300 3257
rect 4907 3231 4923 3237
rect 5047 3237 5093 3243
rect 6047 3237 6153 3243
rect 3567 3197 3633 3203
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 2737 3107 2743 3123
rect 2727 3097 2743 3107
rect 2727 3093 2740 3097
rect 3847 3057 3913 3063
rect 4467 3037 4533 3043
rect 4620 3043 4633 3047
rect 4617 3033 4633 3043
rect 727 3017 783 3023
rect 777 2967 783 3017
rect 3767 3017 3793 3023
rect 4447 3017 4473 3023
rect 3877 2997 3913 3003
rect 3877 2967 3883 2997
rect 4340 3003 4353 3007
rect 4337 2993 4353 3003
rect 777 2957 793 2967
rect 780 2953 793 2957
rect 3867 2957 3883 2967
rect 4337 2967 4343 2993
rect 4337 2957 4353 2967
rect 3867 2953 3880 2957
rect 4340 2953 4353 2957
rect 4617 2947 4623 3033
rect 5807 3017 5853 3023
rect 6127 3017 6153 3023
rect 6167 3017 6193 3023
rect 4640 3003 4653 3007
rect 4637 2993 4653 3003
rect 4907 3003 4920 3007
rect 5820 3003 5833 3007
rect 4907 2993 4923 3003
rect 4637 2967 4643 2993
rect 4637 2957 4653 2967
rect 4640 2953 4653 2957
rect 4027 2937 4073 2943
rect 4167 2937 4193 2943
rect 4917 2946 4923 2993
rect 5817 2993 5833 3003
rect 5980 3003 5993 3007
rect 5977 2993 5993 3003
rect 5817 2963 5823 2993
rect 5977 2967 5983 2993
rect 5817 2957 5843 2963
rect 5977 2957 5993 2967
rect 5837 2943 5843 2957
rect 5980 2953 5993 2957
rect 5837 2937 5893 2943
rect 6243 2878 6303 3382
rect 6210 2862 6303 2878
rect 2087 2837 2133 2843
rect 4347 2837 4393 2843
rect 5027 2817 5093 2823
rect 767 2797 853 2803
rect 4487 2797 4553 2803
rect 1200 2783 1213 2787
rect 1197 2773 1213 2783
rect 1327 2783 1340 2787
rect 4100 2783 4113 2787
rect 1327 2773 1343 2783
rect 1197 2747 1203 2773
rect 1337 2747 1343 2773
rect 1197 2737 1213 2747
rect 1200 2733 1213 2737
rect 1327 2737 1343 2747
rect 4097 2773 4113 2783
rect 4227 2783 4240 2787
rect 4333 2783 4347 2792
rect 4227 2773 4243 2783
rect 4333 2780 4373 2783
rect 4337 2777 4373 2780
rect 5240 2783 5253 2787
rect 5237 2773 5253 2783
rect 5380 2783 5393 2787
rect 5377 2773 5393 2783
rect 4097 2747 4103 2773
rect 4237 2747 4243 2773
rect 4097 2737 4113 2747
rect 1327 2733 1340 2737
rect 4100 2733 4113 2737
rect 4237 2737 4253 2747
rect 4240 2733 4253 2737
rect 5237 2743 5243 2773
rect 5377 2746 5383 2773
rect 5477 2747 5483 2793
rect 5500 2783 5513 2787
rect 5207 2737 5243 2743
rect 5467 2737 5483 2747
rect 5497 2773 5513 2783
rect 5627 2783 5640 2787
rect 5780 2783 5793 2787
rect 5627 2773 5643 2783
rect 5497 2747 5503 2773
rect 5637 2747 5643 2773
rect 5777 2773 5793 2783
rect 5777 2747 5783 2773
rect 5497 2737 5513 2747
rect 5467 2733 5480 2737
rect 5500 2733 5513 2737
rect 5637 2737 5653 2747
rect 5640 2733 5653 2737
rect 5767 2737 5783 2747
rect 5767 2733 5780 2737
rect 1827 2717 1873 2723
rect 3927 2717 3973 2723
rect 4067 2717 4153 2723
rect 4487 2717 4533 2723
rect 4787 2717 4813 2723
rect 4907 2717 4933 2723
rect 5587 2717 5693 2723
rect 6007 2717 6173 2723
rect 4527 2697 4573 2703
rect -63 2602 30 2618
rect 807 2613 810 2627
rect -63 2098 -3 2602
rect 4807 2577 4833 2583
rect 4120 2523 4133 2527
rect 4117 2513 4133 2523
rect 1327 2497 1363 2503
rect 1200 2483 1213 2487
rect 1197 2473 1213 2483
rect 1197 2447 1203 2473
rect 1187 2437 1203 2447
rect 1357 2443 1363 2497
rect 2107 2497 2133 2503
rect 3647 2497 3733 2503
rect 3807 2497 3833 2503
rect 1467 2483 1480 2487
rect 3540 2483 3553 2487
rect 1467 2473 1483 2483
rect 1337 2437 1363 2443
rect 1187 2433 1200 2437
rect 1337 2423 1343 2437
rect 1477 2427 1483 2473
rect 3537 2473 3553 2483
rect 3537 2447 3543 2473
rect 4117 2447 4123 2513
rect 5380 2503 5393 2507
rect 4227 2497 4263 2503
rect 4257 2447 4263 2497
rect 5377 2493 5393 2503
rect 5467 2497 5503 2503
rect 4487 2483 4500 2487
rect 4487 2473 4503 2483
rect 4667 2483 4680 2487
rect 5377 2483 5383 2493
rect 4667 2473 4683 2483
rect 4497 2447 4503 2473
rect 3537 2437 3553 2447
rect 3540 2433 3553 2437
rect 4117 2437 4133 2447
rect 4120 2433 4133 2437
rect 4257 2437 4273 2447
rect 4260 2433 4273 2437
rect 4487 2437 4503 2447
rect 4677 2447 4683 2473
rect 5357 2477 5383 2483
rect 5357 2447 5363 2477
rect 4677 2437 4693 2447
rect 4487 2433 4500 2437
rect 4680 2433 4693 2437
rect 5357 2437 5373 2447
rect 5360 2433 5373 2437
rect 5497 2443 5503 2497
rect 5987 2497 6073 2503
rect 5807 2477 5833 2483
rect 5497 2437 5523 2443
rect 1307 2417 1343 2423
rect 2107 2417 2133 2423
rect 4807 2417 4873 2423
rect 5517 2423 5523 2437
rect 5517 2417 5553 2423
rect 6243 2358 6303 2862
rect 6210 2342 6303 2358
rect 5907 2317 5933 2323
rect 2087 2277 2113 2283
rect 3657 2277 3693 2283
rect 900 2263 913 2267
rect 897 2253 913 2263
rect 1167 2263 1180 2267
rect 2080 2263 2093 2267
rect 1167 2253 1183 2263
rect 897 2227 903 2253
rect 1177 2227 1183 2253
rect 897 2217 913 2227
rect 900 2213 913 2217
rect 1167 2217 1183 2227
rect 2077 2253 2093 2263
rect 2367 2263 2380 2267
rect 2367 2253 2383 2263
rect 2547 2263 2560 2267
rect 2800 2263 2813 2267
rect 2547 2253 2563 2263
rect 2077 2223 2083 2253
rect 2377 2223 2383 2253
rect 2077 2217 2103 2223
rect 2377 2217 2413 2223
rect 1167 2213 1180 2217
rect 2097 2207 2103 2217
rect 967 2197 1013 2203
rect 1027 2197 1053 2203
rect 2097 2197 2113 2207
rect 2100 2193 2113 2197
rect 2240 2203 2253 2207
rect 2237 2193 2253 2203
rect 2557 2203 2563 2253
rect 2797 2253 2813 2263
rect 3520 2263 3533 2267
rect 3367 2257 3403 2263
rect 2797 2227 2803 2253
rect 2787 2217 2803 2227
rect 3397 2226 3403 2257
rect 3517 2253 3533 2263
rect 3517 2227 3523 2253
rect 3657 2227 3663 2277
rect 3967 2277 4013 2283
rect 4107 2277 4143 2283
rect 2787 2213 2800 2217
rect 3507 2217 3523 2227
rect 3507 2213 3520 2217
rect 3647 2217 3663 2227
rect 4137 2223 4143 2277
rect 4367 2263 4380 2267
rect 4367 2253 4383 2263
rect 4527 2263 4540 2267
rect 4527 2253 4543 2263
rect 4767 2263 4780 2267
rect 4920 2263 4933 2267
rect 4767 2253 4783 2263
rect 4377 2227 4383 2253
rect 4137 2217 4163 2223
rect 3647 2213 3660 2217
rect 2507 2197 2563 2203
rect 2667 2197 2733 2203
rect 3067 2197 3113 2203
rect 4157 2203 4163 2217
rect 4367 2217 4383 2227
rect 4537 2223 4543 2253
rect 4777 2227 4783 2253
rect 4917 2253 4933 2263
rect 5047 2263 5060 2267
rect 5047 2253 5063 2263
rect 4917 2227 4923 2253
rect 5057 2227 5063 2253
rect 5757 2257 5793 2263
rect 5757 2227 5763 2257
rect 4537 2217 4573 2223
rect 4367 2213 4380 2217
rect 4777 2217 4793 2227
rect 4780 2213 4793 2217
rect 4907 2217 4923 2227
rect 4907 2213 4920 2217
rect 5047 2217 5063 2227
rect 5047 2213 5060 2217
rect 5747 2217 5763 2227
rect 5747 2213 5760 2217
rect 4157 2197 4213 2203
rect 5407 2197 5493 2203
rect 2237 2183 2243 2193
rect 2167 2177 2243 2183
rect 4547 2157 4593 2163
rect 2173 2143 2187 2153
rect 2173 2140 2233 2143
rect 2177 2137 2233 2140
rect 4667 2126 4680 2127
rect 4667 2113 4673 2126
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 3787 2017 3813 2023
rect 1147 1977 1213 1983
rect 1227 1977 1253 1983
rect 1897 1977 1953 1983
rect 320 1963 333 1967
rect 317 1953 333 1963
rect 857 1957 913 1963
rect 317 1927 323 1953
rect 317 1917 333 1927
rect 320 1913 333 1917
rect 857 1906 863 1957
rect 1447 1963 1460 1967
rect 1447 1953 1463 1963
rect 1457 1927 1463 1953
rect 1897 1927 1903 1977
rect 2027 1977 2073 1983
rect 2707 1977 2773 1983
rect 3747 1977 3813 1983
rect 4007 1977 4053 1983
rect 4187 1977 4233 1983
rect 2167 1963 2180 1967
rect 2500 1963 2513 1967
rect 2167 1953 2183 1963
rect 2177 1927 2183 1953
rect 1457 1917 1473 1927
rect 1460 1913 1473 1917
rect 1897 1917 1913 1927
rect 1900 1913 1913 1917
rect 2167 1917 2183 1927
rect 2497 1953 2513 1963
rect 3333 1963 3347 1973
rect 5327 1977 5453 1983
rect 5667 1977 5773 1983
rect 5907 1977 6053 1983
rect 3317 1960 3347 1963
rect 3317 1957 3343 1960
rect 3477 1957 3513 1963
rect 2497 1927 2503 1953
rect 2497 1917 2513 1927
rect 2167 1913 2180 1917
rect 2500 1913 2513 1917
rect 3317 1923 3323 1957
rect 3477 1927 3483 1957
rect 3887 1963 3900 1967
rect 4580 1963 4593 1967
rect 3887 1953 3903 1963
rect 3287 1917 3323 1923
rect 3467 1917 3483 1927
rect 3897 1923 3903 1953
rect 4577 1953 4593 1963
rect 5140 1963 5153 1967
rect 5137 1953 5153 1963
rect 4577 1927 4583 1953
rect 5137 1927 5143 1953
rect 3897 1917 3933 1923
rect 3467 1913 3480 1917
rect 4577 1917 4593 1927
rect 4580 1913 4593 1917
rect 5127 1917 5143 1927
rect 5127 1913 5140 1917
rect 907 1897 933 1903
rect 6243 1838 6303 2342
rect 6210 1822 6303 1838
rect 2027 1757 2113 1763
rect 3507 1757 3553 1763
rect 1800 1743 1813 1747
rect 1797 1733 1813 1743
rect 1927 1743 1940 1747
rect 1927 1733 1943 1743
rect 487 1723 500 1727
rect 487 1713 503 1723
rect 497 1707 503 1713
rect 1797 1707 1803 1733
rect 1937 1707 1943 1733
rect 2057 1737 2093 1743
rect 2057 1707 2063 1737
rect 3913 1743 3927 1753
rect 4157 1757 4193 1763
rect 3913 1740 3943 1743
rect 3917 1737 3943 1740
rect 497 1697 513 1707
rect 500 1693 513 1697
rect 1797 1697 1813 1707
rect 1800 1693 1813 1697
rect 1937 1697 1953 1707
rect 1940 1693 1953 1697
rect 2047 1697 2063 1707
rect 3937 1707 3943 1737
rect 4157 1707 4163 1757
rect 5847 1757 5883 1763
rect 4407 1743 4420 1747
rect 4407 1733 4423 1743
rect 4847 1743 4860 1747
rect 4847 1733 4863 1743
rect 5147 1743 5160 1747
rect 5877 1743 5883 1757
rect 5147 1733 5163 1743
rect 5877 1737 5903 1743
rect 3937 1697 3953 1707
rect 2047 1693 2060 1697
rect 3940 1693 3953 1697
rect 4157 1697 4173 1707
rect 4160 1693 4173 1697
rect 4257 1704 4263 1720
rect 4257 1698 4293 1704
rect 4417 1703 4423 1733
rect 4417 1697 4453 1703
rect 1627 1677 1653 1683
rect 2367 1677 2413 1683
rect 4027 1677 4073 1683
rect 4857 1686 4863 1733
rect 5157 1707 5163 1733
rect 5147 1697 5163 1707
rect 5897 1703 5903 1737
rect 5897 1697 5933 1703
rect 5147 1693 5160 1697
rect 5087 1677 5233 1683
rect 5707 1677 5773 1683
rect 5937 1683 5943 1693
rect 5827 1677 5943 1683
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 537 1547 543 1563
rect 527 1537 543 1547
rect 527 1533 540 1537
rect 1607 1457 1633 1463
rect 1827 1457 1893 1463
rect 3947 1457 3993 1463
rect 3020 1443 3033 1447
rect 3017 1433 3033 1443
rect 3153 1443 3167 1453
rect 5927 1457 5953 1463
rect 3420 1443 3433 1447
rect 3137 1440 3167 1443
rect 3137 1437 3163 1440
rect 3017 1407 3023 1433
rect 3137 1407 3143 1437
rect 3417 1433 3433 1443
rect 3540 1443 3553 1447
rect 3537 1433 3553 1443
rect 5847 1443 5860 1447
rect 5847 1433 5863 1443
rect 3417 1407 3423 1433
rect 3017 1397 3033 1407
rect 3020 1393 3033 1397
rect 3137 1397 3153 1407
rect 3140 1393 3153 1397
rect 3407 1397 3423 1407
rect 3537 1407 3543 1433
rect 3537 1397 3553 1407
rect 3407 1393 3420 1397
rect 3540 1393 3553 1397
rect 4327 1377 4413 1383
rect 5147 1377 5213 1383
rect 5857 1383 5863 1433
rect 5827 1377 5863 1383
rect 5547 1357 5573 1363
rect 3267 1337 3313 1343
rect 3787 1337 3813 1343
rect 6243 1318 6303 1822
rect 6210 1302 6303 1318
rect 697 1280 753 1283
rect 693 1277 753 1280
rect 693 1267 707 1277
rect 297 1257 333 1263
rect 297 1243 303 1257
rect 2347 1257 2393 1263
rect 267 1237 303 1243
rect 4407 1237 4453 1243
rect 407 1223 420 1227
rect 580 1223 593 1227
rect 407 1213 423 1223
rect 417 1187 423 1213
rect 407 1177 423 1187
rect 577 1213 593 1223
rect 2020 1223 2033 1227
rect 2017 1213 2033 1223
rect 5340 1223 5353 1227
rect 5337 1213 5353 1223
rect 5587 1223 5600 1227
rect 5587 1213 5603 1223
rect 5900 1223 5913 1227
rect 577 1183 583 1213
rect 1797 1187 1803 1213
rect 2017 1187 2023 1213
rect 557 1180 583 1183
rect 553 1177 583 1180
rect 407 1173 420 1177
rect 553 1167 567 1177
rect 1787 1177 1803 1187
rect 1787 1173 1800 1177
rect 2007 1177 2023 1187
rect 2007 1173 2020 1177
rect 3087 1177 3113 1183
rect 5337 1183 5343 1213
rect 5597 1187 5603 1213
rect 5337 1177 5363 1183
rect 927 1157 993 1163
rect 1107 1157 1133 1163
rect 2907 1157 2953 1163
rect 3027 1157 3113 1163
rect 4707 1157 4773 1163
rect 5287 1157 5333 1163
rect 5357 1143 5363 1177
rect 5587 1177 5603 1187
rect 5587 1173 5600 1177
rect 5777 1163 5783 1218
rect 5897 1213 5913 1223
rect 5897 1187 5903 1213
rect 5897 1177 5913 1187
rect 5900 1173 5913 1177
rect 5721 1157 5783 1163
rect 5247 1137 5363 1143
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 2867 937 2933 943
rect 4187 937 4233 943
rect 4767 937 4813 943
rect 4927 937 5013 943
rect 5027 937 5053 943
rect 5127 937 5173 943
rect 5327 937 5393 943
rect 5407 937 5433 943
rect 307 923 320 927
rect 307 913 323 923
rect 447 923 460 927
rect 447 913 463 923
rect 747 923 760 927
rect 4560 923 4573 927
rect 747 913 763 923
rect 317 887 323 913
rect 457 887 463 913
rect 317 877 333 887
rect 320 873 333 877
rect 447 877 463 887
rect 757 883 763 913
rect 4557 913 4573 923
rect 5527 923 5540 927
rect 5527 913 5543 923
rect 5827 923 5840 927
rect 5827 913 5843 923
rect 4557 887 4563 913
rect 5537 887 5543 913
rect 5837 887 5843 913
rect 757 877 793 883
rect 447 873 460 877
rect 4547 877 4563 887
rect 4547 873 4560 877
rect 4967 880 5003 883
rect 4967 877 5007 880
rect 5537 877 5553 887
rect 4993 867 5007 877
rect 5540 873 5553 877
rect 5837 877 5853 887
rect 5840 873 5853 877
rect 6067 857 6153 863
rect 6243 798 6303 1302
rect 6210 782 6303 798
rect 2447 717 2473 723
rect 1320 703 1333 707
rect 1317 693 1333 703
rect 1980 703 1993 707
rect 1977 693 1993 703
rect 4187 697 4223 703
rect 1317 667 1323 693
rect 1977 667 1983 693
rect 4217 667 4223 697
rect 1317 657 1333 667
rect 1320 653 1333 657
rect 1977 657 1993 667
rect 1980 653 1993 657
rect 4217 657 4233 667
rect 4220 653 4233 657
rect 5947 657 5973 663
rect 847 637 973 643
rect 1387 637 1453 643
rect 1967 637 2013 643
rect 3727 637 3793 643
rect 1927 617 1993 623
rect -63 522 30 538
rect -63 18 -3 522
rect 5847 497 5893 503
rect 227 417 283 423
rect 277 403 283 417
rect 307 417 333 423
rect 387 417 423 423
rect 277 397 313 403
rect 417 403 423 417
rect 417 397 443 403
rect 437 367 443 397
rect 427 357 443 367
rect 577 367 583 453
rect 727 417 773 423
rect 1327 417 1453 423
rect 2427 417 2473 423
rect 2987 417 3093 423
rect 5447 417 5493 423
rect 5697 417 5793 423
rect 2127 403 2140 407
rect 2760 403 2773 407
rect 2127 393 2143 403
rect 577 357 593 367
rect 427 353 440 357
rect 580 353 593 357
rect 1407 337 1493 343
rect 2137 346 2143 393
rect 2757 393 2773 403
rect 2757 367 2763 393
rect 2747 357 2763 367
rect 2747 353 2760 357
rect 3547 337 3673 343
rect 3987 337 4073 343
rect 4747 337 4773 343
rect 5487 337 5553 343
rect 5697 346 5703 417
rect 6007 403 6020 407
rect 6007 393 6023 403
rect 6017 367 6023 393
rect 6017 357 6033 367
rect 6020 353 6033 357
rect 1547 317 1573 323
rect 2587 297 2633 303
rect 6243 278 6303 782
rect 6210 262 6303 278
rect 1507 237 1533 243
rect 2867 197 2893 203
rect 2157 177 2193 183
rect 2157 143 2163 177
rect 2137 140 2163 143
rect 2133 137 2163 140
rect 2133 127 2147 137
rect 3287 137 3313 143
rect 3927 137 3953 143
rect 907 117 973 123
rect 1647 117 1733 123
rect 2907 117 2973 123
rect 5047 117 5153 123
rect 1907 97 1933 103
rect 4027 97 4053 103
rect -63 2 30 18
rect 6243 2 6303 262
<< m2contact >>
rect 2813 6173 2827 6187
rect 2833 6173 2847 6187
rect 2053 6133 2067 6147
rect 2193 6133 2207 6147
rect 2613 6133 2627 6147
rect 2673 6133 2687 6147
rect 2993 6113 3007 6127
rect 5313 6113 5327 6127
rect 5353 6113 5367 6127
rect 2013 6073 2027 6087
rect 2953 6073 2967 6087
rect 1973 6053 1987 6067
rect 3733 6053 3747 6067
rect 3833 6051 3847 6065
rect 3873 6053 3887 6067
rect 3933 6053 3947 6067
rect 5573 6053 5587 6067
rect 5653 6053 5667 6067
rect 3373 6013 3387 6027
rect 3413 6013 3427 6027
rect 2313 5933 2327 5947
rect 2373 5933 2387 5947
rect 1973 5913 1987 5927
rect 2013 5913 2027 5927
rect 3533 5893 3547 5907
rect 3953 5893 3967 5907
rect 3993 5893 4007 5907
rect 5013 5893 5027 5907
rect 5153 5893 5167 5907
rect 513 5833 527 5847
rect 613 5833 627 5847
rect 2153 5833 2167 5847
rect 2193 5833 2207 5847
rect 3413 5833 3427 5847
rect 4633 5833 4647 5847
rect 4693 5833 4707 5847
rect 5093 5833 5107 5847
rect 5933 5893 5947 5907
rect 6033 5893 6047 5907
rect 5933 5853 5947 5867
rect 5173 5832 5187 5846
rect 6013 5831 6027 5845
rect 6133 5833 6147 5847
rect 73 5613 87 5627
rect 113 5614 127 5628
rect 173 5613 187 5627
rect 233 5613 247 5627
rect 3213 5613 3227 5627
rect 453 5593 467 5607
rect 893 5593 907 5607
rect 1353 5593 1367 5607
rect 1493 5593 1507 5607
rect 893 5553 907 5567
rect 1293 5553 1307 5567
rect 473 5533 487 5547
rect 613 5533 627 5547
rect 673 5533 687 5547
rect 1413 5533 1427 5547
rect 2733 5593 2747 5607
rect 3153 5593 3167 5607
rect 2673 5553 2687 5567
rect 3153 5553 3167 5567
rect 4093 5593 4107 5607
rect 5673 5593 5687 5607
rect 5713 5593 5727 5607
rect 4093 5553 4107 5567
rect 2233 5533 2247 5547
rect 2333 5533 2347 5547
rect 3293 5533 3307 5547
rect 3513 5531 3527 5545
rect 3553 5533 3567 5547
rect 373 5393 387 5407
rect 733 5393 747 5407
rect 1413 5394 1427 5408
rect 1613 5393 1627 5407
rect 1653 5393 1667 5407
rect 693 5333 707 5347
rect 1953 5373 1967 5387
rect 1373 5333 1387 5347
rect 1953 5333 1967 5347
rect 2013 5373 2027 5387
rect 2553 5373 2567 5387
rect 2593 5373 2607 5387
rect 3233 5393 3247 5407
rect 3473 5393 3487 5407
rect 3553 5394 3567 5408
rect 4073 5393 4087 5407
rect 4953 5393 4967 5407
rect 5013 5393 5027 5407
rect 6113 5393 6127 5407
rect 6193 5393 6207 5407
rect 53 5313 67 5327
rect 93 5313 107 5327
rect 373 5313 387 5327
rect 1613 5311 1627 5325
rect 1653 5313 1667 5327
rect 1813 5313 1827 5327
rect 1873 5313 1887 5327
rect 3133 5333 3147 5347
rect 3373 5373 3387 5387
rect 3533 5373 3547 5387
rect 3373 5333 3387 5347
rect 3473 5333 3487 5347
rect 4173 5373 4187 5387
rect 4093 5333 4107 5347
rect 4493 5373 4507 5387
rect 4233 5333 4247 5347
rect 4453 5333 4467 5347
rect 2053 5313 2067 5327
rect 3393 5313 3407 5327
rect 3413 5313 3427 5327
rect 3473 5312 3487 5326
rect 3553 5313 3567 5327
rect 3633 5313 3647 5327
rect 3693 5313 3707 5327
rect 4193 5312 4207 5326
rect 4253 5313 4267 5327
rect 1653 5292 1667 5306
rect 1693 5293 1707 5307
rect 4573 5293 4587 5307
rect 4633 5293 4647 5307
rect 3473 5252 3487 5266
rect 3533 5253 3547 5267
rect 953 5133 967 5147
rect 993 5113 1007 5127
rect 4313 5113 4327 5127
rect 4353 5113 4367 5127
rect 4693 5113 4707 5127
rect 4733 5113 4747 5127
rect 5493 5113 5507 5127
rect 5613 5113 5627 5127
rect 1073 5093 1087 5107
rect 1113 5093 1127 5107
rect 1333 5093 1347 5107
rect 1573 5093 1587 5107
rect 1713 5093 1727 5107
rect 1813 5093 1827 5107
rect 313 5033 327 5047
rect 1373 5033 1387 5047
rect 1813 5033 1827 5047
rect 1933 5033 1947 5047
rect 593 5013 607 5027
rect 673 5013 687 5027
rect 773 5013 787 5027
rect 1853 5013 1867 5027
rect 1993 5093 2007 5107
rect 2073 5093 2087 5107
rect 2613 5093 2627 5107
rect 3133 5093 3147 5107
rect 3213 5093 3227 5107
rect 3293 5093 3307 5107
rect 4773 5093 4787 5107
rect 4833 5093 4847 5107
rect 2273 5073 2287 5087
rect 2113 5033 2127 5047
rect 2913 5073 2927 5087
rect 5533 5092 5547 5106
rect 5613 5093 5627 5107
rect 6113 5093 6127 5107
rect 3713 5073 3727 5087
rect 3813 5073 3827 5087
rect 2253 5032 2267 5046
rect 2593 5033 2607 5047
rect 2913 5033 2927 5047
rect 3273 5033 3287 5047
rect 3653 5033 3667 5047
rect 3993 5073 4007 5087
rect 4173 5073 4187 5087
rect 5293 5073 5307 5087
rect 3813 5033 3827 5047
rect 3933 5033 3947 5047
rect 4153 5033 4167 5047
rect 5233 5033 5247 5047
rect 6153 5033 6167 5047
rect 333 4993 347 5007
rect 1933 5012 1947 5026
rect 2213 5013 2227 5027
rect 2313 5011 2327 5025
rect 5373 5013 5387 5027
rect 5433 5013 5447 5027
rect 833 4993 847 5007
rect 1913 4973 1927 4987
rect 1953 4973 1967 4987
rect 5233 4912 5247 4926
rect 5273 4913 5287 4927
rect 213 4893 227 4907
rect 313 4893 327 4907
rect 5673 4873 5687 4887
rect 5713 4872 5727 4886
rect 1613 4853 1627 4867
rect 3333 4853 3347 4867
rect 3793 4853 3807 4867
rect 4233 4853 4247 4867
rect 4313 4853 4327 4867
rect 4613 4853 4627 4867
rect 5113 4853 5127 4867
rect 5373 4853 5387 4867
rect 5513 4853 5527 4867
rect 5813 4853 5827 4867
rect 1613 4813 1627 4827
rect 3053 4813 3067 4827
rect 3333 4813 3347 4827
rect 3793 4813 3807 4827
rect 4093 4813 4107 4827
rect 4233 4813 4247 4827
rect 4313 4813 4327 4827
rect 4573 4813 4587 4827
rect 353 4793 367 4807
rect 413 4793 427 4807
rect 853 4793 867 4807
rect 933 4793 947 4807
rect 753 4779 767 4793
rect 813 4779 827 4793
rect 1393 4791 1407 4805
rect 1493 4793 1507 4807
rect 2173 4793 2187 4807
rect 2233 4793 2247 4807
rect 2393 4793 2407 4807
rect 2513 4793 2527 4807
rect 2573 4793 2587 4807
rect 2613 4793 2627 4807
rect 2993 4793 3007 4807
rect 3033 4793 3047 4807
rect 4133 4793 4147 4807
rect 4193 4793 4207 4807
rect 4253 4793 4267 4807
rect 5013 4793 5027 4807
rect 5373 4813 5387 4827
rect 5573 4813 5587 4827
rect 5813 4813 5827 4827
rect 5453 4793 5467 4807
rect 5553 4793 5567 4807
rect 5633 4793 5647 4807
rect 5773 4793 5787 4807
rect 5873 4793 5887 4807
rect 3053 4773 3067 4787
rect 1273 4673 1287 4687
rect 1993 4673 2007 4687
rect 3413 4673 3427 4687
rect 5913 4593 5927 4607
rect 5973 4593 5987 4607
rect 493 4573 507 4587
rect 1253 4573 1267 4587
rect 1293 4573 1307 4587
rect 2833 4573 2847 4587
rect 2893 4573 2907 4587
rect 3793 4573 3807 4587
rect 3873 4574 3887 4588
rect 3913 4573 3927 4587
rect 4793 4573 4807 4587
rect 4833 4573 4847 4587
rect 5533 4573 5547 4587
rect 5593 4574 5607 4588
rect 5633 4573 5647 4587
rect 5893 4573 5907 4587
rect 373 4553 387 4567
rect 373 4513 387 4527
rect 453 4513 467 4527
rect 733 4553 747 4567
rect 4253 4553 4267 4567
rect 4593 4553 4607 4567
rect 4653 4553 4667 4567
rect 5433 4553 5447 4567
rect 5833 4553 5847 4567
rect 3393 4513 3407 4527
rect 3433 4513 3447 4527
rect 4213 4513 4227 4527
rect 753 4492 767 4506
rect 2693 4493 2707 4507
rect 2753 4493 2767 4507
rect 3753 4493 3767 4507
rect 3833 4493 3847 4507
rect 3953 4493 3967 4507
rect 4033 4493 4047 4507
rect 4713 4493 4727 4507
rect 4813 4493 4827 4507
rect 4853 4493 4867 4507
rect 5353 4493 5367 4507
rect 5793 4513 5807 4527
rect 5933 4513 5947 4527
rect 2793 4393 2807 4407
rect 2833 4393 2847 4407
rect 6153 4393 6167 4407
rect 6213 4393 6227 4407
rect 3773 4373 3787 4387
rect 3813 4373 3827 4387
rect 5953 4373 5967 4387
rect 6013 4373 6027 4387
rect 2273 4353 2287 4367
rect 2313 4353 2327 4367
rect 3173 4353 3187 4367
rect 3793 4353 3807 4367
rect 3833 4353 3847 4367
rect 5953 4353 5967 4367
rect 3033 4293 3047 4307
rect 3073 4293 3087 4307
rect 4933 4333 4947 4347
rect 5073 4333 5087 4347
rect 5113 4333 5127 4347
rect 5633 4333 5647 4347
rect 5773 4333 5787 4347
rect 4893 4293 4907 4307
rect 5633 4293 5647 4307
rect 5733 4293 5747 4307
rect 6193 4353 6207 4367
rect 6033 4293 6047 4307
rect 6133 4293 6147 4307
rect 493 4273 507 4287
rect 533 4273 547 4287
rect 1253 4273 1267 4287
rect 1333 4273 1347 4287
rect 3213 4273 3227 4287
rect 4193 4273 4207 4287
rect 4253 4273 4267 4287
rect 4533 4273 4547 4287
rect 4613 4273 4627 4287
rect 4693 4273 4707 4287
rect 5713 4273 5727 4287
rect 5773 4273 5787 4287
rect 5953 4273 5967 4287
rect 6073 4273 6087 4287
rect 5313 4232 5327 4246
rect 5353 4233 5367 4247
rect 3053 4212 3067 4226
rect 3093 4213 3107 4227
rect 1593 4153 1607 4167
rect 1733 4153 1747 4167
rect 2873 4153 2887 4167
rect 3533 4153 3547 4167
rect 3693 4152 3707 4166
rect 773 4093 787 4107
rect 813 4093 827 4107
rect 6173 4093 6187 4107
rect 4493 4073 4507 4087
rect 4573 4073 4587 4087
rect 6113 4073 6127 4087
rect 1153 4053 1167 4067
rect 1213 4053 1227 4067
rect 2613 4054 2627 4068
rect 233 4033 247 4047
rect 1173 4033 1187 4047
rect 173 3993 187 4007
rect 1013 3987 1027 4001
rect 1073 3973 1087 3987
rect 2053 4033 2067 4047
rect 2133 4033 2147 4047
rect 2433 4033 2447 4047
rect 2553 4033 2567 4047
rect 2713 4053 2727 4067
rect 2753 4053 2767 4067
rect 2773 4053 2787 4067
rect 4393 4053 4407 4067
rect 4853 4053 4867 4067
rect 5093 4053 5107 4067
rect 5153 4053 5167 4067
rect 5753 4053 5767 4067
rect 5853 4053 5867 4067
rect 1713 3993 1727 4007
rect 1193 3972 1207 3986
rect 1673 3973 1687 3987
rect 1733 3973 1747 3987
rect 2013 3993 2027 4007
rect 2133 3993 2147 4007
rect 2393 3993 2407 4007
rect 2533 3993 2547 4007
rect 2873 4033 2887 4047
rect 3593 4033 3607 4047
rect 3693 4033 3707 4047
rect 2733 3993 2747 4007
rect 2873 3993 2887 4007
rect 3533 3992 3547 4006
rect 3733 3993 3747 4007
rect 4953 4033 4967 4047
rect 4993 4033 5007 4047
rect 5133 4033 5147 4047
rect 5313 4033 5327 4047
rect 4813 3993 4827 4007
rect 5093 3993 5107 4007
rect 6153 4033 6167 4047
rect 5333 3992 5347 4006
rect 6093 3993 6107 4007
rect 2613 3973 2627 3987
rect 2693 3973 2707 3987
rect 4413 3972 4427 3986
rect 733 3952 747 3966
rect 773 3953 787 3967
rect 1013 3953 1027 3967
rect 1053 3953 1067 3967
rect 1753 3953 1767 3967
rect 833 3853 847 3867
rect 4933 3853 4947 3867
rect 433 3833 447 3847
rect 493 3833 507 3847
rect 273 3813 287 3827
rect 713 3813 727 3827
rect 313 3773 327 3787
rect 673 3773 687 3787
rect 5033 3833 5047 3847
rect 5293 3833 5307 3847
rect 6053 3834 6067 3848
rect 953 3813 967 3827
rect 1413 3813 1427 3827
rect 1973 3813 1987 3827
rect 2173 3813 2187 3827
rect 853 3773 867 3787
rect 1453 3793 1467 3807
rect 1413 3773 1427 3787
rect 373 3753 387 3767
rect 493 3753 507 3767
rect 1013 3753 1027 3767
rect 1073 3753 1087 3767
rect 1153 3752 1167 3766
rect 1393 3751 1407 3765
rect 2333 3813 2347 3827
rect 2433 3813 2447 3827
rect 2033 3773 2047 3787
rect 2173 3773 2187 3787
rect 2273 3773 2287 3787
rect 2433 3773 2447 3787
rect 2613 3813 2627 3827
rect 3633 3813 3647 3827
rect 3873 3813 3887 3827
rect 4973 3813 4987 3827
rect 5133 3813 5147 3827
rect 5233 3813 5247 3827
rect 5533 3813 5547 3827
rect 2413 3751 2427 3765
rect 2493 3753 2507 3767
rect 2533 3753 2547 3767
rect 3593 3773 3607 3787
rect 3853 3773 3867 3787
rect 4973 3773 4987 3787
rect 5133 3773 5147 3787
rect 5573 3773 5587 3787
rect 6153 3772 6167 3786
rect 3973 3753 3987 3767
rect 4013 3753 4027 3767
rect 4293 3751 4307 3765
rect 4333 3753 4347 3767
rect 4493 3753 4507 3767
rect 4533 3753 4547 3767
rect 5393 3753 5407 3767
rect 5473 3753 5487 3767
rect 493 3633 507 3647
rect 1953 3633 1967 3647
rect 3933 3633 3947 3647
rect 3233 3573 3247 3587
rect 3293 3573 3307 3587
rect 4573 3553 4587 3567
rect 4693 3553 4707 3567
rect 673 3533 687 3547
rect 1453 3533 1467 3547
rect 613 3513 627 3527
rect 833 3513 847 3527
rect 933 3513 947 3527
rect 673 3473 687 3487
rect 833 3473 847 3487
rect 933 3473 947 3487
rect 1113 3513 1127 3527
rect 1173 3513 1187 3527
rect 1413 3513 1427 3527
rect 1113 3473 1127 3487
rect 1173 3473 1187 3487
rect 1413 3473 1427 3487
rect 4573 3532 4587 3546
rect 4493 3513 4507 3527
rect 4773 3533 4787 3547
rect 4793 3513 4807 3527
rect 1473 3473 1487 3487
rect 4493 3473 4507 3487
rect 4633 3473 4647 3487
rect 4813 3472 4827 3486
rect 633 3453 647 3467
rect 1033 3453 1047 3467
rect 1093 3452 1107 3466
rect 4793 3452 4807 3466
rect 5873 3533 5887 3547
rect 4913 3453 4927 3467
rect 5033 3453 5047 3467
rect 5073 3453 5087 3467
rect 5233 3513 5247 3527
rect 5473 3513 5487 3527
rect 5673 3513 5687 3527
rect 5773 3513 5787 3527
rect 5513 3473 5527 3487
rect 5613 3473 5627 3487
rect 5773 3473 5787 3487
rect 6073 3533 6087 3547
rect 5953 3473 5967 3487
rect 6113 3473 6127 3487
rect 6033 3453 6047 3467
rect 6073 3453 6087 3467
rect 3793 3353 3807 3367
rect 3853 3353 3867 3367
rect 1413 3313 1427 3327
rect 1273 3293 1287 3307
rect 1373 3293 1387 3307
rect 1253 3272 1267 3286
rect 1373 3253 1387 3267
rect 1353 3233 1367 3247
rect 4433 3293 4447 3307
rect 4933 3293 4947 3307
rect 5033 3293 5047 3307
rect 3833 3253 3847 3267
rect 4433 3253 4447 3267
rect 3873 3231 3887 3245
rect 4893 3226 4907 3240
rect 5333 3293 5347 3307
rect 5073 3253 5087 3267
rect 5273 3253 5287 3267
rect 5033 3233 5047 3247
rect 5093 3233 5107 3247
rect 6033 3233 6047 3247
rect 6153 3233 6167 3247
rect 3553 3193 3567 3207
rect 3633 3193 3647 3207
rect 793 3113 807 3127
rect 3313 3113 3327 3127
rect 3473 3113 3487 3127
rect 2713 3093 2727 3107
rect 3833 3053 3847 3067
rect 3913 3053 3927 3067
rect 4453 3033 4467 3047
rect 4533 3033 4547 3047
rect 4633 3033 4647 3047
rect 713 3013 727 3027
rect 3753 3013 3767 3027
rect 3793 3013 3807 3027
rect 4433 3014 4447 3028
rect 4473 3012 4487 3026
rect 3913 2993 3927 3007
rect 4353 2993 4367 3007
rect 793 2953 807 2967
rect 3853 2953 3867 2967
rect 4353 2953 4367 2967
rect 5793 3013 5807 3027
rect 5853 3013 5867 3027
rect 6113 3013 6127 3027
rect 6153 3014 6167 3028
rect 6193 3013 6207 3027
rect 4653 2993 4667 3007
rect 4893 2993 4907 3007
rect 4653 2953 4667 2967
rect 4013 2933 4027 2947
rect 4073 2933 4087 2947
rect 4153 2933 4167 2947
rect 4193 2933 4207 2947
rect 4613 2933 4627 2947
rect 5833 2993 5847 3007
rect 5993 2993 6007 3007
rect 4913 2932 4927 2946
rect 5993 2953 6007 2967
rect 5893 2933 5907 2947
rect 2073 2833 2087 2847
rect 2133 2833 2147 2847
rect 4333 2833 4347 2847
rect 4393 2833 4407 2847
rect 5013 2813 5027 2827
rect 5093 2813 5107 2827
rect 753 2792 767 2806
rect 853 2793 867 2807
rect 4333 2792 4347 2806
rect 4473 2793 4487 2807
rect 4553 2793 4567 2807
rect 5473 2793 5487 2807
rect 1213 2773 1227 2787
rect 1313 2773 1327 2787
rect 1213 2733 1227 2747
rect 1313 2733 1327 2747
rect 4113 2773 4127 2787
rect 4213 2773 4227 2787
rect 4373 2773 4387 2787
rect 5253 2773 5267 2787
rect 5393 2773 5407 2787
rect 4113 2733 4127 2747
rect 4253 2733 4267 2747
rect 5193 2733 5207 2747
rect 5373 2732 5387 2746
rect 5453 2733 5467 2747
rect 5513 2773 5527 2787
rect 5613 2773 5627 2787
rect 5793 2773 5807 2787
rect 5513 2733 5527 2747
rect 5653 2733 5667 2747
rect 5753 2733 5767 2747
rect 1813 2713 1827 2727
rect 1873 2713 1887 2727
rect 3913 2713 3927 2727
rect 3973 2713 3987 2727
rect 4053 2713 4067 2727
rect 4153 2713 4167 2727
rect 4473 2713 4487 2727
rect 4533 2713 4547 2727
rect 4773 2713 4787 2727
rect 4813 2713 4827 2727
rect 4893 2713 4907 2727
rect 4933 2713 4947 2727
rect 5573 2713 5587 2727
rect 5693 2713 5707 2727
rect 5993 2713 6007 2727
rect 6173 2713 6187 2727
rect 4513 2693 4527 2707
rect 4573 2693 4587 2707
rect 793 2613 807 2627
rect 333 2593 347 2607
rect 1113 2593 1127 2607
rect 1633 2593 1647 2607
rect 2033 2593 2047 2607
rect 2373 2593 2387 2607
rect 4793 2572 4807 2586
rect 4833 2573 4847 2587
rect 4133 2513 4147 2527
rect 1313 2494 1327 2508
rect 1213 2473 1227 2487
rect 1173 2433 1187 2447
rect 2093 2493 2107 2507
rect 2133 2493 2147 2507
rect 3633 2493 3647 2507
rect 3733 2494 3747 2508
rect 3793 2493 3807 2507
rect 3833 2493 3847 2507
rect 1453 2473 1467 2487
rect 1293 2413 1307 2427
rect 3553 2473 3567 2487
rect 4213 2493 4227 2507
rect 5393 2493 5407 2507
rect 5453 2494 5467 2508
rect 4473 2473 4487 2487
rect 4653 2473 4667 2487
rect 3553 2433 3567 2447
rect 4133 2433 4147 2447
rect 4273 2433 4287 2447
rect 4473 2433 4487 2447
rect 4693 2433 4707 2447
rect 5373 2433 5387 2447
rect 5973 2493 5987 2507
rect 6073 2493 6087 2507
rect 5793 2473 5807 2487
rect 5833 2473 5847 2487
rect 1473 2413 1487 2427
rect 2093 2413 2107 2427
rect 2133 2413 2147 2427
rect 4793 2413 4807 2427
rect 4873 2413 4887 2427
rect 5553 2413 5567 2427
rect 5893 2313 5907 2327
rect 5933 2313 5947 2327
rect 2073 2273 2087 2287
rect 2113 2273 2127 2287
rect 913 2253 927 2267
rect 1153 2253 1167 2267
rect 913 2213 927 2227
rect 1153 2213 1167 2227
rect 2093 2253 2107 2267
rect 2353 2253 2367 2267
rect 2533 2253 2547 2267
rect 2413 2213 2427 2227
rect 953 2193 967 2207
rect 1013 2193 1027 2207
rect 1053 2193 1067 2207
rect 2113 2193 2127 2207
rect 2253 2193 2267 2207
rect 2493 2193 2507 2207
rect 2813 2253 2827 2267
rect 3353 2253 3367 2267
rect 2773 2213 2787 2227
rect 3533 2253 3547 2267
rect 3693 2273 3707 2287
rect 3953 2273 3967 2287
rect 4013 2273 4027 2287
rect 4093 2273 4107 2287
rect 3393 2212 3407 2226
rect 3493 2213 3507 2227
rect 3633 2213 3647 2227
rect 4353 2253 4367 2267
rect 4513 2253 4527 2267
rect 4753 2253 4767 2267
rect 2653 2193 2667 2207
rect 2733 2193 2747 2207
rect 3053 2193 3067 2207
rect 3113 2193 3127 2207
rect 4353 2213 4367 2227
rect 4933 2253 4947 2267
rect 5033 2253 5047 2267
rect 5793 2253 5807 2267
rect 4573 2213 4587 2227
rect 4793 2213 4807 2227
rect 4893 2213 4907 2227
rect 5033 2213 5047 2227
rect 5733 2213 5747 2227
rect 4213 2193 4227 2207
rect 5393 2193 5407 2207
rect 5493 2193 5507 2207
rect 2153 2173 2167 2187
rect 2173 2153 2187 2167
rect 4533 2153 4547 2167
rect 4593 2153 4607 2167
rect 2233 2133 2247 2147
rect 4653 2113 4667 2127
rect 4673 2112 4687 2126
rect 113 2073 127 2087
rect 1073 2073 1087 2087
rect 3773 2012 3787 2026
rect 3813 2013 3827 2027
rect 1133 1973 1147 1987
rect 1213 1973 1227 1987
rect 1253 1973 1267 1987
rect 333 1953 347 1967
rect 333 1913 347 1927
rect 913 1953 927 1967
rect 1433 1953 1447 1967
rect 1953 1973 1967 1987
rect 2013 1973 2027 1987
rect 2073 1973 2087 1987
rect 2693 1973 2707 1987
rect 2773 1973 2787 1987
rect 3333 1973 3347 1987
rect 3733 1973 3747 1987
rect 3813 1973 3827 1987
rect 3993 1974 4007 1988
rect 4053 1973 4067 1987
rect 4173 1973 4187 1987
rect 4233 1973 4247 1987
rect 2153 1953 2167 1967
rect 1473 1913 1487 1927
rect 1913 1913 1927 1927
rect 2153 1913 2167 1927
rect 2513 1953 2527 1967
rect 5313 1972 5327 1986
rect 5453 1973 5467 1987
rect 5653 1973 5667 1987
rect 5773 1973 5787 1987
rect 5893 1973 5907 1987
rect 6053 1973 6067 1987
rect 2513 1913 2527 1927
rect 3273 1913 3287 1927
rect 3513 1953 3527 1967
rect 3873 1953 3887 1967
rect 3453 1913 3467 1927
rect 4593 1953 4607 1967
rect 5153 1953 5167 1967
rect 3933 1913 3947 1927
rect 4593 1913 4607 1927
rect 5113 1913 5127 1927
rect 853 1892 867 1906
rect 893 1893 907 1907
rect 933 1893 947 1907
rect 2013 1753 2027 1767
rect 2113 1753 2127 1767
rect 3493 1753 3507 1767
rect 3553 1753 3567 1767
rect 3913 1753 3927 1767
rect 1813 1733 1827 1747
rect 1913 1733 1927 1747
rect 473 1713 487 1727
rect 2093 1733 2107 1747
rect 513 1693 527 1707
rect 1813 1693 1827 1707
rect 1953 1693 1967 1707
rect 2033 1693 2047 1707
rect 4193 1753 4207 1767
rect 5833 1752 5847 1766
rect 4253 1720 4267 1734
rect 4393 1733 4407 1747
rect 4833 1733 4847 1747
rect 5133 1733 5147 1747
rect 3953 1693 3967 1707
rect 4173 1693 4187 1707
rect 4293 1693 4307 1707
rect 4453 1693 4467 1707
rect 1613 1673 1627 1687
rect 1653 1673 1667 1687
rect 2353 1673 2367 1687
rect 2413 1673 2427 1687
rect 4013 1673 4027 1687
rect 4073 1673 4087 1687
rect 5133 1693 5147 1707
rect 5933 1693 5947 1707
rect 4853 1672 4867 1686
rect 5073 1673 5087 1687
rect 5233 1673 5247 1687
rect 5693 1673 5707 1687
rect 5773 1673 5787 1687
rect 5813 1671 5827 1685
rect 1253 1553 1267 1567
rect 513 1533 527 1547
rect 1593 1453 1607 1467
rect 1633 1453 1647 1467
rect 1813 1452 1827 1466
rect 1893 1453 1907 1467
rect 3153 1453 3167 1467
rect 3933 1453 3947 1467
rect 3993 1453 4007 1467
rect 3033 1433 3047 1447
rect 5913 1452 5927 1466
rect 5953 1454 5967 1468
rect 3433 1433 3447 1447
rect 3553 1433 3567 1447
rect 5833 1433 5847 1447
rect 3033 1393 3047 1407
rect 3153 1393 3167 1407
rect 3393 1393 3407 1407
rect 3553 1393 3567 1407
rect 4313 1373 4327 1387
rect 4413 1373 4427 1387
rect 5133 1373 5147 1387
rect 5213 1373 5227 1387
rect 5813 1373 5827 1387
rect 5533 1353 5547 1367
rect 5573 1353 5587 1367
rect 3253 1333 3267 1347
rect 3313 1333 3327 1347
rect 3773 1333 3787 1347
rect 3813 1333 3827 1347
rect 753 1273 767 1287
rect 253 1234 267 1248
rect 333 1253 347 1267
rect 693 1253 707 1267
rect 2333 1253 2347 1267
rect 2393 1253 2407 1267
rect 4393 1233 4407 1247
rect 4453 1233 4467 1247
rect 393 1213 407 1227
rect 393 1173 407 1187
rect 593 1213 607 1227
rect 1793 1213 1807 1227
rect 2033 1213 2047 1227
rect 5353 1213 5367 1227
rect 5573 1213 5587 1227
rect 5773 1218 5787 1232
rect 1773 1173 1787 1187
rect 1993 1173 2007 1187
rect 3073 1173 3087 1187
rect 3113 1173 3127 1187
rect 553 1153 567 1167
rect 913 1153 927 1167
rect 993 1153 1007 1167
rect 1093 1153 1107 1167
rect 1133 1153 1147 1167
rect 2893 1153 2907 1167
rect 2953 1153 2967 1167
rect 3013 1153 3027 1167
rect 3113 1152 3127 1166
rect 4693 1153 4707 1167
rect 4773 1153 4787 1167
rect 5273 1151 5287 1165
rect 5333 1153 5347 1167
rect 5233 1133 5247 1147
rect 5573 1173 5587 1187
rect 5707 1153 5721 1167
rect 5913 1213 5927 1227
rect 5913 1173 5927 1187
rect 2853 933 2867 947
rect 2933 933 2947 947
rect 4173 933 4187 947
rect 4233 933 4247 947
rect 4753 934 4767 948
rect 4813 933 4827 947
rect 4913 933 4927 947
rect 5013 934 5027 948
rect 5053 933 5067 947
rect 5113 933 5127 947
rect 5173 933 5187 947
rect 5313 933 5327 947
rect 5393 932 5407 946
rect 5433 934 5447 948
rect 293 913 307 927
rect 433 913 447 927
rect 733 913 747 927
rect 333 873 347 887
rect 433 873 447 887
rect 4573 913 4587 927
rect 5513 913 5527 927
rect 5813 913 5827 927
rect 793 873 807 887
rect 4533 873 4547 887
rect 4953 873 4967 887
rect 5553 873 5567 887
rect 5853 873 5867 887
rect 4993 853 5007 867
rect 6053 853 6067 867
rect 6153 853 6167 867
rect 2433 713 2447 727
rect 2473 713 2487 727
rect 1333 693 1347 707
rect 1993 693 2007 707
rect 4173 693 4187 707
rect 1333 653 1347 667
rect 1993 653 2007 667
rect 4233 653 4247 667
rect 5933 653 5947 667
rect 5973 653 5987 667
rect 833 633 847 647
rect 973 633 987 647
rect 1373 633 1387 647
rect 1453 633 1467 647
rect 1953 633 1967 647
rect 2013 633 2027 647
rect 3713 633 3727 647
rect 3793 633 3807 647
rect 1913 613 1927 627
rect 1993 613 2007 627
rect 5833 493 5847 507
rect 5893 493 5907 507
rect 573 453 587 467
rect 213 414 227 428
rect 293 413 307 427
rect 333 413 347 427
rect 373 413 387 427
rect 313 392 327 406
rect 413 353 427 367
rect 713 413 727 427
rect 773 414 787 428
rect 1313 413 1327 427
rect 1453 413 1467 427
rect 2413 413 2427 427
rect 2473 413 2487 427
rect 2973 413 2987 427
rect 3093 413 3107 427
rect 5433 413 5447 427
rect 5493 413 5507 427
rect 2113 393 2127 407
rect 593 353 607 367
rect 1393 333 1407 347
rect 1493 333 1507 347
rect 2773 393 2787 407
rect 2733 353 2747 367
rect 2133 332 2147 346
rect 3533 333 3547 347
rect 3673 333 3687 347
rect 3973 333 3987 347
rect 4073 333 4087 347
rect 4733 333 4747 347
rect 4773 333 4787 347
rect 5473 333 5487 347
rect 5553 333 5567 347
rect 5793 414 5807 428
rect 5993 393 6007 407
rect 6033 353 6047 367
rect 5693 332 5707 346
rect 1533 313 1547 327
rect 1573 313 1587 327
rect 2573 293 2587 307
rect 2633 293 2647 307
rect 1493 233 1507 247
rect 1533 233 1547 247
rect 2853 193 2867 207
rect 2893 193 2907 207
rect 2193 173 2207 187
rect 3273 133 3287 147
rect 3313 133 3327 147
rect 3913 133 3927 147
rect 3953 133 3967 147
rect 893 113 907 127
rect 973 113 987 127
rect 1633 113 1647 127
rect 1733 113 1747 127
rect 2133 113 2147 127
rect 2893 113 2907 127
rect 2973 113 2987 127
rect 5033 113 5047 127
rect 5153 113 5167 127
rect 1893 93 1907 107
rect 1933 93 1947 107
rect 4013 93 4027 107
rect 4053 93 4067 107
<< metal2 >>
rect 96 5947 103 6083
rect 136 6080 143 6083
rect 133 6067 147 6080
rect 256 5947 263 6083
rect 316 6007 323 6133
rect 353 6107 367 6110
rect 376 6074 384 6083
rect 416 6074 423 6193
rect 496 6116 503 6153
rect 336 6047 343 6073
rect 376 6067 423 6074
rect 16 5866 23 5933
rect 16 5566 23 5852
rect 36 5667 43 5893
rect 156 5866 163 5893
rect 116 5628 123 5852
rect 176 5643 183 5933
rect 316 5866 323 5953
rect 376 5947 383 6067
rect 436 5866 443 5892
rect 276 5827 283 5863
rect 456 5863 463 6053
rect 476 6047 483 6083
rect 516 6043 523 6073
rect 536 6067 543 6303
rect 576 6116 583 6153
rect 616 6116 623 6213
rect 516 6036 543 6043
rect 536 5908 543 6036
rect 596 5967 603 6083
rect 656 6023 663 6114
rect 676 6083 683 6153
rect 773 6126 823 6133
rect 773 6120 787 6126
rect 776 6116 783 6120
rect 676 6076 703 6083
rect 636 6016 663 6023
rect 636 5927 643 6016
rect 456 5856 483 5863
rect 516 5860 523 5863
rect 376 5647 383 5833
rect 396 5827 403 5852
rect 156 5636 183 5643
rect 73 5600 87 5613
rect 156 5607 163 5636
rect 76 5596 83 5600
rect 56 5327 63 5453
rect 116 5388 123 5533
rect 136 5527 143 5563
rect 156 5408 163 5553
rect 176 5527 183 5613
rect 233 5600 247 5613
rect 236 5596 243 5600
rect 396 5596 403 5653
rect 440 5603 453 5607
rect 436 5596 453 5603
rect 96 5340 103 5343
rect 56 5027 63 5273
rect 76 5087 83 5333
rect 93 5327 107 5340
rect 196 5287 203 5552
rect 316 5487 323 5594
rect 440 5593 453 5596
rect 476 5563 483 5856
rect 513 5847 527 5860
rect 556 5747 563 5863
rect 596 5843 603 5913
rect 656 5896 663 5993
rect 596 5836 613 5843
rect 496 5607 503 5713
rect 536 5596 543 5633
rect 576 5608 583 5753
rect 96 5076 103 5173
rect 116 4856 123 5043
rect 136 4867 143 5013
rect 16 3547 23 4593
rect 36 4567 43 4854
rect 56 4348 63 4613
rect 76 4527 83 4793
rect 96 4627 103 4823
rect 156 4807 163 5033
rect 176 4987 183 5173
rect 216 5103 223 5413
rect 336 5346 343 5533
rect 376 5523 383 5563
rect 416 5527 423 5563
rect 456 5556 483 5563
rect 376 5516 403 5523
rect 376 5407 383 5493
rect 396 5487 403 5516
rect 436 5387 443 5413
rect 296 5307 303 5343
rect 376 5340 383 5343
rect 216 5096 243 5103
rect 236 5088 243 5096
rect 316 5047 323 5074
rect 196 4907 203 5033
rect 216 4907 223 5043
rect 256 4987 263 5043
rect 336 5023 343 5332
rect 373 5327 387 5340
rect 456 5343 463 5556
rect 476 5467 483 5533
rect 496 5523 503 5553
rect 516 5543 523 5563
rect 556 5560 563 5563
rect 553 5547 567 5560
rect 516 5540 543 5543
rect 516 5536 547 5540
rect 533 5527 547 5536
rect 496 5516 523 5523
rect 516 5376 523 5516
rect 553 5380 567 5393
rect 556 5376 563 5380
rect 456 5336 483 5343
rect 316 5016 343 5023
rect 316 4907 323 5016
rect 347 5003 360 5007
rect 347 5000 363 5003
rect 347 4993 367 5000
rect 353 4987 367 4993
rect 416 4907 423 5003
rect 476 4967 483 5336
rect 496 5287 503 5343
rect 316 4856 323 4893
rect 436 4883 443 4953
rect 416 4876 443 4883
rect 156 4556 163 4593
rect 176 4467 183 4554
rect 56 3567 63 4073
rect 116 4063 123 4303
rect 176 4287 183 4334
rect 196 4087 203 4823
rect 236 4523 243 4645
rect 236 4516 263 4523
rect 236 4367 243 4516
rect 276 4507 283 4564
rect 336 4567 343 4823
rect 356 4527 363 4793
rect 396 4747 403 4854
rect 416 4807 423 4876
rect 476 4856 483 4913
rect 496 4863 503 5213
rect 536 5167 543 5332
rect 596 5307 603 5553
rect 616 5547 623 5833
rect 696 5727 703 6076
rect 716 5987 723 6083
rect 756 6080 763 6083
rect 753 6067 767 6080
rect 776 6007 783 6053
rect 733 5900 747 5913
rect 736 5896 743 5900
rect 776 5896 783 5993
rect 816 5987 823 6126
rect 836 6027 843 6193
rect 896 6128 903 6213
rect 876 5987 883 6083
rect 716 5608 723 5813
rect 636 5563 643 5594
rect 636 5556 663 5563
rect 656 5527 663 5556
rect 696 5547 703 5563
rect 687 5536 703 5547
rect 687 5533 700 5536
rect 716 5447 723 5533
rect 536 5076 543 5113
rect 576 5076 583 5153
rect 596 5147 603 5293
rect 616 5187 623 5333
rect 636 5307 643 5343
rect 716 5346 723 5433
rect 736 5407 743 5553
rect 756 5547 763 5733
rect 776 5523 783 5633
rect 796 5607 803 5913
rect 816 5747 823 5973
rect 916 5866 923 6083
rect 876 5827 883 5863
rect 896 5607 903 5713
rect 956 5647 963 5853
rect 976 5767 983 6303
rect 1076 6116 1083 6193
rect 1216 6167 1223 6193
rect 1216 6116 1223 6153
rect 1136 6067 1143 6114
rect 1296 6116 1323 6123
rect 1196 6080 1203 6083
rect 1056 5936 1063 6013
rect 996 5896 1023 5903
rect 996 5803 1003 5896
rect 1136 5863 1143 5893
rect 1116 5856 1143 5863
rect 996 5796 1023 5803
rect 976 5667 983 5753
rect 996 5608 1003 5633
rect 807 5556 823 5563
rect 756 5516 783 5523
rect 756 5383 763 5516
rect 796 5407 803 5553
rect 856 5483 863 5553
rect 876 5527 883 5593
rect 896 5527 903 5553
rect 847 5476 863 5483
rect 736 5376 763 5383
rect 796 5376 803 5393
rect 836 5376 843 5473
rect 696 5307 703 5333
rect 596 5040 603 5043
rect 556 5023 563 5032
rect 536 5016 563 5023
rect 593 5027 607 5040
rect 536 4867 543 5016
rect 636 4947 643 5033
rect 656 5007 663 5113
rect 676 5027 683 5073
rect 556 4887 563 4913
rect 496 4856 523 4863
rect 516 4627 523 4856
rect 576 4856 583 4893
rect 373 4567 387 4573
rect 507 4573 513 4587
rect 413 4560 427 4573
rect 500 4566 520 4567
rect 416 4556 423 4560
rect 507 4563 520 4566
rect 507 4556 523 4563
rect 573 4560 587 4573
rect 576 4556 583 4560
rect 507 4553 520 4556
rect 276 4383 283 4493
rect 296 4407 303 4523
rect 440 4523 453 4527
rect 376 4427 383 4513
rect 396 4467 403 4523
rect 436 4516 453 4523
rect 440 4513 453 4516
rect 476 4487 483 4533
rect 596 4526 603 4553
rect 276 4376 303 4383
rect 236 4336 243 4353
rect 96 4056 123 4063
rect 96 3947 103 4056
rect 196 4007 203 4034
rect 116 4000 123 4003
rect 113 3987 127 4000
rect 136 3667 143 3993
rect 176 3823 183 3993
rect 216 3883 223 4053
rect 236 4047 243 4193
rect 256 4127 263 4303
rect 296 4087 303 4376
rect 336 4336 343 4393
rect 496 4348 503 4513
rect 616 4487 623 4812
rect 656 4747 663 4953
rect 696 4856 703 5293
rect 716 5287 723 5332
rect 736 5107 743 5376
rect 756 5107 763 5233
rect 876 5227 883 5492
rect 916 5407 923 5533
rect 936 5447 943 5563
rect 976 5527 983 5563
rect 1016 5527 1023 5796
rect 1156 5767 1163 6072
rect 1193 6067 1207 6080
rect 1276 6086 1283 6113
rect 1256 5947 1263 6073
rect 1296 6027 1303 6116
rect 1376 5967 1383 6043
rect 1176 5727 1183 5933
rect 1256 5896 1263 5933
rect 1316 5866 1323 5893
rect 1276 5767 1283 5863
rect 1036 5547 1043 5693
rect 1196 5607 1203 5653
rect 1296 5603 1303 5773
rect 1276 5596 1303 5603
rect 1173 5563 1187 5573
rect 1156 5560 1187 5563
rect 1156 5556 1183 5560
rect 936 5376 943 5412
rect 976 5247 983 5513
rect 1116 5467 1123 5523
rect 996 5207 1003 5374
rect 1136 5207 1143 5473
rect 1176 5383 1183 5533
rect 1156 5376 1183 5383
rect 1196 5376 1203 5593
rect 1316 5587 1323 5733
rect 1256 5543 1263 5563
rect 1236 5536 1263 5543
rect 1236 5388 1243 5536
rect 1156 5346 1163 5376
rect 1256 5347 1263 5513
rect 1296 5427 1303 5553
rect 1313 5380 1327 5393
rect 1336 5383 1343 5953
rect 1416 5896 1423 5933
rect 1436 5927 1443 6153
rect 1536 6128 1543 6153
rect 1696 6116 1743 6123
rect 1596 6086 1603 6114
rect 1516 5967 1523 6083
rect 1556 6080 1563 6083
rect 1553 6067 1567 6080
rect 1596 6007 1603 6072
rect 1576 5908 1583 5953
rect 1356 5607 1363 5633
rect 1436 5596 1443 5852
rect 1516 5727 1523 5863
rect 1556 5827 1563 5863
rect 1616 5727 1623 6053
rect 1736 6027 1743 6116
rect 1756 6087 1763 6114
rect 1636 5863 1643 5894
rect 1636 5856 1653 5863
rect 1716 5827 1723 5933
rect 1776 5908 1783 6053
rect 1816 5967 1823 6083
rect 1827 5956 1843 5963
rect 1496 5607 1503 5653
rect 1476 5567 1483 5594
rect 1516 5596 1523 5713
rect 1556 5596 1563 5653
rect 1416 5547 1423 5563
rect 1576 5560 1583 5563
rect 1573 5547 1587 5560
rect 1376 5387 1383 5433
rect 1416 5408 1423 5533
rect 1316 5376 1323 5380
rect 1336 5376 1363 5383
rect 1216 5307 1223 5343
rect 1356 5346 1363 5376
rect 1456 5376 1463 5413
rect 1296 5267 1303 5332
rect 953 5127 967 5133
rect 776 5076 803 5083
rect 736 4967 743 5013
rect 773 5007 787 5013
rect 796 4987 803 5076
rect 836 5007 843 5113
rect 776 4907 783 4972
rect 816 4907 823 4993
rect 856 4963 863 5033
rect 856 4956 873 4963
rect 716 4820 723 4823
rect 713 4807 727 4820
rect 756 4793 763 4812
rect 776 4807 783 4893
rect 876 4856 883 4953
rect 896 4867 903 5043
rect 936 5027 943 5043
rect 927 5016 943 5027
rect 927 5013 940 5016
rect 916 4947 923 4992
rect 956 4987 963 5033
rect 936 4976 953 4983
rect 816 4820 823 4823
rect 856 4820 863 4823
rect 636 4526 643 4613
rect 736 4567 743 4733
rect 756 4527 763 4613
rect 796 4568 803 4813
rect 813 4807 827 4820
rect 853 4807 867 4820
rect 576 4348 583 4473
rect 616 4336 623 4373
rect 696 4336 703 4473
rect 356 4247 363 4303
rect 396 4300 403 4303
rect 393 4287 407 4300
rect 273 4040 287 4053
rect 276 4036 283 4040
rect 207 3876 223 3883
rect 156 3816 183 3823
rect 196 3816 203 3873
rect 256 3843 263 4003
rect 296 3947 303 4003
rect 356 3967 363 4034
rect 376 3947 383 4113
rect 396 4047 403 4233
rect 436 4167 443 4333
rect 536 4287 543 4334
rect 496 4007 503 4273
rect 596 4127 603 4303
rect 536 4036 543 4073
rect 636 4027 643 4273
rect 416 3927 423 3992
rect 436 3907 443 3953
rect 396 3847 403 3873
rect 256 3840 283 3843
rect 256 3836 287 3840
rect 156 3767 163 3816
rect 273 3827 287 3836
rect 216 3780 223 3783
rect 176 3707 183 3773
rect 213 3767 227 3780
rect 256 3747 263 3783
rect 96 3627 103 3653
rect 296 3647 303 3813
rect 336 3780 343 3783
rect 376 3780 383 3783
rect 316 3647 323 3773
rect 333 3767 347 3780
rect 373 3767 387 3780
rect 16 2788 23 3493
rect 36 3023 43 3293
rect 56 3247 63 3493
rect 76 3383 83 3503
rect 96 3407 103 3613
rect 196 3496 203 3633
rect 76 3376 103 3383
rect 76 3067 83 3353
rect 96 3347 103 3376
rect 136 3308 143 3393
rect 196 3287 203 3393
rect 336 3387 343 3533
rect 376 3500 383 3503
rect 373 3487 387 3500
rect 396 3407 403 3633
rect 416 3547 423 3814
rect 436 3647 443 3833
rect 493 3820 507 3833
rect 536 3828 543 3933
rect 556 3847 563 4003
rect 596 3947 603 4003
rect 496 3816 503 3820
rect 456 3527 463 3693
rect 476 3687 483 3772
rect 516 3767 523 3783
rect 507 3757 523 3767
rect 507 3753 520 3757
rect 496 3663 503 3732
rect 476 3656 503 3663
rect 453 3503 467 3513
rect 436 3500 467 3503
rect 436 3496 463 3500
rect 416 3447 423 3493
rect 476 3487 483 3656
rect 436 3407 443 3473
rect 476 3307 483 3433
rect 496 3347 503 3633
rect 556 3587 563 3783
rect 576 3727 583 3773
rect 596 3767 603 3833
rect 616 3827 623 3993
rect 656 3987 663 4293
rect 716 4147 723 4303
rect 756 4247 763 4492
rect 876 4467 883 4573
rect 916 4563 923 4912
rect 936 4807 943 4976
rect 976 4927 983 5133
rect 1007 5113 1013 5127
rect 1036 5076 1043 5153
rect 1076 5107 1083 5193
rect 1073 5080 1087 5093
rect 1076 5076 1083 5080
rect 1016 4947 1023 5043
rect 1056 4887 1063 5032
rect 1116 4907 1123 5093
rect 1216 5087 1223 5133
rect 1136 5046 1143 5073
rect 1236 5046 1243 5113
rect 1296 5076 1303 5153
rect 1333 5087 1347 5093
rect 1316 5007 1323 5032
rect 1076 4823 1083 4893
rect 1176 4856 1183 4893
rect 1356 4868 1363 5332
rect 1376 5247 1383 5333
rect 1436 5307 1443 5343
rect 1496 5327 1503 5413
rect 1556 5407 1563 5513
rect 1596 5427 1603 5473
rect 1616 5407 1623 5713
rect 1656 5608 1663 5693
rect 1676 5507 1683 5563
rect 1736 5547 1743 5853
rect 1756 5727 1763 5833
rect 1756 5527 1763 5653
rect 1816 5643 1823 5863
rect 1836 5667 1843 5956
rect 1856 5787 1863 6083
rect 1816 5640 1843 5643
rect 1816 5636 1847 5640
rect 1833 5627 1847 5636
rect 1856 5607 1863 5773
rect 1876 5563 1883 6303
rect 2053 6120 2067 6133
rect 2093 6120 2107 6133
rect 2056 6116 2063 6120
rect 2096 6116 2103 6120
rect 1936 6047 1943 6083
rect 1996 6086 2003 6113
rect 1986 6073 1987 6080
rect 1973 6067 1987 6073
rect 2027 6083 2040 6087
rect 2027 6076 2043 6083
rect 2027 6073 2040 6076
rect 1896 5907 1903 6013
rect 1936 6007 1943 6033
rect 1996 5927 2003 6072
rect 2036 5967 2043 6053
rect 2013 5927 2027 5933
rect 1933 5900 1947 5913
rect 1973 5900 1987 5913
rect 1936 5896 1943 5900
rect 1976 5896 1983 5900
rect 2136 5896 2143 6033
rect 2156 5947 2163 6153
rect 2196 6147 2203 6173
rect 2196 6116 2203 6133
rect 2313 6120 2327 6133
rect 2316 6116 2323 6120
rect 2276 6087 2283 6114
rect 2216 5987 2223 6083
rect 2336 6027 2343 6083
rect 2376 6047 2383 6083
rect 2416 6047 2423 6193
rect 2456 6128 2463 6233
rect 2573 6120 2587 6133
rect 2613 6120 2627 6133
rect 2576 6116 2583 6120
rect 2616 6116 2623 6120
rect 2536 6087 2543 6114
rect 2676 6087 2683 6133
rect 2756 6116 2763 6193
rect 2807 6173 2813 6187
rect 2833 6167 2847 6173
rect 2816 6087 2823 6133
rect 2636 6047 2643 6083
rect 2736 6063 2743 6072
rect 2736 6056 2763 6063
rect 2676 5947 2683 5973
rect 2256 5936 2313 5943
rect 2256 5927 2263 5936
rect 2387 5943 2400 5947
rect 2387 5940 2403 5943
rect 2387 5933 2407 5940
rect 2393 5927 2407 5933
rect 2247 5913 2263 5927
rect 2287 5923 2300 5927
rect 2287 5913 2303 5923
rect 1956 5687 1963 5863
rect 1996 5807 2003 5863
rect 2056 5807 2063 5894
rect 2296 5896 2303 5913
rect 2513 5900 2527 5913
rect 2696 5908 2703 5953
rect 2516 5896 2523 5900
rect 2156 5860 2163 5863
rect 2153 5847 2167 5860
rect 2196 5847 2203 5893
rect 2336 5867 2343 5894
rect 2236 5807 2243 5863
rect 2536 5860 2543 5863
rect 1836 5507 1843 5563
rect 1856 5556 1883 5563
rect 1856 5483 1863 5556
rect 1836 5476 1863 5483
rect 1516 5376 1563 5383
rect 1436 5076 1443 5153
rect 1456 5147 1463 5233
rect 1516 5167 1523 5376
rect 1656 5327 1663 5393
rect 1676 5327 1683 5413
rect 1756 5376 1763 5413
rect 1796 5376 1803 5453
rect 1536 5207 1543 5293
rect 1573 5080 1587 5093
rect 1616 5083 1623 5311
rect 1696 5307 1703 5333
rect 1576 5076 1583 5080
rect 1616 5076 1643 5083
rect 1416 5040 1423 5043
rect 1373 5027 1387 5033
rect 1413 5027 1427 5040
rect 1496 5007 1503 5074
rect 1636 5003 1643 5076
rect 1616 4996 1643 5003
rect 1376 4856 1383 4973
rect 1416 4887 1423 4913
rect 1416 4856 1423 4873
rect 1056 4816 1083 4823
rect 1096 4687 1103 4853
rect 1476 4826 1483 4853
rect 896 4556 923 4563
rect 936 4556 943 4613
rect 976 4556 983 4593
rect 1096 4588 1103 4673
rect 1136 4567 1143 4793
rect 1156 4707 1163 4823
rect 1276 4820 1283 4823
rect 1273 4807 1287 4820
rect 1176 4607 1183 4713
rect 1273 4667 1287 4673
rect 896 4487 903 4556
rect 956 4447 963 4523
rect 1007 4520 1023 4523
rect 1007 4516 1027 4520
rect 1013 4507 1027 4516
rect 776 4107 783 4433
rect 816 4336 823 4413
rect 896 4307 903 4393
rect 976 4343 983 4433
rect 967 4336 983 4343
rect 996 4306 1003 4333
rect 676 4047 683 4073
rect 716 4036 723 4093
rect 687 4003 700 4007
rect 687 3996 703 4003
rect 736 4000 743 4003
rect 687 3993 700 3996
rect 676 3823 683 3993
rect 733 3987 747 4000
rect 696 3847 703 3973
rect 776 3967 783 4072
rect 733 3947 747 3952
rect 816 3947 823 4093
rect 836 4036 843 4153
rect 896 4036 923 4043
rect 856 3967 863 4003
rect 716 3887 723 3913
rect 916 3907 923 4036
rect 936 3987 943 4233
rect 956 4047 963 4133
rect 976 4036 983 4073
rect 1016 4043 1023 4433
rect 1036 4387 1043 4553
rect 1076 4467 1083 4523
rect 1156 4467 1163 4573
rect 1253 4560 1267 4573
rect 1256 4556 1263 4560
rect 1136 4456 1153 4463
rect 1096 4336 1103 4373
rect 1136 4267 1143 4456
rect 1236 4407 1243 4523
rect 1296 4507 1303 4573
rect 1356 4568 1363 4613
rect 1396 4556 1403 4791
rect 1436 4767 1443 4823
rect 1496 4807 1503 4893
rect 1616 4867 1623 4996
rect 1656 4907 1663 5292
rect 1736 5247 1743 5343
rect 1776 5247 1783 5343
rect 1807 5313 1813 5327
rect 1836 5287 1843 5476
rect 1856 5387 1863 5433
rect 1876 5423 1883 5453
rect 1896 5447 1903 5613
rect 2016 5556 2033 5563
rect 1953 5523 1967 5533
rect 1953 5520 1983 5523
rect 1956 5516 1983 5520
rect 1916 5467 1923 5493
rect 1876 5416 1903 5423
rect 1896 5376 1903 5416
rect 1956 5387 1963 5493
rect 1976 5467 1983 5493
rect 1876 5327 1883 5343
rect 1876 5287 1883 5313
rect 1676 5087 1683 5213
rect 1696 5147 1703 5213
rect 1713 5088 1727 5093
rect 1756 5076 1763 5113
rect 1736 5007 1743 5043
rect 1796 5027 1803 5273
rect 1813 5088 1827 5093
rect 1896 5088 1903 5313
rect 1956 5267 1963 5333
rect 1936 5047 1943 5073
rect 1727 4996 1743 5007
rect 1727 4993 1740 4996
rect 1693 4860 1707 4873
rect 1696 4856 1703 4860
rect 1536 4820 1543 4823
rect 1533 4807 1547 4820
rect 1613 4807 1627 4813
rect 1636 4767 1643 4853
rect 1416 4587 1423 4693
rect 1196 4336 1203 4393
rect 1156 4163 1163 4293
rect 1176 4187 1183 4303
rect 1216 4207 1223 4303
rect 1256 4300 1263 4303
rect 1253 4287 1267 4300
rect 1296 4267 1303 4292
rect 1316 4227 1323 4554
rect 1496 4543 1503 4653
rect 1596 4568 1603 4613
rect 1476 4536 1503 4543
rect 1376 4520 1383 4523
rect 1336 4348 1343 4512
rect 1373 4507 1387 4520
rect 1333 4267 1347 4273
rect 1376 4207 1383 4292
rect 1396 4267 1403 4373
rect 1416 4348 1423 4513
rect 1456 4427 1463 4533
rect 1156 4156 1183 4163
rect 1016 4036 1043 4043
rect 1096 4036 1103 4093
rect 1156 4067 1163 4093
rect 996 4001 1027 4003
rect 996 3994 1013 4001
rect 956 3907 963 3993
rect 816 3843 823 3873
rect 836 3867 843 3893
rect 816 3836 843 3843
rect 656 3816 683 3823
rect 673 3767 687 3773
rect 576 3716 593 3727
rect 580 3713 593 3716
rect 596 3607 603 3673
rect 616 3527 623 3633
rect 636 3483 643 3733
rect 656 3627 663 3693
rect 676 3547 683 3673
rect 696 3547 703 3833
rect 727 3823 740 3827
rect 727 3816 743 3823
rect 727 3813 740 3816
rect 796 3776 823 3783
rect 756 3747 763 3772
rect 716 3587 723 3653
rect 756 3647 763 3712
rect 796 3603 803 3713
rect 816 3703 823 3776
rect 836 3727 843 3836
rect 856 3827 863 3853
rect 956 3827 963 3853
rect 856 3747 863 3773
rect 816 3696 843 3703
rect 796 3596 823 3603
rect 667 3516 703 3523
rect 616 3476 643 3483
rect 596 3407 603 3472
rect 216 3276 243 3283
rect 96 3260 103 3263
rect 93 3247 107 3260
rect 236 3247 243 3276
rect 176 3240 183 3243
rect 173 3227 187 3240
rect 316 3223 323 3273
rect 496 3283 503 3333
rect 476 3276 503 3283
rect 516 3283 523 3393
rect 596 3308 603 3393
rect 596 3283 603 3294
rect 516 3276 543 3283
rect 576 3276 603 3283
rect 476 3227 483 3276
rect 316 3216 343 3223
rect 336 3127 343 3216
rect 536 3187 543 3276
rect 496 3127 503 3173
rect 36 3016 63 3023
rect 36 2907 43 2994
rect 56 2847 63 3016
rect 156 2980 163 2983
rect 153 2966 167 2980
rect 36 1887 43 2053
rect 56 1967 63 2793
rect 116 2776 123 2952
rect 136 2483 143 2653
rect 196 2607 203 3053
rect 216 2887 223 2983
rect 256 2807 263 3113
rect 496 2887 503 3113
rect 556 3016 563 3233
rect 256 2776 283 2783
rect 216 2740 223 2743
rect 213 2727 227 2740
rect 276 2647 283 2776
rect 127 2476 143 2483
rect 233 2480 247 2493
rect 236 2476 243 2480
rect 136 2223 143 2476
rect 116 2216 143 2223
rect 113 2067 127 2073
rect 16 1756 33 1763
rect 16 708 23 1756
rect 36 1716 43 1753
rect 56 1723 63 1913
rect 76 1767 83 1923
rect 56 1716 83 1723
rect 96 1716 103 1813
rect 136 1726 143 1993
rect 156 1922 163 2413
rect 196 1987 203 2353
rect 256 2223 263 2253
rect 236 2216 263 2223
rect 256 2027 263 2216
rect 276 2167 283 2573
rect 296 2507 303 2873
rect 336 2687 343 2743
rect 333 2607 347 2613
rect 376 2587 383 2743
rect 416 2503 423 2733
rect 436 2627 443 2793
rect 476 2776 483 2833
rect 516 2807 523 2983
rect 516 2707 523 2743
rect 536 2687 543 2813
rect 596 2783 603 2833
rect 616 2827 623 3476
rect 636 3367 643 3453
rect 656 3447 663 3513
rect 676 3423 683 3473
rect 656 3416 683 3423
rect 656 3207 663 3416
rect 716 3367 723 3483
rect 736 3296 743 3433
rect 756 3327 763 3483
rect 776 3307 783 3473
rect 796 3467 803 3573
rect 816 3487 823 3596
rect 836 3527 843 3696
rect 876 3647 883 3783
rect 916 3627 923 3693
rect 856 3567 863 3593
rect 853 3520 867 3532
rect 856 3516 863 3520
rect 936 3527 943 3733
rect 956 3667 963 3772
rect 976 3587 983 3973
rect 1007 3953 1013 3967
rect 1036 3887 1043 4036
rect 1176 4047 1183 4156
rect 1196 4007 1203 4113
rect 1076 4000 1083 4003
rect 1073 3987 1087 4000
rect 1116 3983 1123 4003
rect 1216 4006 1223 4053
rect 1256 4036 1263 4073
rect 1096 3976 1123 3983
rect 1096 3963 1103 3976
rect 1067 3956 1103 3963
rect 1036 3876 1053 3887
rect 1040 3873 1053 3876
rect 996 3856 1033 3863
rect 996 3827 1003 3856
rect 1013 3820 1027 3833
rect 1016 3816 1023 3820
rect 1096 3827 1103 3933
rect 996 3687 1003 3773
rect 1016 3647 1023 3753
rect 1036 3727 1043 3783
rect 1076 3780 1083 3783
rect 1073 3767 1087 3780
rect 1096 3623 1103 3773
rect 1116 3747 1123 3953
rect 1196 3947 1203 3972
rect 1136 3767 1143 3873
rect 1156 3787 1163 3933
rect 1196 3816 1203 3853
rect 1236 3843 1243 4032
rect 1316 4000 1323 4003
rect 1313 3990 1327 4000
rect 1356 3990 1363 4113
rect 1436 4087 1443 4393
rect 1476 4336 1483 4453
rect 1496 4367 1503 4473
rect 1736 4447 1743 4973
rect 1756 4687 1763 5013
rect 1776 4887 1783 4933
rect 1796 4907 1803 4953
rect 1816 4856 1823 5033
rect 1856 4868 1863 5013
rect 1876 4887 1883 5043
rect 1956 5046 1963 5213
rect 1796 4820 1803 4823
rect 1776 4707 1783 4812
rect 1793 4807 1807 4820
rect 1836 4787 1843 4823
rect 1916 4783 1923 4973
rect 1936 4823 1943 5012
rect 1956 4987 1963 5032
rect 1976 4987 1983 5374
rect 1996 5307 2003 5473
rect 2036 5447 2043 5552
rect 2013 5387 2027 5393
rect 2036 5376 2043 5433
rect 2076 5376 2083 5633
rect 2096 5608 2103 5673
rect 2107 5596 2123 5603
rect 2096 5407 2103 5594
rect 2236 5547 2243 5693
rect 2176 5427 2183 5523
rect 2256 5507 2263 5773
rect 2276 5587 2283 5852
rect 2533 5847 2547 5860
rect 2336 5647 2343 5813
rect 2313 5600 2327 5613
rect 2316 5596 2323 5600
rect 2456 5596 2463 5833
rect 2516 5663 2523 5713
rect 2496 5656 2523 5663
rect 2496 5596 2503 5656
rect 2416 5567 2423 5594
rect 2336 5560 2343 5563
rect 2333 5547 2347 5560
rect 2056 5340 2063 5343
rect 2053 5327 2067 5340
rect 2096 5287 2103 5343
rect 1996 5107 2003 5153
rect 2036 5107 2043 5253
rect 1996 5076 2003 5093
rect 2056 5076 2063 5193
rect 2076 5107 2083 5273
rect 2113 5247 2127 5253
rect 2107 5240 2127 5247
rect 2107 5236 2123 5240
rect 2107 5233 2120 5236
rect 2176 5207 2183 5332
rect 2196 5207 2203 5293
rect 2127 5180 2163 5183
rect 2127 5176 2167 5180
rect 2153 5167 2167 5176
rect 2036 4868 2043 4993
rect 2076 4947 2083 5072
rect 2096 5047 2103 5113
rect 2156 5076 2163 5113
rect 2096 4856 2103 4933
rect 2116 4887 2123 5033
rect 2136 4856 2143 5043
rect 2213 5027 2227 5033
rect 1936 4816 1963 4823
rect 1896 4776 1923 4783
rect 1796 4687 1803 4713
rect 1496 4296 1523 4303
rect 1313 3983 1363 3990
rect 1376 3927 1383 4073
rect 1236 3836 1263 3843
rect 1256 3783 1263 3836
rect 1176 3767 1183 3783
rect 1236 3776 1263 3783
rect 1160 3766 1183 3767
rect 1136 3667 1143 3753
rect 1167 3756 1183 3766
rect 1167 3753 1180 3756
rect 1076 3616 1103 3623
rect 1053 3520 1067 3533
rect 1076 3527 1083 3616
rect 1056 3516 1063 3520
rect 836 3447 843 3473
rect 876 3447 883 3483
rect 916 3447 923 3483
rect 936 3387 943 3473
rect 956 3387 963 3514
rect 1096 3487 1103 3593
rect 1176 3527 1183 3633
rect 1127 3523 1140 3527
rect 1127 3516 1143 3523
rect 1127 3513 1140 3516
rect 1036 3480 1043 3483
rect 1033 3467 1047 3480
rect 1033 3447 1047 3453
rect 836 3307 843 3373
rect 807 3283 820 3287
rect 807 3276 823 3283
rect 807 3273 820 3276
rect 716 3107 723 3263
rect 776 3240 783 3243
rect 676 3008 683 3093
rect 756 3023 763 3233
rect 773 3227 787 3240
rect 776 3147 783 3213
rect 796 3127 803 3233
rect 836 3127 843 3253
rect 756 3016 783 3023
rect 713 3000 727 3013
rect 716 2996 723 3000
rect 656 2907 663 2963
rect 756 2827 763 2993
rect 576 2776 603 2783
rect 416 2496 443 2503
rect 436 2476 443 2496
rect 456 2487 463 2633
rect 316 2227 323 2474
rect 516 2463 523 2493
rect 516 2456 543 2463
rect 376 2440 383 2443
rect 373 2427 387 2440
rect 416 2327 423 2443
rect 456 2307 463 2433
rect 576 2427 583 2776
rect 656 2746 663 2813
rect 740 2806 760 2807
rect 740 2803 753 2806
rect 736 2793 753 2803
rect 736 2776 743 2793
rect 776 2787 783 3016
rect 856 2996 863 3053
rect 876 3027 883 3073
rect 896 3016 903 3133
rect 916 3027 923 3113
rect 936 3047 943 3173
rect 793 2947 807 2953
rect 936 2963 943 2983
rect 916 2956 943 2963
rect 876 2847 883 2953
rect 896 2867 903 2953
rect 636 2736 653 2743
rect 756 2627 763 2743
rect 796 2627 803 2813
rect 836 2787 843 2833
rect 916 2827 923 2956
rect 853 2780 867 2793
rect 856 2776 863 2780
rect 816 2567 823 2773
rect 916 2746 923 2792
rect 716 2456 723 2533
rect 876 2508 883 2693
rect 376 2256 423 2263
rect 416 2248 423 2256
rect 473 2240 487 2253
rect 516 2246 523 2293
rect 756 2287 763 2353
rect 816 2267 823 2493
rect 916 2463 923 2732
rect 936 2687 943 2933
rect 956 2807 963 3153
rect 1076 3143 1083 3453
rect 1096 3403 1103 3452
rect 1116 3427 1123 3473
rect 1096 3396 1163 3403
rect 1136 3167 1143 3373
rect 1156 3367 1163 3396
rect 1176 3347 1183 3473
rect 1196 3427 1203 3533
rect 1216 3527 1223 3713
rect 1276 3647 1283 3913
rect 1376 3816 1383 3873
rect 1413 3827 1427 3833
rect 1256 3516 1263 3553
rect 1296 3547 1303 3813
rect 1287 3533 1303 3547
rect 1293 3506 1307 3513
rect 1156 3283 1163 3313
rect 1156 3276 1173 3283
rect 1156 3187 1163 3233
rect 1056 3136 1083 3143
rect 1056 3043 1063 3136
rect 1036 3036 1063 3043
rect 1036 2987 1043 3036
rect 1056 2976 1063 3013
rect 1033 2783 1047 2793
rect 1016 2780 1047 2783
rect 1016 2776 1043 2780
rect 956 2707 963 2733
rect 996 2727 1003 2743
rect 996 2716 1013 2727
rect 1000 2713 1013 2716
rect 996 2476 1003 2693
rect 1016 2507 1023 2633
rect 1056 2587 1063 2853
rect 1076 2746 1083 2793
rect 1076 2627 1083 2732
rect 1036 2476 1043 2553
rect 896 2456 923 2463
rect 836 2247 843 2413
rect 856 2327 863 2433
rect 476 2236 483 2240
rect 196 1976 213 1987
rect 236 1956 243 1993
rect 156 1915 224 1922
rect 316 1827 323 2013
rect 336 1967 343 2053
rect 376 1956 383 1993
rect 396 1967 403 2153
rect 456 2067 463 2233
rect 756 2236 783 2243
rect 756 2107 763 2236
rect 856 2206 863 2253
rect 416 1923 423 1943
rect 456 1943 463 2013
rect 456 1936 483 1943
rect 336 1847 343 1913
rect 356 1903 363 1923
rect 396 1916 423 1923
rect 396 1903 403 1916
rect 356 1896 403 1903
rect 36 1347 43 1423
rect 76 1367 83 1716
rect 296 1663 303 1713
rect 276 1656 303 1663
rect 276 1483 283 1656
rect 276 1476 303 1483
rect 16 366 23 493
rect 36 188 43 1333
rect 76 1216 83 1332
rect 116 1227 123 1353
rect 136 1127 143 1453
rect 276 1416 283 1453
rect 296 1427 303 1476
rect 336 1267 343 1313
rect 376 1267 383 1833
rect 396 1716 403 1873
rect 416 1727 423 1916
rect 436 1847 443 1933
rect 476 1727 483 1936
rect 656 1936 663 1973
rect 756 1943 763 2093
rect 816 1976 823 2192
rect 756 1936 783 1943
rect 436 1456 443 1672
rect 216 1216 223 1253
rect 253 1248 267 1253
rect 236 1127 243 1183
rect 216 927 223 1073
rect 156 916 203 923
rect 96 880 103 883
rect 76 807 83 873
rect 93 867 107 880
rect 196 867 203 916
rect 296 927 303 993
rect 256 880 263 883
rect 156 666 163 853
rect 216 747 223 873
rect 253 867 267 880
rect 116 447 123 663
rect 56 -24 63 433
rect 93 400 107 413
rect 96 396 103 400
rect 156 367 163 652
rect 207 414 213 427
rect 200 413 220 414
rect 256 396 263 493
rect 316 427 323 1253
rect 396 1227 403 1373
rect 416 1207 423 1393
rect 476 1307 483 1692
rect 496 1407 503 1933
rect 556 1736 563 1833
rect 596 1736 603 1833
rect 516 1607 523 1693
rect 536 1667 543 1703
rect 636 1686 643 1773
rect 516 1427 523 1533
rect 556 1436 563 1533
rect 596 1447 603 1553
rect 636 1487 643 1672
rect 656 1667 663 1813
rect 676 1747 683 1833
rect 756 1807 763 1853
rect 716 1736 723 1793
rect 776 1787 783 1913
rect 836 1907 843 1933
rect 856 1927 863 2192
rect 836 1748 843 1893
rect 856 1763 863 1892
rect 876 1827 883 2373
rect 896 1907 903 2456
rect 1016 2327 1023 2443
rect 927 2263 940 2267
rect 927 2256 943 2263
rect 976 2256 983 2313
rect 1016 2267 1023 2292
rect 927 2253 940 2256
rect 916 1967 923 2213
rect 953 2207 967 2212
rect 996 2027 1003 2173
rect 1016 2007 1023 2193
rect 1036 2187 1043 2413
rect 1076 2307 1083 2513
rect 1096 2427 1103 2573
rect 1116 2487 1123 2593
rect 1176 2527 1183 2833
rect 1196 2788 1203 3413
rect 1216 3363 1223 3473
rect 1236 3383 1243 3483
rect 1236 3376 1263 3383
rect 1216 3356 1243 3363
rect 1216 3167 1223 3333
rect 1216 3027 1223 3093
rect 1236 3067 1243 3356
rect 1256 3307 1263 3376
rect 1316 3327 1323 3473
rect 1336 3467 1343 3593
rect 1356 3527 1363 3783
rect 1376 3687 1383 3753
rect 1396 3667 1403 3751
rect 1416 3527 1423 3773
rect 1436 3727 1443 3853
rect 1456 3807 1463 4173
rect 1476 3848 1483 4073
rect 1496 3867 1503 4173
rect 1516 4127 1523 4296
rect 1536 4087 1543 4353
rect 1556 4243 1563 4413
rect 1576 4387 1583 4413
rect 1636 4367 1643 4433
rect 1633 4340 1647 4353
rect 1676 4347 1683 4393
rect 1636 4336 1643 4340
rect 1696 4327 1703 4433
rect 1756 4423 1763 4533
rect 1776 4507 1783 4543
rect 1796 4427 1803 4633
rect 1816 4487 1823 4533
rect 1836 4447 1843 4543
rect 1856 4427 1863 4753
rect 1876 4527 1883 4593
rect 1896 4487 1903 4776
rect 2016 4763 2023 4823
rect 2036 4787 2043 4854
rect 2056 4767 2063 4812
rect 2176 4767 2183 4793
rect 2016 4756 2053 4763
rect 2196 4747 2203 4933
rect 2236 4887 2243 5074
rect 2256 5067 2263 5493
rect 2516 5487 2523 5552
rect 2556 5507 2563 5633
rect 2596 5608 2603 5893
rect 2636 5863 2643 5894
rect 2636 5856 2663 5863
rect 2633 5600 2647 5613
rect 2636 5596 2643 5600
rect 2496 5376 2503 5433
rect 2656 5427 2663 5563
rect 2540 5383 2553 5387
rect 2536 5376 2553 5383
rect 2276 5346 2283 5373
rect 2356 5267 2363 5343
rect 2287 5083 2300 5087
rect 2287 5076 2303 5083
rect 2336 5076 2343 5113
rect 2287 5073 2300 5076
rect 2396 5087 2403 5343
rect 2416 5127 2423 5333
rect 2436 5227 2443 5374
rect 2540 5373 2553 5376
rect 2456 5336 2473 5343
rect 2456 5287 2463 5336
rect 2516 5340 2523 5343
rect 2513 5327 2527 5340
rect 2576 5327 2583 5413
rect 2676 5403 2683 5553
rect 2696 5547 2703 5613
rect 2736 5607 2743 5973
rect 2756 5967 2763 6056
rect 2776 6047 2783 6083
rect 2836 6047 2843 6114
rect 2936 6067 2943 6083
rect 2776 5947 2783 5973
rect 2773 5900 2787 5912
rect 2776 5896 2783 5900
rect 2796 5847 2803 5863
rect 2836 5860 2843 5863
rect 2833 5847 2847 5860
rect 2796 5663 2803 5833
rect 2876 5827 2883 6033
rect 2916 5867 2923 6033
rect 2936 5947 2943 6053
rect 2956 6047 2963 6073
rect 2976 5967 2983 6114
rect 3007 6123 3020 6127
rect 3007 6116 3023 6123
rect 3007 6113 3020 6116
rect 3096 6027 3103 6193
rect 3156 6116 3163 6153
rect 3316 6128 3323 6153
rect 3356 6116 3363 6193
rect 3436 6116 3443 6193
rect 3136 6080 3143 6083
rect 3133 6067 3147 6080
rect 3176 6027 3183 6083
rect 3136 5927 3143 5953
rect 3133 5900 3147 5913
rect 3136 5896 3143 5900
rect 3016 5843 3023 5863
rect 3036 5847 3043 5894
rect 3116 5860 3123 5863
rect 3113 5847 3127 5860
rect 2996 5836 3023 5843
rect 2996 5827 3003 5836
rect 2796 5656 2813 5663
rect 2716 5563 2723 5594
rect 2816 5596 2823 5653
rect 2716 5556 2733 5563
rect 2676 5396 2703 5403
rect 2696 5376 2703 5396
rect 2716 5387 2723 5493
rect 2596 5346 2603 5373
rect 2456 5088 2463 5233
rect 2476 5207 2483 5253
rect 2496 5167 2503 5213
rect 2516 5143 2523 5193
rect 2496 5136 2523 5143
rect 2407 5076 2423 5083
rect 2256 4856 2263 5032
rect 2236 4820 2243 4823
rect 2233 4807 2247 4820
rect 1936 4556 1943 4693
rect 1996 4567 2003 4673
rect 2016 4523 2023 4653
rect 2076 4627 2083 4653
rect 2056 4556 2063 4593
rect 2096 4556 2103 4693
rect 2116 4687 2123 4713
rect 2156 4627 2163 4673
rect 2176 4587 2183 4633
rect 2147 4583 2160 4587
rect 2147 4576 2163 4583
rect 2147 4573 2160 4576
rect 2016 4516 2043 4523
rect 2036 4503 2043 4516
rect 2116 4516 2143 4523
rect 1987 4496 2023 4503
rect 2036 4496 2063 4503
rect 1736 4416 1763 4423
rect 1736 4347 1743 4416
rect 1716 4316 1743 4323
rect 1556 4236 1573 4243
rect 1556 3967 1563 4003
rect 1576 3987 1583 4233
rect 1576 3807 1583 3973
rect 1596 3796 1603 4153
rect 1616 4147 1623 4303
rect 1676 4247 1683 4283
rect 1696 4223 1703 4273
rect 1676 4216 1703 4223
rect 1636 4048 1643 4073
rect 1676 4048 1683 4216
rect 1696 4167 1703 4193
rect 1736 4167 1743 4316
rect 1816 4287 1823 4313
rect 1696 4043 1703 4153
rect 1696 4036 1723 4043
rect 1716 4007 1723 4036
rect 1816 4036 1823 4073
rect 1836 4067 1843 4323
rect 1656 3987 1663 4003
rect 1656 3976 1673 3987
rect 1660 3973 1673 3976
rect 1456 3707 1463 3772
rect 1513 3766 1527 3772
rect 1476 3683 1483 3753
rect 1456 3680 1483 3683
rect 1456 3676 1487 3680
rect 1287 3303 1300 3307
rect 1287 3296 1303 3303
rect 1336 3296 1343 3413
rect 1356 3383 1363 3473
rect 1376 3407 1383 3483
rect 1356 3376 1383 3383
rect 1376 3307 1383 3376
rect 1287 3293 1300 3296
rect 1256 3243 1263 3272
rect 1356 3260 1363 3263
rect 1256 3236 1283 3243
rect 1216 2787 1223 2973
rect 1236 2887 1243 2983
rect 1256 2847 1263 3153
rect 1276 3027 1283 3236
rect 1296 3107 1303 3233
rect 1316 3087 1323 3252
rect 1353 3247 1367 3260
rect 1373 3247 1387 3253
rect 1336 3187 1343 3233
rect 1296 2947 1303 2983
rect 1116 2367 1123 2433
rect 1116 2268 1123 2313
rect 1176 2303 1183 2433
rect 1156 2296 1183 2303
rect 1156 2267 1163 2296
rect 1053 2207 1067 2212
rect 1136 2167 1143 2223
rect 1073 2087 1087 2093
rect 1156 2047 1163 2213
rect 936 1956 943 1993
rect 973 1960 987 1973
rect 976 1956 983 1960
rect 956 1920 963 1923
rect 953 1907 967 1920
rect 856 1756 883 1763
rect 876 1736 883 1756
rect 736 1696 763 1703
rect 756 1647 763 1696
rect 656 1467 663 1593
rect 616 1420 623 1423
rect 613 1407 627 1420
rect 656 1423 663 1453
rect 656 1416 683 1423
rect 356 1180 363 1183
rect 336 1127 343 1173
rect 353 1167 367 1180
rect 436 1183 443 1253
rect 473 1220 487 1233
rect 476 1216 483 1220
rect 556 1227 563 1273
rect 416 1180 443 1183
rect 413 1176 443 1180
rect 336 1087 343 1113
rect 356 916 363 1053
rect 396 1007 403 1173
rect 413 1167 427 1176
rect 536 1180 543 1183
rect 533 1167 547 1180
rect 426 1160 427 1167
rect 553 1167 567 1172
rect 436 927 443 1153
rect 576 923 583 1392
rect 636 1327 643 1413
rect 693 1267 707 1273
rect 596 1240 663 1243
rect 593 1236 663 1240
rect 593 1227 607 1236
rect 656 1216 663 1236
rect 596 1127 603 1173
rect 636 1127 643 1183
rect 576 916 603 923
rect 376 880 383 883
rect 336 427 343 873
rect 373 867 387 880
rect 416 827 423 883
rect 433 867 447 873
rect 456 847 463 914
rect 536 880 543 883
rect 356 708 363 793
rect 496 708 503 872
rect 533 867 547 880
rect 576 747 583 873
rect 536 696 543 733
rect 396 627 403 663
rect 456 627 463 694
rect 596 663 603 916
rect 656 916 663 1153
rect 676 1147 683 1183
rect 716 1167 723 1633
rect 776 1567 783 1733
rect 816 1547 823 1703
rect 856 1416 863 1703
rect 896 1627 903 1703
rect 936 1703 943 1893
rect 1056 1887 1063 1954
rect 956 1747 963 1872
rect 976 1736 983 1833
rect 936 1696 963 1703
rect 916 1667 923 1693
rect 956 1387 963 1696
rect 996 1547 1003 1703
rect 1013 1460 1027 1473
rect 1016 1456 1023 1460
rect 767 1273 773 1287
rect 736 1228 743 1253
rect 793 1220 807 1233
rect 796 1216 803 1220
rect 856 1187 863 1293
rect 896 1216 903 1313
rect 1056 1307 1063 1653
rect 1076 1587 1083 2013
rect 1096 1967 1103 2033
rect 1133 1960 1147 1973
rect 1136 1956 1143 1960
rect 1176 1956 1183 2273
rect 1196 2268 1203 2774
rect 1233 2780 1247 2793
rect 1236 2776 1243 2780
rect 1316 2787 1323 3013
rect 1336 2827 1343 3173
rect 1396 2947 1403 3453
rect 1416 3327 1423 3473
rect 1436 3303 1443 3653
rect 1456 3627 1463 3676
rect 1473 3667 1487 3676
rect 1453 3547 1467 3553
rect 1476 3523 1483 3632
rect 1496 3627 1503 3733
rect 1456 3516 1483 3523
rect 1456 3323 1463 3516
rect 1556 3527 1563 3673
rect 1476 3447 1483 3473
rect 1536 3480 1543 3483
rect 1533 3467 1547 3480
rect 1456 3316 1483 3323
rect 1416 3296 1443 3303
rect 1476 3296 1483 3316
rect 1516 3307 1523 3433
rect 1556 3403 1563 3473
rect 1536 3396 1563 3403
rect 1536 3367 1543 3396
rect 1416 3127 1423 3296
rect 1536 3266 1543 3353
rect 1576 3303 1583 3693
rect 1596 3587 1603 3653
rect 1616 3647 1623 3953
rect 1696 3947 1703 3993
rect 1736 3987 1743 4034
rect 1836 3967 1843 4003
rect 1756 3907 1763 3953
rect 1716 3800 1723 3803
rect 1713 3787 1727 3800
rect 1856 3787 1863 3992
rect 1876 3967 1883 4113
rect 1976 4107 1983 4413
rect 1996 4407 2003 4473
rect 2016 4387 2023 4496
rect 2016 4316 2023 4373
rect 2036 4307 2043 4353
rect 2056 4347 2063 4496
rect 2136 4447 2143 4516
rect 2076 4316 2103 4323
rect 1996 4127 2003 4213
rect 1896 3947 1903 4053
rect 1876 3807 1883 3932
rect 1916 3907 1923 3993
rect 1936 3967 1943 4003
rect 1976 3967 1983 4003
rect 1896 3863 1903 3893
rect 1896 3856 1923 3863
rect 1896 3796 1903 3833
rect 1633 3520 1647 3533
rect 1636 3516 1643 3520
rect 1616 3480 1623 3483
rect 1613 3467 1627 3480
rect 1656 3427 1663 3483
rect 1696 3447 1703 3673
rect 1916 3667 1923 3856
rect 1976 3827 1983 3893
rect 1967 3796 1983 3803
rect 1976 3687 1983 3796
rect 1753 3520 1767 3533
rect 1756 3516 1763 3520
rect 1796 3516 1803 3553
rect 1816 3527 1823 3613
rect 1556 3296 1603 3303
rect 1456 3260 1463 3263
rect 1453 3247 1467 3260
rect 1456 2986 1463 3113
rect 1556 3107 1563 3296
rect 1716 3303 1723 3513
rect 1696 3296 1723 3303
rect 1616 3260 1623 3263
rect 1576 3087 1583 3253
rect 1613 3247 1627 3260
rect 1696 3107 1703 3296
rect 1816 3263 1823 3433
rect 1776 3207 1783 3263
rect 1796 3256 1823 3263
rect 1776 3127 1783 3193
rect 1596 3007 1603 3093
rect 1416 2976 1443 2983
rect 1436 2927 1443 2976
rect 1616 2983 1623 3033
rect 1596 2976 1623 2983
rect 1436 2887 1443 2913
rect 1436 2807 1443 2873
rect 1216 2487 1223 2733
rect 1256 2707 1263 2743
rect 1296 2707 1303 2743
rect 1236 2607 1243 2633
rect 1276 2476 1283 2533
rect 1316 2508 1323 2733
rect 1256 2367 1263 2443
rect 1296 2440 1303 2443
rect 1293 2427 1307 2440
rect 1276 2256 1283 2293
rect 1216 2220 1223 2223
rect 1213 2207 1227 2220
rect 1196 1967 1203 2093
rect 1256 2087 1263 2223
rect 1316 2167 1323 2253
rect 1336 2207 1343 2313
rect 1356 2267 1363 2773
rect 1376 2527 1383 2743
rect 1396 2507 1403 2673
rect 1436 2587 1443 2753
rect 1456 2567 1463 2972
rect 1476 2707 1483 2813
rect 1536 2747 1543 2773
rect 1516 2667 1523 2743
rect 1456 2487 1463 2513
rect 1376 2387 1383 2473
rect 1476 2443 1483 2573
rect 1436 2436 1483 2443
rect 1416 2387 1423 2413
rect 1396 2256 1403 2333
rect 1456 2307 1463 2413
rect 1376 2187 1383 2223
rect 1416 2220 1423 2223
rect 1413 2207 1427 2220
rect 1267 1983 1280 1987
rect 1267 1973 1283 1983
rect 1116 1748 1123 1923
rect 1216 1823 1223 1973
rect 1276 1956 1283 1973
rect 1376 1963 1383 2152
rect 1356 1956 1383 1963
rect 1336 1926 1343 1953
rect 1256 1847 1263 1923
rect 1216 1816 1243 1823
rect 1096 1736 1113 1743
rect 1096 1706 1103 1736
rect 1156 1736 1163 1773
rect 1216 1706 1223 1793
rect 1236 1747 1243 1816
rect 1316 1736 1323 1793
rect 1336 1747 1343 1912
rect 1356 1807 1363 1956
rect 1436 1967 1443 2133
rect 1456 2067 1463 2253
rect 1476 2107 1483 2413
rect 1496 2407 1503 2633
rect 1516 2627 1523 2653
rect 1536 2488 1543 2712
rect 1556 2527 1563 2833
rect 1656 2743 1663 2793
rect 1636 2736 1663 2743
rect 1676 2727 1683 2853
rect 1696 2827 1703 3053
rect 1736 3027 1743 3093
rect 1753 3020 1767 3033
rect 1796 3027 1803 3256
rect 1816 3047 1823 3133
rect 1836 3067 1843 3653
rect 1953 3627 1967 3633
rect 1856 3347 1863 3553
rect 1876 3447 1883 3573
rect 1876 3323 1883 3433
rect 1856 3316 1883 3323
rect 1856 3296 1863 3316
rect 1956 3287 1963 3513
rect 1976 3267 1983 3534
rect 1996 3387 2003 3833
rect 2016 3787 2023 3993
rect 2036 3967 2043 4272
rect 2056 4047 2063 4213
rect 2076 4048 2083 4253
rect 2096 4227 2103 4316
rect 2116 4036 2123 4073
rect 2136 4047 2143 4373
rect 2176 4363 2183 4453
rect 2196 4427 2203 4493
rect 2216 4467 2223 4773
rect 2276 4747 2283 4823
rect 2296 4767 2303 4812
rect 2316 4687 2323 5011
rect 2356 5007 2363 5043
rect 2416 4943 2423 5076
rect 2496 5076 2503 5136
rect 2536 5076 2543 5173
rect 2576 5167 2583 5233
rect 2416 4936 2443 4943
rect 2376 4856 2383 4893
rect 2416 4856 2423 4913
rect 2436 4867 2443 4936
rect 2356 4787 2363 4823
rect 2396 4820 2403 4823
rect 2393 4807 2407 4820
rect 2456 4607 2463 4993
rect 2476 4967 2483 5043
rect 2576 5046 2583 5093
rect 2596 5087 2603 5332
rect 2676 5307 2683 5343
rect 2613 5080 2627 5093
rect 2616 5076 2623 5080
rect 2656 5076 2663 5193
rect 2516 4868 2523 4933
rect 2536 4887 2543 4913
rect 2556 4856 2563 5033
rect 2536 4807 2543 4823
rect 2576 4820 2583 4823
rect 2573 4807 2587 4820
rect 2527 4797 2543 4807
rect 2527 4793 2540 4797
rect 2476 4583 2483 4633
rect 2456 4576 2483 4583
rect 2456 4443 2463 4576
rect 2516 4547 2523 4772
rect 2556 4687 2563 4793
rect 2436 4436 2463 4443
rect 2380 4423 2393 4427
rect 2376 4413 2393 4423
rect 2156 4356 2183 4363
rect 2216 4356 2273 4363
rect 2116 3823 2123 3973
rect 2136 3847 2143 3993
rect 2116 3816 2143 3823
rect 2036 3663 2043 3773
rect 2096 3780 2103 3783
rect 2056 3687 2063 3772
rect 2093 3767 2107 3780
rect 2136 3727 2143 3816
rect 2027 3656 2043 3663
rect 2016 3516 2023 3653
rect 2116 3547 2123 3613
rect 1996 3260 2003 3263
rect 1896 3147 1903 3252
rect 1993 3247 2007 3260
rect 2036 3247 2043 3373
rect 2056 3367 2063 3472
rect 2076 3127 2083 3493
rect 2156 3347 2163 4356
rect 2216 4336 2223 4356
rect 2296 4327 2303 4353
rect 2176 4007 2183 4093
rect 2196 4047 2203 4213
rect 2236 4167 2243 4292
rect 2316 4183 2323 4353
rect 2376 4336 2383 4413
rect 2436 4387 2443 4436
rect 2476 4427 2483 4533
rect 2496 4407 2503 4543
rect 2536 4536 2563 4543
rect 2476 4348 2483 4373
rect 2516 4347 2523 4512
rect 2356 4227 2363 4303
rect 2316 4176 2343 4183
rect 2176 3827 2183 3972
rect 2216 3816 2223 3933
rect 2256 3828 2263 3993
rect 2276 3967 2283 4173
rect 2336 4036 2343 4176
rect 2316 4000 2323 4003
rect 2313 3987 2327 4000
rect 2356 3967 2363 4003
rect 2416 4003 2423 4273
rect 2496 4227 2503 4303
rect 2536 4287 2543 4536
rect 2576 4367 2583 4593
rect 2596 4527 2603 5033
rect 2716 5007 2723 5333
rect 2736 4967 2743 5552
rect 2756 5487 2763 5563
rect 2796 5560 2803 5563
rect 2793 5547 2807 5560
rect 2836 5388 2843 5453
rect 2856 5407 2863 5693
rect 2916 5596 2923 5733
rect 2976 5566 2983 5633
rect 2876 5556 2893 5563
rect 2776 5347 2783 5374
rect 2796 5307 2803 5343
rect 2776 5076 2783 5233
rect 2796 5227 2803 5293
rect 2876 5287 2883 5556
rect 2996 5547 3003 5813
rect 3036 5596 3043 5693
rect 3076 5596 3083 5673
rect 3116 5567 3123 5594
rect 3136 5567 3143 5793
rect 3176 5787 3183 5933
rect 3196 5903 3203 6053
rect 3236 5967 3243 6114
rect 3296 5967 3303 6083
rect 3196 5896 3223 5903
rect 3336 5863 3343 6083
rect 3396 6027 3403 6114
rect 3360 6023 3373 6027
rect 3356 6013 3373 6023
rect 3356 5887 3363 6013
rect 3413 6007 3427 6013
rect 3556 6007 3563 6193
rect 3596 6027 3603 6083
rect 3636 6076 3663 6083
rect 3393 5900 3407 5913
rect 3396 5896 3403 5900
rect 3496 5866 3503 5973
rect 3533 5907 3547 5913
rect 3516 5867 3523 5894
rect 3616 5896 3623 5973
rect 3656 5967 3663 6076
rect 3316 5856 3343 5863
rect 3416 5860 3423 5863
rect 3413 5847 3427 5860
rect 3556 5767 3563 5863
rect 3596 5843 3603 5852
rect 3576 5836 3603 5843
rect 3156 5607 3163 5713
rect 3176 5647 3183 5733
rect 3213 5600 3227 5613
rect 3216 5596 3223 5600
rect 2876 5247 2883 5273
rect 2816 5076 2823 5113
rect 2836 5107 2843 5213
rect 2876 5027 2883 5173
rect 2896 5088 2903 5393
rect 2936 5376 2943 5473
rect 2976 5376 2983 5433
rect 3036 5343 3043 5533
rect 3156 5527 3163 5553
rect 3236 5543 3243 5563
rect 3216 5536 3243 5543
rect 2956 5307 2963 5332
rect 2916 5087 2923 5273
rect 2936 5247 2943 5293
rect 2996 5287 3003 5343
rect 3016 5336 3043 5343
rect 2896 5046 2903 5074
rect 2976 5076 2983 5113
rect 2996 5087 3003 5133
rect 2956 5040 2963 5043
rect 2676 4856 2683 4893
rect 2616 4807 2623 4853
rect 2636 4767 2643 4793
rect 2656 4787 2663 4823
rect 2616 4568 2623 4733
rect 2696 4647 2703 4773
rect 2696 4587 2703 4633
rect 2693 4560 2707 4573
rect 2696 4556 2703 4560
rect 2616 4427 2623 4554
rect 2676 4427 2683 4473
rect 2696 4467 2703 4493
rect 2736 4487 2743 4953
rect 2756 4767 2763 4873
rect 2796 4747 2803 4812
rect 2836 4787 2843 4823
rect 2896 4743 2903 4893
rect 2916 4867 2923 5033
rect 2953 5027 2967 5040
rect 3016 5007 3023 5336
rect 3076 5307 3083 5343
rect 3116 5340 3123 5343
rect 3113 5327 3127 5340
rect 3056 5076 3063 5113
rect 3116 5076 3123 5233
rect 3136 5147 3143 5333
rect 3156 5327 3163 5473
rect 3216 5407 3223 5536
rect 3236 5407 3243 5513
rect 3276 5467 3283 5594
rect 3293 5547 3307 5553
rect 3256 5427 3263 5453
rect 3236 5376 3243 5393
rect 3176 5323 3183 5373
rect 3216 5340 3223 5343
rect 3213 5327 3227 5340
rect 3176 5316 3203 5323
rect 3156 5267 3163 5313
rect 3036 4947 3043 5073
rect 3076 4967 3083 5043
rect 3136 4907 3143 5093
rect 2996 4856 3003 4893
rect 2936 4793 2953 4807
rect 2896 4736 2913 4743
rect 2816 4627 2823 4673
rect 2836 4667 2843 4713
rect 2796 4556 2803 4593
rect 2833 4560 2847 4573
rect 2836 4556 2843 4560
rect 2753 4507 2767 4513
rect 2896 4487 2903 4573
rect 2656 4303 2663 4413
rect 2736 4336 2743 4413
rect 2756 4407 2763 4433
rect 2776 4336 2783 4413
rect 2796 4407 2803 4473
rect 2816 4407 2823 4453
rect 2676 4306 2683 4333
rect 2576 4300 2583 4303
rect 2573 4287 2587 4300
rect 2616 4267 2623 4303
rect 2636 4296 2663 4303
rect 2436 4047 2443 4193
rect 2456 4036 2463 4133
rect 2616 4068 2623 4213
rect 2636 4207 2643 4296
rect 2656 4227 2663 4273
rect 2756 4267 2763 4303
rect 2667 4216 2683 4223
rect 2567 4033 2573 4047
rect 2656 4036 2663 4073
rect 2676 4047 2683 4216
rect 2416 3996 2443 4003
rect 2393 3983 2407 3993
rect 2376 3980 2407 3983
rect 2376 3976 2403 3980
rect 2176 3747 2183 3773
rect 2236 3780 2243 3783
rect 2233 3767 2247 3780
rect 2276 3707 2283 3773
rect 2296 3627 2303 3853
rect 2316 3707 2323 3873
rect 2336 3827 2343 3933
rect 2376 3887 2383 3976
rect 2396 3816 2403 3853
rect 2436 3827 2443 3996
rect 2520 4003 2533 4007
rect 2516 3993 2533 4003
rect 2553 4003 2567 4012
rect 2553 4000 2583 4003
rect 2556 3996 2583 4000
rect 2516 3947 2523 3993
rect 2576 3983 2583 3996
rect 2696 3987 2703 4153
rect 2736 4087 2743 4193
rect 2756 4107 2763 4253
rect 2756 4067 2763 4093
rect 2796 4087 2803 4233
rect 2816 4147 2823 4313
rect 2836 4303 2843 4393
rect 2893 4340 2907 4353
rect 2896 4336 2903 4340
rect 2836 4296 2863 4303
rect 2836 4067 2843 4273
rect 2916 4223 2923 4733
rect 2936 4247 2943 4793
rect 2976 4787 2983 4812
rect 3036 4807 3043 4853
rect 3056 4827 3063 4893
rect 2996 4763 3003 4793
rect 2967 4756 3003 4763
rect 3053 4763 3067 4773
rect 3136 4767 3143 4823
rect 3053 4760 3083 4763
rect 3056 4756 3083 4760
rect 2956 4556 2963 4693
rect 2996 4667 3003 4693
rect 3016 4568 3023 4633
rect 3036 4627 3043 4713
rect 3036 4527 3043 4613
rect 2956 4227 2963 4493
rect 2976 4487 2983 4523
rect 2980 4443 2993 4447
rect 2976 4440 2993 4443
rect 2973 4433 2993 4440
rect 2973 4427 2987 4433
rect 2996 4336 3003 4393
rect 3016 4300 3023 4303
rect 3013 4287 3027 4300
rect 2916 4216 2943 4223
rect 2576 3976 2603 3983
rect 2376 3762 2383 3783
rect 2456 3786 2463 3813
rect 2376 3755 2413 3762
rect 2376 3667 2383 3755
rect 2436 3667 2443 3773
rect 2496 3780 2503 3783
rect 2493 3767 2507 3780
rect 2536 3767 2543 3783
rect 2516 3756 2533 3763
rect 2236 3507 2243 3533
rect 2256 3496 2263 3613
rect 2116 3260 2123 3263
rect 2113 3247 2127 3260
rect 2256 3247 2263 3263
rect 2296 3247 2303 3333
rect 1756 3016 1763 3020
rect 1816 3016 1823 3033
rect 1696 2707 1703 2792
rect 1716 2607 1723 2983
rect 1736 2787 1743 2973
rect 1796 2847 1803 2973
rect 1836 2867 1843 2953
rect 1836 2807 1843 2853
rect 1773 2780 1787 2793
rect 1856 2787 1863 2983
rect 1876 2803 1883 2973
rect 1876 2796 1903 2803
rect 1776 2776 1783 2780
rect 1896 2776 1903 2796
rect 1933 2780 1947 2793
rect 1936 2776 1943 2780
rect 1756 2667 1763 2743
rect 1813 2707 1827 2713
rect 1647 2593 1653 2607
rect 1556 2440 1563 2443
rect 1553 2427 1567 2440
rect 1516 2327 1523 2413
rect 1536 2327 1543 2333
rect 1536 2313 1553 2327
rect 1536 2256 1543 2313
rect 1616 2268 1623 2553
rect 1816 2476 1823 2573
rect 1836 2488 1843 2772
rect 1876 2740 1883 2743
rect 1856 2687 1863 2732
rect 1873 2727 1887 2740
rect 1916 2707 1923 2743
rect 1916 2667 1923 2693
rect 1976 2647 1983 2773
rect 1716 2446 1723 2473
rect 1856 2367 1863 2513
rect 1876 2447 1883 2533
rect 1976 2476 1983 2573
rect 1996 2487 2003 2813
rect 2036 2803 2043 2873
rect 2016 2796 2043 2803
rect 2016 2776 2023 2796
rect 2036 2607 2043 2633
rect 1916 2407 1923 2443
rect 1516 1983 1523 2223
rect 1576 2187 1583 2253
rect 1636 2147 1643 2223
rect 1676 2127 1683 2273
rect 1696 2207 1703 2353
rect 1736 2256 1743 2353
rect 1496 1976 1523 1983
rect 1496 1956 1503 1976
rect 1536 1956 1543 1993
rect 1576 1967 1583 2013
rect 1396 1887 1403 1923
rect 1456 1887 1463 1953
rect 1476 1847 1483 1913
rect 1516 1887 1523 1923
rect 1367 1796 1383 1803
rect 1096 1647 1103 1692
rect 1296 1667 1303 1703
rect 1176 1436 1243 1443
rect 1136 1400 1143 1403
rect 1133 1387 1147 1400
rect 736 927 743 1113
rect 616 867 623 914
rect 756 887 763 1173
rect 776 1147 783 1183
rect 916 1180 923 1183
rect 913 1167 927 1180
rect 996 1167 1003 1233
rect 1036 1216 1043 1273
rect 1136 1247 1143 1273
rect 1096 1180 1103 1183
rect 873 920 887 933
rect 876 916 883 920
rect 676 863 683 883
rect 656 856 683 863
rect 656 696 663 856
rect 576 656 603 663
rect 576 467 583 656
rect 236 227 243 363
rect 296 188 303 413
rect 320 406 340 407
rect 327 403 340 406
rect 327 396 343 403
rect 373 400 387 413
rect 376 396 383 400
rect 327 393 340 396
rect 356 327 363 363
rect 416 147 423 353
rect 436 188 443 413
rect 456 366 463 393
rect 576 366 583 432
rect 596 407 603 633
rect 676 587 683 663
rect 736 627 743 813
rect 776 707 783 914
rect 796 787 803 873
rect 816 847 823 883
rect 856 880 863 883
rect 853 867 867 880
rect 916 707 923 1033
rect 936 827 943 873
rect 956 787 963 883
rect 996 880 1003 883
rect 993 867 1007 880
rect 1056 847 1063 1172
rect 1093 1167 1107 1180
rect 1136 1167 1143 1233
rect 1216 1216 1223 1313
rect 1196 1180 1203 1183
rect 1193 1167 1207 1180
rect 1076 867 1083 993
rect 1096 883 1103 1113
rect 1096 876 1123 883
rect 996 747 1003 813
rect 1156 807 1163 843
rect 956 696 963 733
rect 996 696 1003 733
rect 1176 707 1183 833
rect 796 660 803 663
rect 836 660 843 663
rect 793 647 807 660
rect 833 647 847 660
rect 676 396 683 453
rect 787 416 823 423
rect 496 188 503 213
rect 536 147 543 363
rect 136 -24 143 143
rect 216 -24 223 143
rect 336 -24 343 143
rect 576 107 583 352
rect 596 176 603 353
rect 656 227 663 363
rect 716 227 723 413
rect 816 396 823 416
rect 736 327 743 393
rect 856 267 863 453
rect 876 447 883 693
rect 936 660 943 663
rect 933 647 947 660
rect 976 647 983 663
rect 1036 647 1043 694
rect 1196 666 1203 773
rect 1236 763 1243 1436
rect 1256 1427 1263 1553
rect 1336 1501 1343 1693
rect 1356 1507 1363 1772
rect 1376 1743 1383 1796
rect 1376 1736 1403 1743
rect 1436 1736 1443 1813
rect 1476 1736 1483 1833
rect 1496 1743 1503 1813
rect 1516 1767 1523 1873
rect 1556 1743 1563 1923
rect 1596 1827 1603 2053
rect 1696 1956 1703 2053
rect 1736 1926 1743 2133
rect 1756 2023 1763 2223
rect 1796 2047 1803 2333
rect 1833 2283 1847 2293
rect 1816 2280 1847 2283
rect 1816 2276 1843 2280
rect 1816 2147 1823 2276
rect 1876 2256 1883 2313
rect 1936 2283 1943 2393
rect 1956 2347 1963 2443
rect 1996 2387 2003 2433
rect 2016 2307 2023 2553
rect 2036 2487 2043 2513
rect 2056 2507 2063 2743
rect 2076 2627 2083 2833
rect 2096 2726 2103 2853
rect 2116 2707 2123 3113
rect 2136 2847 2143 2973
rect 2156 2947 2163 2983
rect 2156 2827 2163 2933
rect 2176 2867 2183 3033
rect 2216 2980 2223 2983
rect 2213 2967 2227 2980
rect 2236 2963 2243 3173
rect 2256 3027 2263 3233
rect 2336 3127 2343 3393
rect 2396 3187 2403 3653
rect 2416 3567 2423 3613
rect 2456 3607 2463 3673
rect 2416 3267 2423 3453
rect 2436 3387 2443 3503
rect 2456 3427 2463 3593
rect 2516 3503 2523 3756
rect 2496 3496 2523 3503
rect 2496 3427 2503 3496
rect 2273 3020 2287 3033
rect 2276 3016 2283 3020
rect 2416 2983 2423 3033
rect 2436 3007 2443 3294
rect 2456 3087 2463 3333
rect 2476 3260 2483 3263
rect 2473 3247 2487 3260
rect 2536 3187 2543 3693
rect 2556 3307 2563 3773
rect 2227 2956 2243 2963
rect 2253 2760 2267 2773
rect 2256 2756 2263 2760
rect 2096 2507 2103 2593
rect 2136 2567 2143 2733
rect 2056 2476 2063 2493
rect 2096 2476 2103 2493
rect 2076 2407 2083 2443
rect 2136 2427 2143 2493
rect 2156 2487 2163 2653
rect 2176 2647 2183 2743
rect 2276 2687 2283 2953
rect 2296 2907 2303 2973
rect 2316 2947 2323 2983
rect 2416 2976 2443 2983
rect 2556 2827 2563 2873
rect 2376 2760 2383 2763
rect 2356 2703 2363 2753
rect 2373 2747 2387 2760
rect 2356 2696 2383 2703
rect 2376 2607 2383 2696
rect 2516 2647 2523 2793
rect 2556 2756 2563 2813
rect 2576 2747 2583 3853
rect 2596 3787 2603 3976
rect 2616 3927 2623 3973
rect 2656 3907 2663 3973
rect 2616 3827 2623 3892
rect 2696 3828 2703 3952
rect 2636 3767 2643 3783
rect 2647 3756 2663 3763
rect 2596 3483 2603 3633
rect 2656 3528 2663 3756
rect 2676 3547 2683 3783
rect 2696 3523 2703 3733
rect 2716 3587 2723 4053
rect 2773 4040 2787 4053
rect 2776 4036 2783 4040
rect 2736 3963 2743 3993
rect 2756 3967 2763 4003
rect 2736 3956 2752 3963
rect 2736 3867 2743 3893
rect 2776 3887 2783 3953
rect 2796 3907 2803 4003
rect 2776 3847 2783 3873
rect 2836 3827 2843 3993
rect 2856 3967 2863 4073
rect 2876 4047 2883 4153
rect 2896 4036 2903 4093
rect 2936 4048 2943 4216
rect 2873 3983 2887 3993
rect 2873 3980 2903 3983
rect 2876 3976 2903 3980
rect 2876 3807 2883 3933
rect 2896 3796 2903 3976
rect 2736 3687 2743 3773
rect 2796 3727 2803 3753
rect 2816 3687 2823 3783
rect 2856 3707 2863 3763
rect 2876 3623 2883 3753
rect 2896 3627 2903 3673
rect 2916 3647 2923 3953
rect 2976 3947 2983 4034
rect 2996 4007 3003 4233
rect 3036 4067 3043 4293
rect 3056 4247 3063 4733
rect 3076 4587 3083 4756
rect 3156 4747 3163 5253
rect 3176 5187 3183 5293
rect 3196 5287 3203 5316
rect 3196 5088 3203 5133
rect 3216 5107 3223 5173
rect 3296 5107 3303 5343
rect 3316 5083 3323 5233
rect 3336 5227 3343 5374
rect 3336 5127 3343 5213
rect 3356 5187 3363 5513
rect 3376 5387 3383 5563
rect 3416 5503 3423 5753
rect 3436 5527 3443 5673
rect 3556 5667 3563 5753
rect 3576 5643 3583 5836
rect 3636 5727 3643 5813
rect 3656 5787 3663 5953
rect 3556 5636 3583 5643
rect 3476 5527 3483 5563
rect 3556 5547 3563 5636
rect 3636 5607 3643 5713
rect 3620 5563 3633 5567
rect 3616 5556 3633 5563
rect 3620 5553 3633 5556
rect 3656 5547 3663 5653
rect 3676 5647 3683 6153
rect 3736 6080 3743 6083
rect 3733 6067 3747 6080
rect 3776 5967 3783 6133
rect 3813 6120 3827 6133
rect 3816 6116 3823 6120
rect 3856 6116 3863 6233
rect 3976 6163 3983 6303
rect 4116 6167 4123 6303
rect 3956 6156 3983 6163
rect 3876 6080 3883 6083
rect 3873 6067 3887 6080
rect 3847 6055 3873 6062
rect 3856 5896 3863 5973
rect 3896 5896 3903 6053
rect 3916 6007 3923 6073
rect 3936 6067 3943 6113
rect 3956 6087 3963 6156
rect 4116 6116 4123 6153
rect 4156 6116 4163 6153
rect 4216 6086 4223 6113
rect 4316 6087 4323 6153
rect 3696 5856 3723 5863
rect 3696 5827 3703 5856
rect 3756 5687 3763 5863
rect 3776 5767 3783 5833
rect 3816 5727 3823 5893
rect 3876 5860 3883 5863
rect 3873 5847 3887 5860
rect 3776 5667 3783 5713
rect 3756 5627 3763 5652
rect 3816 5647 3823 5713
rect 3716 5560 3723 5563
rect 3416 5496 3443 5503
rect 3396 5376 3403 5433
rect 3436 5376 3443 5496
rect 3473 5407 3487 5413
rect 3460 5343 3473 5347
rect 3416 5340 3423 5343
rect 3356 5103 3363 5173
rect 3376 5143 3383 5333
rect 3413 5327 3427 5340
rect 3456 5336 3473 5343
rect 3460 5333 3473 5336
rect 3396 5267 3403 5313
rect 3436 5247 3443 5313
rect 3476 5287 3483 5312
rect 3467 5266 3480 5267
rect 3467 5253 3473 5266
rect 3436 5147 3443 5173
rect 3376 5136 3393 5143
rect 3307 5076 3323 5083
rect 3336 5096 3363 5103
rect 3336 5076 3343 5096
rect 3376 5083 3383 5112
rect 3396 5107 3403 5133
rect 3376 5076 3403 5083
rect 3456 5076 3463 5153
rect 3476 5127 3483 5232
rect 3496 5207 3503 5453
rect 3516 5187 3523 5531
rect 3676 5467 3683 5553
rect 3713 5547 3727 5560
rect 3696 5467 3703 5513
rect 3756 5507 3763 5553
rect 3536 5387 3543 5413
rect 3567 5394 3573 5407
rect 3560 5393 3580 5394
rect 3613 5380 3627 5393
rect 3616 5376 3623 5380
rect 3736 5376 3743 5413
rect 3556 5340 3563 5343
rect 3553 5327 3567 5340
rect 3636 5340 3643 5343
rect 3633 5327 3647 5340
rect 3616 5316 3633 5323
rect 3533 5247 3547 5253
rect 3296 5047 3303 5072
rect 3260 5043 3273 5047
rect 3176 4727 3183 4854
rect 3196 4847 3203 5013
rect 3216 4947 3223 5043
rect 3256 5036 3273 5043
rect 3260 5033 3273 5036
rect 3316 4827 3323 5013
rect 3356 4967 3363 5043
rect 3396 5043 3403 5076
rect 3396 5036 3423 5043
rect 3436 5040 3443 5043
rect 3376 4987 3383 5033
rect 3336 4867 3343 4913
rect 3416 4907 3423 5036
rect 3433 5027 3447 5040
rect 3476 5007 3483 5043
rect 3236 4787 3243 4823
rect 3276 4727 3283 4823
rect 3347 4823 3360 4827
rect 3476 4826 3483 4972
rect 3536 4947 3543 5153
rect 3516 4856 3523 4913
rect 3556 4868 3563 5173
rect 3596 5147 3603 5273
rect 3596 5076 3603 5133
rect 3616 5127 3623 5316
rect 3656 5287 3663 5332
rect 3633 5080 3647 5093
rect 3656 5087 3663 5233
rect 3676 5183 3683 5374
rect 3696 5267 3703 5313
rect 3716 5280 3723 5343
rect 3756 5307 3763 5332
rect 3776 5280 3783 5632
rect 3833 5600 3847 5613
rect 3836 5596 3843 5600
rect 3876 5596 3883 5633
rect 3896 5607 3903 5773
rect 3916 5747 3923 5813
rect 3796 5343 3803 5513
rect 3816 5447 3823 5563
rect 3916 5563 3923 5733
rect 3936 5707 3943 5753
rect 3956 5687 3963 5893
rect 3976 5847 3983 6033
rect 3996 5907 4003 6072
rect 4036 5908 4043 5933
rect 4076 5896 4083 5993
rect 4196 5896 4203 5933
rect 4216 5927 4223 6072
rect 4276 5987 4283 6083
rect 4316 6047 4323 6073
rect 4016 5727 4023 5863
rect 3936 5608 3943 5653
rect 4016 5596 4023 5653
rect 4056 5607 4063 5863
rect 3896 5556 3923 5563
rect 3896 5527 3903 5556
rect 3936 5403 3943 5594
rect 3996 5507 4003 5563
rect 4036 5543 4043 5563
rect 4016 5536 4043 5543
rect 4016 5467 4023 5536
rect 3927 5396 3943 5403
rect 3796 5336 3823 5343
rect 3716 5273 3783 5280
rect 3716 5247 3723 5273
rect 3676 5176 3703 5183
rect 3636 5076 3643 5080
rect 3656 4967 3663 5033
rect 3676 4987 3683 5073
rect 3696 4883 3703 5176
rect 3716 5087 3723 5193
rect 3736 5147 3743 5213
rect 3727 5083 3740 5087
rect 3727 5076 3743 5083
rect 3776 5076 3783 5113
rect 3796 5107 3803 5213
rect 3816 5087 3823 5336
rect 3727 5073 3740 5076
rect 3800 5044 3813 5047
rect 3716 4903 3723 5033
rect 3756 4947 3763 5043
rect 3796 5033 3813 5044
rect 3716 4896 3743 4903
rect 3696 4876 3723 4883
rect 3347 4816 3363 4823
rect 3347 4813 3360 4816
rect 3436 4787 3443 4823
rect 3476 4767 3483 4812
rect 3136 4556 3143 4613
rect 3176 4568 3183 4653
rect 3076 4307 3083 4513
rect 3116 4487 3123 4523
rect 3176 4507 3183 4554
rect 3216 4520 3223 4523
rect 3196 4447 3203 4513
rect 3213 4507 3227 4520
rect 3276 4507 3283 4713
rect 3316 4627 3323 4733
rect 3576 4687 3583 4823
rect 3596 4787 3603 4813
rect 3616 4747 3623 4854
rect 3380 4523 3393 4527
rect 3336 4487 3343 4523
rect 3376 4516 3393 4523
rect 3380 4513 3393 4516
rect 3416 4507 3423 4673
rect 3436 4527 3443 4633
rect 3476 4627 3483 4653
rect 3456 4563 3463 4593
rect 3456 4556 3483 4563
rect 3516 4556 3523 4653
rect 3173 4347 3187 4353
rect 3116 4227 3123 4303
rect 3107 4213 3113 4227
rect 3056 4087 3063 4212
rect 3056 4036 3063 4073
rect 3016 3967 3023 4003
rect 3076 3947 3083 4213
rect 3096 4127 3103 4153
rect 3096 3967 3103 4023
rect 3076 3946 3100 3947
rect 3076 3936 3093 3946
rect 3080 3933 3093 3936
rect 3116 3907 3123 4013
rect 3136 3927 3143 4272
rect 3156 4207 3163 4303
rect 3156 4016 3183 4023
rect 3016 3783 3023 3803
rect 2996 3776 3023 3783
rect 2996 3747 3003 3776
rect 3016 3703 3023 3753
rect 3156 3747 3163 3993
rect 3176 3987 3183 4016
rect 3176 3803 3183 3973
rect 3196 3847 3203 4353
rect 3236 4336 3243 4433
rect 3273 4340 3287 4353
rect 3276 4336 3283 4340
rect 3356 4327 3363 4353
rect 3376 4316 3383 4493
rect 3496 4467 3503 4523
rect 3576 4467 3583 4673
rect 3596 4487 3603 4593
rect 3616 4556 3623 4733
rect 3213 4287 3227 4292
rect 3256 4227 3263 4303
rect 3316 4207 3323 4233
rect 3396 4167 3403 4353
rect 3496 4167 3503 4273
rect 3636 4227 3643 4453
rect 3656 4447 3663 4523
rect 3676 4383 3683 4753
rect 3716 4627 3723 4876
rect 3736 4583 3743 4896
rect 3796 4867 3803 5033
rect 3816 4868 3823 5012
rect 3816 4827 3823 4854
rect 3756 4767 3763 4823
rect 3796 4687 3803 4813
rect 3836 4787 3843 5253
rect 3896 5247 3903 5373
rect 3916 5347 3923 5393
rect 3973 5380 3987 5393
rect 3976 5376 3983 5380
rect 4016 5376 4023 5413
rect 3996 5307 4003 5343
rect 3896 5076 3903 5113
rect 3936 5087 3943 5193
rect 3920 5043 3933 5047
rect 3856 4987 3863 5033
rect 3876 4963 3883 5043
rect 3916 5036 3933 5043
rect 3920 5033 3933 5036
rect 3956 5027 3963 5153
rect 3976 5107 3983 5273
rect 3976 5047 3983 5093
rect 4007 5083 4020 5087
rect 4056 5083 4063 5453
rect 4076 5407 4083 5673
rect 4116 5667 4123 5894
rect 4256 5866 4263 5913
rect 4216 5827 4223 5863
rect 4107 5603 4120 5607
rect 4107 5596 4123 5603
rect 4107 5593 4120 5596
rect 4096 5427 4103 5553
rect 4156 5467 4163 5533
rect 4196 5527 4203 5594
rect 4176 5387 4183 5433
rect 4076 5346 4083 5372
rect 4196 5347 4203 5453
rect 4096 5127 4103 5333
rect 4116 5287 4123 5343
rect 4136 5227 4143 5253
rect 4007 5076 4023 5083
rect 4056 5076 4073 5083
rect 4007 5073 4020 5076
rect 4176 5087 4183 5173
rect 4196 5147 4203 5312
rect 4216 5187 4223 5613
rect 4256 5608 4263 5653
rect 4276 5627 4283 5933
rect 4336 5896 4343 5933
rect 4296 5727 4303 5793
rect 4316 5787 4323 5863
rect 4356 5603 4363 6302
rect 4416 6123 4423 6303
rect 4616 6207 4623 6303
rect 4416 6116 4443 6123
rect 4436 5927 4443 6116
rect 4556 6116 4563 6153
rect 4596 6087 4603 6114
rect 4496 6027 4503 6083
rect 4536 5987 4543 6072
rect 4396 5647 4403 5913
rect 4453 5900 4467 5913
rect 4456 5896 4463 5900
rect 4536 5863 4543 5973
rect 4596 5927 4603 6073
rect 4616 5903 4623 6193
rect 4656 6116 4663 6173
rect 5247 6156 5273 6163
rect 4716 6047 4723 6083
rect 4756 6047 4763 6153
rect 4796 6116 4803 6153
rect 4927 6116 4943 6123
rect 4596 5896 4623 5903
rect 4436 5827 4443 5863
rect 4536 5856 4563 5863
rect 4636 5847 4643 6033
rect 4816 5987 4823 6072
rect 4656 5847 4663 5933
rect 4716 5896 4723 5973
rect 4856 5896 4863 5993
rect 4916 5927 4923 6114
rect 4696 5847 4703 5863
rect 4696 5647 4703 5833
rect 4736 5787 4743 5863
rect 4336 5596 4363 5603
rect 4276 5467 4283 5563
rect 4336 5547 4343 5596
rect 4396 5527 4403 5553
rect 4436 5507 4443 5563
rect 4256 5340 4263 5343
rect 4296 5340 4303 5343
rect 4233 5327 4247 5333
rect 4253 5327 4267 5340
rect 4293 5327 4307 5340
rect 4376 5287 4383 5493
rect 4456 5407 4463 5633
rect 4696 5596 4723 5603
rect 4413 5380 4427 5393
rect 4416 5376 4423 5380
rect 4256 5167 4263 5273
rect 4036 5040 4043 5043
rect 4033 5027 4047 5040
rect 4046 5020 4047 5027
rect 3856 4956 3883 4963
rect 3856 4907 3863 4956
rect 3856 4727 3863 4893
rect 3916 4856 3923 4913
rect 3696 4576 3743 4583
rect 3696 4407 3703 4576
rect 3793 4560 3807 4573
rect 3796 4556 3803 4560
rect 3676 4376 3703 4383
rect 3653 4323 3667 4333
rect 3653 4320 3683 4323
rect 3656 4316 3683 4320
rect 3696 4187 3703 4376
rect 3716 4327 3723 4473
rect 3756 4447 3763 4493
rect 3776 4463 3783 4523
rect 3836 4507 3843 4673
rect 3876 4588 3883 4823
rect 3896 4687 3903 4793
rect 3936 4767 3943 4823
rect 3913 4560 3927 4573
rect 3956 4567 3963 4973
rect 3976 4587 3983 4953
rect 3996 4807 4003 5013
rect 4056 4927 4063 5013
rect 4076 4907 4083 5074
rect 4056 4820 4063 4823
rect 4053 4807 4067 4820
rect 4076 4803 4083 4872
rect 4096 4827 4103 4893
rect 4116 4887 4123 4973
rect 4136 4856 4143 4913
rect 4156 4887 4163 5033
rect 4176 4927 4183 5052
rect 4196 4987 4203 5112
rect 4273 5080 4287 5093
rect 4276 5076 4283 5080
rect 4176 4856 4183 4892
rect 4236 4867 4243 5043
rect 4296 4856 4303 5133
rect 4313 5107 4327 5113
rect 4316 4967 4323 5072
rect 4336 4947 4343 5253
rect 4416 5247 4423 5313
rect 4367 5113 4373 5127
rect 4396 5103 4403 5153
rect 4376 5096 4403 5103
rect 4376 5088 4383 5096
rect 4416 5076 4423 5233
rect 4436 5207 4443 5343
rect 4456 5067 4463 5333
rect 4396 5027 4403 5043
rect 4396 4987 4403 5013
rect 4313 4867 4327 4873
rect 4476 4863 4483 5513
rect 4496 5387 4503 5413
rect 4516 5340 4523 5343
rect 4513 5327 4527 5340
rect 4556 5287 4563 5343
rect 4576 5307 4583 5333
rect 4596 5263 4603 5493
rect 4636 5487 4643 5594
rect 4656 5527 4663 5552
rect 4616 5387 4623 5453
rect 4676 5376 4683 5473
rect 4696 5427 4703 5513
rect 4716 5387 4723 5596
rect 4616 5346 4623 5373
rect 4736 5343 4743 5713
rect 4776 5667 4783 5893
rect 4916 5866 4923 5913
rect 4956 5896 4963 6072
rect 4993 5900 5007 5913
rect 5016 5907 5023 6153
rect 5136 6116 5143 6153
rect 5196 6087 5203 6153
rect 5300 6123 5313 6127
rect 5296 6116 5313 6123
rect 5300 6113 5313 6116
rect 5536 6116 5543 6173
rect 5636 6116 5643 6173
rect 5676 6128 5683 6153
rect 5156 5987 5163 6083
rect 5336 6086 5343 6113
rect 5167 5976 5183 5983
rect 4996 5896 5003 5900
rect 5036 5867 5043 5913
rect 5073 5900 5087 5913
rect 5076 5896 5083 5900
rect 5153 5907 5167 5913
rect 5176 5867 5183 5976
rect 5236 5927 5243 6083
rect 5256 5927 5263 5973
rect 4836 5860 4843 5863
rect 4833 5847 4847 5860
rect 5096 5860 5103 5863
rect 4816 5608 4823 5633
rect 4796 5376 4803 5433
rect 4836 5376 4843 5733
rect 4876 5623 4883 5852
rect 5093 5847 5107 5860
rect 4856 5616 4883 5623
rect 4856 5527 4863 5616
rect 4936 5596 4943 5653
rect 5073 5600 5087 5613
rect 5176 5608 5183 5832
rect 5196 5627 5203 5913
rect 5253 5900 5267 5913
rect 5256 5896 5263 5900
rect 5336 5866 5343 6072
rect 5356 6007 5363 6113
rect 5396 5896 5403 5993
rect 5416 5927 5423 6083
rect 5456 6047 5463 6114
rect 5573 6047 5587 6053
rect 5556 5896 5563 5933
rect 5476 5866 5483 5893
rect 5236 5747 5243 5863
rect 5256 5703 5263 5773
rect 5276 5727 5283 5863
rect 5576 5787 5583 5863
rect 5256 5696 5283 5703
rect 5207 5616 5223 5623
rect 5076 5596 5083 5600
rect 4876 5566 4883 5593
rect 4856 5407 4863 5513
rect 4976 5507 4983 5594
rect 5216 5596 5223 5616
rect 5116 5566 5123 5593
rect 5016 5447 5023 5563
rect 4616 5287 4623 5332
rect 4696 5307 4703 5343
rect 4716 5336 4743 5343
rect 4647 5293 4653 5307
rect 4596 5256 4623 5263
rect 4516 5167 4523 5213
rect 4536 5076 4543 5113
rect 4573 5080 4587 5093
rect 4576 5076 4583 5080
rect 4616 5047 4623 5256
rect 4716 5227 4723 5336
rect 4516 4987 4523 5043
rect 4636 5027 4643 5173
rect 4736 5127 4743 5233
rect 4756 5187 4763 5332
rect 4776 5287 4783 5343
rect 4696 5076 4703 5113
rect 4556 4947 4563 4973
rect 4456 4856 4483 4863
rect 4516 4856 4523 4893
rect 4156 4820 4163 4823
rect 4196 4820 4203 4823
rect 4153 4807 4167 4820
rect 4076 4796 4103 4803
rect 3916 4556 3923 4560
rect 3776 4456 3803 4463
rect 3736 4316 3743 4373
rect 3756 4207 3763 4433
rect 3796 4407 3803 4456
rect 3816 4387 3823 4453
rect 3876 4403 3883 4493
rect 3896 4427 3903 4523
rect 3936 4507 3943 4523
rect 3976 4507 3983 4573
rect 3936 4496 3953 4507
rect 3940 4493 3953 4496
rect 3876 4396 3903 4403
rect 3776 4347 3783 4373
rect 3333 4020 3347 4033
rect 3336 4016 3343 4020
rect 3436 3987 3443 4153
rect 3496 4056 3503 4153
rect 3536 4027 3543 4153
rect 3176 3796 3193 3803
rect 3016 3696 3043 3703
rect 3036 3683 3043 3696
rect 3036 3676 3063 3683
rect 2856 3616 2883 3623
rect 2736 3567 2743 3613
rect 2676 3516 2703 3523
rect 2796 3516 2803 3573
rect 2596 3476 2623 3483
rect 2596 3147 2603 3413
rect 2616 3296 2623 3476
rect 2656 3207 2663 3263
rect 2676 3167 2683 3516
rect 2696 3347 2703 3493
rect 2756 3427 2763 3483
rect 2756 3367 2763 3413
rect 2776 3347 2783 3433
rect 2796 3407 2803 3453
rect 2596 2847 2603 2973
rect 2616 2887 2623 2983
rect 2616 2756 2623 2852
rect 2176 2476 2183 2533
rect 2216 2476 2223 2533
rect 2276 2446 2283 2493
rect 2316 2476 2323 2593
rect 2516 2527 2523 2633
rect 2636 2607 2643 3153
rect 2656 2976 2673 2983
rect 2396 2516 2413 2523
rect 1916 2276 1943 2283
rect 1916 2223 1923 2276
rect 1896 2216 1923 2223
rect 1876 2067 1883 2153
rect 1756 2016 1803 2023
rect 1756 1996 1773 2003
rect 1496 1736 1523 1743
rect 1456 1667 1463 1703
rect 1516 1667 1523 1736
rect 1536 1736 1563 1743
rect 1277 1494 1343 1501
rect 1277 1404 1284 1494
rect 1396 1443 1403 1533
rect 1536 1507 1543 1736
rect 1636 1747 1643 1912
rect 1676 1887 1683 1923
rect 1567 1703 1580 1707
rect 1567 1696 1583 1703
rect 1616 1700 1623 1703
rect 1567 1693 1580 1696
rect 1613 1687 1627 1700
rect 1376 1436 1403 1443
rect 1256 928 1263 1313
rect 1316 1287 1323 1363
rect 1396 1347 1403 1436
rect 1436 1403 1443 1493
rect 1436 1396 1463 1403
rect 1436 1267 1443 1396
rect 1576 1387 1583 1653
rect 1296 1180 1303 1183
rect 1293 1167 1307 1180
rect 1336 1127 1343 1183
rect 1376 1167 1383 1253
rect 1456 1216 1463 1333
rect 1496 1327 1503 1363
rect 1496 1216 1503 1253
rect 1576 1216 1583 1373
rect 1596 1243 1603 1453
rect 1616 1448 1623 1493
rect 1636 1467 1643 1693
rect 1656 1687 1663 1793
rect 1736 1763 1743 1833
rect 1756 1807 1763 1996
rect 1776 1956 1783 1993
rect 1796 1987 1803 2016
rect 1836 1963 1843 2053
rect 1836 1956 1863 1963
rect 1736 1756 1763 1763
rect 1756 1736 1763 1756
rect 1796 1706 1803 1893
rect 1856 1887 1863 1956
rect 1876 1787 1883 2053
rect 1956 2047 1963 2213
rect 1976 2187 1983 2223
rect 1976 2107 1983 2173
rect 1996 2147 2003 2193
rect 2016 2167 2023 2223
rect 2020 2143 2033 2147
rect 2016 2133 2033 2143
rect 2016 2087 2023 2133
rect 1896 1926 1903 2013
rect 1916 1967 1923 2033
rect 1956 1987 1963 2033
rect 2016 1987 2023 2033
rect 2036 2007 2043 2112
rect 2056 2047 2063 2253
rect 2076 2067 2083 2273
rect 2096 2267 2103 2413
rect 2116 2287 2123 2393
rect 2176 2267 2183 2353
rect 2216 2307 2223 2413
rect 2236 2347 2243 2443
rect 2336 2407 2343 2443
rect 2216 2296 2233 2307
rect 2220 2293 2233 2296
rect 2276 2256 2283 2353
rect 2356 2267 2363 2333
rect 2116 2220 2123 2223
rect 1956 1956 1963 1973
rect 1813 1747 1827 1753
rect 1836 1736 1843 1773
rect 1916 1747 1923 1913
rect 1936 1847 1943 1923
rect 1976 1887 1983 1923
rect 2016 1767 2023 1913
rect 1696 1700 1703 1703
rect 1656 1487 1663 1673
rect 1627 1436 1643 1443
rect 1676 1436 1683 1693
rect 1693 1687 1707 1700
rect 1616 1267 1623 1393
rect 1656 1363 1663 1403
rect 1636 1356 1663 1363
rect 1596 1236 1623 1243
rect 1616 1216 1623 1236
rect 1636 1227 1643 1356
rect 1396 1186 1403 1213
rect 1476 1180 1483 1183
rect 1473 1167 1487 1180
rect 1536 1047 1543 1213
rect 1296 916 1303 953
rect 1336 916 1343 973
rect 1396 886 1403 973
rect 1216 756 1243 763
rect 976 607 983 633
rect 1076 607 1083 663
rect 1116 627 1123 663
rect 896 360 903 363
rect 893 347 907 360
rect 936 287 943 363
rect 796 146 803 213
rect 996 203 1003 493
rect 1016 347 1023 593
rect 1216 430 1223 756
rect 1236 696 1243 733
rect 1296 667 1303 733
rect 1316 507 1323 883
rect 1336 707 1343 833
rect 1356 827 1363 883
rect 1396 696 1403 733
rect 1456 666 1463 773
rect 1536 747 1543 873
rect 1556 847 1563 883
rect 1376 660 1383 663
rect 1336 443 1343 653
rect 1373 647 1387 660
rect 1416 527 1423 652
rect 1453 647 1467 652
rect 1536 527 1543 663
rect 1136 423 1223 430
rect 1316 436 1343 443
rect 1316 427 1323 436
rect 1036 327 1043 353
rect 1076 267 1083 363
rect 1116 287 1123 353
rect 833 180 847 193
rect 976 196 1003 203
rect 836 176 843 180
rect 636 -24 643 143
rect 756 107 763 143
rect 856 107 863 143
rect 896 140 903 143
rect 893 127 907 140
rect 976 127 983 196
rect 1036 176 1043 213
rect 1096 146 1103 213
rect 996 107 1003 143
rect 756 47 763 93
rect 1056 47 1063 143
rect 1136 -24 1143 423
rect 1316 396 1323 413
rect 1356 396 1363 453
rect 1216 176 1223 313
rect 1236 307 1243 393
rect 1416 366 1423 413
rect 1453 400 1467 413
rect 1456 396 1463 400
rect 1496 396 1503 433
rect 1576 427 1583 753
rect 1636 696 1643 733
rect 1656 727 1663 1333
rect 1716 1267 1723 1533
rect 1816 1487 1823 1693
rect 1896 1587 1903 1703
rect 1776 1436 1783 1473
rect 1813 1440 1827 1452
rect 1856 1447 1863 1573
rect 1936 1547 1943 1753
rect 1993 1740 2007 1753
rect 2036 1747 2043 1993
rect 2096 1987 2103 2213
rect 2113 2207 2127 2220
rect 2113 2187 2127 2193
rect 2140 2183 2153 2187
rect 2136 2173 2153 2183
rect 2136 2163 2143 2173
rect 2116 2156 2143 2163
rect 2116 2107 2123 2156
rect 2173 2147 2187 2153
rect 2176 2067 2183 2112
rect 2196 2107 2203 2173
rect 2216 2167 2223 2253
rect 2256 2220 2263 2223
rect 2253 2207 2267 2220
rect 2247 2133 2253 2147
rect 2073 1960 2087 1973
rect 2076 1956 2083 1960
rect 2156 1967 2163 2053
rect 2176 1947 2183 2013
rect 2140 1923 2153 1927
rect 2136 1916 2153 1923
rect 2140 1913 2153 1916
rect 1996 1736 2003 1740
rect 1816 1436 1823 1440
rect 1876 1406 1883 1473
rect 1956 1467 1963 1693
rect 2020 1703 2033 1707
rect 2016 1696 2033 1703
rect 2020 1693 2033 1696
rect 2056 1647 2063 1833
rect 1907 1453 1913 1467
rect 1967 1456 1983 1463
rect 1896 1436 1923 1443
rect 1976 1436 1983 1456
rect 1676 867 1683 1253
rect 1756 1216 1763 1253
rect 1796 1227 1803 1403
rect 1836 1400 1843 1403
rect 1833 1387 1847 1400
rect 1896 1347 1903 1436
rect 1996 1267 2003 1473
rect 2016 1407 2023 1613
rect 2036 1367 2043 1453
rect 2076 1436 2083 1893
rect 2176 1847 2183 1912
rect 2196 1827 2203 2013
rect 2276 1956 2283 2053
rect 2296 1963 2303 2223
rect 2336 2216 2363 2223
rect 2356 2107 2363 2216
rect 2376 2167 2383 2453
rect 2396 2226 2403 2516
rect 2416 2476 2423 2513
rect 2456 2268 2463 2432
rect 2496 2256 2503 2373
rect 2536 2267 2543 2533
rect 2596 2476 2603 2573
rect 2636 2488 2643 2513
rect 2656 2487 2663 2976
rect 2696 2963 2703 3293
rect 2736 3260 2743 3263
rect 2733 3247 2747 3260
rect 2776 3207 2783 3263
rect 2816 3127 2823 3533
rect 2856 3467 2863 3616
rect 2916 3516 2923 3573
rect 2936 3547 2943 3573
rect 2896 3467 2903 3483
rect 2856 3347 2863 3373
rect 2896 3367 2903 3453
rect 2896 3296 2903 3332
rect 2936 3296 2943 3353
rect 2836 3263 2843 3293
rect 2996 3283 3003 3653
rect 3016 3387 3023 3593
rect 3036 3407 3043 3633
rect 3056 3516 3063 3676
rect 3176 3647 3183 3753
rect 3216 3647 3223 3913
rect 3236 3807 3243 3833
rect 3256 3803 3263 3893
rect 3256 3796 3283 3803
rect 3236 3667 3243 3753
rect 3176 3607 3183 3633
rect 3220 3583 3233 3587
rect 3216 3573 3233 3583
rect 3216 3516 3223 3573
rect 2976 3276 3023 3283
rect 3036 3276 3043 3393
rect 3096 3387 3103 3483
rect 3116 3467 3123 3514
rect 3176 3427 3183 3483
rect 3236 3407 3243 3514
rect 3256 3447 3263 3733
rect 3276 3707 3283 3796
rect 3276 3587 3283 3693
rect 3296 3687 3303 3913
rect 3316 3627 3323 3814
rect 3336 3587 3343 3772
rect 3356 3727 3363 3873
rect 3307 3573 3313 3587
rect 3336 3516 3343 3573
rect 3376 3548 3383 3613
rect 3396 3607 3403 3653
rect 3416 3627 3423 3783
rect 3056 3287 3063 3373
rect 2836 3256 2883 3263
rect 2836 3107 2843 3233
rect 2916 3207 2923 3263
rect 2676 2956 2703 2963
rect 2676 2447 2683 2956
rect 2716 2947 2723 3093
rect 2736 2788 2743 3053
rect 2756 3047 2763 3093
rect 2756 2996 2783 3003
rect 2756 2827 2763 2996
rect 2836 2963 2843 3093
rect 2896 2986 2903 3173
rect 3016 3167 3023 3276
rect 3076 3143 3083 3333
rect 3316 3227 3323 3433
rect 3396 3303 3403 3473
rect 3396 3296 3423 3303
rect 3416 3246 3423 3296
rect 3436 3263 3443 3952
rect 3456 3907 3463 3933
rect 3536 3863 3543 3992
rect 3556 3947 3563 4033
rect 3576 3967 3583 4093
rect 3596 4047 3603 4173
rect 3696 4047 3703 4152
rect 3776 4063 3783 4093
rect 3796 4087 3803 4353
rect 3833 4348 3847 4353
rect 3856 4267 3863 4303
rect 3816 4063 3823 4113
rect 3776 4056 3823 4063
rect 3836 4056 3843 4153
rect 3856 4107 3863 4193
rect 3753 4040 3767 4053
rect 3756 4036 3763 4040
rect 3796 4036 3803 4056
rect 3716 4007 3723 4034
rect 3616 4000 3623 4003
rect 3527 3856 3543 3863
rect 3596 3863 3603 3993
rect 3613 3987 3627 4000
rect 3616 3907 3623 3952
rect 3656 3947 3663 4003
rect 3696 3867 3703 3893
rect 3736 3887 3743 3993
rect 3853 4003 3867 4013
rect 3836 4000 3867 4003
rect 3836 3996 3863 4000
rect 3596 3856 3623 3863
rect 3516 3816 3523 3853
rect 3476 3647 3483 3813
rect 3580 3783 3593 3787
rect 3576 3776 3593 3783
rect 3580 3773 3593 3776
rect 3536 3747 3543 3772
rect 3616 3747 3623 3856
rect 3633 3827 3647 3833
rect 3776 3816 3783 3893
rect 3816 3816 3823 3993
rect 3836 3927 3843 3996
rect 3876 3943 3883 4023
rect 3896 3987 3903 4396
rect 3916 4347 3923 4493
rect 3976 4336 3983 4413
rect 3996 4407 4003 4753
rect 4056 4607 4063 4653
rect 4056 4556 4063 4593
rect 4096 4523 4103 4796
rect 4193 4807 4207 4820
rect 4233 4807 4247 4813
rect 4276 4807 4283 4823
rect 4267 4796 4283 4807
rect 4267 4793 4280 4796
rect 4116 4647 4123 4793
rect 4136 4767 4143 4793
rect 4316 4747 4323 4813
rect 4416 4767 4423 4823
rect 4033 4507 4047 4512
rect 4076 4516 4103 4523
rect 4116 4523 4123 4633
rect 4196 4556 4203 4653
rect 4256 4567 4263 4733
rect 4236 4527 4243 4554
rect 4316 4556 4323 4693
rect 4116 4516 4143 4523
rect 4056 4306 4063 4393
rect 3916 4167 3923 4293
rect 3996 4267 4003 4303
rect 4076 4207 4083 4516
rect 4136 4336 4143 4516
rect 4116 4283 4123 4303
rect 4116 4276 4143 4283
rect 4136 4227 4143 4276
rect 4156 4247 4163 4303
rect 4196 4287 4203 4334
rect 4216 4267 4223 4513
rect 4296 4467 4303 4523
rect 4293 4340 4307 4353
rect 4296 4336 4303 4340
rect 4336 4306 4343 4413
rect 4356 4387 4363 4713
rect 4376 4527 4383 4673
rect 4436 4667 4443 4813
rect 4456 4727 4463 4856
rect 4416 4556 4423 4633
rect 4496 4607 4503 4823
rect 4536 4767 4543 4823
rect 4576 4647 4583 4813
rect 4356 4287 4363 4352
rect 4413 4340 4427 4353
rect 4456 4347 4463 4473
rect 4516 4427 4523 4613
rect 4596 4567 4603 4933
rect 4676 4907 4683 5043
rect 4716 5007 4723 5043
rect 4613 4867 4627 4873
rect 4696 4856 4703 4953
rect 4636 4707 4643 4812
rect 4676 4787 4683 4823
rect 4636 4587 4643 4693
rect 4716 4627 4723 4813
rect 4736 4767 4743 4873
rect 4756 4867 4763 5033
rect 4776 5007 4783 5093
rect 4796 4887 4803 5173
rect 4816 5127 4823 5343
rect 4896 5287 4903 5433
rect 5016 5407 5023 5433
rect 4953 5380 4967 5393
rect 4956 5376 4963 5380
rect 5053 5380 5067 5393
rect 5056 5376 5063 5380
rect 4916 5307 4923 5333
rect 4936 5247 4943 5343
rect 4836 5107 4843 5133
rect 4936 5047 4943 5074
rect 4767 4856 4783 4863
rect 4733 4560 4747 4573
rect 4756 4567 4763 4813
rect 4816 4823 4823 4953
rect 4836 4867 4843 5043
rect 4856 4867 4863 5013
rect 4876 5007 4883 5043
rect 4896 4856 4903 4893
rect 4816 4816 4843 4823
rect 4793 4567 4807 4573
rect 4736 4556 4743 4560
rect 4616 4526 4623 4553
rect 4416 4336 4423 4340
rect 3976 4027 3983 4073
rect 3993 4020 4007 4033
rect 3996 4016 4003 4020
rect 3856 3936 3883 3943
rect 3856 3887 3863 3936
rect 3873 3827 3887 3833
rect 3696 3747 3703 3783
rect 3556 3607 3563 3693
rect 3736 3667 3743 3793
rect 3840 3783 3853 3787
rect 3836 3776 3853 3783
rect 3840 3773 3853 3776
rect 3796 3727 3803 3772
rect 3876 3727 3883 3792
rect 3533 3563 3547 3573
rect 3516 3560 3547 3563
rect 3516 3556 3543 3560
rect 3516 3507 3523 3556
rect 3676 3527 3683 3633
rect 3533 3500 3547 3513
rect 3536 3496 3543 3500
rect 3736 3503 3743 3653
rect 3776 3607 3783 3653
rect 3716 3496 3743 3503
rect 3693 3483 3707 3493
rect 3693 3480 3723 3483
rect 3696 3476 3723 3480
rect 3493 3300 3507 3313
rect 3496 3296 3503 3300
rect 3536 3296 3543 3373
rect 3436 3256 3463 3263
rect 3076 3136 3103 3143
rect 2816 2956 2843 2963
rect 2816 2867 2823 2956
rect 2856 2827 2863 2983
rect 2876 2776 2883 2933
rect 2896 2927 2903 2972
rect 2916 2887 2923 2983
rect 2736 2476 2743 2593
rect 2776 2587 2783 2773
rect 2816 2667 2823 2693
rect 2416 2187 2423 2213
rect 2516 2220 2523 2223
rect 2376 2027 2383 2153
rect 2436 2027 2443 2212
rect 2456 2107 2463 2193
rect 2476 2087 2483 2212
rect 2513 2207 2527 2220
rect 2556 2207 2563 2433
rect 2576 2407 2583 2443
rect 2616 2407 2623 2443
rect 2636 2267 2643 2293
rect 2296 1956 2323 1963
rect 2096 1747 2103 1813
rect 2113 1748 2127 1753
rect 2153 1740 2167 1753
rect 2156 1736 2163 1740
rect 2196 1736 2203 1792
rect 2316 1767 2323 1956
rect 2336 1956 2363 1963
rect 2236 1706 2243 1753
rect 2336 1736 2343 1956
rect 2396 1706 2403 1833
rect 2416 1747 2423 1883
rect 2476 1847 2483 2033
rect 2496 1887 2503 2193
rect 2516 1967 2523 2172
rect 2536 1968 2543 2013
rect 2596 1963 2603 2193
rect 2616 1987 2623 2223
rect 2636 2007 2643 2213
rect 2656 2207 2663 2293
rect 2716 2268 2723 2393
rect 2776 2387 2783 2432
rect 2816 2267 2823 2653
rect 2836 2446 2843 2732
rect 2956 2707 2963 3113
rect 3096 2976 3103 3136
rect 3196 3067 3203 3113
rect 2976 2776 2983 2813
rect 2876 2476 2883 2513
rect 2956 2467 2963 2672
rect 3036 2527 3043 2774
rect 3056 2607 3063 2873
rect 3196 2803 3203 3053
rect 3316 2987 3323 3113
rect 3356 2927 3363 3053
rect 3376 3028 3383 3232
rect 3176 2796 3203 2803
rect 3036 2476 3043 2513
rect 2856 2307 2863 2313
rect 2847 2293 2863 2307
rect 2896 2303 2903 2443
rect 2956 2303 2963 2453
rect 3016 2327 3023 2443
rect 3096 2387 3103 2732
rect 3116 2446 3123 2553
rect 3176 2476 3183 2796
rect 3236 2788 3243 2913
rect 3336 2788 3343 2893
rect 3376 2827 3383 2963
rect 3436 2947 3443 3153
rect 3456 3087 3463 3256
rect 3476 3127 3483 3231
rect 3516 3187 3523 3252
rect 3556 3127 3563 3193
rect 3436 2776 3443 2933
rect 3256 2488 3263 2743
rect 3356 2687 3363 2743
rect 3476 2740 3483 2743
rect 3473 2727 3487 2740
rect 3496 2687 3503 3033
rect 3556 2996 3563 3053
rect 3576 2907 3583 3393
rect 3676 3227 3683 3263
rect 3556 2896 3573 2903
rect 3316 2307 3323 2443
rect 2896 2296 2923 2303
rect 2856 2256 2863 2293
rect 2893 2260 2907 2273
rect 2916 2267 2923 2296
rect 2936 2296 2963 2303
rect 2896 2256 2903 2260
rect 2696 2187 2703 2223
rect 2736 2220 2743 2223
rect 2733 2207 2747 2220
rect 2776 2167 2783 2213
rect 2596 1956 2623 1963
rect 2656 1956 2663 2153
rect 2693 1968 2707 1973
rect 2516 1867 2523 1913
rect 2476 1787 2483 1812
rect 2556 1807 2563 1912
rect 2616 1776 2623 1956
rect 2453 1740 2467 1753
rect 2456 1736 2463 1740
rect 2736 1743 2743 1993
rect 2776 1987 2783 2153
rect 2796 2127 2803 2253
rect 2876 2187 2883 2223
rect 2796 1956 2803 2073
rect 2876 1927 2883 2173
rect 2936 2047 2943 2296
rect 3347 2296 3363 2303
rect 2956 2087 2963 2273
rect 2993 2260 3007 2273
rect 2996 2256 3003 2260
rect 3036 2256 3043 2293
rect 3156 2256 3163 2293
rect 3016 2127 3023 2223
rect 3056 2220 3063 2223
rect 3053 2207 3067 2220
rect 2956 1956 2963 1993
rect 2656 1736 2683 1743
rect 2096 1487 2103 1693
rect 2136 1627 2143 1703
rect 2356 1700 2363 1703
rect 2316 1627 2323 1692
rect 2353 1687 2367 1700
rect 2436 1687 2443 1703
rect 2427 1676 2443 1687
rect 2427 1673 2440 1676
rect 2136 1587 2143 1613
rect 2113 1440 2127 1453
rect 2116 1436 2123 1440
rect 2236 1436 2243 1473
rect 2276 1436 2283 1533
rect 2316 1407 2323 1433
rect 1736 987 1743 1183
rect 1793 1183 1807 1192
rect 1916 1186 1923 1253
rect 1793 1180 1843 1183
rect 1796 1176 1843 1180
rect 1776 1127 1783 1173
rect 1980 1183 1993 1187
rect 1976 1176 1993 1183
rect 1980 1173 1993 1176
rect 2016 1186 2023 1273
rect 2047 1223 2060 1227
rect 2047 1216 2063 1223
rect 2096 1216 2103 1353
rect 2136 1227 2143 1403
rect 2047 1213 2060 1216
rect 1796 967 1803 1153
rect 2116 1067 2123 1183
rect 2156 1147 2163 1193
rect 2176 983 2183 1392
rect 2216 1243 2223 1403
rect 2196 1236 2223 1243
rect 2196 1007 2203 1236
rect 2256 1216 2263 1333
rect 2336 1267 2343 1513
rect 2376 1436 2383 1513
rect 2496 1443 2503 1733
rect 2536 1696 2563 1703
rect 2536 1547 2543 1696
rect 2676 1667 2683 1736
rect 2716 1736 2743 1743
rect 2776 1736 2783 1853
rect 2816 1827 2823 1923
rect 2716 1706 2723 1736
rect 2876 1703 2883 1873
rect 3016 1823 3023 2033
rect 3056 1956 3063 2033
rect 3096 1987 3103 2254
rect 3176 2220 3183 2223
rect 3113 2207 3127 2213
rect 3173 2207 3187 2220
rect 3187 2196 3203 2203
rect 3116 1963 3123 2113
rect 3096 1956 3123 1963
rect 2996 1816 3023 1823
rect 2716 1527 2723 1692
rect 2796 1627 2803 1703
rect 2876 1696 2903 1703
rect 2476 1436 2503 1443
rect 2436 1400 2443 1403
rect 2433 1387 2447 1400
rect 2436 1347 2443 1373
rect 2167 976 2183 983
rect 1796 923 1803 953
rect 1776 916 1803 923
rect 1776 886 1783 916
rect 1896 916 1903 973
rect 1736 880 1743 883
rect 1733 867 1747 880
rect 1936 883 1943 914
rect 1716 856 1733 863
rect 1676 827 1683 853
rect 1676 696 1683 753
rect 1716 707 1723 856
rect 1776 743 1783 872
rect 1876 827 1883 883
rect 1936 876 1963 883
rect 1956 803 1963 876
rect 1956 796 1983 803
rect 1776 736 1803 743
rect 1596 587 1603 693
rect 1656 660 1663 663
rect 1653 647 1667 660
rect 1736 447 1743 713
rect 1796 696 1803 736
rect 1893 700 1907 713
rect 1896 696 1903 700
rect 1776 660 1783 663
rect 1773 647 1787 660
rect 1816 408 1823 593
rect 1836 527 1843 693
rect 1876 647 1883 663
rect 1656 396 1703 403
rect 1553 363 1567 373
rect 1696 367 1703 396
rect 1536 360 1567 363
rect 1536 356 1563 360
rect 1296 227 1303 352
rect 1396 307 1403 333
rect 1316 176 1323 253
rect 1416 176 1423 213
rect 1436 207 1443 293
rect 1496 247 1503 333
rect 1516 267 1523 352
rect 1536 327 1543 356
rect 1636 360 1643 363
rect 1633 347 1647 360
rect 1516 227 1523 253
rect 1256 147 1263 174
rect 1536 183 1543 233
rect 1516 176 1543 183
rect 1556 176 1563 213
rect 1576 207 1583 313
rect 1696 307 1703 353
rect 1716 347 1723 394
rect 1756 267 1763 363
rect 1796 327 1803 363
rect 1196 107 1203 143
rect 1496 87 1503 173
rect 1516 146 1523 176
rect 1856 176 1863 393
rect 1876 207 1883 633
rect 1916 627 1923 663
rect 1956 647 1963 713
rect 1976 647 1983 796
rect 1996 707 2003 872
rect 2076 827 2083 914
rect 2096 887 2103 933
rect 2156 916 2163 973
rect 2116 708 2123 833
rect 2136 807 2143 883
rect 2176 847 2183 883
rect 2216 803 2223 1133
rect 2236 847 2243 1153
rect 2276 1147 2283 1183
rect 2356 1167 2363 1214
rect 2273 920 2287 933
rect 2276 916 2283 920
rect 2316 916 2323 1093
rect 2376 883 2383 1293
rect 2476 1287 2483 1436
rect 2796 1436 2803 1533
rect 2816 1487 2823 1553
rect 2836 1527 2843 1653
rect 2956 1627 2963 1703
rect 2976 1647 2983 1734
rect 2996 1607 3003 1816
rect 3076 1807 3083 1923
rect 2836 1436 2843 1513
rect 2736 1407 2743 1434
rect 2516 1347 2523 1403
rect 2527 1336 2543 1343
rect 2396 1067 2403 1253
rect 2436 1216 2443 1273
rect 2536 1186 2543 1336
rect 2556 1228 2563 1403
rect 2636 1400 2643 1403
rect 2616 1228 2623 1393
rect 2633 1387 2647 1400
rect 2456 1167 2463 1183
rect 2556 1167 2563 1214
rect 2596 1180 2603 1183
rect 2593 1167 2607 1180
rect 2436 916 2443 1133
rect 2456 927 2463 1153
rect 2656 1047 2663 1273
rect 2676 1227 2683 1403
rect 2876 1406 2883 1473
rect 2936 1436 2943 1493
rect 3016 1448 3023 1793
rect 3116 1703 3123 1813
rect 3136 1748 3143 2053
rect 3156 1926 3163 1973
rect 3196 1968 3203 2196
rect 3216 2007 3223 2223
rect 3236 1956 3243 1993
rect 3256 1987 3263 2293
rect 3336 2256 3343 2293
rect 3356 2267 3363 2296
rect 3376 2268 3383 2573
rect 3396 2423 3403 2673
rect 3476 2483 3483 2553
rect 3476 2476 3503 2483
rect 3396 2416 3423 2423
rect 3416 2263 3423 2416
rect 3436 2407 3443 2443
rect 3496 2347 3503 2476
rect 3516 2307 3523 2433
rect 3396 2260 3423 2263
rect 3393 2256 3423 2260
rect 3456 2256 3463 2293
rect 3356 2067 3363 2213
rect 3376 2007 3383 2254
rect 3393 2247 3407 2256
rect 3480 2223 3493 2227
rect 3260 1923 3273 1927
rect 3256 1916 3273 1923
rect 3260 1913 3273 1916
rect 3196 1736 3203 1773
rect 3296 1743 3303 1973
rect 3316 1926 3323 1993
rect 3396 1983 3403 2212
rect 3436 2203 3443 2223
rect 3476 2216 3493 2223
rect 3480 2213 3493 2216
rect 3436 2196 3463 2203
rect 3333 1967 3347 1973
rect 3376 1976 3403 1983
rect 3376 1956 3383 1976
rect 3416 1956 3423 2073
rect 3456 2027 3463 2196
rect 3396 1847 3403 1923
rect 3476 1926 3483 1953
rect 3276 1736 3303 1743
rect 3036 1507 3043 1703
rect 3096 1696 3123 1703
rect 3096 1447 3103 1633
rect 3016 1406 3023 1434
rect 3047 1443 3060 1447
rect 3047 1436 3063 1443
rect 3047 1433 3060 1436
rect 2816 1400 2823 1403
rect 2813 1387 2827 1400
rect 2716 1216 2723 1333
rect 2756 1216 2763 1293
rect 2696 1147 2703 1172
rect 2736 1107 2743 1172
rect 2656 987 2663 1033
rect 2207 796 2223 803
rect 2016 660 2023 663
rect 1996 627 2003 653
rect 2013 647 2027 660
rect 1916 396 1923 453
rect 1996 367 2003 613
rect 2056 396 2063 453
rect 2116 407 2123 694
rect 2136 666 2143 793
rect 2196 696 2203 793
rect 2296 787 2303 883
rect 2336 876 2383 883
rect 2406 873 2407 880
rect 2393 863 2407 873
rect 2376 860 2407 863
rect 2376 856 2403 860
rect 2176 660 2183 663
rect 2173 647 2187 660
rect 2216 627 2223 663
rect 2016 367 2023 394
rect 1896 227 1903 353
rect 2076 360 2083 363
rect 2073 347 2087 360
rect 2136 363 2143 613
rect 2216 396 2223 553
rect 2256 467 2263 694
rect 2356 607 2363 753
rect 2376 667 2383 856
rect 2416 827 2423 872
rect 2476 727 2483 973
rect 2516 916 2523 973
rect 2676 943 2683 993
rect 2656 936 2683 943
rect 2553 920 2567 933
rect 2556 916 2563 920
rect 2596 807 2603 933
rect 2656 928 2663 936
rect 2693 920 2707 933
rect 2696 916 2703 920
rect 2576 796 2593 803
rect 2433 700 2447 713
rect 2436 696 2443 700
rect 2576 707 2583 796
rect 2476 627 2483 692
rect 2276 403 2283 473
rect 2316 427 2323 573
rect 2256 396 2283 403
rect 2127 356 2143 363
rect 1916 187 1923 253
rect 2076 176 2083 253
rect 2116 176 2123 353
rect 2133 327 2147 332
rect 1616 107 1623 143
rect 1736 140 1743 143
rect 1733 127 1747 140
rect 1636 83 1643 113
rect 1896 107 1903 153
rect 1976 123 1983 132
rect 1956 116 1983 123
rect 2133 127 2147 132
rect 1956 107 1963 116
rect 1947 96 1963 107
rect 1947 93 1960 96
rect 2156 87 2163 394
rect 2316 366 2323 413
rect 2376 396 2383 473
rect 2476 427 2483 613
rect 2596 587 2603 713
rect 2616 708 2623 913
rect 2676 847 2683 883
rect 2413 400 2427 413
rect 2456 416 2473 423
rect 2416 396 2423 400
rect 2196 263 2203 363
rect 2356 327 2363 363
rect 2176 256 2203 263
rect 2176 227 2183 256
rect 2200 223 2213 227
rect 2196 213 2213 223
rect 2196 187 2203 213
rect 2213 180 2227 192
rect 2216 176 2223 180
rect 2256 176 2263 273
rect 2176 146 2183 173
rect 2336 146 2343 233
rect 2393 180 2407 193
rect 2396 176 2403 180
rect 2436 176 2443 213
rect 2456 183 2463 416
rect 2516 396 2523 513
rect 2496 207 2503 363
rect 2536 327 2543 363
rect 2596 307 2603 453
rect 2636 447 2643 833
rect 2656 767 2663 813
rect 2676 708 2683 733
rect 2736 687 2743 933
rect 2756 867 2763 1033
rect 2796 947 2803 1253
rect 2816 1007 2823 1273
rect 2856 1147 2863 1183
rect 2896 1180 2903 1183
rect 2893 1167 2907 1180
rect 2936 1143 2943 1373
rect 2956 1287 2963 1403
rect 3036 1327 3043 1393
rect 3116 1367 3123 1696
rect 2996 1216 3003 1253
rect 3053 1243 3067 1253
rect 3036 1240 3067 1243
rect 3036 1236 3063 1240
rect 3036 1216 3043 1236
rect 2956 1167 2963 1213
rect 3016 1180 3023 1183
rect 3013 1167 3027 1180
rect 3096 1186 3103 1313
rect 3116 1187 3123 1273
rect 3136 1247 3143 1513
rect 3216 1507 3223 1692
rect 3276 1687 3283 1736
rect 3456 1743 3463 1913
rect 3496 1807 3503 1973
rect 3516 1967 3523 2272
rect 3536 2267 3543 2793
rect 3556 2487 3563 2896
rect 3596 2823 3603 3093
rect 3576 2816 3603 2823
rect 3576 2776 3583 2816
rect 3616 2807 3623 3213
rect 3647 3193 3653 3207
rect 3636 2966 3643 3073
rect 3656 3008 3663 3073
rect 3676 3067 3683 3213
rect 3716 3163 3723 3476
rect 3736 3407 3743 3453
rect 3776 3403 3783 3503
rect 3796 3427 3803 3692
rect 3816 3527 3823 3673
rect 3896 3547 3903 3973
rect 4136 3923 4143 4213
rect 4176 4083 4183 4193
rect 4196 4107 4203 4173
rect 4176 4076 4203 4083
rect 4116 3916 4143 3923
rect 4036 3887 4043 3913
rect 3953 3820 3967 3833
rect 3956 3816 3963 3820
rect 4016 3807 4023 3833
rect 4036 3787 4043 3873
rect 4096 3816 4103 3853
rect 4116 3847 4123 3916
rect 4136 3827 4143 3893
rect 3976 3780 3983 3783
rect 3973 3767 3987 3780
rect 3936 3587 3943 3633
rect 3756 3396 3783 3403
rect 3756 3308 3763 3396
rect 3796 3307 3803 3353
rect 3776 3187 3783 3263
rect 3696 3156 3723 3163
rect 3696 3047 3703 3156
rect 3796 3027 3803 3253
rect 3816 3127 3823 3472
rect 3836 3387 3843 3533
rect 3916 3516 3943 3523
rect 3856 3467 3863 3513
rect 3856 3367 3863 3393
rect 3876 3367 3883 3413
rect 3916 3367 3923 3453
rect 3836 3267 3843 3352
rect 3936 3347 3943 3516
rect 3956 3407 3963 3713
rect 3996 3703 4003 3772
rect 3976 3696 4003 3703
rect 3976 3467 3983 3696
rect 4016 3587 4023 3753
rect 3856 3167 3863 3293
rect 3856 3127 3863 3153
rect 3596 2503 3603 2693
rect 3616 2567 3623 2743
rect 3636 2667 3643 2952
rect 3716 2827 3723 2933
rect 3736 2788 3743 2873
rect 3756 2803 3763 3013
rect 3796 2996 3803 3013
rect 3836 2996 3843 3053
rect 3856 3007 3863 3113
rect 3756 2796 3783 2803
rect 3656 2736 3703 2743
rect 3656 2607 3663 2736
rect 3756 2727 3763 2743
rect 3636 2507 3643 2533
rect 3676 2527 3683 2633
rect 3596 2496 3623 2503
rect 3616 2476 3623 2496
rect 3676 2446 3683 2513
rect 3696 2467 3703 2713
rect 3756 2587 3763 2713
rect 3776 2627 3783 2796
rect 3796 2523 3803 2893
rect 3856 2867 3863 2953
rect 3876 2943 3883 3231
rect 3896 2963 3903 3073
rect 3916 3067 3923 3233
rect 3936 3227 3943 3263
rect 3956 3247 3963 3353
rect 3976 3267 3983 3432
rect 3996 3387 4003 3553
rect 4016 3516 4023 3573
rect 4016 3343 4023 3453
rect 4056 3427 4063 3483
rect 3996 3336 4023 3343
rect 3996 3263 4003 3336
rect 4076 3296 4083 3733
rect 4116 3723 4123 3783
rect 4096 3716 4123 3723
rect 4096 3647 4103 3716
rect 4136 3687 4143 3773
rect 4156 3707 4163 3993
rect 4176 3907 4183 4023
rect 4196 3883 4203 4076
rect 4256 4048 4263 4273
rect 4236 4020 4243 4023
rect 4233 4007 4247 4020
rect 4176 3876 4203 3883
rect 4176 3827 4183 3876
rect 4216 3828 4223 3853
rect 4256 3783 4263 4034
rect 4276 4007 4283 4173
rect 4296 3967 4303 4273
rect 4336 4127 4343 4173
rect 4396 4067 4403 4303
rect 4336 3887 4343 4003
rect 4313 3820 4327 3833
rect 4316 3816 4323 3820
rect 4356 3816 4363 3913
rect 4096 3487 4103 3633
rect 4136 3523 4143 3593
rect 4176 3547 4183 3673
rect 4196 3627 4203 3783
rect 4236 3776 4263 3783
rect 4116 3516 4143 3523
rect 4196 3516 4203 3553
rect 4116 3447 4123 3516
rect 4176 3427 4183 3483
rect 3996 3256 4023 3263
rect 4016 3123 4023 3256
rect 4056 3187 4063 3263
rect 4096 3227 4103 3263
rect 4076 3216 4093 3223
rect 3996 3116 4023 3123
rect 4036 3176 4053 3183
rect 3927 3003 3940 3007
rect 3927 2996 3943 3003
rect 3927 2993 3940 2996
rect 3896 2956 3923 2963
rect 3876 2936 3903 2943
rect 3776 2516 3803 2523
rect 3747 2494 3753 2507
rect 3740 2493 3753 2494
rect 3776 2476 3783 2516
rect 3793 2487 3807 2493
rect 3556 2367 3563 2433
rect 3596 2323 3603 2443
rect 3576 2316 3603 2323
rect 3576 2287 3583 2316
rect 3596 2256 3603 2293
rect 3616 2287 3623 2353
rect 3636 2263 3643 2333
rect 3656 2327 3663 2393
rect 3676 2267 3683 2373
rect 3696 2327 3703 2453
rect 3756 2367 3763 2443
rect 3816 2387 3823 2813
rect 3896 2776 3903 2936
rect 3836 2707 3843 2773
rect 3836 2507 3843 2613
rect 3856 2607 3863 2743
rect 3916 2727 3923 2956
rect 3956 2927 3963 2952
rect 3976 2847 3983 2933
rect 3996 2907 4003 3116
rect 4016 2947 4023 3013
rect 4036 3007 4043 3176
rect 4076 3023 4083 3216
rect 4096 3047 4103 3153
rect 4116 3087 4123 3252
rect 4136 3127 4143 3293
rect 4156 3227 4163 3393
rect 4176 3307 4183 3413
rect 4216 3407 4223 3514
rect 4236 3327 4243 3776
rect 4336 3780 4343 3783
rect 4333 3767 4347 3780
rect 4293 3747 4307 3751
rect 4316 3567 4323 3713
rect 4396 3607 4403 4032
rect 4416 4003 4423 4273
rect 4456 4036 4463 4213
rect 4476 4087 4483 4393
rect 4536 4367 4543 4433
rect 4536 4300 4543 4303
rect 4496 4087 4503 4293
rect 4533 4287 4547 4300
rect 4616 4287 4623 4512
rect 4636 4487 4643 4533
rect 4656 4363 4663 4553
rect 4716 4520 4723 4523
rect 4713 4507 4727 4520
rect 4816 4507 4823 4773
rect 4836 4587 4843 4816
rect 4876 4787 4883 4823
rect 4876 4568 4883 4713
rect 4896 4607 4903 4753
rect 4916 4556 4923 4633
rect 4936 4587 4943 5033
rect 4956 5007 4963 5153
rect 4976 5107 4983 5313
rect 4996 5187 5003 5373
rect 5036 5307 5043 5343
rect 5076 5336 5103 5343
rect 5036 5107 5043 5293
rect 5096 5287 5103 5336
rect 4976 5076 5003 5083
rect 5056 5076 5063 5193
rect 4976 4983 4983 5076
rect 4956 4976 4983 4983
rect 4956 4727 4963 4976
rect 5076 4967 5083 5033
rect 5096 4987 5103 5273
rect 5116 5167 5123 5453
rect 5136 5287 5143 5573
rect 5196 5507 5203 5563
rect 5236 5527 5243 5563
rect 5236 5516 5253 5527
rect 5240 5513 5253 5516
rect 5236 5447 5243 5493
rect 5236 5376 5243 5433
rect 5276 5382 5283 5696
rect 5356 5596 5363 5713
rect 5396 5566 5403 5753
rect 5616 5747 5623 6072
rect 5653 6067 5667 6072
rect 5696 5987 5703 6083
rect 5756 6007 5763 6173
rect 5796 6116 5803 6153
rect 5896 6027 5903 6113
rect 5676 5896 5683 5933
rect 5696 5787 5703 5863
rect 5416 5563 5423 5653
rect 5456 5623 5463 5673
rect 5456 5616 5483 5623
rect 5476 5596 5483 5616
rect 5516 5596 5523 5653
rect 5556 5566 5563 5693
rect 5736 5633 5743 5853
rect 5756 5783 5763 5972
rect 5933 5907 5947 5913
rect 5956 5896 5963 5993
rect 5976 5947 5983 6083
rect 5996 5908 6003 5973
rect 6036 5907 6043 6073
rect 6056 5987 6063 6113
rect 6196 6086 6203 6153
rect 5776 5807 5783 5893
rect 5916 5866 5923 5893
rect 5796 5787 5803 5853
rect 5756 5776 5783 5783
rect 5696 5626 5743 5633
rect 5660 5603 5673 5607
rect 5656 5596 5673 5603
rect 5660 5593 5673 5596
rect 5416 5556 5463 5563
rect 5596 5527 5603 5563
rect 5256 5375 5283 5382
rect 5176 5340 5183 5343
rect 5173 5327 5187 5340
rect 5216 5287 5223 5343
rect 5156 5147 5163 5233
rect 5116 5007 5123 5093
rect 5176 5076 5183 5133
rect 5216 5076 5223 5113
rect 5256 5043 5263 5375
rect 5316 5203 5323 5433
rect 5376 5376 5383 5473
rect 5416 5388 5423 5513
rect 5436 5367 5443 5493
rect 5456 5347 5463 5473
rect 5516 5407 5523 5473
rect 5416 5340 5463 5347
rect 5396 5247 5403 5332
rect 5296 5196 5323 5203
rect 5276 5067 5283 5153
rect 5296 5087 5303 5196
rect 5316 5076 5323 5173
rect 5416 5147 5423 5340
rect 5436 5227 5443 5313
rect 5496 5287 5503 5343
rect 5456 5207 5463 5233
rect 5516 5187 5523 5273
rect 5536 5127 5543 5333
rect 5556 5143 5563 5493
rect 5636 5407 5643 5563
rect 5696 5527 5703 5626
rect 5776 5608 5783 5776
rect 5816 5605 5823 5733
rect 5836 5647 5843 5863
rect 5816 5598 5843 5605
rect 5816 5597 5823 5598
rect 5716 5566 5723 5593
rect 5676 5516 5693 5523
rect 5626 5393 5627 5400
rect 5613 5380 5627 5393
rect 5616 5376 5623 5380
rect 5656 5376 5663 5433
rect 5676 5387 5683 5516
rect 5716 5467 5723 5552
rect 5796 5507 5803 5563
rect 5596 5207 5603 5343
rect 5576 5196 5593 5203
rect 5576 5167 5583 5196
rect 5556 5136 5583 5143
rect 5496 5076 5503 5113
rect 5533 5088 5547 5092
rect 5256 5036 5283 5043
rect 5236 4947 5243 5033
rect 4996 4856 5003 4933
rect 5096 4907 5103 4933
rect 5227 4926 5240 4927
rect 5227 4913 5233 4926
rect 5096 4826 5103 4893
rect 5116 4867 5123 4913
rect 5153 4860 5167 4873
rect 5156 4856 5163 4860
rect 5236 4826 5243 4892
rect 5016 4820 5023 4823
rect 5013 4807 5027 4820
rect 5136 4727 5143 4823
rect 4836 4527 4843 4552
rect 4836 4447 4843 4513
rect 4656 4356 4683 4363
rect 4676 4348 4683 4356
rect 4696 4300 4703 4303
rect 4693 4287 4707 4300
rect 4536 4006 4543 4073
rect 4416 3996 4433 4003
rect 4416 3727 4423 3972
rect 4436 3827 4443 3992
rect 4473 3820 4487 3833
rect 4516 3828 4523 3953
rect 4476 3816 4483 3820
rect 4556 3807 4563 4253
rect 4456 3727 4463 3783
rect 4496 3780 4503 3783
rect 4493 3767 4507 3780
rect 4316 3516 4323 3553
rect 4193 3300 4207 3313
rect 4196 3296 4203 3300
rect 4236 3296 4283 3303
rect 4336 3296 4343 3373
rect 4356 3367 4363 3533
rect 4376 3407 4383 3553
rect 4476 3516 4483 3753
rect 4496 3527 4503 3732
rect 4396 3407 4403 3473
rect 4416 3467 4423 3483
rect 4216 3107 4223 3263
rect 4276 3067 4283 3296
rect 4396 3266 4403 3293
rect 4356 3243 4363 3263
rect 4336 3236 4363 3243
rect 4336 3147 4343 3236
rect 4416 3204 4423 3453
rect 4456 3367 4463 3483
rect 4493 3467 4507 3473
rect 4516 3427 4523 3653
rect 4536 3527 4543 3753
rect 4576 3567 4583 4073
rect 4596 4036 4603 4233
rect 4636 4167 4643 4213
rect 4656 4187 4663 4253
rect 4636 3847 4643 3992
rect 4593 3820 4607 3833
rect 4596 3816 4603 3820
rect 4636 3687 4643 3783
rect 4573 3520 4587 3532
rect 4613 3520 4627 3533
rect 4636 3527 4643 3613
rect 4576 3516 4583 3520
rect 4616 3516 4623 3520
rect 4436 3307 4443 3333
rect 4367 3197 4423 3204
rect 4056 3016 4083 3023
rect 4056 2996 4063 3016
rect 4256 2996 4263 3033
rect 4076 2960 4083 2963
rect 3936 2687 3943 2833
rect 3876 2587 3883 2673
rect 3836 2480 3863 2483
rect 3833 2476 3863 2480
rect 3916 2476 3923 2533
rect 3833 2467 3847 2476
rect 3716 2303 3723 2353
rect 3696 2300 3723 2303
rect 3693 2296 3723 2300
rect 3693 2287 3707 2296
rect 3756 2268 3763 2313
rect 3636 2256 3663 2263
rect 3536 2087 3543 2113
rect 3536 1956 3543 2073
rect 3556 2007 3563 2193
rect 3576 1968 3583 2153
rect 3616 1927 3623 2223
rect 3636 1967 3643 2213
rect 3656 2107 3663 2256
rect 3676 1987 3683 2153
rect 3696 2127 3703 2212
rect 3736 2167 3743 2223
rect 3776 2203 3783 2223
rect 3756 2196 3783 2203
rect 3756 2167 3763 2196
rect 3796 2183 3803 2213
rect 3776 2176 3803 2183
rect 3756 2107 3763 2153
rect 3676 1956 3683 1973
rect 3716 1956 3723 2053
rect 3776 2047 3783 2176
rect 3736 1987 3743 2033
rect 3816 2027 3823 2373
rect 3836 2087 3843 2293
rect 3896 2287 3903 2443
rect 3936 2387 3943 2473
rect 3936 2307 3943 2373
rect 3893 2260 3907 2273
rect 3896 2256 3903 2260
rect 3936 2256 3943 2293
rect 3956 2287 3963 2793
rect 4016 2776 4023 2833
rect 4036 2807 4043 2953
rect 4073 2947 4087 2960
rect 3976 2740 3983 2743
rect 3973 2727 3987 2740
rect 4056 2727 4063 2933
rect 3976 2447 3983 2633
rect 3996 2487 4003 2653
rect 4016 2567 4023 2713
rect 4056 2643 4063 2713
rect 4076 2667 4083 2933
rect 4116 2867 4123 2963
rect 4153 2947 4167 2953
rect 4176 2927 4183 2973
rect 4316 2967 4323 2994
rect 4207 2943 4220 2947
rect 4207 2933 4223 2943
rect 4196 2887 4203 2912
rect 4156 2823 4163 2873
rect 4216 2843 4223 2933
rect 4236 2867 4243 2963
rect 4276 2887 4283 2963
rect 4336 2907 4343 3053
rect 4356 3007 4363 3193
rect 4396 2996 4403 3153
rect 4436 3028 4443 3253
rect 4496 3243 4503 3263
rect 4536 3247 4543 3473
rect 4556 3427 4563 3483
rect 4573 3300 4587 3313
rect 4576 3296 4583 3300
rect 4616 3296 4623 3393
rect 4636 3387 4643 3473
rect 4656 3407 4663 4073
rect 4676 4007 4683 4133
rect 4736 4048 4743 4213
rect 4756 4087 4763 4353
rect 4856 4336 4863 4493
rect 4896 4343 4903 4523
rect 4936 4487 4943 4523
rect 4936 4347 4943 4433
rect 4896 4336 4923 4343
rect 4776 4147 4783 4333
rect 4876 4227 4883 4303
rect 4916 4306 4923 4336
rect 4956 4343 4963 4512
rect 4976 4367 4983 4573
rect 4996 4447 5003 4613
rect 5096 4467 5103 4673
rect 4956 4336 4983 4343
rect 5016 4336 5023 4373
rect 5116 4347 5123 4633
rect 5156 4568 5163 4773
rect 5236 4568 5243 4812
rect 5256 4527 5263 4973
rect 5276 4967 5283 5036
rect 5376 5040 5383 5043
rect 5373 5027 5387 5040
rect 5287 4913 5293 4927
rect 5356 4923 5363 5013
rect 5336 4920 5363 4923
rect 5333 4916 5363 4920
rect 5316 4856 5323 4913
rect 5333 4907 5347 4916
rect 5346 4900 5347 4907
rect 5356 4868 5363 4893
rect 5376 4867 5383 4953
rect 5416 4907 5423 5033
rect 5436 5027 5443 5073
rect 5476 5040 5483 5043
rect 5473 5027 5487 5040
rect 5176 4520 5183 4523
rect 5173 4507 5187 4520
rect 5176 4348 5183 4453
rect 4896 4267 4903 4293
rect 4776 4036 4783 4093
rect 4676 3643 4683 3793
rect 4696 3663 4703 4033
rect 4796 4000 4803 4003
rect 4793 3987 4807 4000
rect 4836 4006 4843 4133
rect 4936 4067 4943 4312
rect 5076 4306 5083 4333
rect 5036 4300 5043 4303
rect 5033 4287 5047 4300
rect 5096 4147 5103 4334
rect 4853 4048 4867 4053
rect 4936 4033 4953 4047
rect 4696 3656 4723 3663
rect 4676 3636 4703 3643
rect 4676 3587 4683 3613
rect 4696 3607 4703 3636
rect 4676 3447 4683 3573
rect 4696 3527 4703 3553
rect 4716 3516 4723 3656
rect 4756 3528 4763 3772
rect 4776 3547 4783 3673
rect 4796 3583 4803 3853
rect 4816 3787 4823 3993
rect 4876 4000 4883 4003
rect 4836 3828 4843 3992
rect 4873 3987 4887 4000
rect 4916 3967 4923 4003
rect 4976 3987 4983 4053
rect 5056 4036 5063 4093
rect 5093 4047 5107 4053
rect 4956 3976 4973 3983
rect 4847 3816 4863 3823
rect 4896 3816 4903 3853
rect 4933 3847 4947 3853
rect 4836 3667 4843 3713
rect 4796 3576 4823 3583
rect 4796 3527 4803 3553
rect 4816 3507 4823 3576
rect 4696 3427 4703 3473
rect 4656 3303 4663 3353
rect 4696 3308 4703 3353
rect 4736 3308 4743 3433
rect 4776 3427 4783 3483
rect 4807 3486 4820 3487
rect 4807 3473 4813 3486
rect 4796 3323 4803 3452
rect 4776 3316 4803 3323
rect 4656 3296 4683 3303
rect 4476 3236 4503 3243
rect 4456 3107 4463 3173
rect 4456 3047 4463 3072
rect 4476 3043 4483 3236
rect 4536 3127 4543 3153
rect 4467 3036 4483 3043
rect 4367 2963 4380 2967
rect 4367 2956 4383 2963
rect 4367 2953 4380 2956
rect 4356 2927 4363 2953
rect 4296 2863 4303 2893
rect 4276 2856 4303 2863
rect 4216 2836 4243 2843
rect 4136 2816 4163 2823
rect 4096 2787 4103 2813
rect 4136 2787 4143 2816
rect 4127 2776 4143 2787
rect 4127 2773 4140 2776
rect 4216 2787 4223 2813
rect 4156 2740 4163 2743
rect 4116 2703 4123 2733
rect 4153 2727 4167 2740
rect 4116 2696 4143 2703
rect 4036 2636 4063 2643
rect 4036 2488 4043 2636
rect 4056 2527 4063 2613
rect 4076 2476 4083 2533
rect 4136 2527 4143 2696
rect 4156 2507 4163 2653
rect 4176 2603 4183 2673
rect 4176 2596 4203 2603
rect 4176 2476 4183 2573
rect 4196 2507 4203 2596
rect 4216 2527 4223 2693
rect 4196 2496 4213 2507
rect 4200 2493 4213 2496
rect 4236 2483 4243 2836
rect 4256 2787 4263 2813
rect 4276 2807 4283 2856
rect 4396 2847 4403 2893
rect 4333 2827 4347 2833
rect 4333 2787 4347 2792
rect 4356 2746 4363 2833
rect 4387 2773 4393 2787
rect 4436 2776 4443 2933
rect 4456 2907 4463 2953
rect 4476 2947 4483 3012
rect 4496 2927 4503 2993
rect 4496 2847 4503 2913
rect 4473 2780 4487 2793
rect 4516 2787 4523 3033
rect 4536 2996 4543 3033
rect 4556 3027 4563 3213
rect 4596 3147 4603 3263
rect 4676 3227 4683 3296
rect 4616 2987 4623 3053
rect 4636 3047 4643 3133
rect 4556 2867 4563 2933
rect 4576 2847 4583 2963
rect 4613 2947 4627 2952
rect 4636 2907 4643 3012
rect 4656 3007 4663 3033
rect 4696 3008 4703 3233
rect 4716 3047 4723 3263
rect 4756 3187 4763 3253
rect 4776 3147 4783 3316
rect 4816 3296 4823 3353
rect 4836 3327 4843 3653
rect 4856 3587 4863 3693
rect 4893 3520 4907 3533
rect 4956 3528 4963 3976
rect 4976 3827 4983 3933
rect 4996 3847 5003 4033
rect 5076 3907 5083 4003
rect 5096 3967 5103 3993
rect 5047 3843 5060 3847
rect 5047 3833 5063 3843
rect 5013 3820 5027 3833
rect 5016 3816 5023 3820
rect 5056 3816 5063 3833
rect 4987 3783 5000 3787
rect 4987 3773 5003 3783
rect 4996 3687 5003 3773
rect 5096 3767 5103 3953
rect 4896 3516 4903 3520
rect 4967 3516 4983 3523
rect 4876 3387 4883 3483
rect 4916 3480 4923 3483
rect 4913 3467 4927 3480
rect 4976 3467 4983 3516
rect 4856 3296 4863 3353
rect 4896 3307 4903 3453
rect 4916 3266 4923 3313
rect 4936 3307 4943 3373
rect 4976 3308 4983 3393
rect 5016 3327 5023 3593
rect 5036 3507 5043 3751
rect 5116 3607 5123 4293
rect 5156 4187 5163 4303
rect 5216 4227 5223 4523
rect 5276 4487 5283 4813
rect 5296 4787 5303 4823
rect 5316 4627 5323 4693
rect 5336 4647 5343 4812
rect 5316 4556 5323 4613
rect 5356 4556 5363 4753
rect 5376 4707 5383 4813
rect 5336 4447 5343 4523
rect 5396 4507 5403 4873
rect 5476 4856 5483 4893
rect 5516 4867 5523 4893
rect 5536 4826 5543 4953
rect 5576 4903 5583 5136
rect 5616 5127 5623 5293
rect 5676 5287 5683 5333
rect 5696 5327 5703 5413
rect 5716 5343 5723 5373
rect 5836 5347 5843 5598
rect 5856 5387 5863 5793
rect 5876 5767 5883 5863
rect 5916 5707 5923 5852
rect 5936 5827 5943 5853
rect 5976 5647 5983 5863
rect 5913 5600 5927 5613
rect 5916 5596 5923 5600
rect 5956 5596 5963 5633
rect 5896 5527 5903 5563
rect 5716 5336 5743 5343
rect 5627 5093 5633 5107
rect 5656 5076 5663 5113
rect 5716 5043 5723 5313
rect 5736 5207 5743 5336
rect 5776 5267 5783 5332
rect 5816 5247 5823 5343
rect 5876 5327 5883 5473
rect 5973 5380 5987 5393
rect 5996 5387 6003 5552
rect 5976 5376 5983 5380
rect 5916 5247 5923 5343
rect 5956 5287 5963 5343
rect 6016 5346 6023 5831
rect 6056 5807 6063 5913
rect 6153 5900 6167 5913
rect 6156 5896 6163 5900
rect 6096 5827 6103 5863
rect 6136 5860 6143 5863
rect 6133 5847 6147 5860
rect 6036 5596 6043 5633
rect 6096 5603 6103 5653
rect 6096 5596 6123 5603
rect 6076 5407 6083 5563
rect 6116 5407 6123 5596
rect 6136 5487 6143 5793
rect 6196 5767 6203 6072
rect 6196 5527 6203 5753
rect 6216 5627 6223 6013
rect 5836 5076 5843 5173
rect 5996 5167 6003 5333
rect 6036 5307 6043 5393
rect 6073 5380 6087 5393
rect 6113 5380 6127 5393
rect 6076 5376 6083 5380
rect 6116 5376 6123 5380
rect 5936 5076 5943 5153
rect 5613 4983 5627 4993
rect 5676 4987 5683 5043
rect 5696 5036 5723 5043
rect 5613 4980 5643 4983
rect 5616 4976 5643 4980
rect 5556 4896 5583 4903
rect 5456 4820 5463 4823
rect 5453 4807 5467 4820
rect 5556 4807 5563 4896
rect 5616 4856 5623 4953
rect 5636 4947 5643 4976
rect 5673 4887 5687 4893
rect 5653 4860 5667 4873
rect 5656 4856 5663 4860
rect 5587 4823 5600 4827
rect 5587 4816 5603 4823
rect 5636 4820 5643 4823
rect 5587 4813 5600 4816
rect 5633 4807 5647 4820
rect 5696 4807 5703 5036
rect 5716 4907 5723 4933
rect 5736 4887 5743 5074
rect 5756 4927 5763 4993
rect 5713 4863 5727 4872
rect 5713 4860 5743 4863
rect 5716 4856 5743 4860
rect 5816 4867 5823 5032
rect 5800 4824 5813 4827
rect 5756 4820 5763 4823
rect 5436 4567 5443 4653
rect 5533 4567 5547 4573
rect 5576 4563 5583 4613
rect 5596 4588 5603 4793
rect 5556 4556 5583 4563
rect 5376 4496 5393 4503
rect 5133 4047 5147 4053
rect 5153 4040 5167 4053
rect 5193 4040 5207 4053
rect 5216 4047 5223 4133
rect 5156 4036 5163 4040
rect 5196 4036 5203 4040
rect 5136 3827 5143 3993
rect 5176 3907 5183 4003
rect 5216 3843 5223 3993
rect 5196 3836 5223 3843
rect 5196 3828 5203 3836
rect 5236 3827 5243 4373
rect 5276 4247 5283 4303
rect 5316 4267 5323 4303
rect 5356 4247 5363 4493
rect 5376 4287 5383 4496
rect 5416 4487 5423 4553
rect 5416 4368 5423 4473
rect 5476 4387 5483 4523
rect 5536 4423 5543 4453
rect 5556 4447 5563 4556
rect 5633 4560 5647 4573
rect 5636 4556 5643 4560
rect 5536 4416 5563 4423
rect 5453 4340 5467 4353
rect 5556 4363 5563 4416
rect 5576 4363 5583 4413
rect 5596 4387 5603 4493
rect 5616 4487 5623 4523
rect 5656 4487 5663 4523
rect 5676 4367 5683 4513
rect 5696 4467 5703 4772
rect 5716 4563 5723 4813
rect 5753 4807 5767 4820
rect 5796 4813 5813 4824
rect 5756 4583 5763 4693
rect 5776 4647 5783 4793
rect 5796 4767 5803 4813
rect 5836 4803 5843 4993
rect 5856 4927 5863 4993
rect 5876 4903 5883 4933
rect 5856 4896 5883 4903
rect 5856 4867 5863 4896
rect 5896 4856 5903 4953
rect 5916 4887 5923 5043
rect 5936 4887 5943 4993
rect 5956 4967 5963 5043
rect 5936 4856 5943 4873
rect 5876 4820 5883 4823
rect 5827 4796 5843 4803
rect 5816 4747 5823 4792
rect 5800 4683 5813 4687
rect 5796 4673 5813 4683
rect 5796 4587 5803 4673
rect 5856 4627 5863 4813
rect 5873 4807 5887 4820
rect 5887 4800 5903 4803
rect 5887 4796 5907 4800
rect 5893 4787 5907 4796
rect 5876 4727 5883 4772
rect 5916 4663 5923 4812
rect 5896 4656 5923 4663
rect 5756 4576 5783 4583
rect 5716 4556 5743 4563
rect 5776 4556 5783 4576
rect 5836 4567 5843 4593
rect 5896 4587 5903 4656
rect 5796 4487 5803 4513
rect 5816 4467 5823 4554
rect 5916 4556 5923 4593
rect 5936 4567 5943 4733
rect 5556 4356 5583 4363
rect 5456 4336 5463 4340
rect 5556 4336 5563 4356
rect 5633 4347 5647 4353
rect 5436 4283 5443 4303
rect 5416 4276 5443 4283
rect 5316 4047 5323 4232
rect 5336 4027 5343 4213
rect 5296 4000 5303 4003
rect 5293 3987 5307 4000
rect 5336 3967 5343 3992
rect 5356 3867 5363 4053
rect 5376 4047 5383 4252
rect 5396 4036 5403 4233
rect 5416 4207 5423 4276
rect 5436 4036 5443 4213
rect 5456 4107 5463 4273
rect 5516 4227 5523 4313
rect 5616 4227 5623 4334
rect 5696 4336 5703 4432
rect 5756 4347 5763 4453
rect 5856 4387 5863 4523
rect 5787 4343 5800 4347
rect 5787 4336 5803 4343
rect 5787 4333 5800 4336
rect 5876 4347 5883 4493
rect 5896 4427 5903 4523
rect 5616 4067 5623 4093
rect 5616 4036 5623 4053
rect 5636 4043 5643 4293
rect 5676 4207 5683 4303
rect 5716 4300 5723 4303
rect 5713 4287 5727 4300
rect 5756 4306 5763 4333
rect 5676 4107 5683 4193
rect 5736 4103 5743 4293
rect 5776 4247 5783 4273
rect 5816 4107 5823 4303
rect 5856 4227 5863 4303
rect 5736 4096 5763 4103
rect 5636 4036 5663 4043
rect 5256 3786 5263 3833
rect 5136 3707 5143 3773
rect 5176 3687 5183 3783
rect 5053 3520 5067 3533
rect 5113 3520 5127 3533
rect 5056 3516 5063 3520
rect 5116 3516 5123 3520
rect 5036 3467 5043 3493
rect 5156 3480 5163 3483
rect 5076 3407 5083 3453
rect 5136 3447 5143 3472
rect 5153 3467 5167 3480
rect 5020 3303 5033 3307
rect 5016 3296 5033 3303
rect 5020 3293 5033 3296
rect 4836 3227 4843 3263
rect 4816 2996 4823 3053
rect 4853 3000 4867 3013
rect 4896 3007 4903 3226
rect 4856 2996 4863 3000
rect 4476 2776 4483 2780
rect 4256 2587 4263 2733
rect 4316 2627 4323 2673
rect 4236 2476 4263 2483
rect 4296 2476 4303 2533
rect 3976 2287 3983 2412
rect 4036 2387 4043 2413
rect 4056 2367 4063 2443
rect 3856 2216 3873 2223
rect 3767 2026 3780 2027
rect 3767 2013 3773 2026
rect 3796 1967 3803 1993
rect 3813 1960 3827 1973
rect 3816 1956 3823 1960
rect 3856 1956 3863 2216
rect 3896 2127 3903 2173
rect 3916 2107 3923 2223
rect 3956 2187 3963 2223
rect 3876 1967 3883 2053
rect 3936 1963 3943 2113
rect 3916 1956 3943 1963
rect 3956 1956 3963 2173
rect 3976 1987 3983 2153
rect 3996 1988 4003 2293
rect 4016 2047 4023 2273
rect 4076 2256 4083 2333
rect 4096 2287 4103 2353
rect 4116 2307 4123 2473
rect 4147 2443 4160 2447
rect 4147 2436 4163 2443
rect 4147 2433 4160 2436
rect 4036 2216 4063 2223
rect 4036 2167 4043 2216
rect 4096 2187 4103 2223
rect 4096 2107 4103 2152
rect 4116 2127 4123 2213
rect 4136 2127 4143 2293
rect 4156 2267 4163 2353
rect 4196 2256 4203 2443
rect 4236 2256 4243 2293
rect 4256 2267 4263 2476
rect 4376 2443 4383 2752
rect 4416 2607 4423 2743
rect 4456 2707 4463 2743
rect 4496 2740 4503 2743
rect 4493 2727 4507 2740
rect 4536 2727 4543 2833
rect 4553 2787 4567 2793
rect 4596 2776 4603 2813
rect 4636 2787 4643 2853
rect 4656 2807 4663 2953
rect 4676 2783 4683 2952
rect 4716 2907 4723 2963
rect 4776 2927 4783 2994
rect 4916 2967 4923 3073
rect 4936 3063 4943 3253
rect 4956 3187 4963 3263
rect 4936 3056 4963 3063
rect 4776 2847 4783 2892
rect 4796 2867 4803 2953
rect 4656 2776 4683 2783
rect 4693 2780 4707 2793
rect 4696 2776 4703 2780
rect 4416 2488 4423 2572
rect 4456 2488 4463 2593
rect 4476 2487 4483 2713
rect 4576 2707 4583 2732
rect 4613 2727 4627 2732
rect 4607 2713 4627 2727
rect 4500 2703 4513 2707
rect 4496 2693 4513 2703
rect 4496 2527 4503 2693
rect 4276 2367 4283 2433
rect 4316 2327 4323 2443
rect 4356 2436 4383 2443
rect 4156 2216 4183 2223
rect 4216 2220 4223 2223
rect 4027 2036 4043 2043
rect 3556 1767 3563 1912
rect 3436 1736 3463 1743
rect 3493 1740 3507 1753
rect 3496 1736 3503 1740
rect 3336 1700 3343 1703
rect 3153 1448 3167 1453
rect 3196 1436 3203 1473
rect 3276 1406 3283 1493
rect 3156 1267 3163 1393
rect 3216 1383 3223 1403
rect 3196 1376 3223 1383
rect 3196 1287 3203 1376
rect 3173 1220 3187 1233
rect 3176 1216 3183 1220
rect 2927 1136 2943 1143
rect 2853 920 2867 933
rect 2856 916 2863 920
rect 2916 923 2923 1133
rect 2947 943 2960 947
rect 2947 933 2963 943
rect 2916 916 2943 923
rect 2956 916 2963 933
rect 3016 916 3043 923
rect 2736 663 2743 673
rect 2656 487 2663 663
rect 2716 656 2743 663
rect 2756 647 2763 853
rect 2796 787 2803 883
rect 2896 847 2903 914
rect 2916 827 2923 893
rect 2856 696 2863 733
rect 2796 627 2803 663
rect 2676 396 2683 513
rect 2616 327 2623 394
rect 2633 307 2647 313
rect 2576 227 2583 293
rect 2656 267 2663 363
rect 2696 343 2703 352
rect 2696 336 2713 343
rect 2676 247 2683 313
rect 2487 196 2503 207
rect 2487 193 2500 196
rect 2456 176 2483 183
rect 2476 146 2483 176
rect 2593 180 2607 193
rect 2596 176 2603 180
rect 2676 176 2683 212
rect 2716 176 2723 333
rect 2736 227 2743 353
rect 2756 207 2763 433
rect 2776 407 2783 553
rect 2836 447 2843 663
rect 2856 423 2863 453
rect 2836 416 2863 423
rect 2836 396 2843 416
rect 2776 327 2783 353
rect 2816 327 2823 363
rect 2856 207 2863 363
rect 2767 196 2783 203
rect 2276 136 2333 143
rect 2496 107 2503 173
rect 2576 140 2583 143
rect 2573 127 2587 140
rect 2776 143 2783 196
rect 2876 183 2883 353
rect 2896 347 2903 433
rect 2916 408 2923 773
rect 2936 767 2943 916
rect 2996 880 3003 883
rect 2993 867 3007 880
rect 3036 847 3043 916
rect 3076 907 3083 1173
rect 3216 1183 3223 1353
rect 3256 1307 3263 1333
rect 3276 1247 3283 1392
rect 3296 1327 3303 1693
rect 3333 1687 3347 1700
rect 3416 1667 3423 1734
rect 3316 1447 3323 1613
rect 3356 1436 3363 1473
rect 3436 1447 3443 1736
rect 3476 1436 3483 1553
rect 3376 1367 3383 1403
rect 3316 1307 3323 1333
rect 3256 1236 3273 1243
rect 3136 1167 3143 1183
rect 3196 1176 3223 1183
rect 3120 1166 3143 1167
rect 3127 1156 3143 1166
rect 3127 1153 3140 1156
rect 3216 1147 3223 1176
rect 3176 916 3183 1093
rect 3236 1087 3243 1213
rect 3256 1186 3263 1236
rect 3316 1216 3323 1253
rect 3336 1147 3343 1183
rect 3376 1047 3383 1332
rect 3396 1007 3403 1393
rect 3456 1347 3463 1392
rect 3496 1367 3503 1403
rect 3436 1216 3443 1273
rect 3416 1087 3423 1183
rect 3156 880 3163 883
rect 3153 867 3167 880
rect 3016 836 3033 843
rect 3016 807 3023 836
rect 2993 700 3007 713
rect 2996 696 3003 700
rect 3056 666 3063 793
rect 3216 727 3223 993
rect 3233 923 3247 933
rect 3233 920 3263 923
rect 3236 916 3263 920
rect 3496 916 3503 1193
rect 3516 923 3523 1373
rect 3536 1167 3543 1753
rect 3616 1736 3623 1793
rect 3596 1667 3603 1703
rect 3656 1527 3663 1833
rect 3696 1767 3703 1923
rect 3736 1867 3743 1923
rect 3720 1783 3733 1787
rect 3716 1773 3733 1783
rect 3716 1748 3723 1773
rect 3756 1748 3763 1873
rect 3776 1847 3783 1953
rect 3836 1867 3843 1923
rect 3876 1867 3883 1893
rect 3676 1467 3683 1733
rect 3736 1587 3743 1703
rect 3796 1663 3803 1793
rect 3836 1736 3843 1773
rect 3896 1767 3903 1953
rect 3916 1807 3923 1956
rect 3976 1920 3983 1923
rect 3933 1907 3947 1913
rect 3973 1907 3987 1920
rect 4016 1867 4023 1913
rect 4036 1887 4043 2036
rect 4116 1983 4123 2113
rect 4156 2027 4163 2216
rect 4213 2207 4227 2220
rect 4196 2107 4203 2173
rect 4096 1976 4123 1983
rect 3913 1747 3927 1753
rect 3776 1656 3803 1663
rect 3756 1567 3763 1593
rect 3567 1443 3580 1447
rect 3567 1436 3583 1443
rect 3567 1433 3580 1436
rect 3756 1436 3763 1553
rect 3776 1448 3783 1656
rect 3936 1607 3943 1753
rect 3996 1736 4003 1793
rect 3956 1627 3963 1693
rect 4013 1687 4027 1693
rect 4036 1647 4043 1773
rect 4056 1747 4063 1973
rect 4096 1956 4103 1976
rect 4133 1960 4147 1973
rect 4156 1967 4163 2013
rect 4136 1956 4143 1960
rect 4176 1867 4183 1973
rect 4076 1807 4083 1853
rect 4096 1736 4103 1773
rect 4156 1727 4163 1833
rect 4176 1747 4183 1853
rect 4196 1767 4203 2072
rect 4256 1983 4263 2213
rect 4276 2087 4283 2273
rect 4316 2256 4323 2292
rect 4336 2287 4343 2353
rect 4356 2267 4363 2436
rect 4436 2367 4443 2443
rect 4496 2446 4503 2513
rect 4473 2427 4487 2433
rect 4356 2187 4363 2213
rect 4247 1976 4263 1983
rect 4236 1956 4243 1973
rect 4276 1956 4283 2033
rect 4316 1967 4323 2173
rect 4376 2167 4383 2293
rect 4396 2207 4403 2313
rect 4496 2256 4503 2313
rect 4516 2267 4523 2633
rect 4596 2547 4603 2713
rect 4616 2607 4623 2693
rect 4656 2667 4663 2776
rect 4796 2746 4803 2813
rect 4756 2687 4763 2732
rect 4816 2727 4823 2933
rect 4836 2907 4843 2963
rect 4876 2927 4883 2952
rect 4916 2787 4923 2932
rect 4776 2647 4783 2713
rect 4796 2607 4803 2653
rect 4836 2647 4843 2733
rect 4833 2587 4847 2593
rect 4787 2586 4800 2587
rect 4787 2573 4793 2586
rect 4593 2480 4607 2493
rect 4596 2476 4603 2480
rect 4636 2476 4643 2533
rect 4656 2487 4663 2573
rect 4536 2226 4543 2433
rect 4676 2427 4683 2493
rect 4716 2476 4723 2533
rect 4756 2476 4763 2553
rect 4696 2407 4703 2433
rect 4816 2443 4823 2573
rect 4856 2567 4863 2743
rect 4896 2740 4903 2743
rect 4893 2727 4907 2740
rect 4936 2727 4943 3033
rect 4956 2847 4963 3056
rect 4976 3008 4983 3133
rect 4996 3047 5003 3263
rect 5033 3247 5047 3253
rect 5056 3127 5063 3313
rect 5076 3307 5083 3333
rect 5196 3303 5203 3693
rect 5216 3327 5223 3772
rect 5236 3587 5243 3653
rect 5236 3527 5243 3573
rect 5276 3547 5283 3853
rect 5293 3827 5307 3833
rect 5313 3820 5327 3833
rect 5316 3816 5323 3820
rect 5336 3527 5343 3772
rect 5376 3687 5383 3783
rect 5393 3767 5407 3773
rect 5416 3548 5423 4003
rect 5516 4003 5523 4034
rect 5516 3996 5543 4003
rect 5436 3727 5443 3953
rect 5456 3827 5463 3992
rect 5496 3816 5503 3993
rect 5536 3827 5543 3996
rect 5556 3947 5563 4003
rect 5596 4000 5603 4003
rect 5593 3987 5607 4000
rect 5636 3816 5643 3993
rect 5656 3867 5663 4036
rect 5736 4036 5743 4073
rect 5756 4067 5763 4096
rect 5773 4040 5787 4053
rect 5776 4036 5783 4040
rect 5716 3967 5723 4003
rect 5756 4000 5763 4003
rect 5753 3987 5767 4000
rect 5456 3667 5463 3773
rect 5476 3767 5483 3783
rect 5356 3483 5363 3533
rect 5476 3527 5483 3753
rect 5516 3687 5523 3783
rect 5460 3523 5473 3527
rect 5456 3516 5473 3523
rect 5460 3513 5473 3516
rect 5316 3476 5363 3483
rect 5187 3296 5203 3303
rect 5076 3127 5083 3253
rect 5107 3243 5120 3247
rect 5107 3233 5123 3243
rect 5007 3036 5023 3043
rect 5016 3023 5023 3036
rect 5016 3016 5043 3023
rect 5036 2996 5043 3016
rect 5056 2966 5063 3013
rect 5076 2887 5083 3033
rect 4976 2776 4983 2813
rect 5016 2776 5023 2813
rect 5036 2787 5043 2813
rect 4776 2436 4823 2443
rect 4436 2187 4443 2223
rect 4476 2220 4483 2223
rect 4473 2207 4487 2220
rect 4216 1736 4223 1793
rect 4256 1748 4263 1923
rect 4296 1887 4303 1912
rect 4076 1700 4083 1703
rect 4073 1687 4087 1700
rect 3556 1287 3563 1393
rect 3636 1367 3643 1403
rect 3676 1347 3683 1432
rect 3736 1400 3743 1403
rect 3733 1387 3747 1400
rect 3676 1307 3683 1333
rect 3776 1307 3783 1333
rect 3693 1283 3707 1293
rect 3796 1287 3803 1513
rect 3816 1347 3823 1473
rect 3856 1436 3863 1473
rect 3876 1367 3883 1403
rect 3676 1280 3707 1283
rect 3676 1276 3703 1280
rect 3576 1180 3583 1183
rect 3573 1167 3587 1180
rect 3616 1087 3623 1183
rect 3656 1107 3663 1273
rect 3676 1186 3683 1276
rect 3516 916 3543 923
rect 3153 700 3167 713
rect 3156 696 3163 700
rect 2976 660 2983 663
rect 2973 647 2987 660
rect 3076 567 3083 693
rect 3136 660 3143 663
rect 3133 647 3147 660
rect 3216 607 3223 713
rect 3236 707 3243 793
rect 3256 727 3263 753
rect 3276 696 3283 833
rect 3316 703 3323 843
rect 3396 708 3403 914
rect 3536 886 3543 916
rect 3476 863 3483 883
rect 3456 856 3483 863
rect 3316 696 3343 703
rect 3296 607 3303 663
rect 2936 396 2943 513
rect 3336 467 3343 696
rect 3436 696 3443 813
rect 3456 707 3463 856
rect 2973 408 2987 413
rect 3093 400 3107 413
rect 3136 408 3143 453
rect 3096 396 3103 400
rect 2856 176 2883 183
rect 2616 87 2623 133
rect 2696 107 2703 143
rect 2736 136 2783 143
rect 2836 107 2843 143
rect 2876 87 2883 133
rect 2896 127 2903 193
rect 2956 176 2963 363
rect 2996 360 3003 363
rect 3076 360 3083 363
rect 2993 347 3007 360
rect 3073 347 3087 360
rect 3176 327 3183 394
rect 3196 367 3203 413
rect 3253 400 3267 413
rect 3256 396 3263 400
rect 3036 146 3043 233
rect 3076 176 3083 293
rect 3116 227 3123 273
rect 3236 227 3243 363
rect 3276 267 3283 363
rect 3336 247 3343 413
rect 3356 287 3363 694
rect 3393 400 3407 413
rect 3456 408 3463 653
rect 3476 627 3483 833
rect 3556 696 3563 1033
rect 3696 928 3703 1253
rect 3836 1147 3843 1273
rect 3936 1247 3943 1453
rect 3956 1347 3963 1473
rect 4036 1467 4043 1493
rect 4007 1463 4020 1467
rect 4007 1453 4023 1463
rect 4016 1436 4023 1453
rect 3976 1307 3983 1373
rect 4076 1247 4083 1593
rect 4096 1406 4103 1673
rect 4116 1587 4123 1703
rect 4136 1436 4143 1553
rect 4176 1436 4183 1693
rect 4196 1587 4203 1703
rect 4276 1527 4283 1813
rect 4336 1787 4343 2033
rect 4356 1967 4363 2013
rect 4396 1956 4403 2172
rect 4396 1747 4403 1873
rect 4436 1827 4443 1973
rect 4476 1956 4483 2193
rect 4516 1956 4523 2153
rect 4536 2107 4543 2153
rect 4556 2047 4563 2253
rect 4576 2167 4583 2213
rect 4636 2187 4643 2212
rect 4593 2167 4607 2173
rect 4496 1867 4503 1923
rect 4296 1587 4303 1693
rect 4336 1627 4343 1673
rect 4356 1647 4363 1703
rect 4316 1448 4323 1513
rect 4236 1436 4263 1443
rect 3816 1136 3833 1143
rect 3616 666 3623 773
rect 3636 727 3643 843
rect 3716 767 3723 973
rect 3776 916 3783 1033
rect 3816 928 3823 1136
rect 3856 1023 3863 1193
rect 3876 1087 3883 1233
rect 3936 1087 3943 1183
rect 3976 1147 3983 1183
rect 3936 1047 3943 1073
rect 3836 1016 3863 1023
rect 3836 987 3843 1016
rect 3856 886 3863 993
rect 3896 916 3903 993
rect 3733 700 3747 713
rect 3756 708 3763 883
rect 3736 696 3743 700
rect 3536 627 3543 663
rect 3396 396 3403 400
rect 3516 396 3523 573
rect 3556 396 3563 453
rect 3456 363 3463 394
rect 3416 356 3463 363
rect 3496 327 3503 363
rect 3536 360 3543 363
rect 3533 347 3547 360
rect 3616 307 3623 613
rect 3636 527 3643 692
rect 3676 660 3683 663
rect 3716 660 3723 663
rect 3673 647 3687 660
rect 3656 636 3673 643
rect 3656 408 3663 636
rect 3713 647 3727 660
rect 3776 647 3783 753
rect 3916 747 3923 883
rect 3916 707 3923 733
rect 3796 647 3803 693
rect 3856 587 3863 663
rect 3936 547 3943 813
rect 3976 807 3983 1053
rect 4016 1007 4023 1214
rect 4036 1183 4043 1233
rect 4096 1216 4103 1313
rect 4036 1180 4063 1183
rect 4036 1176 4067 1180
rect 4053 1167 4067 1176
rect 4116 947 4123 1183
rect 4136 1107 4143 1293
rect 4156 1127 4163 1403
rect 4236 1267 4243 1436
rect 4356 1406 4363 1453
rect 4396 1443 4403 1693
rect 4416 1467 4423 1773
rect 4516 1736 4523 1793
rect 4556 1747 4563 1913
rect 4436 1463 4443 1733
rect 4496 1700 4503 1703
rect 4456 1507 4463 1693
rect 4493 1687 4507 1700
rect 4536 1567 4543 1692
rect 4576 1507 4583 2153
rect 4676 2147 4683 2353
rect 4696 2267 4703 2393
rect 4713 2260 4727 2273
rect 4756 2267 4763 2313
rect 4716 2256 4723 2260
rect 4736 2167 4743 2223
rect 4596 1967 4603 2132
rect 4616 1987 4623 2133
rect 4647 2113 4653 2127
rect 4680 2126 4693 2127
rect 4687 2113 4693 2126
rect 4596 1887 4603 1913
rect 4616 1847 4623 1923
rect 4596 1836 4613 1843
rect 4596 1747 4603 1836
rect 4636 1736 4643 1793
rect 4676 1767 4683 2073
rect 4756 2023 4763 2213
rect 4776 2187 4783 2436
rect 4796 2367 4803 2413
rect 4816 2367 4823 2413
rect 4796 2267 4803 2332
rect 4816 2256 4823 2353
rect 4836 2287 4843 2513
rect 4896 2476 4903 2513
rect 4936 2487 4943 2673
rect 4876 2440 4883 2443
rect 4873 2427 4887 2440
rect 4856 2256 4863 2313
rect 4956 2303 4963 2733
rect 4996 2707 5003 2743
rect 5036 2607 5043 2733
rect 4996 2387 5003 2413
rect 4936 2296 4963 2303
rect 4796 2147 4803 2213
rect 4876 2187 4883 2223
rect 4916 2226 4923 2273
rect 4936 2267 4943 2296
rect 4996 2256 5003 2373
rect 5016 2347 5023 2443
rect 5033 2267 5047 2273
rect 4896 2027 4903 2213
rect 5036 2107 5043 2213
rect 4756 2016 4783 2023
rect 4696 1923 4703 2013
rect 4776 1987 4783 2016
rect 4836 1963 4843 1993
rect 4816 1956 4843 1963
rect 4696 1916 4723 1923
rect 4676 1736 4703 1744
rect 4436 1456 4463 1463
rect 4396 1436 4423 1443
rect 4456 1436 4463 1456
rect 4316 1347 4323 1373
rect 4396 1327 4403 1353
rect 4416 1347 4423 1373
rect 4176 1067 4183 1253
rect 4356 1228 4363 1313
rect 4436 1287 4443 1403
rect 4393 1220 4407 1233
rect 4396 1216 4403 1220
rect 4216 1180 4223 1183
rect 4196 1007 4203 1173
rect 4213 1167 4227 1180
rect 4336 1180 4343 1183
rect 4333 1167 4347 1180
rect 4376 1063 4383 1183
rect 4416 1147 4423 1183
rect 4416 1067 4423 1133
rect 4376 1056 4403 1063
rect 4233 947 4247 953
rect 4173 920 4187 933
rect 4176 916 4183 920
rect 4036 880 4043 883
rect 4033 867 4047 880
rect 4076 807 4083 883
rect 4116 767 4123 893
rect 4256 886 4263 1053
rect 4376 916 4383 1033
rect 4396 923 4403 1056
rect 4456 1047 4463 1233
rect 4516 1216 4523 1473
rect 4536 1243 4543 1493
rect 4536 1236 4563 1243
rect 4556 1216 4563 1236
rect 4476 1087 4483 1213
rect 4536 1180 4543 1183
rect 4533 1167 4547 1180
rect 4396 916 4423 923
rect 4156 767 4163 883
rect 4316 827 4323 883
rect 4416 847 4423 916
rect 3696 396 3703 453
rect 3816 396 3823 453
rect 3916 367 3923 493
rect 4016 467 4023 613
rect 4056 507 4063 693
rect 4076 666 4083 753
rect 4116 696 4123 753
rect 4156 696 4163 732
rect 4176 707 4183 793
rect 4136 587 4143 663
rect 4196 627 4203 773
rect 4367 756 4423 763
rect 4216 666 4223 713
rect 4276 696 4283 753
rect 4313 700 4327 713
rect 4316 696 4323 700
rect 4247 663 4260 667
rect 4247 656 4263 663
rect 4247 653 4260 656
rect 3973 400 3987 413
rect 3976 396 3983 400
rect 4016 396 4023 453
rect 3673 347 3687 352
rect 3716 327 3723 363
rect 3836 360 3843 363
rect 3876 360 3883 363
rect 3833 347 3847 360
rect 3873 347 3887 360
rect 4056 366 4063 453
rect 4133 400 4147 413
rect 4136 396 4143 400
rect 3827 316 3853 323
rect 3956 307 3963 363
rect 4087 336 4133 343
rect 3973 327 3987 333
rect 3986 320 3987 327
rect 3116 176 3123 213
rect 2976 140 2983 143
rect 2973 127 2987 140
rect 3096 107 3103 143
rect 1607 76 1643 83
rect 3176 47 3183 173
rect 3260 143 3273 147
rect 3256 136 3273 143
rect 3260 133 3273 136
rect 3296 87 3303 173
rect 3316 147 3323 213
rect 3396 176 3403 213
rect 3456 143 3463 193
rect 3516 176 3523 273
rect 3656 176 3663 293
rect 3756 146 3763 213
rect 3376 47 3383 143
rect 3416 136 3463 143
rect 3536 124 3544 143
rect 3676 140 3683 143
rect 3673 124 3687 140
rect 3776 124 3783 273
rect 3976 256 4043 263
rect 3796 188 3803 233
rect 3916 147 3923 233
rect 3956 187 3963 253
rect 3976 176 3983 256
rect 4016 176 4023 233
rect 4036 203 4043 256
rect 4036 200 4063 203
rect 4036 196 4067 200
rect 4053 187 4067 196
rect 3536 117 3783 124
rect 3836 87 3843 113
rect 3856 67 3863 143
rect 3936 127 3943 153
rect 3956 107 3963 133
rect 4036 107 4043 143
rect 4056 107 4063 133
rect 4007 93 4013 107
rect 4076 67 4083 293
rect 4116 176 4123 213
rect 4156 207 4163 363
rect 4196 287 4203 433
rect 4236 396 4243 453
rect 4276 396 4283 493
rect 4356 408 4363 713
rect 4376 707 4383 733
rect 4416 696 4423 756
rect 4436 723 4443 933
rect 4493 920 4507 933
rect 4496 916 4503 920
rect 4556 887 4563 1133
rect 4596 987 4603 1363
rect 4676 1267 4683 1673
rect 4696 1487 4703 1736
rect 4616 1087 4623 1253
rect 4716 1247 4723 1853
rect 4736 1703 4743 1793
rect 4776 1736 4783 1773
rect 4836 1747 4843 1933
rect 4856 1707 4863 2013
rect 4876 1907 4883 1954
rect 4876 1807 4883 1893
rect 4936 1887 4943 1923
rect 4996 1887 5003 1993
rect 5056 1983 5063 2833
rect 5076 2747 5083 2833
rect 5096 2827 5103 3212
rect 5116 3147 5123 3233
rect 5136 3187 5143 3263
rect 5136 2996 5143 3073
rect 5156 3027 5163 3253
rect 5176 3227 5183 3294
rect 5216 3207 5223 3263
rect 5216 3167 5223 3193
rect 5176 2996 5183 3033
rect 5196 3007 5203 3073
rect 5276 3067 5283 3253
rect 5296 3047 5303 3313
rect 5316 3266 5323 3373
rect 5336 3307 5343 3476
rect 5376 3367 5383 3473
rect 5396 3447 5403 3483
rect 5436 3427 5443 3472
rect 5496 3403 5503 3593
rect 5516 3527 5523 3673
rect 5536 3516 5543 3653
rect 5556 3647 5563 3814
rect 5576 3627 5583 3773
rect 5616 3527 5623 3783
rect 5636 3707 5643 3733
rect 5656 3707 5663 3783
rect 5600 3483 5613 3487
rect 5556 3480 5563 3483
rect 5513 3467 5527 3473
rect 5553 3467 5567 3480
rect 5596 3476 5613 3483
rect 5600 3473 5613 3476
rect 5636 3427 5643 3514
rect 5496 3396 5523 3403
rect 5456 3296 5483 3303
rect 5133 2780 5147 2793
rect 5136 2776 5143 2780
rect 5176 2776 5183 2853
rect 5156 2740 5163 2743
rect 5116 2647 5123 2732
rect 5153 2727 5167 2740
rect 5147 2696 5173 2703
rect 5196 2667 5203 2733
rect 5156 2476 5163 2573
rect 5196 2487 5203 2613
rect 5076 2427 5083 2474
rect 5116 2256 5123 2353
rect 5136 2347 5143 2443
rect 5156 2227 5163 2413
rect 5216 2287 5223 3033
rect 5336 3023 5343 3272
rect 5476 3207 5483 3296
rect 5496 3247 5503 3373
rect 5516 3367 5523 3396
rect 5556 3296 5563 3333
rect 5636 3307 5643 3413
rect 5516 3187 5523 3293
rect 5616 3227 5623 3263
rect 5336 3016 5363 3023
rect 5236 2927 5243 2994
rect 5256 2903 5263 3013
rect 5316 2907 5323 2963
rect 5256 2896 5283 2903
rect 5236 2667 5243 2853
rect 5256 2787 5263 2873
rect 5276 2827 5283 2896
rect 5293 2780 5307 2793
rect 5296 2776 5303 2780
rect 5336 2776 5343 2933
rect 5356 2787 5363 3016
rect 5376 2907 5383 3053
rect 5376 2767 5383 2793
rect 5396 2787 5403 3093
rect 5416 3007 5423 3133
rect 5433 3000 5447 3013
rect 5436 2996 5443 3000
rect 5476 2996 5483 3153
rect 5636 3127 5643 3253
rect 5656 3183 5663 3553
rect 5676 3527 5683 3633
rect 5696 3567 5703 3853
rect 5756 3816 5763 3952
rect 5816 3907 5823 4034
rect 5836 3824 5843 4113
rect 5856 3903 5863 4053
rect 5876 4036 5883 4293
rect 5896 4267 5903 4413
rect 5936 4367 5943 4513
rect 5956 4387 5963 4753
rect 5976 4707 5983 4873
rect 5976 4607 5983 4633
rect 5996 4607 6003 4913
rect 6016 4867 6023 5113
rect 6096 5076 6103 5153
rect 6116 5107 6123 5173
rect 6156 5107 6163 5393
rect 6036 5007 6043 5073
rect 6116 5007 6123 5043
rect 6036 4907 6043 4993
rect 6096 4856 6103 4953
rect 6016 4767 6023 4793
rect 5976 4567 5983 4593
rect 5996 4556 6003 4593
rect 6016 4583 6023 4693
rect 6036 4647 6043 4823
rect 6076 4820 6083 4823
rect 6073 4807 6087 4820
rect 6016 4576 6043 4583
rect 6036 4556 6043 4576
rect 6016 4520 6023 4523
rect 5973 4503 5987 4513
rect 6013 4507 6027 4520
rect 5973 4500 6003 4503
rect 5976 4496 6003 4500
rect 5936 4357 5953 4367
rect 5940 4353 5953 4357
rect 5936 4227 5943 4303
rect 5953 4267 5967 4273
rect 5976 4187 5983 4293
rect 5996 4227 6003 4496
rect 6096 4467 6103 4554
rect 5856 3896 5883 3903
rect 5796 3817 5843 3824
rect 5716 3516 5723 3693
rect 5776 3683 5783 3783
rect 5776 3676 5803 3683
rect 5776 3527 5783 3593
rect 5676 3347 5683 3473
rect 5696 3407 5703 3483
rect 5736 3447 5743 3483
rect 5736 3387 5743 3433
rect 5693 3323 5707 3333
rect 5676 3320 5707 3323
rect 5673 3316 5703 3320
rect 5673 3307 5687 3316
rect 5756 3296 5763 3453
rect 5776 3347 5783 3473
rect 5796 3447 5803 3676
rect 5816 3667 5823 3772
rect 5816 3547 5823 3653
rect 5836 3547 5843 3817
rect 5856 3747 5863 3873
rect 5876 3827 5883 3896
rect 5896 3887 5903 4003
rect 5893 3820 5907 3833
rect 5896 3816 5903 3820
rect 5856 3516 5863 3633
rect 5876 3547 5883 3773
rect 5916 3707 5923 3783
rect 5927 3696 5943 3703
rect 5896 3607 5903 3653
rect 5936 3486 5943 3696
rect 5956 3667 5963 4133
rect 5996 4047 6003 4153
rect 6016 4067 6023 4373
rect 6076 4367 6083 4453
rect 6096 4336 6103 4373
rect 6116 4367 6123 4793
rect 6136 4727 6143 4854
rect 6156 4767 6163 5033
rect 6176 4967 6183 5074
rect 6196 4687 6203 5393
rect 6216 4607 6223 5613
rect 6136 4347 6143 4593
rect 6156 4407 6163 4523
rect 6076 4300 6083 4303
rect 6036 4036 6043 4293
rect 6073 4287 6087 4300
rect 6073 4040 6087 4053
rect 6096 4043 6103 4233
rect 6116 4147 6123 4292
rect 6136 4247 6143 4293
rect 6113 4087 6127 4093
rect 6076 4036 6083 4040
rect 6096 4036 6123 4043
rect 5976 3947 5983 4033
rect 5996 3927 6003 3993
rect 6016 3847 6023 4003
rect 6056 3848 6063 4003
rect 6076 3907 6083 3973
rect 6096 3827 6103 3993
rect 5976 3816 6023 3823
rect 5976 3647 5983 3816
rect 6036 3780 6043 3783
rect 5996 3727 6003 3773
rect 6033 3767 6047 3780
rect 6076 3687 6083 3783
rect 5996 3516 6003 3553
rect 6076 3547 6083 3673
rect 5793 3343 5807 3353
rect 5793 3340 5823 3343
rect 5796 3336 5823 3340
rect 5656 3176 5683 3183
rect 5556 2996 5563 3093
rect 5456 2947 5463 2963
rect 5456 2807 5463 2933
rect 5476 2807 5483 2853
rect 5413 2780 5427 2793
rect 5416 2776 5423 2780
rect 5316 2707 5323 2743
rect 5296 2476 5303 2513
rect 5276 2440 5283 2443
rect 5236 2347 5243 2433
rect 5273 2427 5287 2440
rect 5256 2327 5263 2373
rect 5316 2367 5323 2443
rect 5256 2283 5263 2313
rect 5356 2287 5363 2733
rect 5376 2647 5383 2732
rect 5456 2687 5463 2733
rect 5376 2487 5383 2593
rect 5436 2587 5443 2673
rect 5476 2647 5483 2772
rect 5396 2507 5403 2553
rect 5416 2476 5423 2513
rect 5456 2508 5463 2633
rect 5373 2427 5387 2433
rect 5396 2367 5403 2443
rect 5236 2276 5263 2283
rect 5176 2087 5183 2273
rect 5236 2256 5243 2276
rect 5256 2187 5263 2223
rect 5036 1976 5063 1983
rect 5036 1956 5043 1976
rect 5056 1867 5063 1912
rect 5096 1827 5103 1923
rect 5113 1907 5127 1913
rect 4736 1696 4764 1703
rect 4916 1700 4923 1703
rect 4913 1687 4927 1700
rect 4776 1267 4783 1363
rect 4720 1223 4733 1227
rect 4716 1216 4733 1223
rect 4720 1213 4733 1216
rect 4616 943 4623 1073
rect 4656 1047 4663 1183
rect 4696 1180 4703 1183
rect 4693 1167 4707 1180
rect 4596 936 4623 943
rect 4596 927 4603 936
rect 4636 928 4643 973
rect 4587 916 4603 927
rect 4587 913 4600 916
rect 4520 883 4533 887
rect 4516 876 4533 883
rect 4520 873 4533 876
rect 4436 716 4463 723
rect 4456 696 4463 716
rect 4436 607 4443 663
rect 4496 627 4503 693
rect 4516 666 4523 753
rect 4676 747 4683 1113
rect 4716 1087 4723 1113
rect 4736 1007 4743 1173
rect 4716 916 4723 973
rect 4756 948 4763 1233
rect 4776 1223 4783 1253
rect 4856 1223 4863 1672
rect 4896 1406 4903 1573
rect 4936 1436 4943 1553
rect 4976 1448 4983 1633
rect 4996 1547 5003 1773
rect 5036 1743 5043 1773
rect 5016 1736 5043 1743
rect 5016 1706 5023 1736
rect 5136 1747 5143 2013
rect 5316 2007 5323 2273
rect 5356 2147 5363 2223
rect 5396 2207 5403 2223
rect 5396 2127 5403 2193
rect 5167 1963 5180 1967
rect 5167 1956 5183 1963
rect 5167 1953 5180 1956
rect 5076 1700 5083 1703
rect 5073 1687 5087 1700
rect 5116 1507 5123 1703
rect 5133 1687 5147 1693
rect 4996 1367 5003 1403
rect 5096 1400 5103 1403
rect 5093 1387 5107 1400
rect 5087 1356 5113 1363
rect 5136 1347 5143 1373
rect 5156 1327 5163 1813
rect 5176 1807 5183 1853
rect 5196 1847 5203 1912
rect 5236 1767 5243 1993
rect 5313 1960 5327 1972
rect 5316 1956 5323 1960
rect 5436 1963 5443 2353
rect 5476 2327 5483 2433
rect 5496 2287 5503 2913
rect 5516 2787 5523 2952
rect 5596 2788 5603 2893
rect 5616 2867 5623 2963
rect 5616 2787 5623 2813
rect 5656 2783 5663 3153
rect 5676 3007 5683 3176
rect 5696 3087 5703 3263
rect 5716 3107 5723 3233
rect 5736 3207 5743 3252
rect 5796 3167 5803 3293
rect 5816 3203 5823 3336
rect 5836 3307 5843 3483
rect 5916 3296 5923 3353
rect 5816 3196 5843 3203
rect 5696 3047 5703 3073
rect 5693 3000 5707 3012
rect 5696 2996 5703 3000
rect 5736 2996 5743 3053
rect 5776 3007 5783 3093
rect 5796 3027 5803 3053
rect 5676 2827 5683 2953
rect 5716 2927 5723 2963
rect 5716 2887 5723 2913
rect 5796 2867 5803 3013
rect 5636 2776 5663 2783
rect 5516 2563 5523 2733
rect 5576 2727 5583 2743
rect 5573 2707 5587 2713
rect 5516 2556 5533 2563
rect 5536 2476 5543 2553
rect 5576 2527 5583 2672
rect 5596 2507 5603 2653
rect 5616 2476 5623 2713
rect 5636 2483 5643 2776
rect 5716 2776 5723 2852
rect 5756 2783 5763 2813
rect 5816 2803 5823 3173
rect 5836 3007 5843 3196
rect 5856 3107 5863 3263
rect 5896 3187 5903 3263
rect 5896 3147 5903 3173
rect 5916 3023 5923 3113
rect 5907 3016 5923 3023
rect 5853 3000 5867 3013
rect 5856 2996 5863 3000
rect 5896 2996 5903 3013
rect 5796 2800 5823 2803
rect 5793 2796 5823 2800
rect 5793 2787 5807 2796
rect 5836 2788 5843 2933
rect 5876 2927 5883 2963
rect 5756 2776 5783 2783
rect 5696 2740 5703 2743
rect 5656 2707 5663 2733
rect 5693 2727 5707 2740
rect 5776 2743 5783 2776
rect 5873 2780 5887 2793
rect 5896 2787 5903 2933
rect 5916 2807 5923 2873
rect 5876 2776 5883 2780
rect 5776 2736 5803 2743
rect 5656 2507 5663 2653
rect 5636 2476 5663 2483
rect 5556 2440 5563 2443
rect 5553 2427 5567 2440
rect 5456 2103 5463 2273
rect 5476 2147 5483 2233
rect 5496 2220 5503 2223
rect 5493 2207 5507 2220
rect 5456 2096 5483 2103
rect 5456 1987 5463 2073
rect 5476 2027 5483 2096
rect 5416 1956 5443 1963
rect 5456 1956 5463 1973
rect 5256 1736 5263 1873
rect 5296 1847 5303 1923
rect 5336 1887 5343 1923
rect 5296 1706 5303 1753
rect 5356 1736 5363 1773
rect 5396 1736 5403 1813
rect 5416 1747 5423 1956
rect 5536 1963 5543 2033
rect 5556 2007 5563 2223
rect 5576 2167 5583 2413
rect 5576 1968 5583 2153
rect 5596 2087 5603 2373
rect 5616 2287 5623 2313
rect 5636 2263 5643 2433
rect 5656 2347 5663 2476
rect 5616 2256 5643 2263
rect 5656 2256 5663 2312
rect 5676 2307 5683 2513
rect 5696 2487 5703 2573
rect 5736 2476 5743 2732
rect 5756 2507 5763 2733
rect 5776 2476 5783 2713
rect 5796 2487 5803 2736
rect 5816 2707 5823 2743
rect 5856 2740 5863 2743
rect 5853 2727 5867 2740
rect 5896 2667 5903 2733
rect 5916 2727 5923 2793
rect 5956 2783 5963 3473
rect 5976 3427 5983 3483
rect 6016 3407 6023 3483
rect 6076 3467 6083 3512
rect 6016 3367 6023 3393
rect 6036 3343 6043 3453
rect 6076 3387 6083 3453
rect 6016 3336 6043 3343
rect 6016 3296 6023 3336
rect 5976 3047 5983 3193
rect 5996 3067 6003 3263
rect 6036 3260 6043 3263
rect 6033 3247 6047 3260
rect 5936 2776 5963 2783
rect 5976 2776 5983 3033
rect 5996 3007 6003 3053
rect 6036 3008 6043 3212
rect 6096 3127 6103 3773
rect 6116 3767 6123 4036
rect 6136 3967 6143 4173
rect 6156 4167 6163 4372
rect 6176 4123 6183 4473
rect 6196 4367 6203 4512
rect 6196 4187 6203 4332
rect 6156 4116 6183 4123
rect 6156 4047 6163 4116
rect 6216 4107 6223 4393
rect 6187 4093 6193 4107
rect 6136 3743 6143 3813
rect 6156 3807 6163 3913
rect 6116 3736 6143 3743
rect 6116 3527 6123 3736
rect 6156 3567 6163 3772
rect 6196 3727 6203 4003
rect 6156 3516 6163 3553
rect 6216 3523 6223 3953
rect 6236 3687 6243 4452
rect 6216 3516 6243 3523
rect 6116 3427 6123 3473
rect 6136 3447 6143 3483
rect 6176 3463 6183 3483
rect 6156 3456 6183 3463
rect 6156 3387 6163 3456
rect 6176 3296 6183 3413
rect 6196 3407 6203 3453
rect 6156 3247 6163 3263
rect 6076 2996 6083 3093
rect 6156 3028 6163 3233
rect 6196 3187 6203 3263
rect 6216 3227 6223 3294
rect 6176 3176 6193 3183
rect 6176 3047 6183 3176
rect 6007 2963 6020 2967
rect 6007 2956 6023 2963
rect 6007 2953 6020 2956
rect 6056 2847 6063 2963
rect 5936 2746 5943 2776
rect 6036 2740 6043 2743
rect 5993 2727 6007 2732
rect 6033 2727 6047 2740
rect 6076 2647 6083 2774
rect 5816 2387 5823 2493
rect 5896 2488 5903 2613
rect 6096 2527 6103 2893
rect 6116 2867 6123 3013
rect 6193 3000 6207 3013
rect 6196 2996 6203 3000
rect 6216 2907 6223 2963
rect 6156 2776 6163 2873
rect 6236 2863 6243 3516
rect 6216 2856 6243 2863
rect 6196 2776 6203 2853
rect 6136 2647 6143 2743
rect 6176 2740 6183 2743
rect 6173 2727 6187 2740
rect 5936 2496 5973 2503
rect 5936 2476 5943 2496
rect 5836 2427 5843 2473
rect 5976 2447 5983 2493
rect 5696 2256 5703 2353
rect 5736 2267 5743 2293
rect 5616 2047 5623 2256
rect 5636 2187 5643 2213
rect 5720 2223 5733 2227
rect 5716 2216 5733 2223
rect 5720 2213 5733 2216
rect 5653 1987 5667 1993
rect 5536 1956 5563 1963
rect 5476 1887 5483 1923
rect 5196 1700 5203 1703
rect 5176 1627 5183 1693
rect 5193 1687 5207 1700
rect 5236 1687 5243 1703
rect 5236 1587 5243 1673
rect 5256 1436 5263 1473
rect 5176 1367 5183 1434
rect 4776 1216 4803 1223
rect 4836 1216 4883 1223
rect 4773 1167 4787 1173
rect 4876 1167 4883 1216
rect 4736 880 4743 883
rect 4733 867 4747 880
rect 4756 696 4763 793
rect 4796 707 4803 1153
rect 4896 1047 4903 1213
rect 4936 1180 4943 1183
rect 4933 1167 4947 1180
rect 4376 396 4383 493
rect 4256 327 4263 363
rect 4296 287 4303 363
rect 4316 247 4323 293
rect 4396 247 4403 363
rect 4436 360 4443 363
rect 4433 347 4447 360
rect 4156 176 4163 193
rect 4393 180 4407 193
rect 4396 176 4403 180
rect 4436 176 4443 213
rect 4476 146 4483 233
rect 4496 227 4503 573
rect 4536 547 4543 613
rect 4616 587 4623 652
rect 4656 567 4663 694
rect 4696 567 4703 663
rect 4736 627 4743 663
rect 4776 660 4783 663
rect 4773 647 4787 660
rect 4596 427 4603 513
rect 4596 396 4603 413
rect 4536 360 4543 363
rect 4533 347 4547 360
rect 4576 307 4583 363
rect 4576 227 4583 293
rect 4536 176 4543 213
rect 4596 203 4603 313
rect 4636 307 4643 453
rect 4656 327 4663 553
rect 4713 400 4727 413
rect 4716 396 4723 400
rect 4696 360 4703 363
rect 4736 360 4743 363
rect 4693 347 4707 360
rect 4733 347 4747 360
rect 4776 347 4783 393
rect 4796 366 4803 653
rect 4816 408 4823 933
rect 4876 916 4883 993
rect 4913 920 4927 933
rect 4936 927 4943 1153
rect 4916 916 4923 920
rect 4956 887 4963 993
rect 5016 948 5023 1213
rect 5036 1186 5043 1253
rect 5196 1247 5203 1373
rect 5216 1347 5223 1373
rect 5236 1307 5243 1403
rect 5296 1387 5303 1692
rect 5376 1607 5383 1703
rect 5336 1436 5343 1573
rect 5376 1436 5383 1593
rect 5416 1443 5423 1693
rect 5436 1567 5443 1813
rect 5496 1736 5503 1893
rect 5516 1807 5523 1923
rect 5536 1736 5543 1813
rect 5556 1747 5563 1956
rect 5656 1956 5663 1973
rect 5596 1763 5603 1923
rect 5696 1767 5703 1973
rect 5736 1956 5743 2213
rect 5756 1987 5763 2333
rect 5776 2187 5783 2353
rect 5876 2347 5883 2443
rect 5896 2343 5903 2413
rect 5916 2367 5923 2443
rect 5896 2336 5923 2343
rect 5796 2267 5803 2333
rect 5836 2256 5843 2333
rect 5880 2324 5893 2327
rect 5876 2313 5893 2324
rect 5876 2256 5883 2313
rect 5896 2267 5903 2292
rect 5856 2220 5863 2223
rect 5853 2207 5867 2220
rect 5776 1987 5783 2033
rect 5773 1960 5787 1973
rect 5776 1956 5783 1960
rect 5796 1867 5803 1923
rect 5576 1756 5603 1763
rect 5476 1683 5483 1703
rect 5476 1676 5503 1683
rect 5496 1507 5503 1676
rect 5516 1607 5523 1703
rect 5416 1436 5443 1443
rect 5496 1436 5503 1493
rect 5556 1463 5563 1693
rect 5536 1456 5563 1463
rect 5176 1236 5193 1243
rect 5116 1127 5123 1183
rect 5156 1107 5163 1193
rect 5176 947 5183 1236
rect 5356 1227 5363 1403
rect 5396 1400 5403 1403
rect 5393 1387 5407 1400
rect 5236 1147 5243 1183
rect 5053 920 5067 933
rect 5056 916 5063 920
rect 4856 703 4863 883
rect 4896 880 4903 883
rect 4893 867 4907 880
rect 4976 867 4983 913
rect 4993 867 5007 872
rect 4836 696 4863 703
rect 4836 607 4843 696
rect 4936 487 4943 733
rect 4976 696 4983 753
rect 5116 727 5123 933
rect 5196 916 5203 953
rect 5176 827 5183 883
rect 5196 807 5203 853
rect 5076 666 5083 713
rect 5176 696 5183 773
rect 5156 660 5163 663
rect 5153 647 5167 660
rect 4916 366 4923 433
rect 5016 396 5023 473
rect 5056 366 5063 473
rect 5116 396 5163 403
rect 4576 196 4603 203
rect 4576 176 4583 196
rect 4616 146 4623 273
rect 4716 247 4723 313
rect 4676 176 4683 233
rect 4756 187 4763 253
rect 4136 87 4143 143
rect 4276 107 4283 132
rect 4476 87 4483 132
rect 4696 67 4703 143
rect 4776 107 4783 333
rect 4796 207 4803 352
rect 4796 146 4803 193
rect 4856 176 4863 253
rect 4876 107 4883 143
rect 4916 67 4923 352
rect 4996 227 5003 363
rect 5056 327 5063 352
rect 4973 180 4987 193
rect 4976 176 4983 180
rect 5076 146 5083 193
rect 5136 176 5143 253
rect 5156 207 5163 396
rect 5176 287 5183 473
rect 5216 423 5223 883
rect 5256 787 5263 1113
rect 5276 927 5283 1151
rect 5316 1127 5323 1214
rect 5373 1220 5387 1233
rect 5376 1216 5383 1220
rect 5336 1167 5343 1193
rect 5356 1087 5363 1153
rect 5396 967 5403 1183
rect 5313 947 5327 953
rect 5436 948 5443 1436
rect 5476 1400 5483 1403
rect 5473 1387 5487 1400
rect 5536 1367 5543 1456
rect 5576 1443 5583 1756
rect 5596 1627 5603 1733
rect 5656 1700 5663 1703
rect 5653 1687 5667 1700
rect 5696 1687 5704 1703
rect 5736 1706 5743 1753
rect 5716 1663 5723 1693
rect 5707 1656 5723 1663
rect 5596 1467 5603 1613
rect 5556 1436 5583 1443
rect 5616 1436 5623 1553
rect 5656 1436 5663 1493
rect 5676 1447 5683 1593
rect 5313 920 5327 933
rect 5456 943 5463 1233
rect 5536 1216 5543 1332
rect 5556 1247 5563 1436
rect 5576 1227 5583 1353
rect 5456 936 5483 943
rect 5316 916 5323 920
rect 5276 843 5283 873
rect 5296 863 5303 883
rect 5296 856 5323 863
rect 5276 836 5303 843
rect 5296 783 5303 836
rect 5316 803 5323 856
rect 5336 827 5343 872
rect 5316 796 5343 803
rect 5296 776 5323 783
rect 5276 708 5283 753
rect 5316 696 5323 776
rect 5336 707 5343 796
rect 5376 703 5383 773
rect 5396 727 5403 932
rect 5476 928 5483 936
rect 5516 927 5523 1183
rect 5596 1186 5603 1403
rect 5696 1403 5703 1652
rect 5676 1396 5703 1403
rect 5576 947 5583 1173
rect 5596 916 5603 953
rect 5616 947 5623 1313
rect 5636 1227 5643 1273
rect 5676 1216 5683 1396
rect 5716 1327 5723 1473
rect 5736 1447 5743 1553
rect 5756 1527 5763 1773
rect 5796 1736 5803 1813
rect 5836 1787 5843 2073
rect 5856 1967 5863 2193
rect 5916 2067 5923 2336
rect 5936 2267 5943 2313
rect 5996 2307 6003 2513
rect 6073 2480 6087 2493
rect 6076 2476 6083 2480
rect 6016 2268 6023 2393
rect 6056 2367 6063 2443
rect 6096 2363 6103 2443
rect 6096 2356 6123 2363
rect 5936 2007 5943 2213
rect 5956 2047 5963 2223
rect 5893 1960 5907 1973
rect 5976 1968 5983 2193
rect 6036 2167 6043 2213
rect 5896 1956 5903 1960
rect 6016 1956 6023 1993
rect 6056 1987 6063 2293
rect 6076 2226 6083 2313
rect 6056 1956 6063 1973
rect 6096 1967 6103 2333
rect 6116 2287 6123 2356
rect 6136 2256 6143 2293
rect 6176 2256 6183 2373
rect 6216 2347 6223 2856
rect 5976 1926 5983 1954
rect 5833 1740 5847 1752
rect 5876 1747 5883 1923
rect 5836 1736 5843 1740
rect 5787 1676 5813 1683
rect 5856 1667 5863 1703
rect 5756 1463 5763 1513
rect 5756 1456 5783 1463
rect 5776 1436 5783 1456
rect 5820 1443 5833 1447
rect 5816 1436 5833 1443
rect 5820 1433 5833 1436
rect 5716 1216 5723 1253
rect 5736 1227 5743 1293
rect 5696 1180 5703 1183
rect 5693 1167 5707 1180
rect 5636 916 5643 953
rect 5356 696 5403 703
rect 5436 696 5443 773
rect 5496 743 5503 883
rect 5496 736 5523 743
rect 5256 660 5263 663
rect 5253 647 5267 660
rect 5216 416 5243 423
rect 5236 396 5243 416
rect 5273 400 5287 413
rect 5276 396 5283 400
rect 5316 367 5323 513
rect 5336 427 5343 653
rect 5356 403 5363 696
rect 5416 607 5423 663
rect 5336 396 5363 403
rect 5396 396 5403 593
rect 5496 427 5503 713
rect 5516 707 5523 736
rect 5536 727 5543 913
rect 5567 883 5580 887
rect 5567 876 5583 883
rect 5567 873 5580 876
rect 5616 847 5623 883
rect 5556 696 5563 773
rect 5536 587 5543 652
rect 5576 487 5583 652
rect 5636 627 5643 853
rect 5676 703 5683 933
rect 5696 887 5703 1073
rect 5756 1047 5763 1333
rect 5816 1327 5823 1373
rect 5776 1267 5783 1293
rect 5816 1216 5823 1313
rect 5836 1247 5843 1393
rect 5856 1307 5863 1632
rect 5876 1447 5883 1693
rect 5896 1467 5903 1853
rect 5916 1487 5923 1773
rect 5996 1736 6003 1853
rect 6076 1748 6083 1923
rect 6116 1787 6123 2053
rect 6216 1984 6223 2293
rect 6176 1977 6223 1984
rect 6056 1736 6073 1743
rect 5936 1667 5943 1693
rect 5976 1627 5983 1703
rect 5936 1467 5943 1573
rect 5956 1468 5963 1513
rect 5913 1440 5927 1452
rect 5996 1447 6003 1553
rect 6056 1547 6063 1736
rect 6176 1706 6183 1977
rect 6096 1527 6103 1703
rect 6136 1448 6143 1703
rect 5916 1436 5923 1440
rect 5896 1400 5903 1403
rect 5856 1216 5863 1293
rect 5876 1223 5883 1393
rect 5893 1387 5907 1400
rect 5936 1383 5943 1403
rect 5916 1376 5943 1383
rect 5916 1327 5923 1376
rect 5916 1227 5923 1292
rect 5876 1216 5903 1223
rect 5836 1180 5843 1183
rect 5833 1167 5847 1180
rect 5836 1127 5843 1153
rect 5896 1067 5903 1216
rect 5936 1216 5943 1333
rect 5976 1287 5983 1393
rect 5996 1367 6003 1433
rect 5976 1216 5983 1273
rect 6056 1223 6063 1392
rect 6076 1247 6083 1373
rect 6096 1367 6103 1403
rect 6136 1247 6143 1434
rect 6156 1387 6163 1513
rect 6036 1216 6063 1223
rect 6073 1220 6087 1233
rect 6076 1216 6083 1220
rect 6036 1186 6043 1216
rect 5916 1147 5923 1173
rect 5956 1127 5963 1183
rect 5716 928 5723 953
rect 5796 916 5803 973
rect 5816 927 5823 953
rect 5656 696 5683 703
rect 5716 696 5723 773
rect 5756 696 5763 853
rect 5776 847 5783 883
rect 5836 867 5843 973
rect 5896 928 5903 1032
rect 5936 916 5943 973
rect 6056 943 6063 1173
rect 6096 1147 6103 1183
rect 6036 936 6063 943
rect 6036 928 6043 936
rect 6076 916 6083 973
rect 6096 927 6103 1053
rect 5867 883 5880 887
rect 5867 876 5883 883
rect 5867 873 5880 876
rect 5816 856 5833 863
rect 5776 747 5783 833
rect 5433 400 5447 413
rect 5436 396 5443 400
rect 5216 287 5223 363
rect 5336 347 5343 396
rect 5376 360 5383 363
rect 5373 347 5387 360
rect 5296 176 5303 273
rect 5416 267 5423 363
rect 5496 347 5503 413
rect 5467 333 5473 347
rect 4956 107 4963 143
rect 5016 127 5023 143
rect 5156 140 5163 143
rect 5153 127 5167 140
rect 5356 143 5363 213
rect 5436 176 5443 213
rect 5476 143 5483 193
rect 5516 167 5523 413
rect 5596 396 5603 593
rect 5656 547 5663 696
rect 5796 666 5803 693
rect 5736 587 5743 663
rect 5796 587 5803 652
rect 5656 396 5663 473
rect 5556 360 5563 363
rect 5616 360 5623 363
rect 5553 347 5567 360
rect 5613 347 5627 360
rect 5676 343 5683 394
rect 5696 367 5703 493
rect 5656 336 5683 343
rect 5576 176 5583 213
rect 5616 176 5623 253
rect 5656 207 5663 336
rect 5696 307 5703 332
rect 5716 327 5723 533
rect 5816 507 5823 856
rect 5856 696 5863 773
rect 5876 747 5883 853
rect 5916 827 5923 883
rect 5896 696 5903 753
rect 5936 707 5943 733
rect 5956 708 5963 773
rect 5976 747 5983 913
rect 5996 787 6003 853
rect 6016 723 6023 883
rect 6056 880 6063 883
rect 6053 867 6067 880
rect 6036 727 6043 853
rect 6056 827 6063 853
rect 5996 716 6023 723
rect 5996 703 6003 716
rect 5976 696 6003 703
rect 5836 507 5843 613
rect 5793 428 5807 433
rect 5836 407 5843 472
rect 5736 307 5743 353
rect 5676 146 5683 233
rect 5716 207 5723 253
rect 5776 247 5783 363
rect 5816 356 5843 363
rect 5773 180 5787 193
rect 5796 187 5803 253
rect 5776 176 5783 180
rect 5316 136 5363 143
rect 5396 140 5403 143
rect 5016 116 5033 127
rect 5020 113 5033 116
rect 5393 127 5407 140
rect 5456 136 5483 143
rect 5556 140 5563 143
rect 5553 127 5567 140
rect 5596 107 5603 143
rect 5816 107 5823 333
rect 5836 307 5843 356
rect 5836 207 5843 233
rect 5856 183 5863 493
rect 5876 347 5883 613
rect 5896 467 5903 493
rect 5936 396 5943 653
rect 5956 627 5963 694
rect 5976 667 5983 696
rect 6056 696 6063 773
rect 6096 703 6103 873
rect 6096 696 6123 703
rect 5976 408 5983 632
rect 5996 407 6003 453
rect 5836 176 5863 183
rect 5896 176 5903 233
rect 5916 207 5923 363
rect 5936 176 5943 333
rect 5836 146 5843 176
rect 5976 67 5983 313
rect 6016 203 6023 633
rect 6036 587 6043 663
rect 6116 467 6123 696
rect 6036 407 6043 433
rect 6056 396 6063 453
rect 6093 400 6107 413
rect 6136 407 6143 1172
rect 6096 396 6103 400
rect 5996 196 6023 203
rect 5996 146 6003 196
rect 6036 176 6043 353
rect 6076 327 6083 363
rect 6156 247 6163 853
rect 6176 427 6183 1692
rect 6196 1667 6203 1733
rect 6196 1406 6203 1533
rect 6196 207 6203 1013
rect 6016 107 6023 143
rect 6076 67 6083 143
rect 6216 107 6223 1952
rect 6236 1627 6243 2833
rect 6236 327 6243 1613
<< m3contact >>
rect 413 6193 427 6207
rect 313 6133 327 6147
rect 113 6114 127 6128
rect 153 6114 167 6128
rect 233 6114 247 6128
rect 273 6114 287 6128
rect 133 6053 147 6067
rect 353 6110 367 6124
rect 333 6073 347 6087
rect 493 6153 507 6167
rect 453 6114 467 6128
rect 333 6033 347 6047
rect 313 5993 327 6007
rect 313 5953 327 5967
rect 13 5933 27 5947
rect 93 5933 107 5947
rect 173 5933 187 5947
rect 253 5933 267 5947
rect 33 5893 47 5907
rect 93 5894 107 5908
rect 153 5893 167 5907
rect 13 5852 27 5866
rect 73 5852 87 5866
rect 113 5852 127 5866
rect 153 5852 167 5866
rect 33 5653 47 5667
rect 213 5894 227 5908
rect 253 5894 267 5908
rect 453 6053 467 6067
rect 373 5933 387 5947
rect 373 5894 387 5908
rect 433 5892 447 5906
rect 233 5852 247 5866
rect 313 5852 327 5866
rect 353 5852 367 5866
rect 393 5852 407 5866
rect 433 5852 447 5866
rect 513 6073 527 6087
rect 473 6033 487 6047
rect 613 6213 627 6227
rect 893 6213 907 6227
rect 573 6153 587 6167
rect 833 6193 847 6207
rect 673 6153 687 6167
rect 653 6114 667 6128
rect 533 6053 547 6067
rect 733 6114 747 6128
rect 593 5953 607 5967
rect 653 5993 667 6007
rect 593 5913 607 5927
rect 633 5913 647 5927
rect 493 5894 507 5908
rect 533 5894 547 5908
rect 373 5833 387 5847
rect 273 5813 287 5827
rect 393 5813 407 5827
rect 393 5653 407 5667
rect 373 5633 387 5647
rect 113 5593 127 5607
rect 153 5593 167 5607
rect 13 5552 27 5566
rect 93 5552 107 5566
rect 113 5533 127 5547
rect 53 5453 67 5467
rect 153 5553 167 5567
rect 133 5513 147 5527
rect 273 5594 287 5608
rect 313 5594 327 5608
rect 193 5552 207 5566
rect 253 5552 267 5566
rect 173 5513 187 5527
rect 153 5394 167 5408
rect 113 5374 127 5388
rect 153 5373 167 5387
rect 73 5333 87 5347
rect 53 5273 67 5287
rect 133 5332 147 5346
rect 633 5852 647 5866
rect 573 5753 587 5767
rect 553 5733 567 5747
rect 493 5713 507 5727
rect 533 5633 547 5647
rect 493 5593 507 5607
rect 573 5594 587 5608
rect 333 5533 347 5547
rect 313 5473 327 5487
rect 213 5413 227 5427
rect 193 5273 207 5287
rect 93 5173 107 5187
rect 173 5173 187 5187
rect 73 5073 87 5087
rect 133 5074 147 5088
rect 53 5013 67 5027
rect 33 4854 47 4868
rect 73 4854 87 4868
rect 153 5033 167 5047
rect 133 5013 147 5027
rect 13 4593 27 4607
rect 133 4853 147 4867
rect 73 4793 87 4807
rect 53 4613 67 4627
rect 33 4553 47 4567
rect 273 5374 287 5388
rect 373 5493 387 5507
rect 413 5513 427 5527
rect 393 5473 407 5487
rect 433 5413 447 5427
rect 393 5374 407 5388
rect 433 5373 447 5387
rect 253 5332 267 5346
rect 332 5332 346 5346
rect 293 5293 307 5307
rect 233 5074 247 5088
rect 273 5074 287 5088
rect 313 5074 327 5088
rect 193 5033 207 5047
rect 173 4973 187 4987
rect 413 5332 427 5346
rect 493 5553 507 5567
rect 593 5553 607 5567
rect 553 5533 567 5547
rect 473 5453 487 5467
rect 533 5513 547 5527
rect 553 5393 567 5407
rect 353 5074 367 5088
rect 453 5032 467 5046
rect 253 4973 267 4987
rect 353 4973 367 4987
rect 533 5332 547 5346
rect 493 5273 507 5287
rect 493 5213 507 5227
rect 433 4953 447 4967
rect 473 4953 487 4967
rect 193 4893 207 4907
rect 413 4893 427 4907
rect 213 4854 227 4868
rect 473 4913 487 4927
rect 353 4854 367 4868
rect 393 4854 407 4868
rect 153 4793 167 4807
rect 93 4613 107 4627
rect 153 4593 167 4607
rect 93 4554 107 4568
rect 173 4554 187 4568
rect 73 4513 87 4527
rect 113 4512 127 4526
rect 173 4453 187 4467
rect 53 4334 67 4348
rect 93 4334 107 4348
rect 133 4334 147 4348
rect 173 4334 187 4348
rect 53 4073 67 4087
rect 173 4273 187 4287
rect 232 4645 246 4659
rect 312 4554 326 4568
rect 333 4553 347 4567
rect 753 6053 767 6067
rect 773 6053 787 6067
rect 773 5993 787 6007
rect 713 5973 727 5987
rect 733 5913 747 5927
rect 893 6114 907 6128
rect 933 6114 947 6128
rect 833 6013 847 6027
rect 813 5973 827 5987
rect 873 5973 887 5987
rect 793 5913 807 5927
rect 753 5852 767 5866
rect 713 5813 727 5827
rect 693 5713 707 5727
rect 753 5733 767 5747
rect 633 5594 647 5608
rect 673 5594 687 5608
rect 713 5594 727 5608
rect 733 5553 747 5567
rect 713 5533 727 5547
rect 653 5513 667 5527
rect 713 5433 727 5447
rect 653 5374 667 5388
rect 613 5333 627 5347
rect 593 5293 607 5307
rect 533 5153 547 5167
rect 573 5153 587 5167
rect 533 5113 547 5127
rect 673 5332 687 5346
rect 773 5633 787 5647
rect 753 5533 767 5547
rect 893 5894 907 5908
rect 933 5894 947 5908
rect 913 5852 927 5866
rect 953 5853 967 5867
rect 873 5813 887 5827
rect 813 5733 827 5747
rect 893 5713 907 5727
rect 793 5593 807 5607
rect 833 5594 847 5608
rect 1073 6193 1087 6207
rect 1213 6193 1227 6207
rect 1033 6114 1047 6128
rect 1213 6153 1227 6167
rect 1433 6153 1447 6167
rect 1533 6153 1547 6167
rect 1133 6114 1147 6128
rect 1173 6114 1187 6128
rect 1053 6072 1067 6086
rect 1093 6072 1107 6086
rect 1273 6113 1287 6127
rect 1153 6072 1167 6086
rect 1133 6053 1147 6067
rect 1053 6013 1067 6027
rect 1133 5893 1147 5907
rect 973 5753 987 5767
rect 973 5653 987 5667
rect 953 5633 967 5647
rect 993 5633 1007 5647
rect 873 5593 887 5607
rect 913 5594 927 5608
rect 953 5594 967 5608
rect 993 5594 1007 5608
rect 793 5553 807 5567
rect 853 5553 867 5567
rect 833 5473 847 5487
rect 913 5533 927 5547
rect 872 5513 886 5527
rect 893 5513 907 5527
rect 873 5492 887 5506
rect 793 5393 807 5407
rect 713 5332 727 5346
rect 633 5293 647 5307
rect 693 5293 707 5307
rect 613 5173 627 5187
rect 593 5133 607 5147
rect 653 5113 667 5127
rect 613 5074 627 5088
rect 553 5032 567 5046
rect 633 5033 647 5047
rect 673 5073 687 5087
rect 653 4993 667 5007
rect 653 4953 667 4967
rect 633 4933 647 4947
rect 553 4913 567 4927
rect 573 4893 587 4907
rect 553 4873 567 4887
rect 453 4812 467 4826
rect 393 4733 407 4747
rect 533 4853 547 4867
rect 553 4812 567 4826
rect 613 4812 627 4826
rect 513 4613 527 4627
rect 373 4573 387 4587
rect 413 4573 427 4587
rect 513 4573 527 4587
rect 573 4573 587 4587
rect 493 4552 507 4566
rect 593 4553 607 4567
rect 473 4533 487 4547
rect 273 4493 287 4507
rect 353 4513 367 4527
rect 493 4513 507 4527
rect 473 4473 487 4487
rect 393 4453 407 4467
rect 373 4413 387 4427
rect 293 4393 307 4407
rect 333 4393 347 4407
rect 233 4353 247 4367
rect 233 4193 247 4207
rect 193 4073 207 4087
rect 213 4053 227 4067
rect 153 4034 167 4048
rect 193 4034 207 4048
rect 133 3993 147 4007
rect 193 3993 207 4007
rect 113 3973 127 3987
rect 93 3933 107 3947
rect 113 3814 127 3828
rect 73 3772 87 3786
rect 193 3873 207 3887
rect 253 4113 267 4127
rect 553 4512 567 4526
rect 593 4512 607 4526
rect 713 5273 727 5287
rect 773 5332 787 5346
rect 813 5332 827 5346
rect 753 5233 767 5247
rect 1233 6072 1247 6086
rect 1253 6073 1267 6087
rect 1193 6053 1207 6067
rect 1273 6072 1287 6086
rect 1413 6072 1427 6086
rect 1293 6013 1307 6027
rect 1333 5953 1347 5967
rect 1373 5953 1387 5967
rect 1173 5933 1187 5947
rect 1253 5933 1267 5947
rect 1153 5753 1167 5767
rect 1213 5894 1227 5908
rect 1313 5893 1327 5907
rect 1233 5852 1247 5866
rect 1313 5852 1327 5866
rect 1293 5773 1307 5787
rect 1273 5753 1287 5767
rect 1173 5713 1187 5727
rect 1033 5693 1047 5707
rect 1193 5653 1207 5667
rect 1053 5594 1067 5608
rect 1193 5593 1207 5607
rect 1233 5594 1247 5608
rect 1313 5733 1327 5747
rect 1173 5573 1187 5587
rect 1033 5533 1047 5547
rect 1173 5533 1187 5547
rect 973 5513 987 5527
rect 1013 5513 1027 5527
rect 933 5433 947 5447
rect 933 5412 947 5426
rect 913 5393 927 5407
rect 913 5332 927 5346
rect 1133 5473 1147 5487
rect 1113 5453 1127 5467
rect 993 5374 1007 5388
rect 1053 5374 1067 5388
rect 1093 5374 1107 5388
rect 973 5233 987 5247
rect 873 5213 887 5227
rect 1033 5332 1047 5346
rect 1073 5332 1087 5346
rect 1313 5573 1327 5587
rect 1253 5513 1267 5527
rect 1233 5374 1247 5388
rect 1293 5413 1307 5427
rect 1313 5393 1327 5407
rect 1413 5933 1427 5947
rect 1373 5894 1387 5908
rect 1533 6114 1547 6128
rect 1593 6114 1607 6128
rect 1653 6114 1667 6128
rect 1593 6072 1607 6086
rect 1673 6072 1687 6086
rect 1553 6053 1567 6067
rect 1613 6053 1627 6067
rect 1593 5993 1607 6007
rect 1513 5953 1527 5967
rect 1573 5953 1587 5967
rect 1433 5913 1447 5927
rect 1533 5894 1547 5908
rect 1573 5894 1587 5908
rect 1393 5852 1407 5866
rect 1433 5852 1447 5866
rect 1353 5633 1367 5647
rect 1393 5594 1407 5608
rect 1553 5813 1567 5827
rect 1753 6114 1767 6128
rect 1793 6114 1807 6128
rect 1833 6114 1847 6128
rect 1753 6073 1767 6087
rect 1773 6053 1787 6067
rect 1733 6013 1747 6027
rect 1713 5933 1727 5947
rect 1633 5894 1647 5908
rect 1693 5894 1707 5908
rect 1653 5852 1667 5866
rect 1813 5953 1827 5967
rect 1773 5894 1787 5908
rect 1733 5853 1747 5867
rect 1713 5813 1727 5827
rect 1513 5713 1527 5727
rect 1613 5713 1627 5727
rect 1493 5653 1507 5667
rect 1473 5594 1487 5608
rect 1553 5653 1567 5667
rect 1373 5552 1387 5566
rect 1473 5553 1487 5567
rect 1533 5552 1547 5566
rect 1573 5533 1587 5547
rect 1373 5433 1387 5447
rect 1553 5513 1567 5527
rect 1453 5413 1467 5427
rect 1493 5413 1507 5427
rect 1153 5332 1167 5346
rect 1253 5333 1267 5347
rect 1373 5373 1387 5387
rect 1413 5373 1427 5387
rect 1293 5332 1307 5346
rect 1353 5332 1367 5346
rect 1213 5293 1227 5307
rect 1293 5253 1307 5267
rect 993 5193 1007 5207
rect 1073 5193 1087 5207
rect 1133 5193 1147 5207
rect 1033 5153 1047 5167
rect 973 5133 987 5147
rect 833 5113 847 5127
rect 953 5113 967 5127
rect 732 5093 746 5107
rect 753 5093 767 5107
rect 713 5074 727 5088
rect 753 5032 767 5046
rect 732 5013 746 5027
rect 773 4993 787 5007
rect 873 5074 887 5088
rect 913 5074 927 5088
rect 853 5033 867 5047
rect 813 4993 827 5007
rect 772 4972 786 4986
rect 793 4973 807 4987
rect 733 4953 747 4967
rect 873 4953 887 4967
rect 773 4893 787 4907
rect 813 4893 827 4907
rect 733 4854 747 4868
rect 673 4812 687 4826
rect 753 4812 767 4826
rect 713 4793 727 4807
rect 833 4854 847 4868
rect 953 5033 967 5047
rect 913 5013 927 5027
rect 913 4992 927 5006
rect 913 4933 927 4947
rect 913 4912 927 4926
rect 893 4853 907 4867
rect 793 4813 807 4827
rect 773 4793 787 4807
rect 653 4733 667 4747
rect 733 4733 747 4747
rect 633 4613 647 4627
rect 693 4554 707 4568
rect 753 4613 767 4627
rect 813 4793 827 4807
rect 873 4573 887 4587
rect 793 4554 807 4568
rect 833 4554 847 4568
rect 633 4512 647 4526
rect 673 4512 687 4526
rect 713 4512 727 4526
rect 753 4513 767 4527
rect 813 4512 827 4526
rect 573 4473 587 4487
rect 613 4473 627 4487
rect 693 4473 707 4487
rect 613 4373 627 4387
rect 373 4334 387 4348
rect 433 4333 447 4347
rect 493 4334 507 4348
rect 533 4334 547 4348
rect 573 4334 587 4348
rect 393 4273 407 4287
rect 353 4233 367 4247
rect 393 4233 407 4247
rect 373 4113 387 4127
rect 293 4073 307 4087
rect 273 4053 287 4067
rect 313 4034 327 4048
rect 353 4034 367 4048
rect 353 3953 367 3967
rect 473 4292 487 4306
rect 433 4153 447 4167
rect 393 4033 407 4047
rect 433 4034 447 4048
rect 653 4293 667 4307
rect 633 4273 647 4287
rect 593 4113 607 4127
rect 533 4073 547 4087
rect 573 4034 587 4048
rect 633 4013 647 4027
rect 413 3992 427 4006
rect 453 3992 467 4006
rect 493 3993 507 4007
rect 293 3933 307 3947
rect 373 3933 387 3947
rect 433 3953 447 3967
rect 413 3913 427 3927
rect 533 3933 547 3947
rect 433 3893 447 3907
rect 393 3873 407 3887
rect 233 3814 247 3828
rect 393 3833 407 3847
rect 293 3813 307 3827
rect 353 3814 367 3828
rect 413 3814 427 3828
rect 173 3773 187 3787
rect 153 3753 167 3767
rect 213 3753 227 3767
rect 253 3733 267 3747
rect 173 3693 187 3707
rect 93 3653 107 3667
rect 133 3653 147 3667
rect 333 3753 347 3767
rect 193 3633 207 3647
rect 292 3633 306 3647
rect 313 3633 327 3647
rect 393 3633 407 3647
rect 93 3613 107 3627
rect 53 3553 67 3567
rect 12 3533 26 3547
rect 33 3534 47 3548
rect 13 3493 27 3507
rect 53 3493 67 3507
rect 33 3293 47 3307
rect 333 3533 347 3547
rect 93 3393 107 3407
rect 133 3393 147 3407
rect 193 3393 207 3407
rect 73 3353 87 3367
rect 53 3233 67 3247
rect 93 3333 107 3347
rect 133 3294 147 3308
rect 373 3473 387 3487
rect 613 3993 627 4007
rect 593 3933 607 3947
rect 553 3833 567 3847
rect 593 3833 607 3847
rect 533 3814 547 3828
rect 473 3772 487 3786
rect 453 3693 467 3707
rect 433 3633 447 3647
rect 413 3533 427 3547
rect 493 3732 507 3746
rect 473 3673 487 3687
rect 453 3513 467 3527
rect 413 3493 427 3507
rect 433 3473 447 3487
rect 473 3473 487 3487
rect 413 3433 427 3447
rect 473 3433 487 3447
rect 393 3393 407 3407
rect 433 3393 447 3407
rect 333 3373 347 3387
rect 573 3773 587 3787
rect 953 4973 967 4987
rect 1013 5113 1027 5127
rect 1293 5153 1307 5167
rect 1213 5133 1227 5147
rect 1053 5032 1067 5046
rect 1013 4933 1027 4947
rect 973 4913 987 4927
rect 993 4893 1007 4907
rect 1133 5073 1147 5087
rect 1173 5074 1187 5088
rect 1233 5113 1247 5127
rect 1213 5073 1227 5087
rect 1333 5073 1347 5087
rect 1133 5032 1147 5046
rect 1193 5032 1207 5046
rect 1233 5032 1247 5046
rect 1313 5032 1327 5046
rect 1313 4993 1327 5007
rect 1073 4893 1087 4907
rect 1113 4893 1127 4907
rect 1173 4893 1187 4907
rect 1053 4873 1067 4887
rect 953 4854 967 4868
rect 1093 4853 1107 4867
rect 1133 4854 1147 4868
rect 1393 5332 1407 5346
rect 1593 5473 1607 5487
rect 1593 5413 1607 5427
rect 1653 5693 1667 5707
rect 1653 5594 1667 5608
rect 1693 5594 1707 5608
rect 1753 5833 1767 5847
rect 1753 5713 1767 5727
rect 1753 5653 1767 5667
rect 1733 5533 1747 5547
rect 1853 5773 1867 5787
rect 1833 5653 1847 5667
rect 1833 5613 1847 5627
rect 1813 5594 1827 5608
rect 1853 5593 1867 5607
rect 1793 5552 1807 5566
rect 2453 6233 2467 6247
rect 3853 6233 3867 6247
rect 2413 6193 2427 6207
rect 2193 6173 2207 6187
rect 2153 6153 2167 6167
rect 1953 6114 1967 6128
rect 1993 6113 2007 6127
rect 2093 6133 2107 6147
rect 1972 6073 1986 6087
rect 1993 6072 2007 6086
rect 2073 6072 2087 6086
rect 1933 6033 1947 6047
rect 1893 6013 1907 6027
rect 1933 5993 1947 6007
rect 2033 6053 2047 6067
rect 2133 6033 2147 6047
rect 2033 5953 2047 5967
rect 2013 5933 2027 5947
rect 1933 5913 1947 5927
rect 1893 5893 1907 5907
rect 1993 5913 2007 5927
rect 2053 5894 2067 5908
rect 2093 5894 2107 5908
rect 2313 6133 2327 6147
rect 2233 6114 2247 6128
rect 2273 6114 2287 6128
rect 2353 6114 2367 6128
rect 2273 6073 2287 6087
rect 2753 6193 2767 6207
rect 3093 6193 3107 6207
rect 3353 6193 3367 6207
rect 3433 6193 3447 6207
rect 3553 6193 3567 6207
rect 2573 6133 2587 6147
rect 2453 6114 2467 6128
rect 2493 6114 2507 6128
rect 2533 6114 2547 6128
rect 2793 6173 2807 6187
rect 2833 6153 2847 6167
rect 2813 6133 2827 6147
rect 2833 6114 2847 6128
rect 2873 6114 2887 6128
rect 2913 6114 2927 6128
rect 2973 6114 2987 6128
rect 2473 6072 2487 6086
rect 2533 6073 2547 6087
rect 2593 6072 2607 6086
rect 2673 6073 2687 6087
rect 2733 6072 2747 6086
rect 2373 6033 2387 6047
rect 2413 6033 2427 6047
rect 2633 6033 2647 6047
rect 2333 6013 2347 6027
rect 2213 5973 2227 5987
rect 2673 5973 2687 5987
rect 2733 5973 2747 5987
rect 2693 5953 2707 5967
rect 2153 5933 2167 5947
rect 2673 5933 2687 5947
rect 2233 5913 2247 5927
rect 2273 5913 2287 5927
rect 2393 5913 2407 5927
rect 2513 5913 2527 5927
rect 1913 5852 1927 5866
rect 2193 5893 2207 5907
rect 2253 5893 2267 5907
rect 2333 5894 2347 5908
rect 2373 5894 2387 5908
rect 2553 5894 2567 5908
rect 2113 5852 2127 5866
rect 2593 5893 2607 5907
rect 2633 5894 2647 5908
rect 2693 5894 2707 5908
rect 2273 5852 2287 5866
rect 2333 5853 2347 5867
rect 2393 5852 2407 5866
rect 2493 5852 2507 5866
rect 1993 5793 2007 5807
rect 2053 5793 2067 5807
rect 2233 5793 2247 5807
rect 2253 5773 2267 5787
rect 2233 5693 2247 5707
rect 1953 5673 1967 5687
rect 2093 5673 2107 5687
rect 2073 5633 2087 5647
rect 1893 5613 1907 5627
rect 1753 5513 1767 5527
rect 1673 5493 1687 5507
rect 1833 5493 1847 5507
rect 1793 5453 1807 5467
rect 1673 5413 1687 5427
rect 1753 5413 1767 5427
rect 1553 5393 1567 5407
rect 1493 5313 1507 5327
rect 1433 5293 1447 5307
rect 1373 5233 1387 5247
rect 1453 5233 1467 5247
rect 1433 5153 1447 5167
rect 1393 5074 1407 5088
rect 1593 5374 1607 5388
rect 1573 5332 1587 5346
rect 1613 5332 1627 5346
rect 1713 5374 1727 5388
rect 1693 5333 1707 5347
rect 1673 5313 1687 5327
rect 1533 5293 1547 5307
rect 1533 5193 1547 5207
rect 1513 5153 1527 5167
rect 1453 5133 1467 5147
rect 1493 5074 1507 5088
rect 1533 5074 1547 5088
rect 1373 5013 1387 5027
rect 1453 5032 1467 5046
rect 1413 5013 1427 5027
rect 1553 5032 1567 5046
rect 1593 5032 1607 5046
rect 1493 4993 1507 5007
rect 1373 4973 1387 4987
rect 1293 4854 1307 4868
rect 1353 4854 1367 4868
rect 1413 4913 1427 4927
rect 1493 4893 1507 4907
rect 1413 4873 1427 4887
rect 1473 4853 1487 4867
rect 1133 4793 1147 4807
rect 1093 4673 1107 4687
rect 933 4613 947 4627
rect 973 4593 987 4607
rect 1093 4574 1107 4588
rect 1393 4812 1407 4826
rect 1273 4793 1287 4807
rect 1173 4713 1187 4727
rect 1153 4693 1167 4707
rect 1273 4653 1287 4667
rect 1353 4613 1367 4627
rect 1173 4593 1187 4607
rect 1153 4573 1167 4587
rect 1033 4553 1047 4567
rect 1093 4553 1107 4567
rect 1133 4553 1147 4567
rect 893 4473 907 4487
rect 873 4453 887 4467
rect 993 4512 1007 4526
rect 1013 4493 1027 4507
rect 773 4433 787 4447
rect 952 4433 966 4447
rect 973 4433 987 4447
rect 1013 4433 1027 4447
rect 753 4233 767 4247
rect 713 4133 727 4147
rect 813 4413 827 4427
rect 893 4393 907 4407
rect 853 4334 867 4348
rect 953 4334 967 4348
rect 993 4333 1007 4347
rect 833 4292 847 4306
rect 893 4293 907 4307
rect 933 4292 947 4306
rect 993 4292 1007 4306
rect 933 4233 947 4247
rect 833 4153 847 4167
rect 713 4093 727 4107
rect 673 4073 687 4087
rect 673 4033 687 4047
rect 773 4072 787 4086
rect 673 3993 687 4007
rect 653 3973 667 3987
rect 613 3813 627 3827
rect 693 3973 707 3987
rect 733 3973 747 3987
rect 853 3953 867 3967
rect 733 3933 747 3947
rect 813 3933 827 3947
rect 713 3913 727 3927
rect 953 4133 967 4147
rect 973 4073 987 4087
rect 953 4033 967 4047
rect 1113 4512 1127 4526
rect 1213 4554 1227 4568
rect 1193 4512 1207 4526
rect 1073 4453 1087 4467
rect 1033 4373 1047 4387
rect 1093 4373 1107 4387
rect 1053 4334 1067 4348
rect 1073 4292 1087 4306
rect 1153 4453 1167 4467
rect 1313 4554 1327 4568
rect 1353 4554 1367 4568
rect 1473 4812 1487 4826
rect 1553 4854 1567 4868
rect 1593 4854 1607 4868
rect 1793 5313 1807 5327
rect 1873 5453 1887 5467
rect 1853 5433 1867 5447
rect 1913 5594 1927 5608
rect 2033 5552 2047 5566
rect 1953 5533 1967 5547
rect 1913 5493 1927 5507
rect 1952 5493 1966 5507
rect 1973 5493 1987 5507
rect 1913 5453 1927 5467
rect 1893 5433 1907 5447
rect 1853 5373 1867 5387
rect 1933 5374 1947 5388
rect 1993 5473 2007 5487
rect 1973 5453 1987 5467
rect 1973 5374 1987 5388
rect 1913 5332 1927 5346
rect 1893 5313 1907 5327
rect 1793 5273 1807 5287
rect 1833 5273 1847 5287
rect 1873 5273 1887 5287
rect 1733 5233 1747 5247
rect 1773 5233 1787 5247
rect 1672 5213 1686 5227
rect 1693 5213 1707 5227
rect 1693 5133 1707 5147
rect 1753 5113 1767 5127
rect 1673 5073 1687 5087
rect 1713 5074 1727 5088
rect 1693 5032 1707 5046
rect 1953 5253 1967 5267
rect 1953 5213 1967 5227
rect 1813 5074 1827 5088
rect 1853 5074 1867 5088
rect 1893 5074 1907 5088
rect 1933 5073 1947 5087
rect 1753 5013 1767 5027
rect 1793 5013 1807 5027
rect 1713 4993 1727 5007
rect 1733 4973 1747 4987
rect 1653 4893 1667 4907
rect 1693 4873 1707 4887
rect 1633 4853 1647 4867
rect 1573 4812 1587 4826
rect 1533 4793 1547 4807
rect 1613 4793 1627 4807
rect 1673 4812 1687 4826
rect 1433 4753 1447 4767
rect 1633 4753 1647 4767
rect 1413 4693 1427 4707
rect 1493 4653 1507 4667
rect 1412 4573 1426 4587
rect 1433 4574 1447 4588
rect 1293 4493 1307 4507
rect 1193 4393 1207 4407
rect 1233 4393 1247 4407
rect 1233 4334 1247 4348
rect 1153 4293 1167 4307
rect 1133 4253 1147 4267
rect 1293 4292 1307 4306
rect 1293 4253 1307 4267
rect 1453 4533 1467 4547
rect 1593 4613 1607 4627
rect 1593 4554 1607 4568
rect 1593 4533 1607 4547
rect 1333 4512 1347 4526
rect 1413 4513 1427 4527
rect 1373 4493 1387 4507
rect 1393 4373 1407 4387
rect 1333 4334 1347 4348
rect 1373 4292 1387 4306
rect 1333 4253 1347 4267
rect 1313 4213 1327 4227
rect 1493 4473 1507 4487
rect 1473 4453 1487 4467
rect 1453 4413 1467 4427
rect 1433 4393 1447 4407
rect 1413 4334 1427 4348
rect 1393 4253 1407 4267
rect 1213 4193 1227 4207
rect 1373 4193 1387 4207
rect 1173 4173 1187 4187
rect 1093 4093 1107 4107
rect 1153 4093 1167 4107
rect 953 3993 967 4007
rect 933 3973 947 3987
rect 973 3973 987 3987
rect 1013 3973 1027 3987
rect 833 3893 847 3907
rect 913 3893 927 3907
rect 953 3893 967 3907
rect 713 3873 727 3887
rect 813 3873 827 3887
rect 693 3833 707 3847
rect 853 3853 867 3867
rect 953 3853 967 3867
rect 633 3772 647 3786
rect 593 3753 607 3767
rect 673 3753 687 3767
rect 633 3733 647 3747
rect 593 3713 607 3727
rect 593 3673 607 3687
rect 613 3633 627 3647
rect 593 3593 607 3607
rect 553 3573 567 3587
rect 533 3514 547 3528
rect 573 3514 587 3528
rect 553 3472 567 3486
rect 593 3472 607 3486
rect 653 3693 667 3707
rect 673 3673 687 3687
rect 653 3613 667 3627
rect 773 3814 787 3828
rect 753 3772 767 3786
rect 753 3733 767 3747
rect 753 3712 767 3726
rect 793 3713 807 3727
rect 713 3653 727 3667
rect 753 3633 767 3647
rect 853 3813 867 3827
rect 893 3814 907 3828
rect 933 3814 947 3828
rect 853 3733 867 3747
rect 833 3713 847 3727
rect 713 3573 727 3587
rect 793 3573 807 3587
rect 693 3533 707 3547
rect 653 3513 667 3527
rect 733 3514 747 3528
rect 513 3393 527 3407
rect 593 3393 607 3407
rect 493 3333 507 3347
rect 473 3293 487 3307
rect 193 3273 207 3287
rect 312 3273 326 3287
rect 93 3233 107 3247
rect 233 3233 247 3247
rect 173 3213 187 3227
rect 333 3272 347 3286
rect 593 3294 607 3308
rect 473 3213 487 3227
rect 553 3233 567 3247
rect 493 3173 507 3187
rect 533 3173 547 3187
rect 253 3113 267 3127
rect 333 3113 347 3127
rect 493 3113 507 3127
rect 73 3053 87 3067
rect 193 3053 207 3067
rect 33 2994 47 3008
rect 33 2893 47 2907
rect 93 2994 107 3008
rect 113 2952 127 2966
rect 153 2952 167 2966
rect 53 2833 67 2847
rect 53 2793 67 2807
rect 13 2774 27 2788
rect 33 2053 47 2067
rect 73 2732 87 2746
rect 133 2653 147 2667
rect 113 2474 127 2488
rect 213 2873 227 2887
rect 393 2974 407 2988
rect 293 2873 307 2887
rect 493 2873 507 2887
rect 253 2793 267 2807
rect 213 2713 227 2727
rect 273 2633 287 2647
rect 193 2593 207 2607
rect 273 2573 287 2587
rect 233 2493 247 2507
rect 153 2413 167 2427
rect 113 2053 127 2067
rect 133 1993 147 2007
rect 53 1953 67 1967
rect 93 1954 107 1968
rect 53 1913 67 1927
rect 33 1873 47 1887
rect 33 1753 47 1767
rect 93 1813 107 1827
rect 73 1753 87 1767
rect 193 2353 207 2367
rect 253 2253 267 2267
rect 473 2833 487 2847
rect 433 2793 447 2807
rect 353 2774 367 2788
rect 393 2774 407 2788
rect 333 2673 347 2687
rect 333 2613 347 2627
rect 413 2733 427 2747
rect 373 2573 387 2587
rect 293 2493 307 2507
rect 593 2833 607 2847
rect 533 2813 547 2827
rect 513 2793 527 2807
rect 513 2693 527 2707
rect 653 3433 667 3447
rect 633 3353 647 3367
rect 733 3433 747 3447
rect 713 3353 727 3367
rect 693 3294 707 3308
rect 773 3473 787 3487
rect 753 3313 767 3327
rect 913 3772 927 3786
rect 953 3772 967 3786
rect 933 3733 947 3747
rect 913 3693 927 3707
rect 873 3633 887 3647
rect 913 3613 927 3627
rect 853 3593 867 3607
rect 853 3553 867 3567
rect 853 3532 867 3546
rect 893 3514 907 3528
rect 953 3653 967 3667
rect 993 3953 1007 3967
rect 1133 4034 1147 4048
rect 1193 4113 1207 4127
rect 1353 4113 1367 4127
rect 1253 4073 1267 4087
rect 1153 3992 1167 4006
rect 1192 3993 1206 4007
rect 1233 4032 1247 4046
rect 1293 4034 1307 4048
rect 1333 4034 1347 4048
rect 1213 3992 1227 4006
rect 1113 3953 1127 3967
rect 1093 3933 1107 3947
rect 1053 3873 1067 3887
rect 1033 3853 1047 3867
rect 1013 3833 1027 3847
rect 993 3813 1007 3827
rect 1053 3814 1067 3828
rect 1093 3813 1107 3827
rect 993 3773 1007 3787
rect 993 3673 1007 3687
rect 1093 3773 1107 3787
rect 1033 3713 1047 3727
rect 1013 3633 1027 3647
rect 1153 3933 1167 3947
rect 1193 3933 1207 3947
rect 1133 3873 1147 3887
rect 1193 3853 1207 3867
rect 1273 3992 1287 4006
rect 1793 4953 1807 4967
rect 1773 4933 1787 4947
rect 1793 4893 1807 4907
rect 1773 4873 1787 4887
rect 1833 5032 1847 5046
rect 1953 5032 1967 5046
rect 1873 4873 1887 4887
rect 1853 4854 1867 4868
rect 1773 4812 1787 4826
rect 1793 4793 1807 4807
rect 1833 4773 1847 4787
rect 2033 5433 2047 5447
rect 2013 5393 2027 5407
rect 2093 5594 2107 5608
rect 2213 5552 2227 5566
rect 2453 5833 2467 5847
rect 2533 5833 2547 5847
rect 2333 5813 2347 5827
rect 2333 5633 2347 5647
rect 2313 5613 2327 5627
rect 2353 5594 2367 5608
rect 2413 5594 2427 5608
rect 2513 5713 2527 5727
rect 2553 5633 2567 5647
rect 2273 5573 2287 5587
rect 2373 5552 2387 5566
rect 2413 5553 2427 5567
rect 2473 5552 2487 5566
rect 2513 5552 2527 5566
rect 2253 5493 2267 5507
rect 2173 5413 2187 5427
rect 2093 5393 2107 5407
rect 2193 5374 2207 5388
rect 1993 5293 2007 5307
rect 2173 5332 2187 5346
rect 2213 5332 2227 5346
rect 2072 5273 2086 5287
rect 2093 5273 2107 5287
rect 2033 5253 2047 5267
rect 1993 5153 2007 5167
rect 2053 5193 2067 5207
rect 2033 5093 2047 5107
rect 2113 5253 2127 5267
rect 2093 5233 2107 5247
rect 2193 5293 2207 5307
rect 2172 5193 2186 5207
rect 2193 5193 2207 5207
rect 2113 5173 2127 5187
rect 2153 5153 2167 5167
rect 2093 5113 2107 5127
rect 2153 5113 2167 5127
rect 2073 5072 2087 5086
rect 2033 5032 2047 5046
rect 2033 4993 2047 5007
rect 1973 4973 1987 4987
rect 2193 5074 2207 5088
rect 2233 5074 2247 5088
rect 2093 5033 2107 5047
rect 2072 4933 2086 4947
rect 2093 4933 2107 4947
rect 1993 4854 2007 4868
rect 2033 4854 2047 4868
rect 2113 4873 2127 4887
rect 2173 5032 2187 5046
rect 2213 5033 2227 5047
rect 2193 4933 2207 4947
rect 1853 4753 1867 4767
rect 1793 4713 1807 4727
rect 1773 4693 1787 4707
rect 1753 4673 1767 4687
rect 1793 4673 1807 4687
rect 1793 4633 1807 4647
rect 1753 4533 1767 4547
rect 1633 4433 1647 4447
rect 1693 4433 1707 4447
rect 1733 4433 1747 4447
rect 1552 4413 1566 4427
rect 1573 4413 1587 4427
rect 1493 4353 1507 4367
rect 1533 4353 1547 4367
rect 1453 4173 1467 4187
rect 1493 4173 1507 4187
rect 1373 4073 1387 4087
rect 1433 4073 1447 4087
rect 1413 4034 1427 4048
rect 1433 3992 1447 4006
rect 1273 3913 1287 3927
rect 1373 3913 1387 3927
rect 1153 3773 1167 3787
rect 1133 3753 1147 3767
rect 1113 3733 1127 3747
rect 1213 3713 1227 3727
rect 1133 3653 1147 3667
rect 1173 3633 1187 3647
rect 973 3573 987 3587
rect 1053 3533 1067 3547
rect 953 3514 967 3528
rect 1013 3514 1027 3528
rect 1093 3593 1107 3607
rect 813 3473 827 3487
rect 793 3453 807 3467
rect 833 3433 847 3447
rect 873 3433 887 3447
rect 913 3433 927 3447
rect 1073 3513 1087 3527
rect 1193 3533 1207 3547
rect 993 3472 1007 3486
rect 1093 3473 1107 3487
rect 1073 3453 1087 3467
rect 1033 3433 1047 3447
rect 833 3373 847 3387
rect 932 3373 946 3387
rect 953 3373 967 3387
rect 773 3293 787 3307
rect 833 3293 847 3307
rect 793 3273 807 3287
rect 933 3272 947 3286
rect 653 3193 667 3207
rect 833 3253 847 3267
rect 753 3233 767 3247
rect 673 3093 687 3107
rect 713 3093 727 3107
rect 793 3233 807 3247
rect 773 3213 787 3227
rect 773 3133 787 3147
rect 933 3173 947 3187
rect 893 3133 907 3147
rect 833 3113 847 3127
rect 873 3073 887 3087
rect 853 3053 867 3067
rect 673 2994 687 3008
rect 753 2993 767 3007
rect 693 2952 707 2966
rect 653 2893 667 2907
rect 613 2813 627 2827
rect 653 2813 667 2827
rect 753 2813 767 2827
rect 533 2673 547 2687
rect 453 2633 467 2647
rect 433 2613 447 2627
rect 313 2474 327 2488
rect 353 2474 367 2488
rect 393 2474 407 2488
rect 513 2493 527 2507
rect 453 2473 467 2487
rect 473 2452 487 2466
rect 373 2413 387 2427
rect 453 2433 467 2447
rect 413 2313 427 2327
rect 813 2994 827 3008
rect 873 3013 887 3027
rect 913 3113 927 3127
rect 953 3153 967 3167
rect 933 3033 947 3047
rect 913 3013 927 3027
rect 833 2952 847 2966
rect 872 2953 886 2967
rect 893 2953 907 2967
rect 793 2933 807 2947
rect 893 2853 907 2867
rect 833 2833 847 2847
rect 873 2833 887 2847
rect 793 2813 807 2827
rect 773 2773 787 2787
rect 653 2732 667 2746
rect 713 2732 727 2746
rect 933 2933 947 2947
rect 913 2813 927 2827
rect 812 2773 826 2787
rect 833 2773 847 2787
rect 913 2792 927 2806
rect 753 2613 767 2627
rect 873 2732 887 2746
rect 913 2732 927 2746
rect 873 2693 887 2707
rect 813 2553 827 2567
rect 713 2533 727 2547
rect 813 2493 827 2507
rect 873 2494 887 2508
rect 573 2413 587 2427
rect 753 2353 767 2367
rect 453 2293 467 2307
rect 513 2293 527 2307
rect 473 2253 487 2267
rect 413 2234 427 2248
rect 453 2233 467 2247
rect 753 2273 767 2287
rect 833 2452 847 2466
rect 1153 3472 1167 3486
rect 1113 3413 1127 3427
rect 1133 3373 1147 3387
rect 1113 3274 1127 3288
rect 1153 3353 1167 3367
rect 1373 3873 1387 3887
rect 1293 3813 1307 3827
rect 1333 3814 1347 3828
rect 1433 3853 1447 3867
rect 1413 3833 1427 3847
rect 1273 3633 1287 3647
rect 1253 3553 1267 3567
rect 1213 3513 1227 3527
rect 1333 3593 1347 3607
rect 1273 3533 1287 3547
rect 1293 3513 1307 3527
rect 1213 3473 1227 3487
rect 1193 3413 1207 3427
rect 1173 3333 1187 3347
rect 1153 3313 1167 3327
rect 1173 3274 1187 3288
rect 1153 3233 1167 3247
rect 1153 3173 1167 3187
rect 1133 3153 1147 3167
rect 1053 3013 1067 3027
rect 1033 2973 1047 2987
rect 1053 2853 1067 2867
rect 953 2793 967 2807
rect 1033 2793 1047 2807
rect 973 2774 987 2788
rect 953 2733 967 2747
rect 1013 2713 1027 2727
rect 953 2693 967 2707
rect 993 2693 1007 2707
rect 933 2673 947 2687
rect 1013 2633 1027 2647
rect 1173 2833 1187 2847
rect 1073 2793 1087 2807
rect 1133 2774 1147 2788
rect 1073 2732 1087 2746
rect 1113 2732 1127 2746
rect 1073 2613 1087 2627
rect 1053 2573 1067 2587
rect 1093 2573 1107 2587
rect 1033 2553 1047 2567
rect 1013 2493 1027 2507
rect 1073 2513 1087 2527
rect 853 2433 867 2447
rect 833 2413 847 2427
rect 813 2253 827 2267
rect 873 2373 887 2387
rect 853 2313 867 2327
rect 853 2253 867 2267
rect 313 2213 327 2227
rect 353 2212 367 2226
rect 273 2153 287 2167
rect 393 2153 407 2167
rect 333 2053 347 2067
rect 253 2013 267 2027
rect 313 2013 327 2027
rect 233 1993 247 2007
rect 213 1973 227 1987
rect 193 1954 207 1968
rect 273 1954 287 1968
rect 253 1912 267 1926
rect 373 1993 387 2007
rect 513 2232 527 2246
rect 653 2232 667 2246
rect 833 2233 847 2247
rect 813 2192 827 2206
rect 853 2192 867 2206
rect 753 2093 767 2107
rect 453 2053 467 2067
rect 453 2013 467 2027
rect 393 1953 407 1967
rect 433 1933 447 1947
rect 653 1973 667 1987
rect 393 1873 407 1887
rect 333 1833 347 1847
rect 373 1833 387 1847
rect 313 1813 327 1827
rect 133 1712 147 1726
rect 272 1712 286 1726
rect 293 1713 307 1727
rect 133 1453 147 1467
rect 273 1453 287 1467
rect 93 1412 107 1426
rect 73 1353 87 1367
rect 113 1353 127 1367
rect 33 1333 47 1347
rect 13 694 27 708
rect 13 493 27 507
rect 13 352 27 366
rect 73 1332 87 1346
rect 113 1213 127 1227
rect 93 1172 107 1186
rect 293 1413 307 1427
rect 333 1313 347 1327
rect 433 1833 447 1847
rect 493 1933 507 1947
rect 833 1933 847 1947
rect 413 1713 427 1727
rect 473 1692 487 1706
rect 433 1672 447 1686
rect 393 1412 407 1426
rect 413 1393 427 1407
rect 393 1373 407 1387
rect 213 1253 227 1267
rect 253 1253 267 1267
rect 313 1253 327 1267
rect 373 1253 387 1267
rect 253 1213 267 1227
rect 193 1172 207 1186
rect 273 1172 287 1186
rect 133 1113 147 1127
rect 233 1113 247 1127
rect 213 1073 227 1087
rect 113 914 127 928
rect 293 993 307 1007
rect 73 873 87 887
rect 133 872 147 886
rect 212 913 226 927
rect 233 914 247 928
rect 273 914 287 928
rect 213 873 227 887
rect 93 853 107 867
rect 153 853 167 867
rect 193 853 207 867
rect 73 793 87 807
rect 73 694 87 708
rect 253 853 267 867
rect 213 733 227 747
rect 253 733 267 747
rect 293 694 307 708
rect 153 652 167 666
rect 193 652 207 666
rect 53 433 67 447
rect 113 433 127 447
rect 33 174 47 188
rect 93 413 107 427
rect 253 493 267 507
rect 193 414 207 428
rect 213 393 227 407
rect 373 1214 387 1228
rect 773 1913 787 1927
rect 753 1853 767 1867
rect 553 1833 567 1847
rect 593 1833 607 1847
rect 673 1833 687 1847
rect 653 1813 667 1827
rect 633 1773 647 1787
rect 573 1692 587 1706
rect 633 1672 647 1686
rect 533 1653 547 1667
rect 513 1593 527 1607
rect 593 1553 607 1567
rect 553 1533 567 1547
rect 713 1793 727 1807
rect 753 1793 767 1807
rect 673 1733 687 1747
rect 853 1913 867 1927
rect 833 1893 847 1907
rect 773 1773 787 1787
rect 973 2432 987 2446
rect 1033 2413 1047 2427
rect 973 2313 987 2327
rect 1013 2313 1027 2327
rect 1013 2292 1027 2306
rect 1013 2253 1027 2267
rect 953 2212 967 2226
rect 993 2212 1007 2226
rect 993 2173 1007 2187
rect 993 2013 1007 2027
rect 1273 3472 1287 3486
rect 1313 3473 1327 3487
rect 1213 3333 1227 3347
rect 1213 3153 1227 3167
rect 1213 3093 1227 3107
rect 1393 3772 1407 3786
rect 1373 3753 1387 3767
rect 1373 3673 1387 3687
rect 1393 3653 1407 3667
rect 1353 3513 1367 3527
rect 1393 3514 1407 3528
rect 1473 4073 1487 4087
rect 1513 4113 1527 4127
rect 1573 4373 1587 4387
rect 1673 4393 1687 4407
rect 1633 4353 1647 4367
rect 1593 4334 1607 4348
rect 1673 4333 1687 4347
rect 1773 4493 1787 4507
rect 1813 4533 1827 4547
rect 1813 4473 1827 4487
rect 1833 4433 1847 4447
rect 1873 4593 1887 4607
rect 1873 4513 1887 4527
rect 2053 4812 2067 4826
rect 2113 4812 2127 4826
rect 2153 4812 2167 4826
rect 2033 4773 2047 4787
rect 2053 4753 2067 4767
rect 2173 4753 2187 4767
rect 2633 5613 2647 5627
rect 2693 5613 2707 5627
rect 2593 5594 2607 5608
rect 2613 5552 2627 5566
rect 2553 5493 2567 5507
rect 2513 5473 2527 5487
rect 2493 5433 2507 5447
rect 2273 5373 2287 5387
rect 2333 5374 2347 5388
rect 2373 5374 2387 5388
rect 2433 5374 2447 5388
rect 2573 5413 2587 5427
rect 2653 5413 2667 5427
rect 2273 5332 2287 5346
rect 2313 5332 2327 5346
rect 2353 5253 2367 5267
rect 2333 5113 2347 5127
rect 2373 5074 2387 5088
rect 2413 5333 2427 5347
rect 2473 5332 2487 5346
rect 2713 5594 2727 5608
rect 2813 6073 2827 6087
rect 2893 6072 2907 6086
rect 2933 6053 2947 6067
rect 2773 6033 2787 6047
rect 2833 6033 2847 6047
rect 2873 6033 2887 6047
rect 2913 6033 2927 6047
rect 2773 5973 2787 5987
rect 2753 5953 2767 5967
rect 2773 5933 2787 5947
rect 2773 5912 2787 5926
rect 2813 5894 2827 5908
rect 2793 5833 2807 5847
rect 2833 5833 2847 5847
rect 2953 6033 2967 6047
rect 3053 6114 3067 6128
rect 3033 6072 3047 6086
rect 3153 6153 3167 6167
rect 3313 6153 3327 6167
rect 3193 6114 3207 6128
rect 3233 6114 3247 6128
rect 3313 6114 3327 6128
rect 3393 6114 3407 6128
rect 3473 6114 3487 6128
rect 3133 6053 3147 6067
rect 3193 6053 3207 6067
rect 3093 6013 3107 6027
rect 3173 6013 3187 6027
rect 2973 5953 2987 5967
rect 3133 5953 3147 5967
rect 2933 5933 2947 5947
rect 3173 5933 3187 5947
rect 3133 5913 3147 5927
rect 2933 5894 2947 5908
rect 2993 5894 3007 5908
rect 3033 5894 3047 5908
rect 2913 5853 2927 5867
rect 2953 5852 2967 5866
rect 3033 5833 3047 5847
rect 3113 5833 3127 5847
rect 2873 5813 2887 5827
rect 2993 5813 3007 5827
rect 2913 5733 2927 5747
rect 2853 5693 2867 5707
rect 2813 5653 2827 5667
rect 2773 5594 2787 5608
rect 2733 5552 2747 5566
rect 2693 5533 2707 5547
rect 2713 5493 2727 5507
rect 2653 5374 2667 5388
rect 2713 5373 2727 5387
rect 2593 5332 2607 5346
rect 2633 5332 2647 5346
rect 2513 5313 2527 5327
rect 2573 5313 2587 5327
rect 2453 5273 2467 5287
rect 2473 5253 2487 5267
rect 2453 5233 2467 5247
rect 2433 5213 2447 5227
rect 2413 5113 2427 5127
rect 2573 5233 2587 5247
rect 2493 5213 2507 5227
rect 2473 5193 2487 5207
rect 2513 5193 2527 5207
rect 2493 5153 2507 5167
rect 2533 5173 2547 5187
rect 2393 5073 2407 5087
rect 2253 5053 2267 5067
rect 2313 5032 2327 5046
rect 2233 4873 2247 4887
rect 2213 4773 2227 4787
rect 2193 4733 2207 4747
rect 2113 4713 2127 4727
rect 1933 4693 1947 4707
rect 2093 4693 2107 4707
rect 1972 4554 1986 4568
rect 2013 4653 2027 4667
rect 2073 4653 2087 4667
rect 1993 4553 2007 4567
rect 1953 4512 1967 4526
rect 2073 4613 2087 4627
rect 2053 4593 2067 4607
rect 2113 4673 2127 4687
rect 2153 4673 2167 4687
rect 2173 4633 2187 4647
rect 2153 4613 2167 4627
rect 2133 4573 2147 4587
rect 2173 4573 2187 4587
rect 2193 4532 2207 4546
rect 1973 4493 1987 4507
rect 2073 4512 2087 4526
rect 1893 4473 1907 4487
rect 1993 4473 2007 4487
rect 1793 4413 1807 4427
rect 1853 4413 1867 4427
rect 1973 4413 1987 4427
rect 1733 4333 1747 4347
rect 1693 4313 1707 4327
rect 1573 4233 1587 4247
rect 1533 4073 1547 4087
rect 1513 4034 1527 4048
rect 1573 3973 1587 3987
rect 1553 3953 1567 3967
rect 1493 3853 1507 3867
rect 1473 3834 1487 3848
rect 1473 3813 1487 3827
rect 1573 3793 1587 3807
rect 1693 4273 1707 4287
rect 1673 4233 1687 4247
rect 1613 4133 1627 4147
rect 1633 4073 1647 4087
rect 1693 4193 1707 4207
rect 1813 4313 1827 4327
rect 1813 4273 1827 4287
rect 1693 4153 1707 4167
rect 1633 4034 1647 4048
rect 1673 4034 1687 4048
rect 1813 4073 1827 4087
rect 1733 4034 1747 4048
rect 1773 4034 1787 4048
rect 1873 4113 1887 4127
rect 1833 4053 1847 4067
rect 1693 3993 1707 4007
rect 1613 3953 1627 3967
rect 1453 3772 1467 3786
rect 1513 3772 1527 3786
rect 1433 3713 1447 3727
rect 1473 3753 1487 3767
rect 1453 3693 1467 3707
rect 1513 3752 1527 3766
rect 1553 3752 1567 3766
rect 1493 3733 1507 3747
rect 1433 3653 1447 3667
rect 1353 3473 1367 3487
rect 1333 3453 1347 3467
rect 1333 3413 1347 3427
rect 1313 3313 1327 3327
rect 1253 3293 1267 3307
rect 1393 3453 1407 3467
rect 1373 3393 1387 3407
rect 1313 3252 1327 3266
rect 1253 3153 1267 3167
rect 1233 3053 1247 3067
rect 1213 3013 1227 3027
rect 1213 2973 1227 2987
rect 1193 2774 1207 2788
rect 1233 2873 1247 2887
rect 1293 3233 1307 3247
rect 1293 3093 1307 3107
rect 1333 3233 1347 3247
rect 1373 3233 1387 3247
rect 1333 3173 1347 3187
rect 1313 3073 1327 3087
rect 1273 3013 1287 3027
rect 1313 3013 1327 3027
rect 1293 2933 1307 2947
rect 1253 2833 1267 2847
rect 1233 2793 1247 2807
rect 1173 2513 1187 2527
rect 1113 2473 1127 2487
rect 1153 2474 1167 2488
rect 1112 2433 1126 2447
rect 1093 2413 1107 2427
rect 1133 2432 1147 2446
rect 1113 2353 1127 2367
rect 1113 2313 1127 2327
rect 1073 2293 1087 2307
rect 1073 2254 1087 2268
rect 1113 2254 1127 2268
rect 1173 2273 1187 2287
rect 1053 2212 1067 2226
rect 1093 2212 1107 2226
rect 1033 2173 1047 2187
rect 1133 2153 1147 2167
rect 1073 2093 1087 2107
rect 1093 2033 1107 2047
rect 1153 2033 1167 2047
rect 1073 2013 1087 2027
rect 933 1993 947 2007
rect 1013 1993 1027 2007
rect 973 1973 987 1987
rect 1013 1954 1027 1968
rect 1053 1954 1067 1968
rect 993 1912 1007 1926
rect 953 1893 967 1907
rect 873 1813 887 1827
rect 773 1733 787 1747
rect 833 1734 847 1748
rect 693 1692 707 1706
rect 653 1653 667 1667
rect 713 1633 727 1647
rect 753 1633 767 1647
rect 653 1593 667 1607
rect 633 1473 647 1487
rect 653 1453 667 1467
rect 593 1433 607 1447
rect 513 1413 527 1427
rect 633 1413 647 1427
rect 493 1393 507 1407
rect 573 1392 587 1406
rect 613 1393 627 1407
rect 473 1293 487 1307
rect 553 1273 567 1287
rect 433 1253 447 1267
rect 413 1193 427 1207
rect 333 1173 347 1187
rect 473 1233 487 1247
rect 513 1214 527 1228
rect 553 1213 567 1227
rect 353 1153 367 1167
rect 333 1113 347 1127
rect 333 1073 347 1087
rect 353 1053 367 1067
rect 493 1172 507 1186
rect 412 1153 426 1167
rect 433 1153 447 1167
rect 533 1153 547 1167
rect 553 1172 567 1186
rect 393 993 407 1007
rect 393 914 407 928
rect 453 914 467 928
rect 513 914 527 928
rect 553 914 567 928
rect 633 1313 647 1327
rect 693 1273 707 1287
rect 613 1214 627 1228
rect 593 1173 607 1187
rect 653 1153 667 1167
rect 593 1113 607 1127
rect 633 1113 647 1127
rect 373 853 387 867
rect 433 853 447 867
rect 493 872 507 886
rect 453 833 467 847
rect 413 813 427 827
rect 353 793 367 807
rect 573 873 587 887
rect 533 853 547 867
rect 533 733 547 747
rect 573 733 587 747
rect 353 694 367 708
rect 413 694 427 708
rect 453 694 467 708
rect 493 694 507 708
rect 513 652 527 666
rect 613 914 627 928
rect 773 1553 787 1567
rect 813 1533 827 1547
rect 913 1693 927 1707
rect 953 1872 967 1886
rect 1053 1873 1067 1887
rect 973 1833 987 1847
rect 953 1733 967 1747
rect 1013 1734 1027 1748
rect 913 1653 927 1667
rect 893 1613 907 1627
rect 1033 1692 1047 1706
rect 1053 1653 1067 1667
rect 993 1533 1007 1547
rect 1013 1473 1027 1487
rect 973 1412 987 1426
rect 953 1373 967 1387
rect 893 1313 907 1327
rect 853 1293 867 1307
rect 773 1273 787 1287
rect 733 1253 747 1267
rect 793 1233 807 1247
rect 733 1214 747 1228
rect 1093 1953 1107 1967
rect 1273 2774 1287 2788
rect 1353 2972 1367 2986
rect 1473 3653 1487 3667
rect 1473 3632 1487 3646
rect 1453 3613 1467 3627
rect 1453 3553 1467 3567
rect 1573 3693 1587 3707
rect 1553 3673 1567 3687
rect 1493 3613 1507 3627
rect 1513 3514 1527 3528
rect 1553 3513 1567 3527
rect 1493 3472 1507 3486
rect 1553 3473 1567 3487
rect 1533 3453 1547 3467
rect 1473 3433 1487 3447
rect 1513 3433 1527 3447
rect 1533 3353 1547 3367
rect 1513 3293 1527 3307
rect 1593 3653 1607 3667
rect 1793 3992 1807 4006
rect 1853 3992 1867 4006
rect 1833 3953 1847 3967
rect 1693 3933 1707 3947
rect 1753 3893 1767 3907
rect 1993 4393 2007 4407
rect 2013 4373 2027 4387
rect 2033 4353 2047 4367
rect 2193 4493 2207 4507
rect 2173 4453 2187 4467
rect 2133 4433 2147 4447
rect 2133 4373 2147 4387
rect 2053 4333 2067 4347
rect 2033 4293 2047 4307
rect 2033 4272 2047 4286
rect 1993 4213 2007 4227
rect 1993 4113 2007 4127
rect 1973 4093 1987 4107
rect 1893 4053 1907 4067
rect 1873 3953 1887 3967
rect 1953 4034 1967 4048
rect 1993 4034 2007 4048
rect 1913 3993 1927 4007
rect 1872 3932 1886 3946
rect 1893 3933 1907 3947
rect 1933 3953 1947 3967
rect 1973 3953 1987 3967
rect 1892 3893 1906 3907
rect 1913 3893 1927 3907
rect 1973 3893 1987 3907
rect 1893 3833 1907 3847
rect 1873 3793 1887 3807
rect 1713 3773 1727 3787
rect 1853 3773 1867 3787
rect 1693 3673 1707 3687
rect 1613 3633 1627 3647
rect 1593 3573 1607 3587
rect 1633 3533 1647 3547
rect 1613 3453 1627 3467
rect 1993 3833 2007 3847
rect 1953 3794 1967 3808
rect 1973 3673 1987 3687
rect 1833 3653 1847 3667
rect 1913 3653 1927 3667
rect 1813 3613 1827 3627
rect 1793 3553 1807 3567
rect 1753 3533 1767 3547
rect 1713 3513 1727 3527
rect 1813 3513 1827 3527
rect 1693 3433 1707 3447
rect 1653 3413 1667 3427
rect 1493 3252 1507 3266
rect 1533 3252 1547 3266
rect 1453 3233 1467 3247
rect 1413 3113 1427 3127
rect 1453 3113 1467 3127
rect 1633 3294 1647 3308
rect 1773 3472 1787 3486
rect 1813 3433 1827 3447
rect 1573 3253 1587 3267
rect 1553 3093 1567 3107
rect 1653 3252 1667 3266
rect 1613 3233 1627 3247
rect 1753 3294 1767 3308
rect 1733 3252 1747 3266
rect 1773 3193 1787 3207
rect 1773 3113 1787 3127
rect 1593 3093 1607 3107
rect 1693 3093 1707 3107
rect 1733 3093 1747 3107
rect 1573 3073 1587 3087
rect 1693 3053 1707 3067
rect 1613 3033 1627 3047
rect 1593 2993 1607 3007
rect 1393 2933 1407 2947
rect 1453 2972 1467 2986
rect 1433 2913 1447 2927
rect 1433 2873 1447 2887
rect 1333 2813 1347 2827
rect 1433 2793 1447 2807
rect 1353 2773 1367 2787
rect 1413 2774 1427 2788
rect 1253 2693 1267 2707
rect 1293 2693 1307 2707
rect 1233 2633 1247 2647
rect 1233 2593 1247 2607
rect 1273 2533 1287 2547
rect 1233 2474 1247 2488
rect 1313 2473 1327 2487
rect 1253 2353 1267 2367
rect 1333 2313 1347 2327
rect 1273 2293 1287 2307
rect 1193 2254 1207 2268
rect 1233 2254 1247 2268
rect 1313 2253 1327 2267
rect 1213 2193 1227 2207
rect 1193 2093 1207 2107
rect 1433 2753 1447 2767
rect 1393 2673 1407 2687
rect 1373 2513 1387 2527
rect 1433 2573 1447 2587
rect 1673 2853 1687 2867
rect 1553 2833 1567 2847
rect 1473 2813 1487 2827
rect 1533 2773 1547 2787
rect 1473 2693 1487 2707
rect 1533 2733 1547 2747
rect 1533 2712 1547 2726
rect 1513 2653 1527 2667
rect 1493 2633 1507 2647
rect 1473 2573 1487 2587
rect 1453 2553 1467 2567
rect 1453 2513 1467 2527
rect 1393 2493 1407 2507
rect 1373 2473 1387 2487
rect 1413 2474 1427 2488
rect 1413 2413 1427 2427
rect 1453 2413 1467 2427
rect 1373 2373 1387 2387
rect 1413 2373 1427 2387
rect 1393 2333 1407 2347
rect 1353 2253 1367 2267
rect 1453 2293 1467 2307
rect 1453 2253 1467 2267
rect 1333 2193 1347 2207
rect 1413 2193 1427 2207
rect 1373 2173 1387 2187
rect 1313 2153 1327 2167
rect 1373 2152 1387 2166
rect 1253 2073 1267 2087
rect 1193 1953 1207 1967
rect 1153 1912 1167 1926
rect 1333 1953 1347 1967
rect 1433 2133 1447 2147
rect 1293 1912 1307 1926
rect 1333 1912 1347 1926
rect 1253 1833 1267 1847
rect 1213 1793 1227 1807
rect 1153 1773 1167 1787
rect 1113 1734 1127 1748
rect 1313 1793 1327 1807
rect 1233 1733 1247 1747
rect 1273 1734 1287 1748
rect 1413 1954 1427 1968
rect 1513 2613 1527 2627
rect 1653 2793 1667 2807
rect 1753 3033 1767 3047
rect 1733 3013 1747 3027
rect 1813 3133 1827 3147
rect 1953 3613 1967 3627
rect 1873 3573 1887 3587
rect 1853 3553 1867 3567
rect 1973 3534 1987 3548
rect 1893 3514 1907 3528
rect 1953 3513 1967 3527
rect 1933 3472 1947 3486
rect 1873 3433 1887 3447
rect 1853 3333 1867 3347
rect 1953 3273 1967 3287
rect 2073 4253 2087 4267
rect 2053 4213 2067 4227
rect 2093 4213 2107 4227
rect 2113 4073 2127 4087
rect 2073 4034 2087 4048
rect 2293 4812 2307 4826
rect 2293 4753 2307 4767
rect 2273 4733 2287 4747
rect 2353 4993 2367 5007
rect 2453 5074 2467 5088
rect 2573 5153 2587 5167
rect 2573 5093 2587 5107
rect 2453 4993 2467 5007
rect 2413 4913 2427 4927
rect 2373 4893 2387 4907
rect 2433 4853 2447 4867
rect 2353 4773 2367 4787
rect 2313 4673 2327 4687
rect 2513 5032 2527 5046
rect 2553 5033 2567 5047
rect 2713 5333 2727 5347
rect 2673 5293 2687 5307
rect 2653 5193 2667 5207
rect 2593 5073 2607 5087
rect 2473 4953 2487 4967
rect 2513 4933 2527 4947
rect 2533 4913 2547 4927
rect 2533 4873 2547 4887
rect 2513 4854 2527 4868
rect 2573 5032 2587 5046
rect 2493 4812 2507 4826
rect 2553 4793 2567 4807
rect 2513 4772 2527 4786
rect 2473 4633 2487 4647
rect 2453 4593 2467 4607
rect 2313 4534 2327 4548
rect 2213 4453 2227 4467
rect 2553 4673 2567 4687
rect 2573 4593 2587 4607
rect 2473 4533 2487 4547
rect 2193 4413 2207 4427
rect 2393 4413 2407 4427
rect 2093 3992 2107 4006
rect 2113 3973 2127 3987
rect 2033 3953 2047 3967
rect 2073 3814 2087 3828
rect 2133 3833 2147 3847
rect 2013 3773 2027 3787
rect 2013 3653 2027 3667
rect 2053 3772 2067 3786
rect 2093 3753 2107 3767
rect 2133 3713 2147 3727
rect 2053 3673 2067 3687
rect 2113 3613 2127 3627
rect 2092 3534 2106 3548
rect 2113 3533 2127 3547
rect 2073 3493 2087 3507
rect 2053 3472 2067 3486
rect 1993 3373 2007 3387
rect 2033 3373 2047 3387
rect 1893 3252 1907 3266
rect 1973 3253 1987 3267
rect 2053 3353 2067 3367
rect 1993 3233 2007 3247
rect 2033 3233 2047 3247
rect 1893 3133 1907 3147
rect 2133 3492 2147 3506
rect 2293 4353 2307 4367
rect 2253 4334 2267 4348
rect 2293 4313 2307 4327
rect 2193 4292 2207 4306
rect 2233 4292 2247 4306
rect 2193 4213 2207 4227
rect 2173 4093 2187 4107
rect 2273 4173 2287 4187
rect 2473 4413 2487 4427
rect 2513 4533 2527 4547
rect 2513 4512 2527 4526
rect 2493 4393 2507 4407
rect 2433 4373 2447 4387
rect 2473 4373 2487 4387
rect 2473 4334 2487 4348
rect 2513 4333 2527 4347
rect 2393 4292 2407 4306
rect 2413 4273 2427 4287
rect 2353 4213 2367 4227
rect 2233 4153 2247 4167
rect 2193 4033 2207 4047
rect 2233 4034 2247 4048
rect 2173 3993 2187 4007
rect 2213 3992 2227 4006
rect 2253 3993 2267 4007
rect 2173 3972 2187 3986
rect 2213 3933 2227 3947
rect 2373 4034 2387 4048
rect 2313 3973 2327 3987
rect 2633 5032 2647 5046
rect 2673 5032 2687 5046
rect 2713 4993 2727 5007
rect 2793 5533 2807 5547
rect 2753 5473 2767 5487
rect 2833 5453 2847 5467
rect 2973 5633 2987 5647
rect 2853 5393 2867 5407
rect 2773 5374 2787 5388
rect 2833 5374 2847 5388
rect 2773 5333 2787 5347
rect 2853 5332 2867 5346
rect 2793 5293 2807 5307
rect 2773 5233 2787 5247
rect 2893 5552 2907 5566
rect 2933 5552 2947 5566
rect 2973 5552 2987 5566
rect 3133 5793 3147 5807
rect 3033 5693 3047 5707
rect 3073 5673 3087 5687
rect 3113 5594 3127 5608
rect 3233 5953 3247 5967
rect 3293 5953 3307 5967
rect 3253 5933 3267 5947
rect 3453 6072 3467 6086
rect 3493 6072 3507 6086
rect 3393 6013 3407 6027
rect 3673 6153 3687 6167
rect 3613 6114 3627 6128
rect 3593 6013 3607 6027
rect 3413 5993 3427 6007
rect 3553 5993 3567 6007
rect 3493 5973 3507 5987
rect 3613 5973 3627 5987
rect 3393 5913 3407 5927
rect 3433 5894 3447 5908
rect 3353 5873 3367 5887
rect 3533 5913 3547 5927
rect 3512 5894 3526 5908
rect 3573 5894 3587 5908
rect 3653 5953 3667 5967
rect 3453 5852 3467 5866
rect 3492 5852 3506 5866
rect 3513 5853 3527 5867
rect 3173 5773 3187 5787
rect 3593 5852 3607 5866
rect 3413 5753 3427 5767
rect 3553 5753 3567 5767
rect 3173 5733 3187 5747
rect 3153 5713 3167 5727
rect 3173 5633 3187 5647
rect 3173 5594 3187 5608
rect 3273 5594 3287 5608
rect 3313 5594 3327 5608
rect 3353 5594 3367 5608
rect 3053 5552 3067 5566
rect 3112 5553 3126 5567
rect 3133 5553 3147 5567
rect 2993 5533 3007 5547
rect 3033 5533 3047 5547
rect 2933 5473 2947 5487
rect 2893 5393 2907 5407
rect 2873 5273 2887 5287
rect 2873 5233 2887 5247
rect 2793 5213 2807 5227
rect 2833 5213 2847 5227
rect 2813 5113 2827 5127
rect 2873 5173 2887 5187
rect 2833 5093 2847 5107
rect 2793 5032 2807 5046
rect 2833 5032 2847 5046
rect 2973 5433 2987 5447
rect 2953 5332 2967 5346
rect 3193 5552 3207 5566
rect 3153 5513 3167 5527
rect 3153 5473 3167 5487
rect 3093 5374 3107 5388
rect 2932 5293 2946 5307
rect 2953 5293 2967 5307
rect 2913 5273 2927 5287
rect 2893 5074 2907 5088
rect 2993 5273 3007 5287
rect 2933 5233 2947 5247
rect 2993 5133 3007 5147
rect 2973 5113 2987 5127
rect 2933 5074 2947 5088
rect 2993 5073 3007 5087
rect 2893 5032 2907 5046
rect 2873 5013 2887 5027
rect 2733 4953 2747 4967
rect 2673 4893 2687 4907
rect 2613 4853 2627 4867
rect 2633 4793 2647 4807
rect 2693 4812 2707 4826
rect 2653 4773 2667 4787
rect 2693 4773 2707 4787
rect 2633 4753 2647 4767
rect 2613 4733 2627 4747
rect 2693 4633 2707 4647
rect 2693 4573 2707 4587
rect 2613 4554 2627 4568
rect 2653 4554 2667 4568
rect 2593 4513 2607 4527
rect 2673 4512 2687 4526
rect 2673 4473 2687 4487
rect 2893 4893 2907 4907
rect 2753 4873 2767 4887
rect 2813 4854 2827 4868
rect 2793 4812 2807 4826
rect 2753 4753 2767 4767
rect 2833 4773 2847 4787
rect 2793 4733 2807 4747
rect 2953 5013 2967 5027
rect 3113 5313 3127 5327
rect 3073 5293 3087 5307
rect 3113 5233 3127 5247
rect 3053 5113 3067 5127
rect 3033 5073 3047 5087
rect 3233 5513 3247 5527
rect 3293 5553 3307 5567
rect 3333 5552 3347 5566
rect 3353 5513 3367 5527
rect 3252 5453 3266 5467
rect 3273 5453 3287 5467
rect 3253 5413 3267 5427
rect 3213 5393 3227 5407
rect 3173 5373 3187 5387
rect 3273 5374 3287 5388
rect 3333 5374 3347 5388
rect 3153 5313 3167 5327
rect 3253 5332 3267 5346
rect 3173 5293 3187 5307
rect 3153 5253 3167 5267
rect 3133 5133 3147 5147
rect 3013 4993 3027 5007
rect 3073 4953 3087 4967
rect 3033 4933 3047 4947
rect 2993 4893 3007 4907
rect 3053 4893 3067 4907
rect 3133 4893 3147 4907
rect 2913 4853 2927 4867
rect 2953 4854 2967 4868
rect 3033 4853 3047 4867
rect 2933 4813 2947 4827
rect 2973 4812 2987 4826
rect 2953 4793 2967 4807
rect 2913 4733 2927 4747
rect 2833 4713 2847 4727
rect 2813 4673 2827 4687
rect 2833 4653 2847 4667
rect 2813 4613 2827 4627
rect 2793 4593 2807 4607
rect 2753 4513 2767 4527
rect 2813 4512 2827 4526
rect 2853 4512 2867 4526
rect 2733 4473 2747 4487
rect 2793 4473 2807 4487
rect 2893 4473 2907 4487
rect 2693 4453 2707 4467
rect 2753 4433 2767 4447
rect 2613 4413 2627 4427
rect 2652 4413 2666 4427
rect 2673 4413 2687 4427
rect 2733 4413 2747 4427
rect 2573 4353 2587 4367
rect 2593 4334 2607 4348
rect 2673 4333 2687 4347
rect 2773 4413 2787 4427
rect 2753 4393 2767 4407
rect 2813 4453 2827 4467
rect 2813 4393 2827 4407
rect 2813 4313 2827 4327
rect 2533 4273 2547 4287
rect 2573 4273 2587 4287
rect 2613 4253 2627 4267
rect 2493 4213 2507 4227
rect 2613 4213 2627 4227
rect 2433 4193 2447 4207
rect 2453 4133 2467 4147
rect 2673 4292 2687 4306
rect 2713 4292 2727 4306
rect 2653 4273 2667 4287
rect 2753 4253 2767 4267
rect 2653 4213 2667 4227
rect 2633 4193 2647 4207
rect 2653 4073 2667 4087
rect 2493 4034 2507 4048
rect 2573 4033 2587 4047
rect 2613 4033 2627 4047
rect 2733 4193 2747 4207
rect 2693 4153 2707 4167
rect 2673 4033 2687 4047
rect 2553 4012 2567 4026
rect 2273 3953 2287 3967
rect 2353 3953 2367 3967
rect 2333 3933 2347 3947
rect 2313 3873 2327 3887
rect 2293 3853 2307 3867
rect 2253 3814 2267 3828
rect 2193 3772 2207 3786
rect 2233 3753 2247 3767
rect 2173 3733 2187 3747
rect 2273 3693 2287 3707
rect 2373 3873 2387 3887
rect 2393 3853 2407 3867
rect 2353 3814 2367 3828
rect 2473 3992 2487 4006
rect 2593 3992 2607 4006
rect 2633 3992 2647 4006
rect 2793 4233 2807 4247
rect 2753 4093 2767 4107
rect 2733 4073 2747 4087
rect 2893 4353 2907 4367
rect 2833 4273 2847 4287
rect 2813 4133 2827 4147
rect 2793 4073 2807 4087
rect 3093 4854 3107 4868
rect 3073 4812 3087 4826
rect 2973 4773 2987 4787
rect 2953 4753 2967 4767
rect 3053 4733 3067 4747
rect 3033 4713 3047 4727
rect 2953 4693 2967 4707
rect 2993 4693 3007 4707
rect 2993 4653 3007 4667
rect 3013 4633 3027 4647
rect 3033 4613 3047 4627
rect 3013 4554 3027 4568
rect 2953 4493 2967 4507
rect 2933 4233 2947 4247
rect 3033 4513 3047 4527
rect 2973 4473 2987 4487
rect 2993 4433 3007 4447
rect 2973 4413 2987 4427
rect 2993 4393 3007 4407
rect 3013 4273 3027 4287
rect 2993 4233 3007 4247
rect 2853 4073 2867 4087
rect 2833 4053 2847 4067
rect 2513 3933 2527 3947
rect 2573 3853 2587 3867
rect 2453 3813 2467 3827
rect 2513 3814 2527 3828
rect 2413 3772 2427 3786
rect 2313 3693 2327 3707
rect 2453 3772 2467 3786
rect 2553 3773 2567 3787
rect 2453 3673 2467 3687
rect 2372 3653 2386 3667
rect 2393 3653 2407 3667
rect 2433 3653 2447 3667
rect 2253 3613 2267 3627
rect 2293 3613 2307 3627
rect 2233 3533 2247 3547
rect 2233 3493 2247 3507
rect 2333 3393 2347 3407
rect 2153 3333 2167 3347
rect 2293 3333 2307 3347
rect 2113 3233 2127 3247
rect 2253 3233 2267 3247
rect 2293 3233 2307 3247
rect 2233 3173 2247 3187
rect 2073 3113 2087 3127
rect 2113 3113 2127 3127
rect 1833 3053 1847 3067
rect 1813 3033 1827 3047
rect 1793 3013 1807 3027
rect 1693 2813 1707 2827
rect 1693 2792 1707 2806
rect 1673 2713 1687 2727
rect 1693 2693 1707 2707
rect 1733 2973 1747 2987
rect 1793 2973 1807 2987
rect 1833 2953 1847 2967
rect 1833 2853 1847 2867
rect 1793 2833 1807 2847
rect 1773 2793 1787 2807
rect 1833 2793 1847 2807
rect 1733 2773 1747 2787
rect 1873 2973 1887 2987
rect 1973 2974 1987 2988
rect 2033 2873 2047 2887
rect 1993 2813 2007 2827
rect 1832 2772 1846 2786
rect 1853 2773 1867 2787
rect 1933 2793 1947 2807
rect 1973 2773 1987 2787
rect 1793 2732 1807 2746
rect 1813 2693 1827 2707
rect 1753 2653 1767 2667
rect 1653 2593 1667 2607
rect 1713 2593 1727 2607
rect 1813 2573 1827 2587
rect 1613 2553 1627 2567
rect 1553 2513 1567 2527
rect 1533 2474 1547 2488
rect 1573 2474 1587 2488
rect 1513 2413 1527 2427
rect 1553 2413 1567 2427
rect 1493 2393 1507 2407
rect 1533 2333 1547 2347
rect 1513 2313 1527 2327
rect 1553 2313 1567 2327
rect 1653 2474 1667 2488
rect 1713 2473 1727 2487
rect 1773 2474 1787 2488
rect 1853 2732 1867 2746
rect 1913 2693 1927 2707
rect 1853 2673 1867 2687
rect 1913 2653 1927 2667
rect 1973 2633 1987 2647
rect 1973 2573 1987 2587
rect 1873 2533 1887 2547
rect 1853 2513 1867 2527
rect 1833 2474 1847 2488
rect 1673 2432 1687 2446
rect 1713 2432 1727 2446
rect 1753 2432 1767 2446
rect 1793 2432 1807 2446
rect 1933 2474 1947 2488
rect 2093 2853 2107 2867
rect 2033 2633 2047 2647
rect 2013 2553 2027 2567
rect 1993 2473 2007 2487
rect 1873 2433 1887 2447
rect 1912 2393 1926 2407
rect 1933 2393 1947 2407
rect 1693 2353 1707 2367
rect 1733 2353 1747 2367
rect 1853 2353 1867 2367
rect 1673 2273 1687 2287
rect 1573 2253 1587 2267
rect 1613 2254 1627 2268
rect 1473 2093 1487 2107
rect 1453 2053 1467 2067
rect 1573 2173 1587 2187
rect 1633 2133 1647 2147
rect 1793 2333 1807 2347
rect 1693 2193 1707 2207
rect 1733 2133 1747 2147
rect 1673 2113 1687 2127
rect 1593 2053 1607 2067
rect 1693 2053 1707 2067
rect 1573 2013 1587 2027
rect 1533 1993 1547 2007
rect 1453 1953 1467 1967
rect 1573 1953 1587 1967
rect 1393 1873 1407 1887
rect 1453 1873 1467 1887
rect 1513 1873 1527 1887
rect 1473 1833 1487 1847
rect 1433 1813 1447 1827
rect 1353 1793 1367 1807
rect 1353 1772 1367 1786
rect 1333 1733 1347 1747
rect 1093 1692 1107 1706
rect 1133 1692 1147 1706
rect 1173 1692 1187 1706
rect 1213 1692 1227 1706
rect 1253 1692 1267 1706
rect 1333 1693 1347 1707
rect 1293 1653 1307 1667
rect 1093 1633 1107 1647
rect 1073 1573 1087 1587
rect 1133 1373 1147 1387
rect 1213 1313 1227 1327
rect 1053 1293 1067 1307
rect 1033 1273 1047 1287
rect 1133 1273 1147 1287
rect 993 1233 1007 1247
rect 933 1214 947 1228
rect 753 1173 767 1187
rect 713 1153 727 1167
rect 673 1133 687 1147
rect 733 1113 747 1127
rect 693 914 707 928
rect 853 1173 867 1187
rect 953 1172 967 1186
rect 1132 1233 1146 1247
rect 1073 1214 1087 1228
rect 1053 1172 1067 1186
rect 773 1133 787 1147
rect 913 1033 927 1047
rect 873 933 887 947
rect 773 914 787 928
rect 833 914 847 928
rect 613 853 627 867
rect 713 872 727 886
rect 753 873 767 887
rect 733 813 747 827
rect 693 694 707 708
rect 393 613 407 627
rect 453 613 467 627
rect 633 652 647 666
rect 593 633 607 647
rect 573 432 587 446
rect 313 413 327 427
rect 433 413 447 427
rect 113 352 127 366
rect 153 353 167 367
rect 193 352 207 366
rect 233 213 247 227
rect 393 352 407 366
rect 353 313 367 327
rect 93 174 107 188
rect 253 174 267 188
rect 293 174 307 188
rect 373 174 387 188
rect 453 393 467 407
rect 513 394 527 408
rect 853 853 867 867
rect 813 833 827 847
rect 793 773 807 787
rect 773 693 787 707
rect 813 694 827 708
rect 973 914 987 928
rect 1013 914 1027 928
rect 933 873 947 887
rect 933 813 947 827
rect 993 853 1007 867
rect 1193 1153 1207 1167
rect 1093 1113 1107 1127
rect 1073 993 1087 1007
rect 1213 914 1227 928
rect 1073 853 1087 867
rect 1053 833 1067 847
rect 993 813 1007 827
rect 953 773 967 787
rect 1173 833 1187 847
rect 1153 793 1167 807
rect 953 733 967 747
rect 993 733 1007 747
rect 873 693 887 707
rect 913 693 927 707
rect 1033 694 1047 708
rect 1093 694 1107 708
rect 1133 694 1147 708
rect 1193 773 1207 787
rect 793 633 807 647
rect 733 613 747 627
rect 673 573 687 587
rect 673 453 687 467
rect 853 453 867 467
rect 593 393 607 407
rect 633 394 647 408
rect 453 352 467 366
rect 493 352 507 366
rect 493 213 507 227
rect 433 174 447 188
rect 493 174 507 188
rect 573 352 587 366
rect 413 133 427 147
rect 473 132 487 146
rect 533 133 547 147
rect 613 352 627 366
rect 733 393 747 407
rect 773 393 787 407
rect 793 352 807 366
rect 733 313 747 327
rect 1173 693 1187 707
rect 1493 1813 1507 1827
rect 1513 1753 1527 1767
rect 1653 1954 1667 1968
rect 1873 2313 1887 2327
rect 1833 2293 1847 2307
rect 1993 2433 2007 2447
rect 1993 2373 2007 2387
rect 1953 2333 1967 2347
rect 2033 2513 2047 2527
rect 2093 2712 2107 2726
rect 2173 3033 2187 3047
rect 2133 2973 2147 2987
rect 2153 2933 2167 2947
rect 2213 2953 2227 2967
rect 2373 3252 2387 3266
rect 2413 3613 2427 3627
rect 2453 3593 2467 3607
rect 2413 3553 2427 3567
rect 2413 3453 2427 3467
rect 2533 3693 2547 3707
rect 2453 3413 2467 3427
rect 2493 3413 2507 3427
rect 2433 3373 2447 3387
rect 2453 3333 2467 3347
rect 2433 3294 2447 3308
rect 2413 3253 2427 3267
rect 2393 3173 2407 3187
rect 2333 3113 2347 3127
rect 2273 3033 2287 3047
rect 2413 3033 2427 3047
rect 2253 3013 2267 3027
rect 2293 2973 2307 2987
rect 2513 3294 2527 3308
rect 2473 3233 2487 3247
rect 2553 3293 2567 3307
rect 2533 3173 2547 3187
rect 2453 3073 2467 3087
rect 2433 2993 2447 3007
rect 2273 2953 2287 2967
rect 2173 2853 2187 2867
rect 2153 2813 2167 2827
rect 2153 2774 2167 2788
rect 2253 2773 2267 2787
rect 2133 2733 2147 2747
rect 2113 2693 2127 2707
rect 2073 2613 2087 2627
rect 2093 2593 2107 2607
rect 2153 2653 2167 2667
rect 2133 2553 2147 2567
rect 2053 2493 2067 2507
rect 2033 2473 2047 2487
rect 2213 2712 2227 2726
rect 2313 2933 2327 2947
rect 2293 2893 2307 2907
rect 2553 2873 2567 2887
rect 2553 2813 2567 2827
rect 2513 2793 2527 2807
rect 2353 2753 2367 2767
rect 2373 2733 2387 2747
rect 2273 2673 2287 2687
rect 2173 2633 2187 2647
rect 2653 3973 2667 3987
rect 2613 3913 2627 3927
rect 2693 3952 2707 3966
rect 2613 3892 2627 3906
rect 2653 3893 2667 3907
rect 2653 3814 2667 3828
rect 2693 3814 2707 3828
rect 2593 3773 2607 3787
rect 2633 3753 2647 3767
rect 2593 3633 2607 3647
rect 2693 3733 2707 3747
rect 2673 3533 2687 3547
rect 2653 3514 2667 3528
rect 2813 4034 2827 4048
rect 2752 3953 2766 3967
rect 2773 3953 2787 3967
rect 2733 3893 2747 3907
rect 2833 3993 2847 4007
rect 2793 3893 2807 3907
rect 2773 3873 2787 3887
rect 2733 3853 2747 3867
rect 2773 3833 2787 3847
rect 2753 3814 2767 3828
rect 2793 3814 2807 3828
rect 2893 4093 2907 4107
rect 2953 4213 2967 4227
rect 2933 4034 2947 4048
rect 2973 4034 2987 4048
rect 2913 3992 2927 4006
rect 2853 3953 2867 3967
rect 2873 3933 2887 3947
rect 2833 3813 2847 3827
rect 2873 3793 2887 3807
rect 2913 3953 2927 3967
rect 2733 3773 2747 3787
rect 2773 3772 2787 3786
rect 2793 3753 2807 3767
rect 2793 3713 2807 3727
rect 2873 3753 2887 3767
rect 2853 3693 2867 3707
rect 2733 3673 2747 3687
rect 2813 3673 2827 3687
rect 2733 3613 2747 3627
rect 2893 3673 2907 3687
rect 3133 4753 3147 4767
rect 3213 5313 3227 5327
rect 3193 5273 3207 5287
rect 3173 5173 3187 5187
rect 3213 5173 3227 5187
rect 3193 5133 3207 5147
rect 3313 5233 3327 5247
rect 3193 5074 3207 5088
rect 3233 5074 3247 5088
rect 3293 5072 3307 5086
rect 3333 5213 3347 5227
rect 3433 5673 3447 5687
rect 3553 5653 3567 5667
rect 3633 5813 3647 5827
rect 3653 5773 3667 5787
rect 3633 5713 3647 5727
rect 3493 5594 3507 5608
rect 3513 5552 3527 5566
rect 3593 5594 3607 5608
rect 3653 5653 3667 5667
rect 3633 5593 3647 5607
rect 3633 5553 3647 5567
rect 3773 6133 3787 6147
rect 3813 6133 3827 6147
rect 3713 6114 3727 6128
rect 3893 6114 3907 6128
rect 3933 6113 3947 6127
rect 3833 6072 3847 6086
rect 3913 6073 3927 6087
rect 3893 6053 3907 6067
rect 3853 5973 3867 5987
rect 3773 5953 3787 5967
rect 3733 5894 3747 5908
rect 3813 5893 3827 5907
rect 4113 6153 4127 6167
rect 4153 6153 4167 6167
rect 4313 6153 4327 6167
rect 4013 6114 4027 6128
rect 4213 6113 4227 6127
rect 4253 6114 4267 6128
rect 3953 6073 3967 6087
rect 3993 6072 4007 6086
rect 4033 6072 4047 6086
rect 4133 6072 4147 6086
rect 4173 6072 4187 6086
rect 4213 6072 4227 6086
rect 3973 6033 3987 6047
rect 3913 5993 3927 6007
rect 3693 5813 3707 5827
rect 3773 5833 3787 5847
rect 3773 5753 3787 5767
rect 3913 5852 3927 5866
rect 3873 5833 3887 5847
rect 3913 5813 3927 5827
rect 3893 5773 3907 5787
rect 3773 5713 3787 5727
rect 3813 5713 3827 5727
rect 3753 5673 3767 5687
rect 3752 5652 3766 5666
rect 3773 5653 3787 5667
rect 3673 5633 3687 5647
rect 3773 5632 3787 5646
rect 3813 5633 3827 5647
rect 3873 5633 3887 5647
rect 3753 5613 3767 5627
rect 3693 5594 3707 5608
rect 3733 5594 3747 5608
rect 3673 5553 3687 5567
rect 3653 5533 3667 5547
rect 3433 5513 3447 5527
rect 3473 5513 3487 5527
rect 3393 5433 3407 5447
rect 3493 5453 3507 5467
rect 3473 5413 3487 5427
rect 3353 5173 3367 5187
rect 3333 5113 3347 5127
rect 3433 5313 3447 5327
rect 3393 5253 3407 5267
rect 3473 5273 3487 5287
rect 3453 5253 3467 5267
rect 3433 5233 3447 5247
rect 3473 5232 3487 5246
rect 3433 5173 3447 5187
rect 3453 5153 3467 5167
rect 3393 5133 3407 5147
rect 3433 5133 3447 5147
rect 3373 5112 3387 5126
rect 3393 5093 3407 5107
rect 3493 5193 3507 5207
rect 3753 5553 3767 5567
rect 3713 5533 3727 5547
rect 3693 5513 3707 5527
rect 3753 5493 3767 5507
rect 3672 5453 3686 5467
rect 3693 5453 3707 5467
rect 3533 5413 3547 5427
rect 3733 5413 3747 5427
rect 3573 5394 3587 5408
rect 3613 5393 3627 5407
rect 3573 5373 3587 5387
rect 3673 5374 3687 5388
rect 3593 5332 3607 5346
rect 3653 5332 3667 5346
rect 3593 5273 3607 5287
rect 3533 5233 3547 5247
rect 3513 5173 3527 5187
rect 3553 5173 3567 5187
rect 3533 5153 3547 5167
rect 3473 5113 3487 5127
rect 3193 5013 3207 5027
rect 3173 4854 3187 4868
rect 3153 4733 3167 4747
rect 3293 5033 3307 5047
rect 3313 5013 3327 5027
rect 3213 4933 3227 4947
rect 3253 4854 3267 4868
rect 3193 4833 3207 4847
rect 3373 5033 3387 5047
rect 3493 5074 3507 5088
rect 3373 4973 3387 4987
rect 3353 4953 3367 4967
rect 3333 4913 3347 4927
rect 3433 5013 3447 5027
rect 3473 4993 3487 5007
rect 3473 4972 3487 4986
rect 3413 4893 3427 4907
rect 3373 4854 3387 4868
rect 3413 4854 3427 4868
rect 3233 4773 3247 4787
rect 3313 4813 3327 4827
rect 3533 4933 3547 4947
rect 3513 4913 3527 4927
rect 3593 5133 3607 5147
rect 3653 5273 3667 5287
rect 3653 5233 3667 5247
rect 3613 5113 3627 5127
rect 3633 5093 3647 5107
rect 3753 5332 3767 5346
rect 3753 5293 3767 5307
rect 3833 5613 3847 5627
rect 3933 5753 3947 5767
rect 3913 5733 3927 5747
rect 3893 5593 3907 5607
rect 3793 5513 3807 5527
rect 3853 5552 3867 5566
rect 3933 5693 3947 5707
rect 4073 5993 4087 6007
rect 4033 5933 4047 5947
rect 4033 5894 4047 5908
rect 4193 5933 4207 5947
rect 4113 5894 4127 5908
rect 4153 5894 4167 5908
rect 4313 6073 4327 6087
rect 4313 6033 4327 6047
rect 4273 5973 4287 5987
rect 4273 5933 4287 5947
rect 4333 5933 4347 5947
rect 4213 5913 4227 5927
rect 4253 5913 4267 5927
rect 3973 5833 3987 5847
rect 4013 5713 4027 5727
rect 3953 5673 3967 5687
rect 3933 5653 3947 5667
rect 4013 5653 4027 5667
rect 3933 5594 3947 5608
rect 3973 5594 3987 5608
rect 4073 5673 4087 5687
rect 3893 5513 3907 5527
rect 3813 5433 3827 5447
rect 3913 5393 3927 5407
rect 4053 5593 4067 5607
rect 3993 5493 4007 5507
rect 4013 5453 4027 5467
rect 4053 5453 4067 5467
rect 4013 5413 4027 5427
rect 3973 5393 3987 5407
rect 3853 5374 3867 5388
rect 3893 5373 3907 5387
rect 3693 5253 3707 5267
rect 3713 5233 3727 5247
rect 3733 5213 3747 5227
rect 3793 5213 3807 5227
rect 3713 5193 3727 5207
rect 3653 5073 3667 5087
rect 3673 5073 3687 5087
rect 3613 5032 3627 5046
rect 3673 4973 3687 4987
rect 3653 4953 3667 4967
rect 3733 5133 3747 5147
rect 3773 5113 3787 5127
rect 3793 5093 3807 5107
rect 3833 5332 3847 5346
rect 3833 5253 3847 5267
rect 3713 5033 3727 5047
rect 3753 4933 3767 4947
rect 3553 4854 3567 4868
rect 3613 4854 3627 4868
rect 3653 4854 3667 4868
rect 3393 4812 3407 4826
rect 3473 4812 3487 4826
rect 3533 4812 3547 4826
rect 3433 4773 3447 4787
rect 3473 4753 3487 4767
rect 3313 4733 3327 4747
rect 3173 4713 3187 4727
rect 3273 4713 3287 4727
rect 3173 4653 3187 4667
rect 3133 4613 3147 4627
rect 3073 4573 3087 4587
rect 3093 4554 3107 4568
rect 3173 4554 3187 4568
rect 3233 4554 3247 4568
rect 3073 4513 3087 4527
rect 3193 4513 3207 4527
rect 3173 4493 3187 4507
rect 3113 4473 3127 4487
rect 3593 4813 3607 4827
rect 3593 4773 3607 4787
rect 3673 4812 3687 4826
rect 3673 4753 3687 4767
rect 3613 4733 3627 4747
rect 3573 4673 3587 4687
rect 3313 4613 3327 4627
rect 3353 4554 3367 4568
rect 3213 4493 3227 4507
rect 3273 4493 3287 4507
rect 3473 4653 3487 4667
rect 3513 4653 3527 4667
rect 3433 4633 3447 4647
rect 3473 4613 3487 4627
rect 3453 4593 3467 4607
rect 3373 4493 3387 4507
rect 3413 4493 3427 4507
rect 3333 4473 3347 4487
rect 3193 4433 3207 4447
rect 3233 4433 3247 4447
rect 3193 4353 3207 4367
rect 3133 4334 3147 4348
rect 3173 4333 3187 4347
rect 3053 4233 3067 4247
rect 3133 4272 3147 4286
rect 3073 4213 3087 4227
rect 3113 4213 3127 4227
rect 3053 4073 3067 4087
rect 3033 4053 3047 4067
rect 2993 3993 3007 4007
rect 3013 3953 3027 3967
rect 3093 4153 3107 4167
rect 3093 4113 3107 4127
rect 3113 4013 3127 4027
rect 3093 3953 3107 3967
rect 2973 3933 2987 3947
rect 3093 3932 3107 3946
rect 3153 4193 3167 4207
rect 3153 3993 3167 4007
rect 3133 3913 3147 3927
rect 3113 3893 3127 3907
rect 3013 3753 3027 3767
rect 2993 3733 3007 3747
rect 3173 3973 3187 3987
rect 3273 4353 3287 4367
rect 3353 4353 3367 4367
rect 3353 4313 3367 4327
rect 3533 4512 3547 4526
rect 3593 4593 3607 4607
rect 3593 4473 3607 4487
rect 3493 4453 3507 4467
rect 3573 4453 3587 4467
rect 3633 4453 3647 4467
rect 3393 4353 3407 4367
rect 3213 4292 3227 4306
rect 3293 4292 3307 4306
rect 3333 4272 3347 4286
rect 3313 4233 3327 4247
rect 3253 4213 3267 4227
rect 3313 4193 3327 4207
rect 3493 4312 3507 4326
rect 3493 4273 3507 4287
rect 3653 4433 3667 4447
rect 3713 4613 3727 4627
rect 3773 4854 3787 4868
rect 3813 5012 3827 5026
rect 3813 4854 3827 4868
rect 3813 4813 3827 4827
rect 3753 4753 3767 4767
rect 3913 5333 3927 5347
rect 3953 5332 3967 5346
rect 3993 5293 4007 5307
rect 3973 5273 3987 5287
rect 3893 5233 3907 5247
rect 3933 5193 3947 5207
rect 3893 5113 3907 5127
rect 3953 5153 3967 5167
rect 3933 5073 3947 5087
rect 3853 5033 3867 5047
rect 3853 4973 3867 4987
rect 3973 5093 3987 5107
rect 4173 5852 4187 5866
rect 4253 5852 4267 5866
rect 4213 5813 4227 5827
rect 4113 5653 4127 5667
rect 4253 5653 4267 5667
rect 4213 5613 4227 5627
rect 4153 5594 4167 5608
rect 4193 5594 4207 5608
rect 4133 5552 4147 5566
rect 4153 5533 4167 5547
rect 4193 5513 4207 5527
rect 4153 5453 4167 5467
rect 4193 5453 4207 5467
rect 4173 5433 4187 5447
rect 4093 5413 4107 5427
rect 4073 5372 4087 5386
rect 4133 5374 4147 5388
rect 4073 5332 4087 5346
rect 4153 5332 4167 5346
rect 4193 5333 4207 5347
rect 4113 5273 4127 5287
rect 4133 5253 4147 5267
rect 4133 5213 4147 5227
rect 4173 5173 4187 5187
rect 4093 5113 4107 5127
rect 4073 5074 4087 5088
rect 4133 5074 4147 5088
rect 4293 5793 4307 5807
rect 4313 5773 4327 5787
rect 4293 5713 4307 5727
rect 4273 5613 4287 5627
rect 4253 5594 4267 5608
rect 4613 6193 4627 6207
rect 4553 6153 4567 6167
rect 4373 6072 4387 6086
rect 4513 6114 4527 6128
rect 4593 6114 4607 6128
rect 4533 6072 4547 6086
rect 4593 6073 4607 6087
rect 4493 6013 4507 6027
rect 4533 5973 4547 5987
rect 4393 5913 4407 5927
rect 4432 5913 4446 5927
rect 4453 5913 4467 5927
rect 4593 5913 4607 5927
rect 4653 6173 4667 6187
rect 5533 6173 5547 6187
rect 5633 6173 5647 6187
rect 5753 6173 5767 6187
rect 4753 6153 4767 6167
rect 4793 6153 4807 6167
rect 5013 6153 5027 6167
rect 5133 6153 5147 6167
rect 5193 6153 5207 6167
rect 5233 6153 5247 6167
rect 5273 6153 5287 6167
rect 4693 6114 4707 6128
rect 4673 6072 4687 6086
rect 4853 6114 4867 6128
rect 4913 6114 4927 6128
rect 4993 6114 5007 6128
rect 4813 6072 4827 6086
rect 4633 6033 4647 6047
rect 4713 6033 4727 6047
rect 4753 6033 4767 6047
rect 4853 5993 4867 6007
rect 4713 5973 4727 5987
rect 4813 5973 4827 5987
rect 4653 5933 4667 5947
rect 4773 5893 4787 5907
rect 4813 5894 4827 5908
rect 4953 6072 4967 6086
rect 4913 5913 4927 5927
rect 4653 5833 4667 5847
rect 4433 5813 4447 5827
rect 4733 5773 4747 5787
rect 4733 5713 4747 5727
rect 4393 5633 4407 5647
rect 4453 5633 4467 5647
rect 4693 5633 4707 5647
rect 4413 5594 4427 5608
rect 4372 5552 4386 5566
rect 4393 5553 4407 5567
rect 4333 5533 4347 5547
rect 4393 5513 4407 5527
rect 4373 5493 4387 5507
rect 4433 5493 4447 5507
rect 4273 5453 4287 5467
rect 4273 5374 4287 5388
rect 4313 5374 4327 5388
rect 4233 5313 4247 5327
rect 4333 5332 4347 5346
rect 4293 5313 4307 5327
rect 4513 5594 4527 5608
rect 4553 5594 4567 5608
rect 4633 5594 4647 5608
rect 4533 5552 4547 5566
rect 4473 5513 4487 5527
rect 4413 5393 4427 5407
rect 4453 5393 4467 5407
rect 4413 5313 4427 5327
rect 4253 5273 4267 5287
rect 4373 5273 4387 5287
rect 4213 5173 4227 5187
rect 4333 5253 4347 5267
rect 4253 5153 4267 5167
rect 4193 5133 4207 5147
rect 4293 5133 4307 5147
rect 4193 5112 4207 5126
rect 3973 5033 3987 5047
rect 3953 5013 3967 5027
rect 3993 5013 4007 5027
rect 4032 5013 4046 5027
rect 4053 5013 4067 5027
rect 3953 4973 3967 4987
rect 3913 4913 3927 4927
rect 3853 4893 3867 4907
rect 3833 4773 3847 4787
rect 3853 4713 3867 4727
rect 3793 4673 3807 4687
rect 3833 4673 3847 4687
rect 3753 4554 3767 4568
rect 3733 4512 3747 4526
rect 3713 4473 3727 4487
rect 3693 4393 3707 4407
rect 3653 4333 3667 4347
rect 3633 4213 3647 4227
rect 3893 4793 3907 4807
rect 3933 4753 3947 4767
rect 3893 4673 3907 4687
rect 3873 4553 3887 4567
rect 3973 4953 3987 4967
rect 4053 4913 4067 4927
rect 4173 5052 4187 5066
rect 4113 5032 4127 5046
rect 4113 4973 4127 4987
rect 4072 4893 4086 4907
rect 4093 4893 4107 4907
rect 4073 4872 4087 4886
rect 4013 4854 4027 4868
rect 3993 4793 4007 4807
rect 4053 4793 4067 4807
rect 4133 4913 4147 4927
rect 4113 4873 4127 4887
rect 4273 5093 4287 5107
rect 4213 5074 4227 5088
rect 4193 4973 4207 4987
rect 4173 4913 4187 4927
rect 4173 4892 4187 4906
rect 4153 4873 4167 4887
rect 4313 5093 4327 5107
rect 4313 5072 4327 5086
rect 4313 4953 4327 4967
rect 4413 5233 4427 5247
rect 4393 5153 4407 5167
rect 4373 5113 4387 5127
rect 4373 5074 4387 5088
rect 4433 5193 4447 5207
rect 4453 5053 4467 5067
rect 4393 5013 4407 5027
rect 4393 4973 4407 4987
rect 4333 4933 4347 4947
rect 4313 4873 4327 4887
rect 4393 4854 4407 4868
rect 4593 5493 4607 5507
rect 4493 5413 4507 5427
rect 4533 5374 4547 5388
rect 4513 5313 4527 5327
rect 4573 5333 4587 5347
rect 4553 5273 4567 5287
rect 4653 5552 4667 5566
rect 4653 5513 4667 5527
rect 4693 5513 4707 5527
rect 4633 5473 4647 5487
rect 4673 5473 4687 5487
rect 4613 5453 4627 5467
rect 4613 5373 4627 5387
rect 4693 5413 4707 5427
rect 4713 5373 4727 5387
rect 4613 5332 4627 5346
rect 4653 5332 4667 5346
rect 4993 5913 5007 5927
rect 5093 6114 5107 6128
rect 5253 6114 5267 6128
rect 5333 6113 5347 6127
rect 5393 6114 5407 6128
rect 5453 6114 5467 6128
rect 5493 6114 5507 6128
rect 5673 6153 5687 6167
rect 5673 6114 5687 6128
rect 5113 6072 5127 6086
rect 5193 6073 5207 6087
rect 5153 5973 5167 5987
rect 5033 5913 5047 5927
rect 5073 5913 5087 5927
rect 5153 5913 5167 5927
rect 5113 5894 5127 5908
rect 5273 6072 5287 6086
rect 5333 6072 5347 6086
rect 5253 5973 5267 5987
rect 5193 5913 5207 5927
rect 5232 5913 5246 5927
rect 5253 5913 5267 5927
rect 4873 5852 4887 5866
rect 4913 5852 4927 5866
rect 4973 5852 4987 5866
rect 5033 5853 5047 5867
rect 4833 5833 4847 5847
rect 4833 5733 4847 5747
rect 4773 5653 4787 5667
rect 4813 5633 4827 5647
rect 4813 5594 4827 5608
rect 4773 5552 4787 5566
rect 4793 5433 4807 5447
rect 5133 5852 5147 5866
rect 5173 5853 5187 5867
rect 4933 5653 4947 5667
rect 4873 5593 4887 5607
rect 5073 5613 5087 5627
rect 4973 5594 4987 5608
rect 5033 5594 5047 5608
rect 5353 5993 5367 6007
rect 5393 5993 5407 6007
rect 5513 6072 5527 6086
rect 5553 6072 5567 6086
rect 5613 6072 5627 6086
rect 5653 6072 5667 6086
rect 5453 6033 5467 6047
rect 5573 6033 5587 6047
rect 5553 5933 5567 5947
rect 5413 5913 5427 5927
rect 5433 5894 5447 5908
rect 5473 5893 5487 5907
rect 5513 5894 5527 5908
rect 5253 5773 5267 5787
rect 5233 5733 5247 5747
rect 5333 5852 5347 5866
rect 5373 5852 5387 5866
rect 5413 5852 5427 5866
rect 5473 5852 5487 5866
rect 5533 5852 5547 5866
rect 5573 5773 5587 5787
rect 5393 5753 5407 5767
rect 5273 5713 5287 5727
rect 5353 5713 5367 5727
rect 5193 5613 5207 5627
rect 4873 5552 4887 5566
rect 4913 5552 4927 5566
rect 4853 5513 4867 5527
rect 5113 5593 5127 5607
rect 5173 5594 5187 5608
rect 5133 5573 5147 5587
rect 4973 5493 4987 5507
rect 5053 5552 5067 5566
rect 5113 5552 5127 5566
rect 5113 5453 5127 5467
rect 4893 5433 4907 5447
rect 5013 5433 5027 5447
rect 4853 5393 4867 5407
rect 4653 5293 4667 5307
rect 4693 5293 4707 5307
rect 4613 5273 4627 5287
rect 4513 5213 4527 5227
rect 4513 5153 4527 5167
rect 4533 5113 4547 5127
rect 4573 5093 4587 5107
rect 4753 5332 4767 5346
rect 4733 5233 4747 5247
rect 4713 5213 4727 5227
rect 4633 5173 4647 5187
rect 4553 5032 4567 5046
rect 4613 5033 4627 5047
rect 4773 5273 4787 5287
rect 4753 5173 4767 5187
rect 4793 5173 4807 5187
rect 4733 5074 4747 5088
rect 4633 5013 4647 5027
rect 4513 4973 4527 4987
rect 4553 4973 4567 4987
rect 4553 4933 4567 4947
rect 4593 4933 4607 4947
rect 4513 4893 4527 4907
rect 3993 4753 4007 4767
rect 3973 4573 3987 4587
rect 3953 4553 3967 4567
rect 3873 4493 3887 4507
rect 3753 4433 3767 4447
rect 3733 4373 3747 4387
rect 3713 4313 3727 4327
rect 3813 4453 3827 4467
rect 3793 4393 3807 4407
rect 3913 4493 3927 4507
rect 3973 4493 3987 4507
rect 3893 4413 3907 4427
rect 3773 4333 3787 4347
rect 3753 4193 3767 4207
rect 3593 4173 3607 4187
rect 3693 4173 3707 4187
rect 3393 4153 3407 4167
rect 3433 4153 3447 4167
rect 3493 4153 3507 4167
rect 3333 4033 3347 4047
rect 3573 4093 3587 4107
rect 3553 4033 3567 4047
rect 3453 4012 3467 4026
rect 3533 4013 3547 4027
rect 3433 3973 3447 3987
rect 3433 3952 3447 3966
rect 3213 3913 3227 3927
rect 3293 3913 3307 3927
rect 3193 3833 3207 3847
rect 3193 3794 3207 3808
rect 3173 3753 3187 3767
rect 3153 3733 3167 3747
rect 2993 3653 3007 3667
rect 2913 3633 2927 3647
rect 2713 3573 2727 3587
rect 2793 3573 2807 3587
rect 2733 3553 2747 3567
rect 2813 3533 2827 3547
rect 2593 3413 2607 3427
rect 2653 3193 2667 3207
rect 2693 3493 2707 3507
rect 2793 3453 2807 3467
rect 2773 3433 2787 3447
rect 2753 3413 2767 3427
rect 2753 3353 2767 3367
rect 2793 3393 2807 3407
rect 2693 3333 2707 3347
rect 2773 3333 2787 3347
rect 2693 3293 2707 3307
rect 2753 3294 2767 3308
rect 2633 3153 2647 3167
rect 2673 3153 2687 3167
rect 2593 3133 2607 3147
rect 2593 2973 2607 2987
rect 2613 2873 2627 2887
rect 2613 2852 2627 2866
rect 2593 2833 2607 2847
rect 2573 2733 2587 2747
rect 2513 2633 2527 2647
rect 2313 2593 2327 2607
rect 2173 2533 2187 2547
rect 2213 2533 2227 2547
rect 2153 2473 2167 2487
rect 2273 2493 2287 2507
rect 2633 2593 2647 2607
rect 2593 2573 2607 2587
rect 2533 2533 2547 2547
rect 2373 2453 2387 2467
rect 2193 2432 2207 2446
rect 2213 2413 2227 2427
rect 2073 2393 2087 2407
rect 2013 2293 2027 2307
rect 1833 2212 1847 2226
rect 1993 2254 2007 2268
rect 2053 2253 2067 2267
rect 1953 2213 1967 2227
rect 1873 2153 1887 2167
rect 1813 2133 1827 2147
rect 1833 2053 1847 2067
rect 1873 2053 1887 2067
rect 1793 2033 1807 2047
rect 1633 1912 1647 1926
rect 1593 1813 1607 1827
rect 1413 1692 1427 1706
rect 1453 1653 1467 1667
rect 1513 1653 1527 1667
rect 1393 1533 1407 1547
rect 1253 1413 1267 1427
rect 1353 1493 1367 1507
rect 1593 1734 1607 1748
rect 1733 1912 1747 1926
rect 1673 1873 1687 1887
rect 1733 1833 1747 1847
rect 1653 1793 1667 1807
rect 1633 1733 1647 1747
rect 1553 1693 1567 1707
rect 1633 1693 1647 1707
rect 1573 1653 1587 1667
rect 1433 1493 1447 1507
rect 1533 1493 1547 1507
rect 1253 1313 1267 1327
rect 1553 1434 1567 1448
rect 1393 1333 1407 1347
rect 1313 1273 1327 1287
rect 1613 1493 1627 1507
rect 1573 1373 1587 1387
rect 1453 1333 1467 1347
rect 1373 1253 1387 1267
rect 1433 1253 1447 1267
rect 1313 1214 1327 1228
rect 1293 1153 1307 1167
rect 1393 1213 1407 1227
rect 1493 1313 1507 1327
rect 1493 1253 1507 1267
rect 1533 1213 1547 1227
rect 1773 1993 1787 2007
rect 1793 1973 1807 1987
rect 1813 1912 1827 1926
rect 1793 1893 1807 1907
rect 1753 1793 1767 1807
rect 1713 1734 1727 1748
rect 1673 1693 1687 1707
rect 1853 1873 1867 1887
rect 1993 2193 2007 2207
rect 1973 2173 1987 2187
rect 2013 2153 2027 2167
rect 1993 2133 2007 2147
rect 2033 2133 2047 2147
rect 1973 2093 1987 2107
rect 2033 2112 2047 2126
rect 2013 2073 2027 2087
rect 1913 2033 1927 2047
rect 1953 2033 1967 2047
rect 2013 2033 2027 2047
rect 1893 2013 1907 2027
rect 2113 2393 2127 2407
rect 2173 2353 2187 2367
rect 2133 2254 2147 2268
rect 2273 2432 2287 2446
rect 2333 2393 2347 2407
rect 2273 2353 2287 2367
rect 2233 2333 2247 2347
rect 2233 2293 2247 2307
rect 2173 2253 2187 2267
rect 2213 2253 2227 2267
rect 2353 2333 2367 2347
rect 2313 2254 2327 2268
rect 2093 2213 2107 2227
rect 2073 2053 2087 2067
rect 2053 2033 2067 2047
rect 2033 1993 2047 2007
rect 1913 1953 1927 1967
rect 1993 1954 2007 1968
rect 1893 1912 1907 1926
rect 1833 1773 1847 1787
rect 1873 1773 1887 1787
rect 1813 1753 1827 1767
rect 1873 1734 1887 1748
rect 2013 1913 2027 1927
rect 1973 1873 1987 1887
rect 1933 1833 1947 1847
rect 1933 1753 1947 1767
rect 1993 1753 2007 1767
rect 1653 1473 1667 1487
rect 1613 1434 1627 1448
rect 1733 1692 1747 1706
rect 1793 1692 1807 1706
rect 1693 1673 1707 1687
rect 1713 1533 1727 1547
rect 1613 1393 1627 1407
rect 1613 1253 1627 1267
rect 1653 1333 1667 1347
rect 1633 1213 1647 1227
rect 1393 1172 1407 1186
rect 1433 1172 1447 1186
rect 1373 1153 1387 1167
rect 1473 1153 1487 1167
rect 1333 1113 1347 1127
rect 1593 1172 1607 1186
rect 1533 1033 1547 1047
rect 1333 973 1347 987
rect 1393 973 1407 987
rect 1293 953 1307 967
rect 1253 914 1267 928
rect 1453 914 1467 928
rect 1573 914 1587 928
rect 1613 914 1627 928
rect 933 633 947 647
rect 1033 633 1047 647
rect 1153 652 1167 666
rect 1193 652 1207 666
rect 1113 613 1127 627
rect 973 593 987 607
rect 1013 593 1027 607
rect 1073 593 1087 607
rect 993 493 1007 507
rect 873 433 887 447
rect 913 394 927 408
rect 953 394 967 408
rect 893 333 907 347
rect 933 273 947 287
rect 853 253 867 267
rect 653 213 667 227
rect 713 213 727 227
rect 793 213 807 227
rect 733 174 747 188
rect 833 193 847 207
rect 1233 733 1247 747
rect 1293 733 1307 747
rect 1253 652 1267 666
rect 1293 653 1307 667
rect 1333 833 1347 847
rect 1393 872 1407 886
rect 1433 872 1447 886
rect 1533 873 1547 887
rect 1353 813 1367 827
rect 1453 773 1467 787
rect 1393 733 1407 747
rect 1353 694 1367 708
rect 1593 872 1607 886
rect 1553 833 1567 847
rect 1573 753 1587 767
rect 1533 733 1547 747
rect 1513 694 1527 708
rect 1313 493 1327 507
rect 1413 652 1427 666
rect 1453 652 1467 666
rect 1493 652 1507 666
rect 1413 513 1427 527
rect 1533 513 1547 527
rect 1353 453 1367 467
rect 1053 394 1067 408
rect 1093 394 1107 408
rect 1033 353 1047 367
rect 1013 333 1027 347
rect 1033 313 1047 327
rect 1113 353 1127 367
rect 1113 273 1127 287
rect 1073 253 1087 267
rect 1033 213 1047 227
rect 1093 213 1107 227
rect 873 174 887 188
rect 573 93 587 107
rect 713 132 727 146
rect 793 132 807 146
rect 753 93 767 107
rect 853 93 867 107
rect 993 93 1007 107
rect 1093 132 1107 146
rect 753 33 767 47
rect 1053 33 1067 47
rect 1173 394 1187 408
rect 1233 393 1247 407
rect 1493 433 1507 447
rect 1413 413 1427 427
rect 1193 352 1207 366
rect 1213 313 1227 327
rect 1173 174 1187 188
rect 1633 733 1647 747
rect 1593 693 1607 707
rect 1853 1692 1867 1706
rect 1853 1573 1867 1587
rect 1893 1573 1907 1587
rect 1773 1473 1787 1487
rect 1813 1473 1827 1487
rect 2153 2212 2167 2226
rect 2113 2173 2127 2187
rect 2193 2173 2207 2187
rect 2173 2133 2187 2147
rect 2173 2112 2187 2126
rect 2113 2093 2127 2107
rect 2213 2153 2227 2167
rect 2253 2133 2267 2147
rect 2193 2093 2207 2107
rect 2152 2053 2166 2067
rect 2173 2053 2187 2067
rect 2273 2053 2287 2067
rect 2093 1973 2107 1987
rect 2113 1954 2127 1968
rect 2172 2013 2186 2027
rect 2193 2013 2207 2027
rect 2173 1933 2187 1947
rect 2093 1912 2107 1926
rect 2173 1912 2187 1926
rect 2073 1893 2087 1907
rect 2053 1833 2067 1847
rect 2033 1733 2047 1747
rect 1933 1533 1947 1547
rect 1873 1473 1887 1487
rect 1853 1433 1867 1447
rect 1973 1692 1987 1706
rect 2053 1633 2067 1647
rect 2013 1613 2027 1627
rect 1993 1473 2007 1487
rect 1913 1453 1927 1467
rect 1953 1453 1967 1467
rect 1673 1253 1687 1267
rect 1713 1253 1727 1267
rect 1753 1253 1767 1267
rect 1713 1214 1727 1228
rect 1873 1392 1887 1406
rect 1833 1373 1847 1387
rect 1933 1392 1947 1406
rect 1893 1333 1907 1347
rect 2033 1453 2047 1467
rect 2013 1393 2027 1407
rect 2173 1833 2187 1847
rect 2233 1954 2247 1968
rect 2413 2513 2427 2527
rect 2513 2513 2527 2527
rect 2473 2474 2487 2488
rect 2453 2432 2467 2446
rect 2493 2373 2507 2387
rect 2453 2254 2467 2268
rect 2633 2513 2647 2527
rect 2632 2474 2646 2488
rect 2673 2972 2687 2986
rect 2733 3233 2747 3247
rect 2773 3193 2787 3207
rect 2893 3613 2907 3627
rect 2912 3573 2926 3587
rect 2933 3573 2947 3587
rect 2933 3533 2947 3547
rect 2953 3514 2967 3528
rect 2933 3472 2947 3486
rect 2853 3453 2867 3467
rect 2893 3453 2907 3467
rect 2853 3373 2867 3387
rect 2893 3353 2907 3367
rect 2933 3353 2947 3367
rect 2853 3333 2867 3347
rect 2893 3332 2907 3346
rect 2833 3293 2847 3307
rect 3033 3633 3047 3647
rect 3013 3593 3027 3607
rect 3253 3893 3267 3907
rect 3233 3833 3247 3847
rect 3233 3793 3247 3807
rect 3233 3753 3247 3767
rect 3253 3733 3267 3747
rect 3233 3653 3247 3667
rect 3173 3633 3187 3647
rect 3213 3633 3227 3647
rect 3173 3593 3187 3607
rect 3113 3514 3127 3528
rect 3233 3514 3247 3528
rect 3033 3393 3047 3407
rect 3013 3373 3027 3387
rect 3113 3453 3127 3467
rect 3173 3413 3187 3427
rect 3273 3693 3287 3707
rect 3353 3873 3367 3887
rect 3313 3814 3327 3828
rect 3293 3673 3307 3687
rect 3333 3772 3347 3786
rect 3313 3613 3327 3627
rect 3373 3814 3387 3828
rect 3353 3713 3367 3727
rect 3393 3653 3407 3667
rect 3373 3613 3387 3627
rect 3272 3573 3286 3587
rect 3313 3573 3327 3587
rect 3333 3573 3347 3587
rect 3293 3514 3307 3528
rect 3413 3613 3427 3627
rect 3393 3593 3407 3607
rect 3373 3534 3387 3548
rect 3413 3492 3427 3506
rect 3313 3472 3327 3486
rect 3393 3473 3407 3487
rect 3253 3433 3267 3447
rect 3313 3433 3327 3447
rect 3233 3393 3247 3407
rect 3053 3373 3067 3387
rect 3093 3373 3107 3387
rect 3073 3333 3087 3347
rect 2833 3233 2847 3247
rect 2813 3113 2827 3127
rect 2913 3193 2927 3207
rect 2892 3173 2906 3187
rect 2753 3093 2767 3107
rect 2833 3093 2847 3107
rect 2653 2473 2667 2487
rect 2733 3053 2747 3067
rect 2713 2933 2727 2947
rect 2753 3033 2767 3047
rect 3053 3273 3067 3287
rect 3013 3153 3027 3167
rect 3213 3272 3227 3286
rect 3333 3274 3347 3288
rect 3453 3933 3467 3947
rect 3453 3893 3467 3907
rect 3513 3853 3527 3867
rect 3633 4034 3647 4048
rect 3673 4034 3687 4048
rect 3773 4093 3787 4107
rect 3753 4053 3767 4067
rect 3833 4334 3847 4348
rect 3853 4253 3867 4267
rect 3853 4193 3867 4207
rect 3833 4153 3847 4167
rect 3813 4113 3827 4127
rect 3793 4073 3807 4087
rect 3853 4093 3867 4107
rect 3713 4034 3727 4048
rect 3853 4013 3867 4027
rect 3593 3993 3607 4007
rect 3573 3953 3587 3967
rect 3553 3933 3567 3947
rect 3613 3973 3627 3987
rect 3613 3952 3627 3966
rect 3713 3993 3727 4007
rect 3653 3933 3667 3947
rect 3613 3893 3627 3907
rect 3693 3893 3707 3907
rect 3773 3992 3787 4006
rect 3813 3993 3827 4007
rect 3773 3893 3787 3907
rect 3733 3873 3747 3887
rect 3473 3813 3487 3827
rect 3553 3814 3567 3828
rect 3533 3772 3547 3786
rect 3693 3853 3707 3867
rect 3633 3833 3647 3847
rect 3673 3814 3687 3828
rect 3973 4413 3987 4427
rect 3913 4333 3927 4347
rect 4053 4653 4067 4667
rect 4053 4593 4067 4607
rect 4033 4512 4047 4526
rect 4113 4793 4127 4807
rect 4153 4793 4167 4807
rect 4233 4793 4247 4807
rect 4133 4753 4147 4767
rect 4373 4812 4387 4826
rect 4433 4813 4447 4827
rect 4413 4753 4427 4767
rect 4253 4733 4267 4747
rect 4313 4733 4327 4747
rect 4193 4653 4207 4667
rect 4113 4633 4127 4647
rect 4153 4554 4167 4568
rect 4233 4554 4247 4568
rect 4353 4713 4367 4727
rect 4313 4693 4327 4707
rect 4273 4554 4287 4568
rect 3993 4393 4007 4407
rect 4053 4393 4067 4407
rect 4013 4334 4027 4348
rect 3913 4293 3927 4307
rect 3953 4292 3967 4306
rect 4053 4292 4067 4306
rect 3993 4253 4007 4267
rect 4173 4512 4187 4526
rect 4233 4513 4247 4527
rect 4193 4334 4207 4348
rect 4293 4453 4307 4467
rect 4333 4413 4347 4427
rect 4293 4353 4307 4367
rect 4253 4334 4267 4348
rect 4373 4673 4387 4687
rect 4553 4854 4567 4868
rect 4453 4713 4467 4727
rect 4433 4653 4447 4667
rect 4413 4633 4427 4647
rect 4533 4753 4547 4767
rect 4573 4633 4587 4647
rect 4513 4613 4527 4627
rect 4493 4593 4507 4607
rect 4453 4554 4467 4568
rect 4373 4513 4387 4527
rect 4433 4512 4447 4526
rect 4453 4473 4467 4487
rect 4353 4373 4367 4387
rect 4353 4352 4367 4366
rect 4413 4353 4427 4367
rect 4273 4292 4287 4306
rect 4333 4292 4347 4306
rect 4553 4554 4567 4568
rect 4753 5033 4767 5047
rect 4713 4993 4727 5007
rect 4693 4953 4707 4967
rect 4673 4893 4687 4907
rect 4613 4873 4627 4887
rect 4653 4854 4667 4868
rect 4733 4873 4747 4887
rect 4633 4812 4647 4826
rect 4713 4813 4727 4827
rect 4673 4773 4687 4787
rect 4633 4693 4647 4707
rect 4773 4993 4787 5007
rect 4853 5332 4867 5346
rect 5053 5393 5067 5407
rect 4993 5373 5007 5387
rect 4913 5333 4927 5347
rect 4913 5293 4927 5307
rect 4893 5273 4907 5287
rect 4973 5313 4987 5327
rect 4933 5233 4947 5247
rect 4953 5153 4967 5167
rect 4833 5133 4847 5147
rect 4813 5113 4827 5127
rect 4853 5074 4867 5088
rect 4893 5074 4907 5088
rect 4933 5074 4947 5088
rect 4813 4953 4827 4967
rect 4793 4873 4807 4887
rect 4753 4853 4767 4867
rect 4753 4813 4767 4827
rect 4733 4753 4747 4767
rect 4713 4613 4727 4627
rect 4633 4573 4647 4587
rect 4733 4573 4747 4587
rect 4613 4553 4627 4567
rect 4673 4554 4687 4568
rect 4793 4812 4807 4827
rect 4853 5013 4867 5027
rect 4933 5033 4947 5047
rect 4873 4993 4887 5007
rect 4893 4893 4907 4907
rect 4832 4853 4846 4867
rect 4853 4853 4867 4867
rect 4813 4773 4827 4787
rect 4753 4553 4767 4567
rect 4793 4553 4807 4567
rect 4633 4533 4647 4547
rect 4573 4512 4587 4526
rect 4613 4512 4627 4526
rect 4533 4433 4547 4447
rect 4513 4413 4527 4427
rect 4473 4393 4487 4407
rect 4453 4333 4467 4347
rect 4293 4273 4307 4287
rect 4353 4273 4367 4287
rect 4213 4253 4227 4267
rect 4153 4233 4167 4247
rect 4133 4213 4147 4227
rect 4073 4193 4087 4207
rect 3913 4153 3927 4167
rect 3973 4073 3987 4087
rect 3993 4033 4007 4047
rect 3973 4013 3987 4027
rect 3893 3973 3907 3987
rect 3833 3913 3847 3927
rect 3853 3873 3867 3887
rect 3873 3833 3887 3847
rect 3733 3793 3747 3807
rect 3653 3772 3667 3786
rect 3533 3733 3547 3747
rect 3613 3733 3627 3747
rect 3693 3733 3707 3747
rect 3553 3693 3567 3707
rect 3473 3633 3487 3647
rect 3873 3792 3887 3806
rect 3793 3772 3807 3786
rect 3793 3713 3807 3727
rect 3873 3713 3887 3727
rect 3793 3692 3807 3706
rect 3733 3653 3747 3667
rect 3773 3653 3787 3667
rect 3673 3633 3687 3647
rect 3553 3593 3567 3607
rect 3533 3573 3547 3587
rect 3533 3513 3547 3527
rect 3673 3513 3687 3527
rect 3513 3493 3527 3507
rect 3693 3493 3707 3507
rect 3773 3593 3787 3607
rect 3573 3393 3587 3407
rect 3533 3373 3547 3387
rect 3493 3313 3507 3327
rect 3373 3232 3387 3246
rect 3413 3232 3427 3246
rect 3313 3213 3327 3227
rect 2953 3113 2967 3127
rect 2813 2853 2827 2867
rect 2893 2972 2907 2986
rect 2873 2933 2887 2947
rect 2753 2813 2767 2827
rect 2853 2813 2867 2827
rect 2733 2774 2747 2788
rect 2773 2773 2787 2787
rect 2893 2913 2907 2927
rect 2913 2873 2927 2887
rect 2713 2732 2727 2746
rect 2733 2593 2747 2607
rect 2833 2732 2847 2746
rect 2813 2693 2827 2707
rect 2813 2653 2827 2667
rect 2773 2573 2787 2587
rect 2793 2474 2807 2488
rect 2553 2433 2567 2447
rect 2393 2212 2407 2226
rect 2433 2212 2447 2226
rect 2473 2212 2487 2226
rect 2413 2173 2427 2187
rect 2373 2153 2387 2167
rect 2353 2093 2367 2107
rect 2453 2193 2467 2207
rect 2453 2093 2467 2107
rect 2673 2433 2687 2447
rect 2773 2432 2787 2446
rect 2573 2393 2587 2407
rect 2613 2393 2627 2407
rect 2713 2393 2727 2407
rect 2632 2293 2646 2307
rect 2653 2293 2667 2307
rect 2593 2254 2607 2268
rect 2633 2253 2647 2267
rect 2513 2193 2527 2207
rect 2553 2193 2567 2207
rect 2593 2193 2607 2207
rect 2473 2073 2487 2087
rect 2473 2033 2487 2047
rect 2373 2013 2387 2027
rect 2433 2013 2447 2027
rect 2253 1912 2267 1926
rect 2093 1813 2107 1827
rect 2193 1813 2207 1827
rect 2193 1792 2207 1806
rect 2113 1734 2127 1748
rect 2153 1753 2167 1767
rect 2233 1753 2247 1767
rect 2313 1753 2327 1767
rect 2093 1693 2107 1707
rect 2293 1734 2307 1748
rect 2453 1912 2467 1926
rect 2393 1833 2407 1847
rect 2513 2172 2527 2186
rect 2533 2013 2547 2027
rect 2533 1954 2547 1968
rect 2573 1954 2587 1968
rect 2633 2213 2647 2227
rect 2773 2373 2787 2387
rect 2713 2254 2727 2268
rect 2753 2254 2767 2268
rect 3193 3113 3207 3127
rect 3193 3053 3207 3067
rect 3053 2873 3067 2887
rect 2973 2813 2987 2827
rect 3033 2774 3047 2788
rect 3013 2732 3027 2746
rect 2953 2693 2967 2707
rect 2953 2672 2967 2686
rect 2873 2513 2887 2527
rect 2913 2474 2927 2488
rect 3253 3014 3267 3028
rect 3353 3053 3367 3067
rect 3213 2972 3227 2986
rect 3313 2973 3327 2987
rect 3433 3153 3447 3167
rect 3373 3014 3387 3028
rect 3413 2994 3427 3008
rect 3233 2913 3247 2927
rect 3353 2913 3367 2927
rect 3113 2774 3127 2788
rect 3093 2732 3107 2746
rect 3053 2593 3067 2607
rect 3033 2513 3047 2527
rect 2993 2474 3007 2488
rect 2953 2453 2967 2467
rect 2833 2432 2847 2446
rect 2853 2313 2867 2327
rect 2833 2293 2847 2307
rect 3053 2432 3067 2446
rect 3113 2553 3127 2567
rect 3333 2893 3347 2907
rect 3473 3252 3487 3266
rect 3513 3252 3527 3266
rect 3473 3231 3487 3245
rect 3513 3173 3527 3187
rect 3553 3113 3567 3127
rect 3453 3073 3467 3087
rect 3553 3053 3567 3067
rect 3493 3033 3507 3047
rect 3433 2933 3447 2947
rect 3373 2813 3387 2827
rect 3233 2774 3247 2788
rect 3333 2774 3347 2788
rect 3193 2732 3207 2746
rect 3473 2713 3487 2727
rect 3513 2952 3527 2966
rect 3653 3294 3667 3308
rect 3633 3252 3647 3266
rect 3613 3213 3627 3227
rect 3673 3213 3687 3227
rect 3593 3093 3607 3107
rect 3533 2793 3547 2807
rect 3353 2673 3367 2687
rect 3393 2673 3407 2687
rect 3493 2673 3507 2687
rect 3373 2573 3387 2587
rect 3213 2474 3227 2488
rect 3253 2474 3267 2488
rect 3293 2474 3307 2488
rect 3333 2474 3347 2488
rect 3113 2432 3127 2446
rect 3153 2432 3167 2446
rect 3193 2432 3207 2446
rect 3093 2373 3107 2387
rect 3013 2313 3027 2327
rect 2793 2253 2807 2267
rect 2893 2273 2907 2287
rect 2913 2253 2927 2267
rect 2693 2173 2707 2187
rect 2653 2153 2667 2167
rect 2773 2153 2787 2167
rect 2633 1993 2647 2007
rect 2613 1973 2627 1987
rect 2733 1993 2747 2007
rect 2493 1873 2507 1887
rect 2553 1912 2567 1926
rect 2513 1853 2527 1867
rect 2473 1833 2487 1847
rect 2473 1812 2487 1826
rect 2553 1793 2567 1807
rect 2473 1773 2487 1787
rect 2693 1954 2707 1968
rect 2673 1912 2687 1926
rect 2453 1753 2467 1767
rect 2413 1733 2427 1747
rect 2493 1733 2507 1747
rect 2833 2212 2847 2226
rect 2873 2173 2887 2187
rect 2793 2113 2807 2127
rect 2793 2073 2807 2087
rect 2833 1954 2847 1968
rect 3033 2293 3047 2307
rect 3153 2293 3167 2307
rect 3253 2293 3267 2307
rect 3312 2293 3326 2307
rect 3333 2293 3347 2307
rect 2953 2273 2967 2287
rect 2993 2273 3007 2287
rect 3093 2254 3107 2268
rect 3193 2254 3207 2268
rect 3013 2113 3027 2127
rect 2953 2073 2967 2087
rect 2933 2033 2947 2047
rect 3013 2033 3027 2047
rect 3053 2033 3067 2047
rect 2953 1993 2967 2007
rect 2773 1912 2787 1926
rect 2773 1853 2787 1867
rect 2173 1692 2187 1706
rect 2233 1692 2247 1706
rect 2313 1692 2327 1706
rect 2393 1692 2407 1706
rect 2133 1613 2147 1627
rect 2313 1613 2327 1627
rect 2133 1573 2147 1587
rect 2273 1533 2287 1547
rect 2093 1473 2107 1487
rect 2233 1473 2247 1487
rect 2113 1453 2127 1467
rect 2333 1513 2347 1527
rect 2373 1513 2387 1527
rect 2313 1433 2327 1447
rect 2093 1392 2107 1406
rect 2033 1353 2047 1367
rect 2093 1353 2107 1367
rect 2013 1273 2027 1287
rect 1913 1253 1927 1267
rect 1993 1253 2007 1267
rect 1853 1214 1867 1228
rect 1793 1192 1807 1206
rect 1953 1214 1967 1228
rect 1873 1172 1887 1186
rect 1913 1172 1927 1186
rect 2173 1392 2187 1406
rect 2133 1213 2147 1227
rect 2153 1193 2167 1207
rect 2013 1172 2027 1186
rect 2073 1172 2087 1186
rect 1793 1153 1807 1167
rect 1773 1113 1787 1127
rect 1733 973 1747 987
rect 2153 1133 2167 1147
rect 2113 1053 2127 1067
rect 1893 973 1907 987
rect 2153 973 2167 987
rect 2253 1392 2267 1406
rect 2313 1393 2327 1407
rect 2253 1333 2267 1347
rect 2413 1434 2427 1448
rect 2873 1913 2887 1927
rect 2933 1912 2947 1926
rect 2873 1873 2887 1887
rect 2813 1813 2827 1827
rect 2813 1734 2827 1748
rect 2713 1692 2727 1706
rect 2753 1692 2767 1706
rect 3113 2213 3127 2227
rect 3173 2193 3187 2207
rect 3113 2113 3127 2127
rect 3093 1973 3107 1987
rect 3133 2053 3147 2067
rect 2913 1734 2927 1748
rect 2973 1734 2987 1748
rect 2673 1653 2687 1667
rect 2533 1533 2547 1547
rect 2833 1653 2847 1667
rect 2793 1613 2807 1627
rect 2813 1553 2827 1567
rect 2793 1533 2807 1547
rect 2713 1513 2727 1527
rect 2393 1392 2407 1406
rect 2433 1373 2447 1387
rect 2433 1333 2447 1347
rect 2373 1293 2387 1307
rect 2313 1214 2327 1228
rect 2353 1214 2367 1228
rect 2213 1172 2227 1186
rect 2233 1153 2247 1167
rect 2213 1133 2227 1147
rect 2193 993 2207 1007
rect 1793 953 1807 967
rect 1713 914 1727 928
rect 1813 914 1827 928
rect 1853 914 1867 928
rect 2093 933 2107 947
rect 1933 914 1947 928
rect 1973 914 1987 928
rect 2013 914 2027 928
rect 2073 914 2087 928
rect 1773 872 1787 886
rect 1833 872 1847 886
rect 1673 853 1687 867
rect 1673 813 1687 827
rect 1673 753 1687 767
rect 1653 713 1667 727
rect 1733 853 1747 867
rect 1873 813 1887 827
rect 1993 872 2007 886
rect 2033 872 2047 886
rect 1733 713 1747 727
rect 1713 693 1727 707
rect 1693 652 1707 666
rect 1653 633 1667 647
rect 1593 573 1607 587
rect 1893 713 1907 727
rect 1953 713 1967 727
rect 1833 693 1847 707
rect 1773 633 1787 647
rect 1813 593 1827 607
rect 1733 433 1747 447
rect 1573 413 1587 427
rect 1873 633 1887 647
rect 1833 513 1847 527
rect 1613 394 1627 408
rect 1553 373 1567 387
rect 1293 352 1307 366
rect 1333 352 1347 366
rect 1413 352 1427 366
rect 1473 352 1487 366
rect 1513 352 1527 366
rect 1713 394 1727 408
rect 1773 394 1787 408
rect 1813 394 1827 408
rect 1233 293 1247 307
rect 1393 293 1407 307
rect 1433 293 1447 307
rect 1313 253 1327 267
rect 1293 213 1307 227
rect 1253 174 1267 188
rect 1413 213 1427 227
rect 1593 352 1607 366
rect 1693 353 1707 367
rect 1633 333 1647 347
rect 1513 253 1527 267
rect 1513 213 1527 227
rect 1433 193 1447 207
rect 1453 174 1467 188
rect 1493 173 1507 187
rect 1553 213 1567 227
rect 1853 393 1867 407
rect 1713 333 1727 347
rect 1693 293 1707 307
rect 1793 313 1807 327
rect 1753 253 1767 267
rect 1573 193 1587 207
rect 1153 132 1167 146
rect 1253 133 1267 147
rect 1293 132 1307 146
rect 1393 132 1407 146
rect 1433 132 1447 146
rect 1193 93 1207 107
rect 1593 174 1607 188
rect 1713 174 1727 188
rect 1753 174 1767 188
rect 2093 873 2107 887
rect 2113 833 2127 847
rect 2073 813 2087 827
rect 2173 833 2187 847
rect 2133 793 2147 807
rect 2193 793 2207 807
rect 2353 1153 2367 1167
rect 2273 1133 2287 1147
rect 2313 1093 2327 1107
rect 2273 933 2287 947
rect 2533 1434 2547 1448
rect 2653 1434 2667 1448
rect 2693 1434 2707 1448
rect 2733 1434 2747 1448
rect 2973 1633 2987 1647
rect 2953 1613 2967 1627
rect 3113 1813 3127 1827
rect 3013 1793 3027 1807
rect 3073 1793 3087 1807
rect 2993 1593 3007 1607
rect 2833 1513 2847 1527
rect 2813 1473 2827 1487
rect 2933 1493 2947 1507
rect 2873 1473 2887 1487
rect 2513 1333 2527 1347
rect 2433 1273 2447 1287
rect 2473 1273 2487 1287
rect 2473 1214 2487 1228
rect 2613 1393 2627 1407
rect 2633 1373 2647 1387
rect 2653 1273 2667 1287
rect 2553 1214 2567 1228
rect 2613 1214 2627 1228
rect 2493 1172 2507 1186
rect 2533 1172 2547 1186
rect 2453 1153 2467 1167
rect 2553 1153 2567 1167
rect 2593 1153 2607 1167
rect 2433 1133 2447 1147
rect 2393 1053 2407 1067
rect 2733 1393 2747 1407
rect 3053 1734 3067 1748
rect 3153 1973 3167 1987
rect 3213 1993 3227 2007
rect 3233 1993 3247 2007
rect 3193 1954 3207 1968
rect 3293 2254 3307 2268
rect 3473 2553 3487 2567
rect 3413 2474 3427 2488
rect 3373 2254 3387 2268
rect 3433 2393 3447 2407
rect 3513 2433 3527 2447
rect 3493 2333 3507 2347
rect 3453 2293 3467 2307
rect 3513 2293 3527 2307
rect 3513 2272 3527 2286
rect 3313 2212 3327 2226
rect 3353 2213 3367 2227
rect 3353 2053 3367 2067
rect 3393 2233 3407 2247
rect 3313 1993 3327 2007
rect 3373 1993 3387 2007
rect 3253 1973 3267 1987
rect 3293 1973 3307 1987
rect 3153 1912 3167 1926
rect 3213 1912 3227 1926
rect 3193 1773 3207 1787
rect 3133 1734 3147 1748
rect 3233 1734 3247 1748
rect 3413 2073 3427 2087
rect 3333 1953 3347 1967
rect 3453 2013 3467 2027
rect 3493 1973 3507 1987
rect 3473 1953 3487 1967
rect 3313 1912 3327 1926
rect 3353 1912 3367 1926
rect 3433 1912 3447 1926
rect 3393 1833 3407 1847
rect 3093 1633 3107 1647
rect 3033 1493 3047 1507
rect 2973 1434 2987 1448
rect 3013 1434 3027 1448
rect 3093 1433 3107 1447
rect 2773 1392 2787 1406
rect 2873 1392 2887 1406
rect 2913 1392 2927 1406
rect 2813 1373 2827 1387
rect 2933 1373 2947 1387
rect 2713 1333 2727 1347
rect 2673 1213 2687 1227
rect 2753 1293 2767 1307
rect 2813 1273 2827 1287
rect 2793 1253 2807 1267
rect 2693 1172 2707 1186
rect 2733 1172 2747 1186
rect 2693 1133 2707 1147
rect 2733 1093 2747 1107
rect 2653 1033 2667 1047
rect 2753 1033 2767 1047
rect 2673 993 2687 1007
rect 2473 973 2487 987
rect 2513 973 2527 987
rect 2653 973 2667 987
rect 2453 913 2467 927
rect 2233 833 2247 847
rect 2033 694 2047 708
rect 2073 694 2087 708
rect 2113 694 2127 708
rect 1973 633 1987 647
rect 2053 652 2067 666
rect 1913 453 1927 467
rect 1953 394 1967 408
rect 2053 453 2067 467
rect 2013 394 2027 408
rect 2093 394 2107 408
rect 2392 873 2406 887
rect 2413 872 2427 886
rect 2293 773 2307 787
rect 2353 753 2367 767
rect 2253 694 2267 708
rect 2293 694 2307 708
rect 2133 652 2147 666
rect 2173 633 2187 647
rect 2133 613 2147 627
rect 2213 613 2227 627
rect 1893 353 1907 367
rect 1933 352 1947 366
rect 1992 353 2006 367
rect 2013 353 2027 367
rect 2113 353 2127 367
rect 2213 553 2227 567
rect 2153 394 2167 408
rect 2313 652 2327 666
rect 2413 813 2427 827
rect 2553 933 2567 947
rect 2593 933 2607 947
rect 2533 872 2547 886
rect 2693 933 2707 947
rect 2733 933 2747 947
rect 2613 913 2627 927
rect 2653 914 2667 928
rect 2473 692 2487 706
rect 2533 694 2547 708
rect 2593 793 2607 807
rect 2593 713 2607 727
rect 2573 693 2587 707
rect 2373 653 2387 667
rect 2413 652 2427 666
rect 2513 652 2527 666
rect 2553 652 2567 666
rect 2473 613 2487 627
rect 2353 593 2367 607
rect 2313 573 2327 587
rect 2273 473 2287 487
rect 2253 453 2267 467
rect 2373 473 2387 487
rect 2313 413 2327 427
rect 2073 333 2087 347
rect 1913 253 1927 267
rect 2073 253 2087 267
rect 1893 213 1907 227
rect 1873 193 1887 207
rect 1913 173 1927 187
rect 1953 174 1967 188
rect 2133 313 2147 327
rect 1893 153 1907 167
rect 1513 132 1527 146
rect 1573 132 1587 146
rect 1693 132 1707 146
rect 1833 132 1847 146
rect 1613 93 1627 107
rect 1493 73 1507 87
rect 1593 73 1607 87
rect 1933 132 1947 146
rect 1973 132 1987 146
rect 2053 132 2067 146
rect 2093 132 2107 146
rect 2133 132 2147 146
rect 2633 833 2647 847
rect 2673 833 2687 847
rect 2613 694 2627 708
rect 2593 573 2607 587
rect 2513 513 2527 527
rect 2233 352 2247 366
rect 2313 352 2327 366
rect 2393 352 2407 366
rect 2353 313 2367 327
rect 2253 273 2267 287
rect 2173 213 2187 227
rect 2213 213 2227 227
rect 2213 192 2227 206
rect 2173 173 2187 187
rect 2333 233 2347 247
rect 2433 213 2447 227
rect 2393 193 2407 207
rect 2593 453 2607 467
rect 2553 394 2567 408
rect 2533 313 2547 327
rect 2653 813 2667 827
rect 2653 753 2667 767
rect 2673 733 2687 747
rect 2673 694 2687 708
rect 2873 1214 2887 1228
rect 2853 1133 2867 1147
rect 2913 1133 2927 1147
rect 3013 1392 3027 1406
rect 3073 1392 3087 1406
rect 3213 1692 3227 1706
rect 3133 1513 3147 1527
rect 3113 1353 3127 1367
rect 3033 1313 3047 1327
rect 3093 1313 3107 1327
rect 2953 1273 2967 1287
rect 2993 1253 3007 1267
rect 3053 1253 3067 1267
rect 2953 1213 2967 1227
rect 3053 1172 3067 1186
rect 3113 1273 3127 1287
rect 3313 1734 3327 1748
rect 3353 1734 3367 1748
rect 3413 1734 3427 1748
rect 3473 1912 3487 1926
rect 3573 2893 3587 2907
rect 3653 3193 3667 3207
rect 3632 3073 3646 3087
rect 3653 3073 3667 3087
rect 3733 3453 3747 3467
rect 3733 3393 3747 3407
rect 3813 3673 3827 3687
rect 4033 3913 4047 3927
rect 4173 4193 4187 4207
rect 4193 4173 4207 4187
rect 4193 4093 4207 4107
rect 4153 3993 4167 4007
rect 4033 3873 4047 3887
rect 3953 3833 3967 3847
rect 4013 3833 4027 3847
rect 4013 3793 4027 3807
rect 4093 3853 4107 3867
rect 4133 3893 4147 3907
rect 4113 3833 4127 3847
rect 4133 3813 4147 3827
rect 3933 3772 3947 3786
rect 3993 3772 4007 3786
rect 4033 3773 4047 3787
rect 4073 3772 4087 3786
rect 3953 3713 3967 3727
rect 3933 3573 3947 3587
rect 3833 3533 3847 3547
rect 3893 3533 3907 3547
rect 3813 3513 3827 3527
rect 3813 3472 3827 3486
rect 3793 3413 3807 3427
rect 3753 3294 3767 3308
rect 3793 3293 3807 3307
rect 3793 3253 3807 3267
rect 3773 3173 3787 3187
rect 3673 3053 3687 3067
rect 3693 3033 3707 3047
rect 3853 3513 3867 3527
rect 3873 3472 3887 3486
rect 3853 3453 3867 3467
rect 3913 3453 3927 3467
rect 3873 3413 3887 3427
rect 3853 3393 3867 3407
rect 3833 3373 3847 3387
rect 3833 3352 3847 3366
rect 3873 3353 3887 3367
rect 3913 3353 3927 3367
rect 4073 3733 4087 3747
rect 4013 3573 4027 3587
rect 3993 3553 4007 3567
rect 3973 3453 3987 3467
rect 3973 3432 3987 3446
rect 3953 3393 3967 3407
rect 3953 3353 3967 3367
rect 3933 3333 3947 3347
rect 3853 3293 3867 3307
rect 3913 3294 3927 3308
rect 3873 3252 3887 3266
rect 3913 3233 3927 3247
rect 3853 3153 3867 3167
rect 3813 3113 3827 3127
rect 3853 3113 3867 3127
rect 3653 2994 3667 3008
rect 3713 2994 3727 3008
rect 3633 2952 3647 2966
rect 3693 2952 3707 2966
rect 3613 2793 3627 2807
rect 3593 2693 3607 2707
rect 3713 2933 3727 2947
rect 3733 2873 3747 2887
rect 3713 2813 3727 2827
rect 3853 2993 3867 3007
rect 3813 2952 3827 2966
rect 3793 2893 3807 2907
rect 3733 2774 3747 2788
rect 3633 2653 3647 2667
rect 3693 2713 3707 2727
rect 3753 2713 3767 2727
rect 3673 2633 3687 2647
rect 3653 2593 3667 2607
rect 3613 2553 3627 2567
rect 3633 2533 3647 2547
rect 3673 2513 3687 2527
rect 3573 2474 3587 2488
rect 3773 2613 3787 2627
rect 3753 2573 3767 2587
rect 3893 3073 3907 3087
rect 4013 3453 4027 3467
rect 3993 3373 4007 3387
rect 4053 3413 4067 3427
rect 3973 3253 3987 3267
rect 4033 3294 4047 3308
rect 4133 3773 4147 3787
rect 4173 3893 4187 3907
rect 4273 4173 4287 4187
rect 4253 4034 4267 4048
rect 4233 3993 4247 4007
rect 4213 3853 4227 3867
rect 4173 3813 4187 3827
rect 4213 3814 4227 3828
rect 4273 3993 4287 4007
rect 4333 4173 4347 4187
rect 4333 4113 4347 4127
rect 4433 4292 4447 4306
rect 4413 4273 4427 4287
rect 4353 4034 4367 4048
rect 4393 4032 4407 4046
rect 4293 3953 4307 3967
rect 4353 3913 4367 3927
rect 4333 3873 4347 3887
rect 4313 3833 4327 3847
rect 4153 3693 4167 3707
rect 4133 3673 4147 3687
rect 4173 3673 4187 3687
rect 4093 3633 4107 3647
rect 4133 3593 4147 3607
rect 4193 3613 4207 3627
rect 4193 3553 4207 3567
rect 4173 3533 4187 3547
rect 4093 3473 4107 3487
rect 4213 3514 4227 3528
rect 4113 3433 4127 3447
rect 4173 3413 4187 3427
rect 4153 3393 4167 3407
rect 4133 3293 4147 3307
rect 3953 3233 3967 3247
rect 3933 3213 3947 3227
rect 4113 3252 4127 3266
rect 3853 2853 3867 2867
rect 3813 2813 3827 2827
rect 3753 2493 3767 2507
rect 3733 2473 3747 2487
rect 3793 2473 3807 2487
rect 3693 2453 3707 2467
rect 3553 2353 3567 2367
rect 3633 2432 3647 2446
rect 3673 2432 3687 2446
rect 3653 2393 3667 2407
rect 3613 2353 3627 2367
rect 3593 2293 3607 2307
rect 3573 2273 3587 2287
rect 3553 2254 3567 2268
rect 3633 2333 3647 2347
rect 3613 2273 3627 2287
rect 3673 2373 3687 2387
rect 3653 2313 3667 2327
rect 3833 2773 3847 2787
rect 3833 2693 3847 2707
rect 3833 2613 3847 2627
rect 3953 2952 3967 2966
rect 3973 2933 3987 2947
rect 3953 2913 3967 2927
rect 4013 3013 4027 3027
rect 4053 3173 4067 3187
rect 4093 3213 4107 3227
rect 4093 3153 4107 3167
rect 4213 3393 4227 3407
rect 4293 3772 4307 3786
rect 4293 3733 4307 3747
rect 4313 3713 4327 3727
rect 4453 4213 4467 4227
rect 4533 4353 4547 4367
rect 4513 4334 4527 4348
rect 4553 4334 4567 4348
rect 4493 4293 4507 4307
rect 4573 4292 4587 4306
rect 4633 4473 4647 4487
rect 4773 4512 4787 4526
rect 4873 4773 4887 4787
rect 4893 4753 4907 4767
rect 4873 4713 4887 4727
rect 4913 4633 4927 4647
rect 4893 4593 4907 4607
rect 4833 4552 4847 4566
rect 4873 4554 4887 4568
rect 5033 5293 5047 5307
rect 4993 5173 5007 5187
rect 5093 5273 5107 5287
rect 5053 5193 5067 5207
rect 4973 5093 4987 5107
rect 5033 5093 5047 5107
rect 4953 4993 4967 5007
rect 5033 5032 5047 5046
rect 5073 5033 5087 5047
rect 5253 5513 5267 5527
rect 5193 5493 5207 5507
rect 5233 5493 5247 5507
rect 5233 5433 5247 5447
rect 5193 5374 5207 5388
rect 5313 5594 5327 5608
rect 5793 6153 5807 6167
rect 6193 6153 6207 6167
rect 5833 6114 5847 6128
rect 5893 6113 5907 6127
rect 5953 6114 5967 6128
rect 5993 6114 6007 6128
rect 6053 6113 6067 6127
rect 6113 6114 6127 6128
rect 5813 6072 5827 6086
rect 5853 6072 5867 6086
rect 5933 6072 5947 6086
rect 5893 6013 5907 6027
rect 5753 5993 5767 6007
rect 5953 5993 5967 6007
rect 5693 5973 5707 5987
rect 5753 5972 5767 5986
rect 5673 5933 5687 5947
rect 5713 5894 5727 5908
rect 5653 5852 5667 5866
rect 5733 5853 5747 5867
rect 5693 5773 5707 5787
rect 5613 5733 5627 5747
rect 5553 5693 5567 5707
rect 5453 5673 5467 5687
rect 5413 5653 5427 5667
rect 5333 5552 5347 5566
rect 5393 5552 5407 5566
rect 5513 5653 5527 5667
rect 5933 5913 5947 5927
rect 5773 5893 5787 5907
rect 5813 5894 5827 5908
rect 5853 5894 5867 5908
rect 5912 5893 5926 5907
rect 6033 6073 6047 6087
rect 5993 5973 6007 5987
rect 5973 5933 5987 5947
rect 5993 5894 6007 5908
rect 6093 6072 6107 6086
rect 6193 6072 6207 6086
rect 6053 5973 6067 5987
rect 6053 5913 6067 5927
rect 6153 5913 6167 5927
rect 5793 5853 5807 5867
rect 5773 5793 5787 5807
rect 5613 5594 5627 5608
rect 5493 5552 5507 5566
rect 5553 5552 5567 5566
rect 5413 5513 5427 5527
rect 5593 5513 5607 5527
rect 5373 5473 5387 5487
rect 5313 5433 5327 5447
rect 5173 5313 5187 5327
rect 5133 5273 5147 5287
rect 5213 5273 5227 5287
rect 5153 5233 5167 5247
rect 5113 5153 5127 5167
rect 5152 5133 5166 5147
rect 5173 5133 5187 5147
rect 5113 5093 5127 5107
rect 5213 5113 5227 5127
rect 5153 5032 5167 5046
rect 5193 5032 5207 5046
rect 5333 5374 5347 5388
rect 5433 5493 5447 5507
rect 5553 5493 5567 5507
rect 5413 5374 5427 5388
rect 5453 5473 5467 5487
rect 5513 5473 5527 5487
rect 5433 5353 5447 5367
rect 5513 5393 5527 5407
rect 5473 5374 5487 5388
rect 5353 5332 5367 5346
rect 5393 5332 5407 5346
rect 5393 5233 5407 5247
rect 5273 5153 5287 5167
rect 5313 5173 5327 5187
rect 5433 5313 5447 5327
rect 5533 5333 5547 5347
rect 5492 5273 5506 5287
rect 5513 5273 5527 5287
rect 5453 5233 5467 5247
rect 5433 5213 5447 5227
rect 5453 5193 5467 5207
rect 5513 5173 5527 5187
rect 5413 5133 5427 5147
rect 5793 5773 5807 5787
rect 5813 5733 5827 5747
rect 5773 5594 5787 5608
rect 5853 5793 5867 5807
rect 5833 5633 5847 5647
rect 5713 5552 5727 5566
rect 5753 5552 5767 5566
rect 5653 5433 5667 5447
rect 5612 5393 5626 5407
rect 5633 5393 5647 5407
rect 5693 5513 5707 5527
rect 5793 5493 5807 5507
rect 5713 5453 5727 5467
rect 5693 5413 5707 5427
rect 5673 5373 5687 5387
rect 5633 5332 5647 5346
rect 5673 5333 5687 5347
rect 5613 5293 5627 5307
rect 5593 5193 5607 5207
rect 5573 5153 5587 5167
rect 5533 5113 5547 5127
rect 5353 5074 5367 5088
rect 5393 5074 5407 5088
rect 5433 5073 5447 5087
rect 5533 5074 5547 5088
rect 5273 5053 5287 5067
rect 5113 4993 5127 5007
rect 5093 4973 5107 4987
rect 5073 4953 5087 4967
rect 5253 4973 5267 4987
rect 4993 4933 5007 4947
rect 5093 4933 5107 4947
rect 5233 4933 5247 4947
rect 5113 4913 5127 4927
rect 5213 4913 5227 4927
rect 5093 4893 5107 4907
rect 5033 4854 5047 4868
rect 5233 4892 5247 4906
rect 5153 4873 5167 4887
rect 5193 4854 5207 4868
rect 5053 4812 5067 4826
rect 5093 4812 5107 4826
rect 5173 4812 5187 4826
rect 5233 4812 5247 4826
rect 5153 4773 5167 4787
rect 4953 4713 4967 4727
rect 5133 4713 5147 4727
rect 5093 4673 5107 4687
rect 4993 4613 5007 4627
rect 4933 4573 4947 4587
rect 4973 4573 4987 4587
rect 4833 4513 4847 4527
rect 4833 4433 4847 4447
rect 4753 4353 4767 4367
rect 4673 4334 4687 4348
rect 4713 4334 4727 4348
rect 4653 4292 4667 4306
rect 4553 4253 4567 4267
rect 4653 4253 4667 4267
rect 4473 4073 4487 4087
rect 4533 4073 4547 4087
rect 4493 4034 4507 4048
rect 4433 3992 4447 4006
rect 4473 3992 4487 4006
rect 4533 3992 4547 4006
rect 4513 3953 4527 3967
rect 4473 3833 4487 3847
rect 4433 3813 4447 3827
rect 4513 3814 4527 3828
rect 4593 4233 4607 4247
rect 4553 3793 4567 3807
rect 4473 3753 4487 3767
rect 4413 3713 4427 3727
rect 4453 3713 4467 3727
rect 4393 3593 4407 3607
rect 4313 3553 4327 3567
rect 4373 3553 4387 3567
rect 4273 3514 4287 3528
rect 4353 3533 4367 3547
rect 4293 3472 4307 3486
rect 4333 3373 4347 3387
rect 4193 3313 4207 3327
rect 4233 3313 4247 3327
rect 4173 3293 4187 3307
rect 4433 3514 4447 3528
rect 4493 3732 4507 3746
rect 4513 3653 4527 3667
rect 4393 3473 4407 3487
rect 4413 3453 4427 3467
rect 4372 3393 4386 3407
rect 4393 3393 4407 3407
rect 4353 3353 4367 3367
rect 4153 3213 4167 3227
rect 4133 3113 4147 3127
rect 4213 3093 4227 3107
rect 4113 3073 4127 3087
rect 4393 3293 4407 3307
rect 4313 3252 4327 3266
rect 4393 3252 4407 3266
rect 4353 3193 4367 3207
rect 4493 3453 4507 3467
rect 4633 4213 4647 4227
rect 4733 4213 4747 4227
rect 4653 4173 4667 4187
rect 4633 4153 4647 4167
rect 4673 4133 4687 4147
rect 4653 4073 4667 4087
rect 4633 3992 4647 4006
rect 4593 3833 4607 3847
rect 4633 3833 4647 3847
rect 4633 3673 4647 3687
rect 4633 3613 4647 3627
rect 4533 3513 4547 3527
rect 4613 3533 4627 3547
rect 4633 3513 4647 3527
rect 4533 3473 4547 3487
rect 4513 3413 4527 3427
rect 4453 3353 4467 3367
rect 4433 3333 4447 3347
rect 4473 3294 4487 3308
rect 4333 3133 4347 3147
rect 4273 3053 4287 3067
rect 4333 3053 4347 3067
rect 4093 3033 4107 3047
rect 4253 3033 4267 3047
rect 4033 2993 4047 3007
rect 4093 2994 4107 3008
rect 4133 2994 4147 3008
rect 4213 2994 4227 3008
rect 4313 2994 4327 3008
rect 4173 2973 4187 2987
rect 4033 2953 4047 2967
rect 3993 2893 4007 2907
rect 3933 2833 3947 2847
rect 3973 2833 3987 2847
rect 4013 2833 4027 2847
rect 3953 2793 3967 2807
rect 3873 2673 3887 2687
rect 3933 2673 3947 2687
rect 3853 2593 3867 2607
rect 3873 2573 3887 2587
rect 3913 2533 3927 2547
rect 3933 2473 3947 2487
rect 3833 2453 3847 2467
rect 3813 2373 3827 2387
rect 3713 2353 3727 2367
rect 3753 2353 3767 2367
rect 3693 2313 3707 2327
rect 3753 2313 3767 2327
rect 3573 2212 3587 2226
rect 3553 2193 3567 2207
rect 3533 2113 3547 2127
rect 3533 2073 3547 2087
rect 3573 2153 3587 2167
rect 3553 1993 3567 2007
rect 3573 1954 3587 1968
rect 3673 2253 3687 2267
rect 3713 2254 3727 2268
rect 3753 2254 3767 2268
rect 3693 2212 3707 2226
rect 3673 2153 3687 2167
rect 3653 2093 3667 2107
rect 3793 2213 3807 2227
rect 3732 2153 3746 2167
rect 3753 2153 3767 2167
rect 3693 2113 3707 2127
rect 3753 2093 3767 2107
rect 3713 2053 3727 2067
rect 3673 1973 3687 1987
rect 3633 1953 3647 1967
rect 3733 2033 3747 2047
rect 3773 2033 3787 2047
rect 3833 2293 3847 2307
rect 3933 2373 3947 2387
rect 3933 2293 3947 2307
rect 3893 2273 3907 2287
rect 4053 2933 4067 2947
rect 4033 2793 4047 2807
rect 4033 2732 4047 2746
rect 4013 2713 4027 2727
rect 3993 2653 4007 2667
rect 3973 2633 3987 2647
rect 4153 2953 4167 2967
rect 4172 2913 4186 2927
rect 4193 2912 4207 2926
rect 4153 2873 4167 2887
rect 4193 2873 4207 2887
rect 4113 2853 4127 2867
rect 4093 2813 4107 2827
rect 4313 2953 4327 2967
rect 4393 3153 4407 3167
rect 4453 3252 4467 3266
rect 4593 3472 4607 3486
rect 4553 3413 4567 3427
rect 4613 3393 4627 3407
rect 4573 3313 4587 3327
rect 4773 4333 4787 4347
rect 4813 4334 4827 4348
rect 4953 4512 4967 4526
rect 4933 4473 4947 4487
rect 4933 4433 4947 4447
rect 4833 4292 4847 4306
rect 5053 4554 5067 4568
rect 5033 4512 5047 4526
rect 5113 4633 5127 4647
rect 5093 4453 5107 4467
rect 4993 4433 5007 4447
rect 5013 4373 5027 4387
rect 4973 4353 4987 4367
rect 5093 4334 5107 4348
rect 5153 4554 5167 4568
rect 5193 4554 5207 4568
rect 5233 4554 5247 4568
rect 5333 5032 5347 5046
rect 5413 5033 5427 5047
rect 5353 5013 5367 5027
rect 5273 4953 5287 4967
rect 5293 4913 5307 4927
rect 5313 4913 5327 4927
rect 5373 4953 5387 4967
rect 5332 4893 5346 4907
rect 5353 4893 5367 4907
rect 5353 4854 5367 4868
rect 5513 5032 5527 5046
rect 5473 5013 5487 5027
rect 5533 4953 5547 4967
rect 5413 4893 5427 4907
rect 5473 4893 5487 4907
rect 5513 4893 5527 4907
rect 5393 4873 5407 4887
rect 5273 4813 5287 4827
rect 5173 4493 5187 4507
rect 5173 4453 5187 4467
rect 4933 4312 4947 4326
rect 4913 4292 4927 4306
rect 4893 4253 4907 4267
rect 4873 4213 4887 4227
rect 4773 4133 4787 4147
rect 4833 4133 4847 4147
rect 4773 4093 4787 4107
rect 4753 4073 4767 4087
rect 4693 4033 4707 4047
rect 4733 4034 4747 4048
rect 4673 3993 4687 4007
rect 4673 3793 4687 3807
rect 4753 3992 4767 4006
rect 4993 4292 5007 4306
rect 5073 4292 5087 4306
rect 5033 4273 5047 4287
rect 5133 4334 5147 4348
rect 5173 4334 5187 4348
rect 5113 4293 5127 4307
rect 5093 4133 5107 4147
rect 5053 4093 5067 4107
rect 4933 4053 4947 4067
rect 4973 4053 4987 4067
rect 4853 4034 4867 4048
rect 4893 4034 4907 4048
rect 4793 3973 4807 3987
rect 4793 3853 4807 3867
rect 4733 3814 4747 3828
rect 4753 3772 4767 3786
rect 4673 3613 4687 3627
rect 4693 3593 4707 3607
rect 4673 3573 4687 3587
rect 4693 3513 4707 3527
rect 4773 3673 4787 3687
rect 4833 3992 4847 4006
rect 4873 3973 4887 3987
rect 5007 4033 5021 4047
rect 5093 4033 5107 4047
rect 4913 3953 4927 3967
rect 4893 3853 4907 3867
rect 4833 3814 4847 3828
rect 4933 3833 4947 3847
rect 4813 3773 4827 3787
rect 4873 3772 4887 3786
rect 4913 3772 4927 3786
rect 4833 3713 4847 3727
rect 4853 3693 4867 3707
rect 4833 3653 4847 3667
rect 4793 3553 4807 3567
rect 4753 3514 4767 3528
rect 4813 3493 4827 3507
rect 4693 3473 4707 3487
rect 4673 3433 4687 3447
rect 4733 3472 4747 3486
rect 4733 3433 4747 3447
rect 4693 3413 4707 3427
rect 4653 3393 4667 3407
rect 4633 3373 4647 3387
rect 4653 3353 4667 3367
rect 4693 3353 4707 3367
rect 4793 3473 4807 3487
rect 4773 3413 4787 3427
rect 4813 3353 4827 3367
rect 4453 3173 4467 3187
rect 4453 3093 4467 3107
rect 4453 3072 4467 3086
rect 4533 3233 4547 3247
rect 4553 3213 4567 3227
rect 4533 3153 4547 3167
rect 4533 3113 4547 3127
rect 4513 3033 4527 3047
rect 4433 2993 4447 3007
rect 4413 2952 4427 2966
rect 4453 2953 4467 2967
rect 4433 2933 4447 2947
rect 4353 2913 4367 2927
rect 4293 2893 4307 2907
rect 4333 2893 4347 2907
rect 4393 2893 4407 2907
rect 4273 2873 4287 2887
rect 4233 2853 4247 2867
rect 4213 2813 4227 2827
rect 4093 2773 4107 2787
rect 4173 2774 4187 2788
rect 4193 2732 4207 2746
rect 4073 2653 4087 2667
rect 4013 2553 4027 2567
rect 4053 2613 4067 2627
rect 4073 2533 4087 2547
rect 4053 2513 4067 2527
rect 3993 2473 4007 2487
rect 4033 2474 4047 2488
rect 4213 2693 4227 2707
rect 4173 2673 4187 2687
rect 4153 2653 4167 2667
rect 4173 2573 4187 2587
rect 4153 2493 4167 2507
rect 4113 2473 4127 2487
rect 4213 2513 4227 2527
rect 4213 2473 4227 2487
rect 4253 2813 4267 2827
rect 4353 2833 4367 2847
rect 4333 2813 4347 2827
rect 4273 2793 4287 2807
rect 4253 2773 4267 2787
rect 4293 2774 4307 2788
rect 4333 2773 4347 2787
rect 4393 2773 4407 2787
rect 4493 2993 4507 3007
rect 4473 2933 4487 2947
rect 4493 2913 4507 2927
rect 4453 2893 4467 2907
rect 4493 2833 4507 2847
rect 4633 3252 4647 3266
rect 4693 3294 4707 3308
rect 4733 3294 4747 3308
rect 4693 3233 4707 3247
rect 4673 3213 4687 3227
rect 4593 3133 4607 3147
rect 4633 3133 4647 3147
rect 4613 3053 4627 3067
rect 4553 3013 4567 3027
rect 4593 2994 4607 3008
rect 4653 3033 4667 3047
rect 4633 3012 4647 3026
rect 4613 2973 4627 2987
rect 4553 2933 4567 2947
rect 4553 2853 4567 2867
rect 4613 2952 4627 2966
rect 4753 3253 4767 3267
rect 4753 3173 4767 3187
rect 4853 3573 4867 3587
rect 4893 3533 4907 3547
rect 4973 3973 4987 3987
rect 4973 3933 4987 3947
rect 5033 3992 5047 4006
rect 5093 3953 5107 3967
rect 5073 3893 5087 3907
rect 4992 3833 5006 3847
rect 5013 3833 5027 3847
rect 5033 3772 5047 3786
rect 5033 3751 5047 3765
rect 5093 3753 5107 3767
rect 4993 3673 5007 3687
rect 5013 3593 5027 3607
rect 4932 3514 4946 3528
rect 4953 3514 4967 3528
rect 4893 3453 4907 3467
rect 4973 3453 4987 3467
rect 4873 3373 4887 3387
rect 4853 3353 4867 3367
rect 4833 3313 4847 3327
rect 4973 3393 4987 3407
rect 4933 3373 4947 3387
rect 4913 3313 4927 3327
rect 4893 3293 4907 3307
rect 5253 4513 5267 4527
rect 5333 4812 5347 4826
rect 5293 4773 5307 4787
rect 5313 4693 5327 4707
rect 5353 4753 5367 4767
rect 5333 4633 5347 4647
rect 5313 4613 5327 4627
rect 5373 4693 5387 4707
rect 5273 4473 5287 4487
rect 5433 4854 5447 4868
rect 5713 5373 5727 5387
rect 5753 5374 5767 5388
rect 5793 5374 5807 5388
rect 5913 5852 5927 5866
rect 5873 5753 5887 5767
rect 5933 5813 5947 5827
rect 5913 5693 5927 5707
rect 6013 5852 6027 5866
rect 5953 5633 5967 5647
rect 5973 5633 5987 5647
rect 5913 5613 5927 5627
rect 5933 5552 5947 5566
rect 5993 5552 6007 5566
rect 5893 5513 5907 5527
rect 5873 5473 5887 5487
rect 5853 5373 5867 5387
rect 5692 5313 5706 5327
rect 5713 5313 5727 5327
rect 5673 5273 5687 5287
rect 5653 5113 5667 5127
rect 5633 5093 5647 5107
rect 5613 5073 5627 5087
rect 5633 5032 5647 5046
rect 5773 5332 5787 5346
rect 5773 5253 5787 5267
rect 5833 5333 5847 5347
rect 5973 5393 5987 5407
rect 5933 5374 5947 5388
rect 5993 5373 6007 5387
rect 5873 5313 5887 5327
rect 5992 5333 6006 5347
rect 6113 5894 6127 5908
rect 6093 5813 6107 5827
rect 6053 5793 6067 5807
rect 6133 5793 6147 5807
rect 6093 5653 6107 5667
rect 6033 5633 6047 5647
rect 6213 6013 6227 6027
rect 6193 5753 6207 5767
rect 6213 5613 6227 5627
rect 6193 5513 6207 5527
rect 6133 5473 6147 5487
rect 6033 5393 6047 5407
rect 6073 5393 6087 5407
rect 5953 5273 5967 5287
rect 5813 5233 5827 5247
rect 5913 5233 5927 5247
rect 5733 5193 5747 5207
rect 5833 5173 5847 5187
rect 5733 5074 5747 5088
rect 5793 5074 5807 5088
rect 6013 5332 6027 5346
rect 6153 5393 6167 5407
rect 6093 5332 6107 5346
rect 6033 5293 6047 5307
rect 6113 5173 6127 5187
rect 5933 5153 5947 5167
rect 5993 5153 6007 5167
rect 6093 5153 6107 5167
rect 6013 5113 6027 5127
rect 5973 5074 5987 5088
rect 5613 4993 5627 5007
rect 5613 4953 5627 4967
rect 5493 4812 5507 4826
rect 5533 4812 5547 4826
rect 5673 4973 5687 4987
rect 5633 4933 5647 4947
rect 5673 4893 5687 4907
rect 5653 4873 5667 4887
rect 5713 4933 5727 4947
rect 5713 4893 5727 4907
rect 5773 5032 5787 5046
rect 5813 5032 5827 5046
rect 5753 4993 5767 5007
rect 5753 4913 5767 4927
rect 5733 4873 5747 4887
rect 5773 4854 5787 4868
rect 5832 4993 5846 5007
rect 5853 4993 5867 5007
rect 5713 4813 5727 4827
rect 5593 4793 5607 4807
rect 5693 4793 5707 4807
rect 5433 4653 5447 4667
rect 5573 4613 5587 4627
rect 5413 4553 5427 4567
rect 5453 4554 5467 4568
rect 5493 4554 5507 4568
rect 5533 4553 5547 4567
rect 5693 4772 5707 4786
rect 5333 4433 5347 4447
rect 5233 4373 5247 4387
rect 5213 4213 5227 4227
rect 5153 4173 5167 4187
rect 5213 4133 5227 4147
rect 5133 4053 5147 4067
rect 5193 4053 5207 4067
rect 5213 4033 5227 4047
rect 5133 3993 5147 4007
rect 5213 3993 5227 4007
rect 5173 3893 5187 3907
rect 5153 3814 5167 3828
rect 5193 3814 5207 3828
rect 5293 4334 5307 4348
rect 5313 4253 5327 4267
rect 5393 4493 5407 4507
rect 5413 4473 5427 4487
rect 5513 4512 5527 4526
rect 5533 4453 5547 4467
rect 5593 4553 5607 4567
rect 5593 4493 5607 4507
rect 5553 4433 5567 4447
rect 5473 4373 5487 4387
rect 5413 4354 5427 4368
rect 5453 4353 5467 4367
rect 5413 4333 5427 4347
rect 5573 4413 5587 4427
rect 5673 4513 5687 4527
rect 5613 4473 5627 4487
rect 5653 4473 5667 4487
rect 5593 4373 5607 4387
rect 5753 4793 5767 4807
rect 5753 4693 5767 4707
rect 5813 4792 5827 4806
rect 5893 4953 5907 4967
rect 5873 4933 5887 4947
rect 5853 4913 5867 4927
rect 5853 4853 5867 4867
rect 5933 4993 5947 5007
rect 5953 4953 5967 4967
rect 5993 4913 6007 4927
rect 5912 4873 5926 4887
rect 5933 4873 5947 4887
rect 5973 4873 5987 4887
rect 5853 4813 5867 4827
rect 5793 4753 5807 4767
rect 5813 4733 5827 4747
rect 5813 4673 5827 4687
rect 5773 4633 5787 4647
rect 5913 4812 5927 4826
rect 5872 4772 5886 4786
rect 5893 4773 5907 4787
rect 5873 4713 5887 4727
rect 5953 4753 5967 4767
rect 5933 4733 5947 4747
rect 5853 4613 5867 4627
rect 5833 4593 5847 4607
rect 5793 4573 5807 4587
rect 5813 4554 5827 4568
rect 5753 4512 5767 4526
rect 5793 4473 5807 4487
rect 5873 4554 5887 4568
rect 5933 4553 5947 4567
rect 5693 4453 5707 4467
rect 5753 4453 5767 4467
rect 5813 4453 5827 4467
rect 5693 4432 5707 4446
rect 5633 4353 5647 4367
rect 5673 4353 5687 4367
rect 5613 4334 5627 4348
rect 5513 4313 5527 4327
rect 5373 4273 5387 4287
rect 5473 4292 5487 4306
rect 5373 4252 5387 4266
rect 5273 4233 5287 4247
rect 5273 4034 5287 4048
rect 5333 4213 5347 4227
rect 5353 4053 5367 4067
rect 5333 4013 5347 4027
rect 5293 3973 5307 3987
rect 5333 3953 5347 3967
rect 5393 4233 5407 4247
rect 5373 4033 5387 4047
rect 5453 4273 5467 4287
rect 5433 4213 5447 4227
rect 5413 4193 5427 4207
rect 5573 4292 5587 4306
rect 5653 4334 5667 4348
rect 5873 4493 5887 4507
rect 5853 4373 5867 4387
rect 5753 4333 5767 4347
rect 5833 4334 5847 4348
rect 5893 4413 5907 4427
rect 5873 4333 5887 4347
rect 5513 4213 5527 4227
rect 5613 4213 5627 4227
rect 5453 4093 5467 4107
rect 5613 4093 5627 4107
rect 5613 4053 5627 4067
rect 5473 4034 5487 4048
rect 5513 4034 5527 4048
rect 5573 4034 5587 4048
rect 5673 4193 5687 4207
rect 5673 4093 5687 4107
rect 5753 4292 5767 4306
rect 5773 4233 5787 4247
rect 5873 4293 5887 4307
rect 5853 4213 5867 4227
rect 5833 4113 5847 4127
rect 5733 4073 5747 4087
rect 5273 3853 5287 3867
rect 5353 3853 5367 3867
rect 5253 3833 5267 3847
rect 5133 3693 5147 3707
rect 5213 3772 5227 3786
rect 5253 3772 5267 3786
rect 5193 3693 5207 3707
rect 5173 3673 5187 3687
rect 5113 3593 5127 3607
rect 5053 3533 5067 3547
rect 5113 3533 5127 3547
rect 5033 3493 5047 3507
rect 5093 3472 5107 3486
rect 5133 3472 5147 3486
rect 5153 3453 5167 3467
rect 5133 3433 5147 3447
rect 5073 3393 5087 3407
rect 5073 3333 5087 3347
rect 5013 3313 5027 3327
rect 5053 3313 5067 3327
rect 4973 3294 4987 3308
rect 4873 3252 4887 3266
rect 4912 3252 4926 3266
rect 4933 3253 4947 3267
rect 4833 3213 4847 3227
rect 4773 3133 4787 3147
rect 4813 3053 4827 3067
rect 4713 3033 4727 3047
rect 4693 2994 4707 3008
rect 4733 2994 4747 3008
rect 4773 2994 4787 3008
rect 4853 3013 4867 3027
rect 4913 3073 4927 3087
rect 4633 2893 4647 2907
rect 4633 2853 4647 2867
rect 4533 2833 4547 2847
rect 4573 2833 4587 2847
rect 4513 2773 4527 2787
rect 4373 2752 4387 2766
rect 4273 2732 4287 2746
rect 4313 2732 4327 2746
rect 4353 2732 4367 2746
rect 4313 2673 4327 2687
rect 4313 2613 4327 2627
rect 4253 2573 4267 2587
rect 4293 2533 4307 2547
rect 3973 2433 3987 2447
rect 4013 2432 4027 2446
rect 3973 2412 3987 2426
rect 4033 2413 4047 2427
rect 4033 2373 4047 2387
rect 4053 2353 4067 2367
rect 4093 2353 4107 2367
rect 4073 2333 4087 2347
rect 3993 2293 4007 2307
rect 3973 2273 3987 2287
rect 3833 2073 3847 2087
rect 3753 2013 3767 2027
rect 3793 1993 3807 2007
rect 3772 1953 3786 1967
rect 3793 1953 3807 1967
rect 3873 2212 3887 2226
rect 3893 2173 3907 2187
rect 3893 2113 3907 2127
rect 3953 2173 3967 2187
rect 3933 2113 3947 2127
rect 3913 2093 3927 2107
rect 3873 2053 3887 2067
rect 3893 1953 3907 1967
rect 3973 2153 3987 2167
rect 4153 2353 4167 2367
rect 4112 2293 4126 2307
rect 4133 2293 4147 2307
rect 4113 2213 4127 2227
rect 4093 2173 4107 2187
rect 4033 2153 4047 2167
rect 4093 2152 4107 2166
rect 4153 2253 4167 2267
rect 4233 2293 4247 2307
rect 4333 2474 4347 2488
rect 4593 2813 4607 2827
rect 4553 2773 4567 2787
rect 4673 2952 4687 2966
rect 4653 2793 4667 2807
rect 4633 2773 4647 2787
rect 4953 3173 4967 3187
rect 4973 3133 4987 3147
rect 4933 3033 4947 3047
rect 4793 2953 4807 2967
rect 4773 2913 4787 2927
rect 4713 2893 4727 2907
rect 4773 2892 4787 2906
rect 4813 2933 4827 2947
rect 4793 2853 4807 2867
rect 4773 2833 4787 2847
rect 4793 2813 4807 2827
rect 4693 2793 4707 2807
rect 4573 2732 4587 2746
rect 4613 2732 4627 2746
rect 4493 2713 4507 2727
rect 4453 2693 4467 2707
rect 4413 2593 4427 2607
rect 4453 2593 4467 2607
rect 4413 2572 4427 2586
rect 4413 2474 4427 2488
rect 4453 2474 4467 2488
rect 4593 2713 4607 2727
rect 4513 2633 4527 2647
rect 4493 2513 4507 2527
rect 4273 2353 4287 2367
rect 4333 2353 4347 2367
rect 4313 2313 4327 2327
rect 4313 2292 4327 2306
rect 4273 2273 4287 2287
rect 4253 2253 4267 2267
rect 4112 2113 4126 2127
rect 4133 2113 4147 2127
rect 4093 2093 4107 2107
rect 4013 2033 4027 2047
rect 3973 1973 3987 1987
rect 3553 1912 3567 1926
rect 3613 1913 3627 1927
rect 3653 1912 3667 1926
rect 3493 1793 3507 1807
rect 3653 1833 3667 1847
rect 3613 1793 3627 1807
rect 3533 1753 3547 1767
rect 3293 1693 3307 1707
rect 3273 1673 3287 1687
rect 3213 1493 3227 1507
rect 3273 1493 3287 1507
rect 3193 1473 3207 1487
rect 3153 1434 3167 1448
rect 3233 1434 3247 1448
rect 3173 1392 3187 1406
rect 3273 1392 3287 1406
rect 3213 1353 3227 1367
rect 3193 1273 3207 1287
rect 3153 1253 3167 1267
rect 3133 1233 3147 1247
rect 3173 1233 3187 1247
rect 2813 993 2827 1007
rect 2793 933 2807 947
rect 2813 914 2827 928
rect 2893 914 2907 928
rect 2753 853 2767 867
rect 2733 673 2747 687
rect 2833 872 2847 886
rect 2913 893 2927 907
rect 2893 833 2907 847
rect 2913 813 2927 827
rect 2793 773 2807 787
rect 2913 773 2927 787
rect 2853 733 2867 747
rect 2813 694 2827 708
rect 2753 633 2767 647
rect 2793 613 2807 627
rect 2773 553 2787 567
rect 2673 513 2687 527
rect 2653 473 2667 487
rect 2633 433 2647 447
rect 2613 394 2627 408
rect 2753 433 2767 447
rect 2713 394 2727 408
rect 2612 313 2626 327
rect 2633 313 2647 327
rect 2593 293 2607 307
rect 2693 352 2707 366
rect 2713 333 2727 347
rect 2673 313 2687 327
rect 2653 253 2667 267
rect 2673 233 2687 247
rect 2573 213 2587 227
rect 2673 212 2687 226
rect 2473 193 2487 207
rect 2593 193 2607 207
rect 2493 173 2507 187
rect 2553 174 2567 188
rect 2733 213 2747 227
rect 2873 652 2887 666
rect 2853 453 2867 467
rect 2833 433 2847 447
rect 2893 433 2907 447
rect 2793 394 2807 408
rect 2773 353 2787 367
rect 2773 313 2787 327
rect 2813 313 2827 327
rect 2873 353 2887 367
rect 2753 193 2767 207
rect 2173 132 2187 146
rect 2233 132 2247 146
rect 2333 132 2347 146
rect 2373 132 2387 146
rect 2413 132 2427 146
rect 2473 132 2487 146
rect 2533 132 2547 146
rect 2613 133 2627 147
rect 2993 853 3007 867
rect 3093 1172 3107 1186
rect 3253 1293 3267 1307
rect 3373 1692 3387 1706
rect 3333 1673 3347 1687
rect 3413 1653 3427 1667
rect 3313 1613 3327 1627
rect 3353 1473 3367 1487
rect 3313 1433 3327 1447
rect 3473 1692 3487 1706
rect 3473 1553 3487 1567
rect 3333 1392 3347 1406
rect 3373 1353 3387 1367
rect 3293 1313 3307 1327
rect 3373 1332 3387 1346
rect 3313 1293 3327 1307
rect 3313 1253 3327 1267
rect 3233 1213 3247 1227
rect 3213 1133 3227 1147
rect 3173 1093 3187 1107
rect 3133 914 3147 928
rect 3273 1233 3287 1247
rect 3253 1172 3267 1186
rect 3293 1172 3307 1186
rect 3333 1133 3347 1147
rect 3233 1073 3247 1087
rect 3373 1033 3387 1047
rect 3453 1392 3467 1406
rect 3513 1373 3527 1387
rect 3493 1353 3507 1367
rect 3453 1333 3467 1347
rect 3433 1273 3447 1287
rect 3493 1193 3507 1207
rect 3473 1172 3487 1186
rect 3413 1073 3427 1087
rect 3213 993 3227 1007
rect 3393 993 3407 1007
rect 3073 893 3087 907
rect 3113 872 3127 886
rect 3153 853 3167 867
rect 3033 833 3047 847
rect 3013 793 3027 807
rect 3053 793 3067 807
rect 2933 753 2947 767
rect 2993 713 3007 727
rect 2953 694 2967 708
rect 3233 933 3247 947
rect 3393 914 3407 928
rect 3453 914 3467 928
rect 3593 1653 3607 1667
rect 3753 1873 3767 1887
rect 3733 1853 3747 1867
rect 3733 1773 3747 1787
rect 3693 1753 3707 1767
rect 3873 1893 3887 1907
rect 3833 1853 3847 1867
rect 3873 1853 3887 1867
rect 3773 1833 3787 1847
rect 3793 1793 3807 1807
rect 3673 1733 3687 1747
rect 3713 1734 3727 1748
rect 3753 1734 3767 1748
rect 3653 1513 3667 1527
rect 3833 1773 3847 1787
rect 3993 1953 4007 1967
rect 3933 1893 3947 1907
rect 4013 1913 4027 1927
rect 3973 1893 3987 1907
rect 4253 2213 4267 2227
rect 4193 2173 4207 2187
rect 4193 2093 4207 2107
rect 4193 2072 4207 2086
rect 4153 2013 4167 2027
rect 4033 1873 4047 1887
rect 4013 1853 4027 1867
rect 3913 1793 3927 1807
rect 3993 1793 4007 1807
rect 3893 1753 3907 1767
rect 3933 1753 3947 1767
rect 3873 1734 3887 1748
rect 3913 1733 3927 1747
rect 3853 1692 3867 1706
rect 3893 1692 3907 1706
rect 3753 1593 3767 1607
rect 3733 1573 3747 1587
rect 3753 1553 3767 1567
rect 3673 1453 3687 1467
rect 3613 1434 3627 1448
rect 3673 1432 3687 1446
rect 3713 1434 3727 1448
rect 4033 1773 4047 1787
rect 3973 1692 3987 1706
rect 4013 1693 4027 1707
rect 4133 1973 4147 1987
rect 4153 1953 4167 1967
rect 4113 1912 4127 1926
rect 4073 1853 4087 1867
rect 4173 1853 4187 1867
rect 4153 1833 4167 1847
rect 4073 1793 4087 1807
rect 4093 1773 4107 1787
rect 4053 1733 4067 1747
rect 4333 2273 4347 2287
rect 4493 2432 4507 2446
rect 4473 2413 4487 2427
rect 4433 2353 4447 2367
rect 4393 2313 4407 2327
rect 4493 2313 4507 2327
rect 4373 2293 4387 2307
rect 4333 2212 4347 2226
rect 4313 2173 4327 2187
rect 4353 2173 4367 2187
rect 4273 2073 4287 2087
rect 4273 2033 4287 2047
rect 4453 2254 4467 2268
rect 4613 2693 4627 2707
rect 4733 2774 4747 2788
rect 4713 2732 4727 2746
rect 4753 2732 4767 2746
rect 4793 2732 4807 2746
rect 4873 2952 4887 2966
rect 4913 2953 4927 2967
rect 4873 2913 4887 2927
rect 4833 2893 4847 2907
rect 4873 2774 4887 2788
rect 4913 2773 4927 2787
rect 4833 2733 4847 2747
rect 4753 2673 4767 2687
rect 4653 2653 4667 2667
rect 4793 2653 4807 2667
rect 4773 2633 4787 2647
rect 4833 2633 4847 2647
rect 4613 2593 4627 2607
rect 4793 2593 4807 2607
rect 4833 2593 4847 2607
rect 4653 2573 4667 2587
rect 4773 2573 4787 2587
rect 4593 2533 4607 2547
rect 4633 2533 4647 2547
rect 4593 2493 4607 2507
rect 4553 2474 4567 2488
rect 4813 2573 4827 2587
rect 4753 2553 4767 2567
rect 4713 2533 4727 2547
rect 4673 2493 4687 2507
rect 4533 2433 4547 2447
rect 4573 2432 4587 2446
rect 4613 2432 4627 2446
rect 4673 2413 4687 2427
rect 4733 2432 4747 2446
rect 5033 3253 5047 3267
rect 5073 3293 5087 3307
rect 5113 3294 5127 3308
rect 5173 3294 5187 3308
rect 5233 3653 5247 3667
rect 5233 3573 5247 3587
rect 5293 3813 5307 3827
rect 5313 3833 5327 3847
rect 5353 3814 5367 3828
rect 5333 3772 5347 3786
rect 5273 3533 5287 3547
rect 5253 3514 5267 3528
rect 5293 3514 5307 3528
rect 5393 3773 5407 3787
rect 5373 3673 5387 3687
rect 5453 3992 5467 4006
rect 5493 3993 5507 4007
rect 5433 3953 5447 3967
rect 5453 3813 5467 3827
rect 5633 3993 5647 4007
rect 5593 3973 5607 3987
rect 5553 3933 5567 3947
rect 5553 3814 5567 3828
rect 5593 3814 5607 3828
rect 5693 4034 5707 4048
rect 5813 4093 5827 4107
rect 5773 4053 5787 4067
rect 5813 4034 5827 4048
rect 5753 3973 5767 3987
rect 5713 3953 5727 3967
rect 5753 3952 5767 3966
rect 5653 3853 5667 3867
rect 5693 3853 5707 3867
rect 5453 3773 5467 3787
rect 5433 3713 5447 3727
rect 5453 3653 5467 3667
rect 5353 3533 5367 3547
rect 5413 3534 5427 3548
rect 5333 3513 5347 3527
rect 5273 3472 5287 3486
rect 5513 3673 5527 3687
rect 5493 3593 5507 3607
rect 5413 3513 5427 3527
rect 5313 3373 5327 3387
rect 5213 3313 5227 3327
rect 5293 3313 5307 3327
rect 5233 3294 5247 3308
rect 5093 3253 5107 3267
rect 5093 3212 5107 3226
rect 5052 3113 5066 3127
rect 5073 3113 5087 3127
rect 4993 3033 5007 3047
rect 5073 3033 5087 3047
rect 4973 2994 4987 3008
rect 5053 3013 5067 3027
rect 5013 2952 5027 2966
rect 5053 2952 5067 2966
rect 5073 2873 5087 2887
rect 4953 2833 4967 2847
rect 5052 2833 5066 2847
rect 5073 2833 5087 2847
rect 4973 2813 4987 2827
rect 5033 2813 5047 2827
rect 5033 2773 5047 2787
rect 4953 2733 4967 2747
rect 4933 2673 4947 2687
rect 4853 2553 4867 2567
rect 4833 2513 4847 2527
rect 4893 2513 4907 2527
rect 4693 2393 4707 2407
rect 4673 2353 4687 2367
rect 4553 2253 4567 2267
rect 4613 2254 4627 2268
rect 4393 2193 4407 2207
rect 4533 2212 4547 2226
rect 4473 2193 4487 2207
rect 4393 2172 4407 2186
rect 4433 2173 4447 2187
rect 4373 2153 4387 2167
rect 4333 2033 4347 2047
rect 4313 1953 4327 1967
rect 4213 1793 4227 1807
rect 4173 1733 4187 1747
rect 4293 1912 4307 1926
rect 4293 1873 4307 1887
rect 4273 1813 4287 1827
rect 4253 1734 4267 1748
rect 4153 1713 4167 1727
rect 4093 1673 4107 1687
rect 4033 1633 4047 1647
rect 3953 1613 3967 1627
rect 3933 1593 3947 1607
rect 4073 1593 4087 1607
rect 3793 1513 3807 1527
rect 3773 1434 3787 1448
rect 3593 1392 3607 1406
rect 3633 1353 3647 1367
rect 3733 1373 3747 1387
rect 3673 1333 3687 1347
rect 3672 1293 3686 1307
rect 3693 1293 3707 1307
rect 3773 1293 3787 1307
rect 3553 1273 3567 1287
rect 3653 1273 3667 1287
rect 4033 1493 4047 1507
rect 3813 1473 3827 1487
rect 3853 1473 3867 1487
rect 3953 1473 3967 1487
rect 3893 1434 3907 1448
rect 3873 1353 3887 1367
rect 3593 1214 3607 1228
rect 3533 1153 3547 1167
rect 3573 1153 3587 1167
rect 3793 1273 3807 1287
rect 3833 1273 3847 1287
rect 3693 1253 3707 1267
rect 3773 1253 3787 1267
rect 3673 1172 3687 1186
rect 3653 1093 3667 1107
rect 3613 1073 3627 1087
rect 3553 1033 3567 1047
rect 3353 872 3367 886
rect 3273 833 3287 847
rect 3233 793 3247 807
rect 3153 713 3167 727
rect 3213 713 3227 727
rect 3073 693 3087 707
rect 3113 694 3127 708
rect 3013 652 3027 666
rect 3053 652 3067 666
rect 2973 633 2987 647
rect 3173 652 3187 666
rect 3133 633 3147 647
rect 3253 753 3267 767
rect 3253 713 3267 727
rect 3233 693 3247 707
rect 3433 872 3447 886
rect 3533 872 3547 886
rect 3433 813 3447 827
rect 3253 652 3267 666
rect 3213 593 3227 607
rect 3293 593 3307 607
rect 3073 553 3087 567
rect 2933 513 2947 527
rect 2913 394 2927 408
rect 3353 694 3367 708
rect 3393 694 3407 708
rect 3473 833 3487 847
rect 3133 453 3147 467
rect 3333 453 3347 467
rect 2973 394 2987 408
rect 3193 413 3207 427
rect 3253 413 3267 427
rect 3333 413 3347 427
rect 3133 394 3147 408
rect 3173 394 3187 408
rect 2893 333 2907 347
rect 2573 113 2587 127
rect 2493 93 2507 107
rect 2873 133 2887 147
rect 2693 93 2707 107
rect 2833 93 2847 107
rect 2993 333 3007 347
rect 3113 352 3127 366
rect 3073 333 3087 347
rect 3293 394 3307 408
rect 3193 353 3207 367
rect 3173 313 3187 327
rect 3073 293 3087 307
rect 3033 233 3047 247
rect 2993 174 3007 188
rect 3113 273 3127 287
rect 3273 253 3287 267
rect 3453 693 3467 707
rect 3413 652 3427 666
rect 3453 653 3467 667
rect 3393 413 3407 427
rect 3813 1214 3827 1228
rect 3713 1172 3727 1186
rect 4033 1453 4047 1467
rect 3993 1392 4007 1406
rect 4033 1392 4047 1406
rect 3973 1373 3987 1387
rect 3953 1333 3967 1347
rect 3973 1293 3987 1307
rect 4113 1573 4127 1587
rect 4133 1553 4147 1567
rect 4233 1692 4247 1706
rect 4193 1573 4207 1587
rect 4353 2013 4367 2027
rect 4353 1953 4367 1967
rect 4433 1973 4447 1987
rect 4373 1912 4387 1926
rect 4393 1873 4407 1887
rect 4333 1773 4347 1787
rect 4333 1734 4347 1748
rect 4373 1734 4387 1748
rect 4513 2153 4527 2167
rect 4533 2093 4547 2107
rect 4593 2212 4607 2226
rect 4633 2212 4647 2226
rect 4593 2173 4607 2187
rect 4633 2173 4647 2187
rect 4573 2153 4587 2167
rect 4553 2033 4567 2047
rect 4532 1912 4546 1926
rect 4553 1913 4567 1927
rect 4493 1853 4507 1867
rect 4433 1813 4447 1827
rect 4513 1793 4527 1807
rect 4413 1773 4427 1787
rect 4313 1692 4327 1706
rect 4333 1673 4347 1687
rect 4393 1693 4407 1707
rect 4353 1633 4367 1647
rect 4333 1613 4347 1627
rect 4293 1573 4307 1587
rect 4273 1513 4287 1527
rect 4313 1513 4327 1527
rect 4353 1453 4367 1467
rect 4093 1392 4107 1406
rect 4093 1313 4107 1327
rect 3873 1233 3887 1247
rect 3933 1233 3947 1247
rect 4033 1233 4047 1247
rect 4073 1233 4087 1247
rect 3853 1193 3867 1207
rect 3773 1033 3787 1047
rect 3713 973 3727 987
rect 3573 914 3587 928
rect 3693 914 3707 928
rect 3673 872 3687 886
rect 3613 773 3627 787
rect 3833 1133 3847 1147
rect 3913 1214 3927 1228
rect 3953 1214 3967 1228
rect 4013 1214 4027 1228
rect 3973 1133 3987 1147
rect 3873 1073 3887 1087
rect 3933 1073 3947 1087
rect 3973 1053 3987 1067
rect 3933 1033 3947 1047
rect 3853 993 3867 1007
rect 3893 993 3907 1007
rect 3833 973 3847 987
rect 3813 914 3827 928
rect 3933 914 3947 928
rect 3713 753 3727 767
rect 3633 713 3647 727
rect 3733 713 3747 727
rect 3633 692 3647 706
rect 3693 694 3707 708
rect 3793 872 3807 886
rect 3853 872 3867 886
rect 3773 753 3787 767
rect 3753 694 3767 708
rect 3573 652 3587 666
rect 3613 652 3627 666
rect 3473 613 3487 627
rect 3533 613 3547 627
rect 3613 613 3627 627
rect 3513 573 3527 587
rect 3453 394 3467 408
rect 3553 453 3567 467
rect 3493 313 3507 327
rect 3633 513 3647 527
rect 3673 633 3687 647
rect 3933 813 3947 827
rect 3913 733 3927 747
rect 3793 693 3807 707
rect 3833 694 3847 708
rect 3873 694 3887 708
rect 3913 693 3927 707
rect 3773 633 3787 647
rect 3893 652 3907 666
rect 3853 573 3867 587
rect 4133 1293 4147 1307
rect 4053 1153 4067 1167
rect 4013 993 4027 1007
rect 4313 1434 4327 1448
rect 4433 1733 4447 1747
rect 4473 1734 4487 1748
rect 4553 1733 4567 1747
rect 4413 1453 4427 1467
rect 4533 1692 4547 1706
rect 4493 1673 4507 1687
rect 4533 1553 4547 1567
rect 4753 2313 4767 2327
rect 4713 2273 4727 2287
rect 4693 2253 4707 2267
rect 4753 2213 4767 2227
rect 4733 2153 4747 2167
rect 4592 2132 4606 2146
rect 4613 2133 4627 2147
rect 4673 2133 4687 2147
rect 4633 2113 4647 2127
rect 4693 2113 4707 2127
rect 4673 2073 4687 2087
rect 4613 1973 4627 1987
rect 4633 1954 4647 1968
rect 4593 1873 4607 1887
rect 4613 1833 4627 1847
rect 4633 1793 4647 1807
rect 4593 1733 4607 1747
rect 4693 2013 4707 2027
rect 4813 2413 4827 2427
rect 4792 2353 4806 2367
rect 4813 2353 4827 2367
rect 4793 2332 4807 2346
rect 4793 2253 4807 2267
rect 4933 2473 4947 2487
rect 4913 2432 4927 2446
rect 4853 2313 4867 2327
rect 4833 2273 4847 2287
rect 5033 2733 5047 2747
rect 4993 2693 5007 2707
rect 5033 2593 5047 2607
rect 4993 2474 5007 2488
rect 4993 2413 5007 2427
rect 4993 2373 5007 2387
rect 4913 2273 4927 2287
rect 4773 2173 4787 2187
rect 4833 2212 4847 2226
rect 4953 2254 4967 2268
rect 5013 2333 5027 2347
rect 5033 2273 5047 2287
rect 4873 2173 4887 2187
rect 4793 2133 4807 2147
rect 4913 2212 4927 2226
rect 4973 2212 4987 2226
rect 5013 2212 5027 2226
rect 5033 2093 5047 2107
rect 4853 2013 4867 2027
rect 4893 2013 4907 2027
rect 4833 1993 4847 2007
rect 4773 1973 4787 1987
rect 4833 1933 4847 1947
rect 4753 1873 4767 1887
rect 4713 1853 4727 1867
rect 4673 1753 4687 1767
rect 4613 1692 4627 1706
rect 4653 1691 4667 1705
rect 4673 1673 4687 1687
rect 4453 1493 4467 1507
rect 4533 1493 4547 1507
rect 4573 1493 4587 1507
rect 4513 1473 4527 1487
rect 4293 1392 4307 1406
rect 4353 1392 4367 1406
rect 4393 1353 4407 1367
rect 4313 1333 4327 1347
rect 4413 1333 4427 1347
rect 4353 1313 4367 1327
rect 4393 1313 4407 1327
rect 4173 1253 4187 1267
rect 4233 1253 4247 1267
rect 4153 1113 4167 1127
rect 4133 1093 4147 1107
rect 4433 1273 4447 1287
rect 4233 1214 4247 1228
rect 4353 1214 4367 1228
rect 4193 1173 4207 1187
rect 4173 1053 4187 1067
rect 4253 1172 4267 1186
rect 4213 1153 4227 1167
rect 4333 1153 4347 1167
rect 4253 1053 4267 1067
rect 4413 1133 4427 1147
rect 4193 993 4207 1007
rect 4233 953 4247 967
rect 4113 933 4127 947
rect 4013 914 4027 928
rect 4053 914 4067 928
rect 4213 914 4227 928
rect 4113 893 4127 907
rect 4033 853 4047 867
rect 3973 793 3987 807
rect 4073 793 4087 807
rect 4373 1033 4387 1047
rect 4333 914 4347 928
rect 4413 1053 4427 1067
rect 4473 1213 4487 1227
rect 4653 1434 4667 1448
rect 4553 1392 4567 1406
rect 4533 1153 4547 1167
rect 4553 1133 4567 1147
rect 4473 1073 4487 1087
rect 4453 1033 4467 1047
rect 4433 933 4447 947
rect 4493 933 4507 947
rect 4193 872 4207 886
rect 4253 872 4267 886
rect 4353 872 4367 886
rect 4413 833 4427 847
rect 4313 813 4327 827
rect 4173 793 4187 807
rect 4073 753 4087 767
rect 4113 753 4127 767
rect 4153 753 4167 767
rect 3993 694 4007 708
rect 4053 693 4067 707
rect 3973 652 3987 666
rect 4013 652 4027 666
rect 4013 613 4027 627
rect 3933 533 3947 547
rect 3913 493 3927 507
rect 3693 453 3707 467
rect 3813 453 3827 467
rect 3653 394 3667 408
rect 3853 394 3867 408
rect 4153 732 4167 746
rect 4193 773 4207 787
rect 4073 652 4087 666
rect 4273 753 4287 767
rect 4353 753 4367 767
rect 4213 713 4227 727
rect 4373 733 4387 747
rect 4313 713 4327 727
rect 4353 713 4367 727
rect 4213 652 4227 666
rect 4293 652 4307 666
rect 4193 613 4207 627
rect 4133 573 4147 587
rect 4053 493 4067 507
rect 4273 493 4287 507
rect 4013 453 4027 467
rect 4053 453 4067 467
rect 4233 453 4247 467
rect 3973 413 3987 427
rect 3673 352 3687 366
rect 3833 333 3847 347
rect 3913 353 3927 367
rect 4193 433 4207 447
rect 4133 413 4147 427
rect 4093 394 4107 408
rect 3873 333 3887 347
rect 3713 313 3727 327
rect 3813 313 3827 327
rect 3853 313 3867 327
rect 3993 352 4007 366
rect 4053 352 4067 366
rect 4113 352 4127 366
rect 4133 333 4147 347
rect 3972 313 3986 327
rect 3613 293 3627 307
rect 3653 293 3667 307
rect 3953 293 3967 307
rect 4073 293 4087 307
rect 3353 273 3367 287
rect 3513 273 3527 287
rect 3333 233 3347 247
rect 3113 213 3127 227
rect 3233 213 3247 227
rect 3313 213 3327 227
rect 3393 213 3407 227
rect 3173 173 3187 187
rect 3233 174 3247 188
rect 3293 173 3307 187
rect 2933 132 2947 146
rect 3033 132 3047 146
rect 3133 132 3147 146
rect 3093 93 3107 107
rect 2153 73 2167 87
rect 2613 73 2627 87
rect 2873 73 2887 87
rect 3213 132 3227 146
rect 3353 174 3367 188
rect 3453 193 3467 207
rect 3553 174 3567 188
rect 3773 273 3787 287
rect 3753 213 3767 227
rect 3693 174 3707 188
rect 3293 73 3307 87
rect 3573 132 3587 146
rect 3713 132 3727 146
rect 3753 132 3767 146
rect 3953 253 3967 267
rect 3793 233 3807 247
rect 3913 233 3927 247
rect 3793 174 3807 188
rect 3833 174 3847 188
rect 3873 174 3887 188
rect 3953 173 3967 187
rect 4013 233 4027 247
rect 4053 173 4067 187
rect 3933 153 3947 167
rect 3813 132 3827 146
rect 3833 113 3847 127
rect 3833 73 3847 87
rect 3933 113 3947 127
rect 3993 132 4007 146
rect 4053 133 4067 147
rect 3953 93 3967 107
rect 3993 93 4007 107
rect 4033 93 4047 107
rect 4113 213 4127 227
rect 4373 693 4387 707
rect 4693 1473 4707 1487
rect 4613 1253 4627 1267
rect 4673 1253 4687 1267
rect 4733 1793 4747 1807
rect 4773 1773 4787 1787
rect 4813 1734 4827 1748
rect 4993 1993 5007 2007
rect 4873 1954 4887 1968
rect 4913 1954 4927 1968
rect 4953 1954 4967 1968
rect 4873 1893 4887 1907
rect 5153 3253 5167 3267
rect 5133 3173 5147 3187
rect 5113 3133 5127 3147
rect 5133 3073 5147 3087
rect 5173 3213 5187 3227
rect 5253 3252 5267 3266
rect 5213 3193 5227 3207
rect 5213 3153 5227 3167
rect 5193 3073 5207 3087
rect 5173 3033 5187 3047
rect 5153 3013 5167 3027
rect 5273 3053 5287 3067
rect 5373 3473 5387 3487
rect 5433 3472 5447 3486
rect 5393 3433 5407 3447
rect 5433 3413 5447 3427
rect 5533 3653 5547 3667
rect 5513 3513 5527 3527
rect 5553 3633 5567 3647
rect 5573 3613 5587 3627
rect 5573 3514 5587 3528
rect 5633 3733 5647 3747
rect 5632 3693 5646 3707
rect 5653 3693 5667 3707
rect 5673 3633 5687 3647
rect 5653 3553 5667 3567
rect 5613 3513 5627 3527
rect 5633 3514 5647 3528
rect 5513 3453 5527 3467
rect 5553 3453 5567 3467
rect 5633 3413 5647 3427
rect 5493 3373 5507 3387
rect 5373 3353 5387 3367
rect 5413 3333 5427 3347
rect 5333 3272 5347 3286
rect 5313 3252 5327 3266
rect 5213 3033 5227 3047
rect 5293 3033 5307 3047
rect 5193 2993 5207 3007
rect 5153 2952 5167 2966
rect 5173 2853 5187 2867
rect 5133 2793 5147 2807
rect 5073 2733 5087 2747
rect 5113 2732 5127 2746
rect 5153 2713 5167 2727
rect 5133 2693 5147 2707
rect 5173 2693 5187 2707
rect 5193 2653 5207 2667
rect 5113 2633 5127 2647
rect 5193 2613 5207 2627
rect 5153 2573 5167 2587
rect 5073 2474 5087 2488
rect 5113 2474 5127 2488
rect 5193 2473 5207 2487
rect 5073 2413 5087 2427
rect 5113 2353 5127 2367
rect 5173 2432 5187 2446
rect 5153 2413 5167 2427
rect 5133 2333 5147 2347
rect 5253 3013 5267 3027
rect 5353 3252 5367 3266
rect 5513 3353 5527 3367
rect 5553 3333 5567 3347
rect 5513 3293 5527 3307
rect 5593 3294 5607 3308
rect 5633 3293 5647 3307
rect 5493 3233 5507 3247
rect 5473 3193 5487 3207
rect 5573 3252 5587 3266
rect 5633 3253 5647 3267
rect 5613 3213 5627 3227
rect 5513 3173 5527 3187
rect 5473 3153 5487 3167
rect 5413 3133 5427 3147
rect 5393 3093 5407 3107
rect 5373 3053 5387 3067
rect 5233 2994 5247 3008
rect 5233 2913 5247 2927
rect 5273 2994 5287 3008
rect 5333 2994 5347 3008
rect 5333 2933 5347 2947
rect 5253 2873 5267 2887
rect 5233 2853 5247 2867
rect 5313 2893 5327 2907
rect 5273 2813 5287 2827
rect 5293 2793 5307 2807
rect 5373 2893 5387 2907
rect 5373 2793 5387 2807
rect 5353 2773 5367 2787
rect 5433 3013 5447 3027
rect 5413 2993 5427 3007
rect 5813 3893 5827 3907
rect 5973 4693 5987 4707
rect 5973 4633 5987 4647
rect 6033 5073 6047 5087
rect 6153 5093 6167 5107
rect 6133 5074 6147 5088
rect 6173 5074 6187 5088
rect 6073 5032 6087 5046
rect 6033 4993 6047 5007
rect 6113 4993 6127 5007
rect 6093 4953 6107 4967
rect 6033 4893 6047 4907
rect 6013 4853 6027 4867
rect 6053 4854 6067 4868
rect 6133 4854 6147 4868
rect 6013 4793 6027 4807
rect 6013 4753 6027 4767
rect 6013 4693 6027 4707
rect 5993 4593 6007 4607
rect 5973 4553 5987 4567
rect 6073 4793 6087 4807
rect 6113 4793 6127 4807
rect 6033 4633 6047 4647
rect 6093 4554 6107 4568
rect 5973 4513 5987 4527
rect 6053 4512 6067 4526
rect 5953 4333 5967 4347
rect 5893 4253 5907 4267
rect 5973 4293 5987 4307
rect 5953 4253 5967 4267
rect 5933 4213 5947 4227
rect 6013 4493 6027 4507
rect 6072 4453 6086 4467
rect 6093 4453 6107 4467
rect 5993 4213 6007 4227
rect 5973 4173 5987 4187
rect 5993 4153 6007 4167
rect 5953 4133 5967 4147
rect 5933 4034 5947 4048
rect 5853 3873 5867 3887
rect 5713 3693 5727 3707
rect 5693 3553 5707 3567
rect 5813 3772 5827 3786
rect 5773 3593 5787 3607
rect 5753 3514 5767 3528
rect 5673 3473 5687 3487
rect 5753 3453 5767 3467
rect 5733 3433 5747 3447
rect 5693 3393 5707 3407
rect 5733 3373 5747 3387
rect 5672 3333 5686 3347
rect 5693 3333 5707 3347
rect 5673 3293 5687 3307
rect 5713 3294 5727 3308
rect 5813 3653 5827 3667
rect 5893 3873 5907 3887
rect 5893 3833 5907 3847
rect 5873 3813 5887 3827
rect 5873 3773 5887 3787
rect 5853 3733 5867 3747
rect 5853 3633 5867 3647
rect 5812 3533 5826 3547
rect 5833 3533 5847 3547
rect 5913 3693 5927 3707
rect 5893 3653 5907 3667
rect 5893 3593 5907 3607
rect 5893 3514 5907 3528
rect 6093 4373 6107 4387
rect 6073 4353 6087 4367
rect 6053 4334 6067 4348
rect 6173 4953 6187 4967
rect 6153 4753 6167 4767
rect 6133 4713 6147 4727
rect 6193 4673 6207 4687
rect 6133 4593 6147 4607
rect 6213 4593 6227 4607
rect 6113 4353 6127 4367
rect 6173 4554 6187 4568
rect 6213 4554 6227 4568
rect 6193 4512 6207 4526
rect 6173 4473 6187 4487
rect 6153 4372 6167 4386
rect 6133 4333 6147 4347
rect 6013 4053 6027 4067
rect 5972 4033 5986 4047
rect 5993 4033 6007 4047
rect 6113 4292 6127 4306
rect 6093 4233 6107 4247
rect 6073 4053 6087 4067
rect 6133 4233 6147 4247
rect 6133 4173 6147 4187
rect 6113 4133 6127 4147
rect 6113 4093 6127 4107
rect 5993 3993 6007 4007
rect 5973 3933 5987 3947
rect 5993 3913 6007 3927
rect 6073 3973 6087 3987
rect 6073 3893 6087 3907
rect 6013 3833 6027 3847
rect 5953 3653 5967 3667
rect 6053 3813 6067 3827
rect 6093 3813 6107 3827
rect 5993 3773 6007 3787
rect 6033 3753 6047 3767
rect 5993 3713 6007 3727
rect 6093 3773 6107 3787
rect 6073 3673 6087 3687
rect 5973 3633 5987 3647
rect 5993 3553 6007 3567
rect 6033 3514 6047 3528
rect 6073 3512 6087 3526
rect 5793 3433 5807 3447
rect 5793 3353 5807 3367
rect 5773 3333 5787 3347
rect 5793 3293 5807 3307
rect 5653 3153 5667 3167
rect 5633 3113 5647 3127
rect 5553 3093 5567 3107
rect 5593 2994 5607 3008
rect 5513 2952 5527 2966
rect 5573 2952 5587 2966
rect 5453 2933 5467 2947
rect 5493 2913 5507 2927
rect 5473 2853 5487 2867
rect 5413 2793 5427 2807
rect 5453 2793 5467 2807
rect 5473 2772 5487 2786
rect 5373 2753 5387 2767
rect 5273 2732 5287 2746
rect 5353 2733 5367 2747
rect 5313 2693 5327 2707
rect 5233 2653 5247 2667
rect 5293 2513 5307 2527
rect 5253 2474 5267 2488
rect 5233 2433 5247 2447
rect 5273 2413 5287 2427
rect 5253 2373 5267 2387
rect 5233 2333 5247 2347
rect 5313 2353 5327 2367
rect 5253 2313 5267 2327
rect 5173 2273 5187 2287
rect 5213 2273 5227 2287
rect 5433 2732 5447 2746
rect 5432 2673 5446 2687
rect 5453 2673 5467 2687
rect 5373 2633 5387 2647
rect 5373 2593 5387 2607
rect 5452 2633 5466 2647
rect 5473 2633 5487 2647
rect 5433 2573 5447 2587
rect 5393 2553 5407 2567
rect 5413 2513 5427 2527
rect 5373 2473 5387 2487
rect 5453 2473 5467 2487
rect 5373 2413 5387 2427
rect 5433 2432 5447 2446
rect 5473 2433 5487 2447
rect 5393 2353 5407 2367
rect 5433 2353 5447 2367
rect 5093 2212 5107 2226
rect 5153 2213 5167 2227
rect 5313 2273 5327 2287
rect 5353 2273 5367 2287
rect 5273 2254 5287 2268
rect 5213 2212 5227 2226
rect 5253 2173 5267 2187
rect 5173 2073 5187 2087
rect 5133 2013 5147 2027
rect 5073 1954 5087 1968
rect 5053 1912 5067 1926
rect 4933 1873 4947 1887
rect 4993 1873 5007 1887
rect 5053 1853 5067 1867
rect 5113 1893 5127 1907
rect 5093 1813 5107 1827
rect 4873 1793 4887 1807
rect 4993 1773 5007 1787
rect 5033 1773 5047 1787
rect 4893 1734 4907 1748
rect 4933 1734 4947 1748
rect 4793 1692 4807 1706
rect 4853 1693 4867 1707
rect 4953 1692 4967 1706
rect 4913 1673 4927 1687
rect 4833 1434 4847 1448
rect 4733 1392 4747 1406
rect 4773 1253 4787 1267
rect 4713 1233 4727 1247
rect 4753 1233 4767 1247
rect 4673 1214 4687 1228
rect 4733 1213 4747 1227
rect 4613 1073 4627 1087
rect 4593 973 4607 987
rect 4733 1173 4747 1187
rect 4673 1113 4687 1127
rect 4713 1113 4727 1127
rect 4653 1033 4667 1047
rect 4633 973 4647 987
rect 4633 914 4647 928
rect 4473 872 4487 886
rect 4553 873 4567 887
rect 4613 872 4627 886
rect 4513 753 4527 767
rect 4493 693 4507 707
rect 4393 652 4407 666
rect 4713 1073 4727 1087
rect 4733 993 4747 1007
rect 4713 973 4727 987
rect 4973 1633 4987 1647
rect 4893 1573 4907 1587
rect 4933 1553 4947 1567
rect 5053 1734 5067 1748
rect 5093 1734 5107 1748
rect 5373 2254 5387 2268
rect 5353 2133 5367 2147
rect 5393 2113 5407 2127
rect 5233 1993 5247 2007
rect 5313 1993 5327 2007
rect 5193 1912 5207 1926
rect 5173 1853 5187 1867
rect 5153 1813 5167 1827
rect 5013 1692 5027 1706
rect 4993 1533 5007 1547
rect 5133 1673 5147 1687
rect 5113 1493 5127 1507
rect 4973 1434 4987 1448
rect 5073 1434 5087 1448
rect 5113 1434 5127 1448
rect 4893 1392 4907 1406
rect 4953 1392 4967 1406
rect 5093 1373 5107 1387
rect 4993 1353 5007 1367
rect 5073 1353 5087 1367
rect 5113 1353 5127 1367
rect 5133 1333 5147 1347
rect 5193 1833 5207 1847
rect 5173 1793 5187 1807
rect 5353 1954 5367 1968
rect 5473 2313 5487 2327
rect 5593 2893 5607 2907
rect 5613 2853 5627 2867
rect 5613 2813 5627 2827
rect 5553 2774 5567 2788
rect 5593 2774 5607 2788
rect 5733 3252 5747 3266
rect 5713 3233 5727 3247
rect 5733 3193 5747 3207
rect 5873 3472 5887 3486
rect 5933 3472 5947 3486
rect 5913 3353 5927 3367
rect 5833 3293 5847 3307
rect 5873 3294 5887 3308
rect 5813 3173 5827 3187
rect 5793 3153 5807 3167
rect 5713 3093 5727 3107
rect 5773 3093 5787 3107
rect 5693 3073 5707 3087
rect 5733 3053 5747 3067
rect 5693 3033 5707 3047
rect 5693 3012 5707 3026
rect 5673 2993 5687 3007
rect 5793 3053 5807 3067
rect 5773 2993 5787 3007
rect 5673 2953 5687 2967
rect 5753 2952 5767 2966
rect 5713 2913 5727 2927
rect 5713 2873 5727 2887
rect 5713 2852 5727 2866
rect 5793 2853 5807 2867
rect 5673 2813 5687 2827
rect 5533 2732 5547 2746
rect 5613 2713 5627 2727
rect 5573 2693 5587 2707
rect 5573 2672 5587 2686
rect 5533 2553 5547 2567
rect 5593 2653 5607 2667
rect 5573 2513 5587 2527
rect 5593 2493 5607 2507
rect 5573 2474 5587 2488
rect 5673 2774 5687 2788
rect 5753 2813 5767 2827
rect 5893 3173 5907 3187
rect 5893 3133 5907 3147
rect 5913 3113 5927 3127
rect 5853 3093 5867 3107
rect 5893 3013 5907 3027
rect 5833 2933 5847 2947
rect 5913 2952 5927 2966
rect 5873 2913 5887 2927
rect 5873 2793 5887 2807
rect 5733 2732 5747 2746
rect 5833 2774 5847 2788
rect 5913 2873 5927 2887
rect 5913 2793 5927 2807
rect 5893 2773 5907 2787
rect 5653 2693 5667 2707
rect 5653 2653 5667 2667
rect 5693 2573 5707 2587
rect 5673 2513 5687 2527
rect 5653 2493 5667 2507
rect 5593 2432 5607 2446
rect 5633 2433 5647 2447
rect 5573 2413 5587 2427
rect 5453 2273 5467 2287
rect 5493 2273 5507 2287
rect 5533 2254 5547 2268
rect 5473 2233 5487 2247
rect 5473 2133 5487 2147
rect 5453 2073 5467 2087
rect 5533 2033 5547 2047
rect 5473 2013 5487 2027
rect 5253 1873 5267 1887
rect 5233 1753 5247 1767
rect 5213 1734 5227 1748
rect 5333 1873 5347 1887
rect 5293 1833 5307 1847
rect 5393 1813 5407 1827
rect 5353 1773 5367 1787
rect 5293 1753 5307 1767
rect 5173 1693 5187 1707
rect 5493 1954 5507 1968
rect 5593 2373 5607 2387
rect 5573 2153 5587 2167
rect 5553 1993 5567 2007
rect 5613 2313 5627 2327
rect 5613 2273 5627 2287
rect 5653 2333 5667 2347
rect 5653 2312 5667 2326
rect 5693 2473 5707 2487
rect 5773 2713 5787 2727
rect 5753 2493 5767 2507
rect 5893 2733 5907 2747
rect 5853 2713 5867 2727
rect 5813 2693 5827 2707
rect 5973 3413 5987 3427
rect 6013 3393 6027 3407
rect 6013 3353 6027 3367
rect 6073 3373 6087 3387
rect 6053 3294 6067 3308
rect 5973 3193 5987 3207
rect 6033 3212 6047 3226
rect 5993 3053 6007 3067
rect 5973 3033 5987 3047
rect 6153 4153 6167 4167
rect 6233 4452 6247 4466
rect 6193 4332 6207 4346
rect 6193 4173 6207 4187
rect 6193 4093 6207 4107
rect 6213 4093 6227 4107
rect 6173 4034 6187 4048
rect 6213 4034 6227 4048
rect 6133 3953 6147 3967
rect 6153 3913 6167 3927
rect 6133 3813 6147 3827
rect 6113 3753 6127 3767
rect 6153 3793 6167 3807
rect 6213 3953 6227 3967
rect 6193 3713 6207 3727
rect 6153 3553 6167 3567
rect 6113 3513 6127 3527
rect 6193 3514 6207 3528
rect 6233 3673 6247 3687
rect 6133 3433 6147 3447
rect 6113 3413 6127 3427
rect 6193 3453 6207 3467
rect 6173 3413 6187 3427
rect 6153 3373 6167 3387
rect 6133 3294 6147 3308
rect 6193 3393 6207 3407
rect 6213 3294 6227 3308
rect 6093 3113 6107 3127
rect 6073 3093 6087 3107
rect 6033 2994 6047 3008
rect 6213 3213 6227 3227
rect 6193 3173 6207 3187
rect 6173 3033 6187 3047
rect 6093 2893 6107 2907
rect 6053 2833 6067 2847
rect 6013 2774 6027 2788
rect 6073 2774 6087 2788
rect 5933 2732 5947 2746
rect 5993 2732 6007 2746
rect 5913 2713 5927 2727
rect 6033 2713 6047 2727
rect 5893 2653 5907 2667
rect 6073 2633 6087 2647
rect 5893 2613 5907 2627
rect 5813 2493 5827 2507
rect 5713 2432 5727 2446
rect 5753 2432 5767 2446
rect 6153 2993 6167 3007
rect 6173 2952 6187 2966
rect 6213 2893 6227 2907
rect 6153 2873 6167 2887
rect 6113 2853 6127 2867
rect 6193 2853 6207 2867
rect 6133 2633 6147 2647
rect 5993 2513 6007 2527
rect 6093 2513 6107 2527
rect 5893 2474 5907 2488
rect 5833 2413 5847 2427
rect 5813 2373 5827 2387
rect 5693 2353 5707 2367
rect 5773 2353 5787 2367
rect 5673 2293 5687 2307
rect 5753 2333 5767 2347
rect 5733 2293 5747 2307
rect 5593 2073 5607 2087
rect 5733 2253 5747 2267
rect 5633 2213 5647 2227
rect 5673 2212 5687 2226
rect 5633 2173 5647 2187
rect 5613 2033 5627 2047
rect 5653 1993 5667 2007
rect 5693 1973 5707 1987
rect 5493 1893 5507 1907
rect 5473 1873 5487 1887
rect 5433 1813 5447 1827
rect 5413 1733 5427 1747
rect 5293 1692 5307 1706
rect 5333 1692 5347 1706
rect 5193 1673 5207 1687
rect 5173 1613 5187 1627
rect 5233 1573 5247 1587
rect 5253 1473 5267 1487
rect 5173 1434 5187 1448
rect 5213 1434 5227 1448
rect 5193 1373 5207 1387
rect 5173 1353 5187 1367
rect 5153 1313 5167 1327
rect 5033 1253 5047 1267
rect 4773 1173 4787 1187
rect 4813 1172 4827 1186
rect 4893 1213 4907 1227
rect 4953 1214 4967 1228
rect 5013 1213 5027 1227
rect 4793 1153 4807 1167
rect 4873 1153 4887 1167
rect 4753 913 4767 927
rect 4733 853 4747 867
rect 4753 793 4767 807
rect 4673 733 4687 747
rect 4553 694 4567 708
rect 4593 694 4607 708
rect 4653 694 4667 708
rect 4713 694 4727 708
rect 4973 1172 4987 1186
rect 4933 1153 4947 1167
rect 4893 1033 4907 1047
rect 4873 993 4887 1007
rect 4513 652 4527 666
rect 4573 652 4587 666
rect 4613 652 4627 666
rect 4493 613 4507 627
rect 4533 613 4547 627
rect 4433 593 4447 607
rect 4493 573 4507 587
rect 4373 493 4387 507
rect 4353 394 4367 408
rect 4413 394 4427 408
rect 4253 313 4267 327
rect 4313 293 4327 307
rect 4193 273 4207 287
rect 4293 273 4307 287
rect 4433 333 4447 347
rect 4313 233 4327 247
rect 4393 233 4407 247
rect 4473 233 4487 247
rect 4433 213 4447 227
rect 4153 193 4167 207
rect 4393 193 4407 207
rect 4253 174 4267 188
rect 4613 573 4627 587
rect 4793 693 4807 707
rect 4793 653 4807 667
rect 4773 633 4787 647
rect 4733 613 4747 627
rect 4653 553 4667 567
rect 4693 553 4707 567
rect 4533 533 4547 547
rect 4593 513 4607 527
rect 4633 453 4647 467
rect 4593 413 4607 427
rect 4553 394 4567 408
rect 4533 333 4547 347
rect 4593 313 4607 327
rect 4573 293 4587 307
rect 4493 213 4507 227
rect 4533 213 4547 227
rect 4573 213 4587 227
rect 4713 413 4727 427
rect 4773 393 4787 407
rect 4693 333 4707 347
rect 4953 993 4967 1007
rect 4933 913 4947 927
rect 5213 1333 5227 1347
rect 5413 1693 5427 1707
rect 5373 1593 5387 1607
rect 5333 1573 5347 1587
rect 5533 1813 5547 1827
rect 5513 1793 5527 1807
rect 5573 1954 5587 1968
rect 5613 1954 5627 1968
rect 5633 1912 5647 1926
rect 5893 2413 5907 2427
rect 5793 2333 5807 2347
rect 5833 2333 5847 2347
rect 5873 2333 5887 2347
rect 5973 2433 5987 2447
rect 5913 2353 5927 2367
rect 5893 2292 5907 2306
rect 5893 2253 5907 2267
rect 5813 2212 5827 2226
rect 5853 2193 5867 2207
rect 5773 2173 5787 2187
rect 5833 2073 5847 2087
rect 5773 2033 5787 2047
rect 5753 1973 5767 1987
rect 5753 1912 5767 1926
rect 5793 1853 5807 1867
rect 5793 1813 5807 1827
rect 5753 1773 5767 1787
rect 5553 1733 5567 1747
rect 5433 1553 5447 1567
rect 5553 1693 5567 1707
rect 5513 1593 5527 1607
rect 5493 1493 5507 1507
rect 5293 1373 5307 1387
rect 5233 1293 5247 1307
rect 5093 1214 5107 1228
rect 5153 1193 5167 1207
rect 5033 1172 5047 1186
rect 5073 1172 5087 1186
rect 5113 1113 5127 1127
rect 5153 1093 5167 1107
rect 5193 1233 5207 1247
rect 5213 1214 5227 1228
rect 5253 1214 5267 1228
rect 5313 1214 5327 1228
rect 5393 1373 5407 1387
rect 5373 1233 5387 1247
rect 5273 1172 5287 1186
rect 5253 1113 5267 1127
rect 5193 953 5207 967
rect 4973 913 4987 927
rect 5013 913 5027 927
rect 4993 872 5007 886
rect 5033 872 5047 886
rect 5073 872 5087 886
rect 4893 853 4907 867
rect 4973 853 4987 867
rect 4973 753 4987 767
rect 4933 733 4947 747
rect 4873 694 4887 708
rect 4893 652 4907 666
rect 4833 593 4847 607
rect 5153 914 5167 928
rect 5193 853 5207 867
rect 5173 813 5187 827
rect 5193 793 5207 807
rect 5173 773 5187 787
rect 5073 713 5087 727
rect 5113 713 5127 727
rect 5013 694 5027 708
rect 5133 694 5147 708
rect 4993 652 5007 666
rect 5033 652 5047 666
rect 5073 652 5087 666
rect 5113 652 5127 666
rect 5153 633 5167 647
rect 4933 473 4947 487
rect 5013 473 5027 487
rect 5053 473 5067 487
rect 5173 473 5187 487
rect 4913 433 4927 447
rect 4813 394 4827 408
rect 4873 394 4887 408
rect 4973 394 4987 408
rect 4793 352 4807 366
rect 4853 352 4867 366
rect 4913 352 4927 366
rect 4953 352 4967 366
rect 4653 313 4667 327
rect 4713 313 4727 327
rect 4633 293 4647 307
rect 4613 273 4627 287
rect 4753 253 4767 267
rect 4673 233 4687 247
rect 4713 233 4727 247
rect 4713 174 4727 188
rect 4753 173 4767 187
rect 4173 132 4187 146
rect 4273 132 4287 146
rect 4373 132 4387 146
rect 4413 132 4427 146
rect 4473 132 4487 146
rect 4513 132 4527 146
rect 4553 132 4567 146
rect 4613 132 4627 146
rect 4273 93 4287 107
rect 4133 73 4147 87
rect 4473 73 4487 87
rect 4733 132 4747 146
rect 4853 253 4867 267
rect 4793 193 4807 207
rect 4793 132 4807 146
rect 4833 132 4847 146
rect 4773 93 4787 107
rect 4873 93 4887 107
rect 5053 352 5067 366
rect 5093 352 5107 366
rect 5053 313 5067 327
rect 5133 253 5147 267
rect 4993 213 5007 227
rect 4973 193 4987 207
rect 5073 193 5087 207
rect 5333 1193 5347 1207
rect 5353 1153 5367 1167
rect 5313 1113 5327 1127
rect 5353 1073 5367 1087
rect 5313 953 5327 967
rect 5393 953 5407 967
rect 5473 1373 5487 1387
rect 5693 1753 5707 1767
rect 5733 1753 5747 1767
rect 5593 1733 5607 1747
rect 5633 1734 5647 1748
rect 5673 1734 5687 1748
rect 5712 1693 5726 1707
rect 5653 1673 5667 1687
rect 5693 1652 5707 1666
rect 5733 1692 5747 1706
rect 5593 1613 5607 1627
rect 5673 1593 5687 1607
rect 5613 1553 5627 1567
rect 5593 1453 5607 1467
rect 5653 1493 5667 1507
rect 5533 1332 5547 1346
rect 5453 1233 5467 1247
rect 5273 913 5287 927
rect 5493 1214 5507 1228
rect 5673 1433 5687 1447
rect 5553 1233 5567 1247
rect 5353 914 5367 928
rect 5273 873 5287 887
rect 5333 872 5347 886
rect 5253 773 5267 787
rect 5333 813 5347 827
rect 5273 753 5287 767
rect 5273 694 5287 708
rect 5373 773 5387 787
rect 5333 693 5347 707
rect 5433 913 5447 927
rect 5473 914 5487 928
rect 5553 1172 5567 1186
rect 5633 1392 5647 1406
rect 5733 1553 5747 1567
rect 5713 1473 5727 1487
rect 5613 1313 5627 1327
rect 5593 1172 5607 1186
rect 5593 953 5607 967
rect 5573 933 5587 947
rect 5533 913 5547 927
rect 5633 1273 5647 1287
rect 5633 1213 5647 1227
rect 6033 2474 6047 2488
rect 6013 2393 6027 2407
rect 5993 2293 6007 2307
rect 6053 2353 6067 2367
rect 6173 2373 6187 2387
rect 6093 2333 6107 2347
rect 6073 2313 6087 2327
rect 6053 2293 6067 2307
rect 5933 2253 5947 2267
rect 5973 2254 5987 2268
rect 6013 2254 6027 2268
rect 5933 2213 5947 2227
rect 5913 2053 5927 2067
rect 5993 2212 6007 2226
rect 6033 2213 6047 2227
rect 5973 2193 5987 2207
rect 5953 2033 5967 2047
rect 5933 1993 5947 2007
rect 5853 1953 5867 1967
rect 6033 2153 6047 2167
rect 6013 1993 6027 2007
rect 5933 1954 5947 1968
rect 5973 1954 5987 1968
rect 6073 2212 6087 2226
rect 6133 2293 6147 2307
rect 6113 2273 6127 2287
rect 6233 2833 6247 2847
rect 6213 2333 6227 2347
rect 6213 2293 6227 2307
rect 6113 2212 6127 2226
rect 6153 2212 6167 2226
rect 6113 2053 6127 2067
rect 6093 1953 6107 1967
rect 5833 1773 5847 1787
rect 5913 1912 5927 1926
rect 5973 1912 5987 1926
rect 6033 1912 6047 1926
rect 5893 1853 5907 1867
rect 5993 1853 6007 1867
rect 5873 1733 5887 1747
rect 5813 1692 5827 1706
rect 5873 1693 5887 1707
rect 5853 1653 5867 1667
rect 5853 1632 5867 1646
rect 5753 1513 5767 1527
rect 5733 1433 5747 1447
rect 5753 1392 5767 1406
rect 5793 1392 5807 1406
rect 5833 1393 5847 1407
rect 5753 1333 5767 1347
rect 5713 1313 5727 1327
rect 5733 1293 5747 1307
rect 5713 1253 5727 1267
rect 5733 1213 5747 1227
rect 5653 1172 5667 1186
rect 5693 1153 5707 1167
rect 5693 1073 5707 1087
rect 5633 953 5647 967
rect 5613 933 5627 947
rect 5673 933 5687 947
rect 5453 872 5467 886
rect 5433 773 5447 787
rect 5393 713 5407 727
rect 5493 713 5507 727
rect 5293 652 5307 666
rect 5333 653 5347 667
rect 5253 633 5267 647
rect 5313 513 5327 527
rect 5273 413 5287 427
rect 5333 413 5347 427
rect 5453 652 5467 666
rect 5393 593 5407 607
rect 5413 593 5427 607
rect 5633 853 5647 867
rect 5613 833 5627 847
rect 5553 773 5567 787
rect 5533 713 5547 727
rect 5513 693 5527 707
rect 5593 694 5607 708
rect 5533 652 5547 666
rect 5573 652 5587 666
rect 5533 573 5547 587
rect 5813 1313 5827 1327
rect 5773 1293 5787 1307
rect 5773 1253 5787 1267
rect 5773 1232 5787 1246
rect 5913 1773 5927 1787
rect 5953 1734 5967 1748
rect 6113 1773 6127 1787
rect 5933 1653 5947 1667
rect 6013 1692 6027 1706
rect 5973 1613 5987 1627
rect 5933 1573 5947 1587
rect 5913 1473 5927 1487
rect 5993 1553 6007 1567
rect 5953 1513 5967 1527
rect 5893 1453 5907 1467
rect 5933 1453 5947 1467
rect 5873 1433 5887 1447
rect 6073 1734 6087 1748
rect 6113 1734 6127 1748
rect 6153 1734 6167 1748
rect 6213 1952 6227 1966
rect 6193 1733 6207 1747
rect 6053 1533 6067 1547
rect 6093 1513 6107 1527
rect 6173 1692 6187 1706
rect 6153 1513 6167 1527
rect 5953 1433 5967 1447
rect 5993 1433 6007 1447
rect 6033 1434 6047 1448
rect 6073 1434 6087 1448
rect 6133 1434 6147 1448
rect 5873 1393 5887 1407
rect 5853 1293 5867 1307
rect 5833 1233 5847 1247
rect 5893 1373 5907 1387
rect 5973 1393 5987 1407
rect 5933 1333 5947 1347
rect 5913 1313 5927 1327
rect 5913 1292 5927 1306
rect 5793 1172 5807 1186
rect 5833 1153 5847 1167
rect 5833 1113 5847 1127
rect 6053 1392 6067 1406
rect 5993 1353 6007 1367
rect 5973 1273 5987 1287
rect 6073 1373 6087 1387
rect 6093 1353 6107 1367
rect 6153 1373 6167 1387
rect 6073 1233 6087 1247
rect 6133 1233 6147 1247
rect 6113 1214 6127 1228
rect 5913 1133 5927 1147
rect 5993 1172 6007 1186
rect 6032 1172 6046 1186
rect 6053 1173 6067 1187
rect 5953 1113 5967 1127
rect 5893 1053 5907 1067
rect 5753 1033 5767 1047
rect 5893 1032 5907 1046
rect 5793 973 5807 987
rect 5833 973 5847 987
rect 5713 953 5727 967
rect 5713 914 5727 928
rect 5753 914 5767 928
rect 5813 953 5827 967
rect 5693 873 5707 887
rect 5733 872 5747 886
rect 5753 853 5767 867
rect 5713 773 5727 787
rect 5933 973 5947 987
rect 5893 914 5907 928
rect 6133 1172 6147 1186
rect 6093 1133 6107 1147
rect 6093 1053 6107 1067
rect 6073 973 6087 987
rect 5973 913 5987 927
rect 6033 914 6047 928
rect 6093 913 6107 927
rect 5773 833 5787 847
rect 5773 733 5787 747
rect 5633 613 5647 627
rect 5593 593 5607 607
rect 5573 473 5587 487
rect 5513 413 5527 427
rect 5253 352 5267 366
rect 5313 353 5327 367
rect 5333 333 5347 347
rect 5373 333 5387 347
rect 5173 273 5187 287
rect 5213 273 5227 287
rect 5293 273 5307 287
rect 5153 193 5167 207
rect 5173 174 5187 188
rect 5453 333 5467 347
rect 5493 333 5507 347
rect 5413 253 5427 267
rect 5353 213 5367 227
rect 5433 213 5447 227
rect 5073 132 5087 146
rect 5113 132 5127 146
rect 5273 132 5287 146
rect 5473 193 5487 207
rect 5793 693 5807 707
rect 5693 652 5707 666
rect 5793 652 5807 666
rect 5733 573 5747 587
rect 5793 573 5807 587
rect 5653 533 5667 547
rect 5713 533 5727 547
rect 5693 493 5707 507
rect 5653 473 5667 487
rect 5673 394 5687 408
rect 5613 333 5627 347
rect 5693 353 5707 367
rect 5613 253 5627 267
rect 5573 213 5587 227
rect 5833 853 5847 867
rect 5873 853 5887 867
rect 5853 773 5867 787
rect 5913 813 5927 827
rect 5953 773 5967 787
rect 5893 753 5907 767
rect 5873 733 5887 747
rect 5933 733 5947 747
rect 5993 853 6007 867
rect 5993 773 6007 787
rect 5973 733 5987 747
rect 6093 873 6107 887
rect 6033 853 6047 867
rect 6053 813 6067 827
rect 6053 773 6067 787
rect 5932 693 5946 707
rect 5953 694 5967 708
rect 6033 713 6047 727
rect 5873 652 5887 666
rect 5913 652 5927 666
rect 5833 613 5847 627
rect 5873 613 5887 627
rect 5813 493 5827 507
rect 5853 493 5867 507
rect 5833 472 5847 486
rect 5793 433 5807 447
rect 5753 394 5767 408
rect 5793 393 5807 407
rect 5833 393 5847 407
rect 5733 353 5747 367
rect 5713 313 5727 327
rect 5693 293 5707 307
rect 5733 293 5747 307
rect 5713 253 5727 267
rect 5673 233 5687 247
rect 5653 193 5667 207
rect 5513 153 5527 167
rect 5813 333 5827 347
rect 5793 253 5807 267
rect 5773 233 5787 247
rect 5713 193 5727 207
rect 5773 193 5787 207
rect 5733 174 5747 188
rect 5793 173 5807 187
rect 5393 113 5407 127
rect 5553 113 5567 127
rect 5633 132 5647 146
rect 5673 132 5687 146
rect 5713 132 5727 146
rect 5753 132 5767 146
rect 5833 293 5847 307
rect 5833 233 5847 247
rect 5833 193 5847 207
rect 5893 453 5907 467
rect 6013 694 6027 708
rect 5973 632 5987 646
rect 6013 633 6027 647
rect 5953 613 5967 627
rect 5993 453 6007 467
rect 5973 394 5987 408
rect 5873 333 5887 347
rect 5893 233 5907 247
rect 5953 352 5967 366
rect 5933 333 5947 347
rect 5913 193 5927 207
rect 5973 313 5987 327
rect 5833 132 5847 146
rect 5873 132 5887 146
rect 5913 132 5927 146
rect 4953 93 4967 107
rect 5593 93 5607 107
rect 5813 93 5827 107
rect 6073 652 6087 666
rect 6033 573 6047 587
rect 6053 453 6067 467
rect 6113 453 6127 467
rect 6033 433 6047 447
rect 6033 393 6047 407
rect 6093 413 6107 427
rect 6133 393 6147 407
rect 6113 352 6127 366
rect 6073 313 6087 327
rect 6193 1653 6207 1667
rect 6193 1533 6207 1547
rect 6193 1392 6207 1406
rect 6193 1013 6207 1027
rect 6173 413 6187 427
rect 6153 233 6167 247
rect 6193 193 6207 207
rect 5993 132 6007 146
rect 6013 93 6027 107
rect 6233 1613 6247 1627
rect 6233 313 6247 327
rect 6213 93 6227 107
rect 3853 53 3867 67
rect 4073 53 4087 67
rect 4693 53 4707 67
rect 4913 53 4927 67
rect 5973 53 5987 67
rect 6073 53 6087 67
rect 3173 33 3187 47
rect 3373 33 3387 47
<< metal3 >>
rect 2467 6236 3853 6244
rect 627 6216 893 6224
rect 427 6196 833 6204
rect 1087 6196 1213 6204
rect 2427 6196 2753 6204
rect 3107 6196 3353 6204
rect 3367 6196 3433 6204
rect 3567 6196 4613 6204
rect 2207 6176 2793 6184
rect 4316 6176 4653 6184
rect 4316 6167 4324 6176
rect 5547 6176 5633 6184
rect 5647 6176 5753 6184
rect 507 6156 573 6164
rect 587 6156 673 6164
rect 1227 6156 1433 6164
rect 1547 6156 2153 6164
rect 2847 6156 2944 6164
rect 236 6136 313 6144
rect 236 6128 244 6136
rect 2107 6136 2313 6144
rect 2327 6136 2573 6144
rect 2587 6136 2813 6144
rect 2936 6144 2944 6156
rect 3167 6156 3313 6164
rect 3687 6156 4113 6164
rect 4167 6156 4313 6164
rect 4567 6156 4753 6164
rect 4807 6156 5013 6164
rect 5027 6156 5133 6164
rect 5207 6156 5233 6164
rect 5287 6156 5673 6164
rect 5807 6156 6193 6164
rect 2936 6136 3004 6144
rect 167 6116 233 6124
rect 116 6084 124 6114
rect 276 6084 284 6114
rect 667 6117 733 6125
rect 947 6116 1033 6124
rect 1047 6117 1133 6125
rect 116 6076 333 6084
rect 356 6064 364 6110
rect 456 6104 464 6114
rect 456 6096 484 6104
rect 476 6084 484 6096
rect 476 6076 513 6084
rect 896 6084 904 6114
rect 816 6076 1053 6084
rect 147 6056 364 6064
rect 467 6056 533 6064
rect 767 6056 773 6064
rect 816 6064 824 6076
rect 1107 6075 1153 6083
rect 1176 6084 1184 6114
rect 1287 6116 1533 6124
rect 1607 6117 1653 6125
rect 1767 6117 1793 6125
rect 1967 6116 1993 6124
rect 1167 6076 1184 6084
rect 1247 6075 1253 6083
rect 1267 6075 1273 6083
rect 1427 6075 1593 6083
rect 1687 6076 1753 6084
rect 1836 6084 1844 6114
rect 2247 6117 2273 6125
rect 2367 6116 2453 6124
rect 2507 6117 2533 6125
rect 2847 6117 2873 6125
rect 2927 6117 2973 6125
rect 1836 6076 1972 6084
rect 2007 6075 2073 6083
rect 2287 6076 2473 6084
rect 2547 6076 2593 6084
rect 2687 6076 2733 6084
rect 2827 6076 2893 6084
rect 2996 6084 3004 6136
rect 3787 6136 3813 6144
rect 3207 6117 3233 6125
rect 3327 6117 3393 6125
rect 3487 6116 3613 6124
rect 3636 6116 3713 6124
rect 3056 6104 3064 6114
rect 3636 6104 3644 6116
rect 3056 6096 3224 6104
rect 2996 6076 3033 6084
rect 3216 6084 3224 6096
rect 3496 6096 3644 6104
rect 3896 6104 3904 6114
rect 3947 6116 4013 6124
rect 4227 6116 4253 6124
rect 4527 6117 4593 6125
rect 4867 6117 4913 6125
rect 5007 6116 5093 6124
rect 5107 6116 5253 6124
rect 4696 6104 4704 6114
rect 5347 6116 5393 6124
rect 5467 6117 5493 6125
rect 5516 6116 5673 6124
rect 3896 6100 3924 6104
rect 3896 6096 3927 6100
rect 3496 6086 3504 6096
rect 3913 6087 3927 6096
rect 4576 6096 4704 6104
rect 3216 6076 3453 6084
rect 3967 6076 3993 6084
rect 4047 6076 4133 6084
rect 4187 6075 4213 6083
rect 4327 6076 4373 6084
rect 4576 6084 4584 6096
rect 4547 6076 4584 6084
rect 4607 6076 4673 6084
rect 4827 6076 4953 6084
rect 5127 6076 5193 6084
rect 5516 6086 5524 6116
rect 5847 6116 5893 6124
rect 5907 6116 5953 6124
rect 6007 6116 6053 6124
rect 6067 6116 6113 6124
rect 5287 6075 5333 6083
rect 5567 6075 5613 6083
rect 5667 6076 5813 6084
rect 5867 6076 5933 6084
rect 5947 6076 6033 6084
rect 6107 6075 6193 6083
rect 787 6056 824 6064
rect 1147 6056 1193 6064
rect 1567 6056 1613 6064
rect 1787 6056 2033 6064
rect 2947 6056 3133 6064
rect 3496 6064 3504 6072
rect 3207 6056 3504 6064
rect 3836 6064 3844 6072
rect 3836 6056 3893 6064
rect 347 6036 473 6044
rect 1947 6036 2133 6044
rect 2387 6036 2413 6044
rect 2647 6036 2773 6044
rect 2787 6036 2833 6044
rect 2847 6036 2873 6044
rect 2927 6036 2953 6044
rect 3987 6036 4313 6044
rect 4647 6036 4713 6044
rect 4727 6036 4753 6044
rect 5467 6036 5573 6044
rect 847 6016 1053 6024
rect 1307 6016 1733 6024
rect 1747 6016 1893 6024
rect 1907 6016 2333 6024
rect 3107 6016 3173 6024
rect 3407 6016 3593 6024
rect 3607 6016 4493 6024
rect 5907 6016 6213 6024
rect 327 5996 384 6004
rect 376 5984 384 5996
rect 667 5996 773 6004
rect 1607 5996 1933 6004
rect 3427 5996 3553 6004
rect 3927 5996 4073 6004
rect 4867 5996 5353 6004
rect 5367 5996 5393 6004
rect 5767 5996 5953 6004
rect 376 5976 713 5984
rect 827 5976 873 5984
rect 1956 5976 2213 5984
rect 327 5956 593 5964
rect 1347 5956 1373 5964
rect 1527 5956 1573 5964
rect 1956 5964 1964 5976
rect 2687 5976 2733 5984
rect 2747 5976 2773 5984
rect 3507 5976 3613 5984
rect 3627 5976 3853 5984
rect 3867 5976 4273 5984
rect 4287 5976 4533 5984
rect 4727 5976 4813 5984
rect 5167 5976 5253 5984
rect 5707 5976 5753 5984
rect 6007 5976 6053 5984
rect 1827 5956 1964 5964
rect 2047 5956 2693 5964
rect 2767 5956 2973 5964
rect 2987 5956 3133 5964
rect 3247 5956 3293 5964
rect 3307 5956 3653 5964
rect 3667 5956 3773 5964
rect 27 5936 93 5944
rect 187 5936 253 5944
rect 336 5936 373 5944
rect 336 5924 344 5936
rect 1187 5936 1253 5944
rect 1427 5936 1713 5944
rect 2027 5936 2124 5944
rect 276 5916 344 5924
rect 47 5896 93 5904
rect 167 5896 213 5904
rect 276 5904 284 5916
rect 607 5916 633 5924
rect 747 5916 793 5924
rect 1377 5916 1433 5924
rect 1377 5908 1385 5916
rect 1947 5916 1993 5924
rect 2116 5924 2124 5936
rect 2167 5936 2673 5944
rect 2273 5927 2287 5936
rect 2787 5936 2933 5944
rect 3187 5936 3253 5944
rect 4047 5936 4193 5944
rect 4287 5936 4333 5944
rect 4347 5936 4653 5944
rect 5567 5936 5673 5944
rect 5687 5936 5973 5944
rect 2116 5916 2233 5924
rect 2407 5916 2513 5924
rect 2636 5916 2773 5924
rect 2636 5908 2644 5916
rect 3147 5916 3393 5924
rect 4227 5916 4253 5924
rect 4407 5916 4432 5924
rect 4467 5916 4593 5924
rect 4927 5916 4993 5924
rect 5047 5916 5073 5924
rect 5207 5916 5232 5924
rect 5267 5916 5413 5924
rect 6067 5916 6153 5924
rect 267 5896 284 5904
rect 236 5876 324 5884
rect 236 5866 244 5876
rect 316 5866 324 5876
rect 27 5855 73 5863
rect 127 5855 153 5863
rect 327 5855 353 5863
rect 376 5847 384 5894
rect 447 5896 493 5904
rect 947 5896 964 5904
rect 407 5855 433 5863
rect 536 5864 544 5894
rect 536 5856 633 5864
rect 896 5864 904 5894
rect 956 5867 964 5896
rect 1147 5896 1213 5904
rect 1327 5896 1373 5904
rect 1396 5896 1533 5904
rect 767 5856 904 5864
rect 1396 5866 1404 5896
rect 1587 5897 1633 5905
rect 1707 5896 1773 5904
rect 1907 5904 1920 5907
rect 1907 5893 1924 5904
rect 2067 5897 2093 5905
rect 2207 5896 2253 5904
rect 2347 5897 2373 5905
rect 2567 5897 2593 5905
rect 2607 5897 2633 5905
rect 2707 5896 2804 5904
rect 1247 5855 1313 5863
rect 1447 5856 1653 5864
rect 1667 5856 1733 5864
rect 1916 5866 1924 5893
rect 2796 5884 2804 5896
rect 2827 5896 2933 5904
rect 3007 5897 3033 5905
rect 3447 5897 3512 5905
rect 3533 5904 3547 5913
rect 3533 5900 3573 5904
rect 3536 5896 3573 5900
rect 3747 5896 3813 5904
rect 3916 5896 4033 5904
rect 2796 5876 3353 5884
rect 2127 5856 2273 5864
rect 2287 5856 2333 5864
rect 2407 5856 2493 5864
rect 2927 5856 2953 5864
rect 3467 5855 3492 5863
rect 3916 5866 3924 5896
rect 4127 5897 4153 5905
rect 4787 5896 4813 5904
rect 5153 5904 5167 5913
rect 5127 5900 5167 5904
rect 5127 5896 5164 5900
rect 5447 5896 5473 5904
rect 5527 5896 5704 5904
rect 5696 5884 5704 5896
rect 5727 5896 5773 5904
rect 5796 5896 5813 5904
rect 5036 5876 5424 5884
rect 5696 5880 5744 5884
rect 5696 5876 5747 5880
rect 5036 5867 5044 5876
rect 3527 5856 3593 5864
rect 4187 5855 4253 5863
rect 4887 5855 4913 5863
rect 4987 5856 5033 5864
rect 5147 5855 5173 5863
rect 5416 5866 5424 5876
rect 5733 5867 5747 5876
rect 5796 5867 5804 5896
rect 5867 5896 5912 5904
rect 5933 5904 5947 5913
rect 5933 5900 5993 5904
rect 5936 5896 5993 5900
rect 5347 5855 5373 5863
rect 5487 5855 5533 5863
rect 5547 5856 5653 5864
rect 5927 5855 6013 5863
rect 6116 5864 6124 5894
rect 6027 5856 6124 5864
rect 1767 5836 2453 5844
rect 2467 5836 2533 5844
rect 2547 5836 2793 5844
rect 2847 5836 3033 5844
rect 3047 5836 3113 5844
rect 3787 5836 3873 5844
rect 3887 5836 3973 5844
rect 4667 5836 4833 5844
rect 287 5816 393 5824
rect 727 5816 873 5824
rect 1567 5816 1713 5824
rect 1727 5816 2333 5824
rect 2887 5816 2993 5824
rect 3647 5816 3684 5824
rect 2007 5796 2053 5804
rect 2067 5796 2233 5804
rect 2247 5796 3133 5804
rect 3676 5804 3684 5816
rect 3707 5816 3913 5824
rect 4227 5816 4433 5824
rect 5947 5816 6093 5824
rect 3676 5796 4293 5804
rect 5787 5796 5853 5804
rect 6067 5796 6133 5804
rect 1307 5776 1853 5784
rect 2267 5776 3173 5784
rect 3667 5776 3893 5784
rect 4327 5776 4733 5784
rect 4747 5776 5253 5784
rect 5587 5776 5693 5784
rect 5707 5776 5793 5784
rect 587 5756 973 5764
rect 1167 5756 1273 5764
rect 1287 5756 3413 5764
rect 3567 5756 3773 5764
rect 4316 5764 4324 5773
rect 3947 5756 4324 5764
rect 5407 5756 5873 5764
rect 5887 5756 6193 5764
rect 567 5736 753 5744
rect 767 5736 813 5744
rect 1327 5736 2913 5744
rect 3187 5736 3664 5744
rect 507 5716 693 5724
rect 907 5716 1173 5724
rect 1527 5716 1613 5724
rect 1627 5716 1753 5724
rect 2527 5716 3153 5724
rect 3167 5716 3633 5724
rect 3656 5724 3664 5736
rect 3927 5736 4833 5744
rect 4847 5736 5233 5744
rect 5627 5736 5813 5744
rect 3656 5716 3773 5724
rect 3827 5716 4013 5724
rect 4307 5716 4733 5724
rect 4747 5716 5273 5724
rect 5287 5716 5353 5724
rect 1047 5696 1653 5704
rect 2516 5704 2524 5713
rect 2247 5696 2524 5704
rect 2867 5696 3033 5704
rect 3047 5696 3933 5704
rect 5567 5696 5913 5704
rect 1967 5676 2093 5684
rect 3087 5676 3433 5684
rect 3447 5676 3753 5684
rect 3767 5676 3953 5684
rect 4087 5676 5453 5684
rect 47 5656 393 5664
rect 987 5656 1193 5664
rect 1507 5656 1553 5664
rect 1767 5656 1833 5664
rect 2827 5656 3553 5664
rect 3667 5656 3752 5664
rect 3787 5656 3933 5664
rect 4027 5656 4113 5664
rect 4127 5656 4253 5664
rect 4787 5656 4933 5664
rect 4947 5656 5413 5664
rect 5527 5656 6093 5664
rect 387 5636 533 5644
rect 547 5636 773 5644
rect 967 5636 993 5644
rect 1367 5636 2073 5644
rect 2347 5636 2553 5644
rect 2987 5636 3173 5644
rect 3687 5636 3773 5644
rect 3827 5636 3873 5644
rect 4407 5636 4453 5644
rect 4707 5636 4813 5644
rect 5847 5636 5953 5644
rect 5967 5636 5973 5644
rect 5987 5636 6033 5644
rect 976 5616 1264 5624
rect 287 5597 313 5605
rect 647 5597 673 5605
rect 27 5555 93 5563
rect 116 5547 124 5593
rect 156 5567 164 5593
rect 496 5567 504 5593
rect 576 5584 584 5594
rect 716 5584 724 5594
rect 847 5596 873 5604
rect 976 5604 984 5616
rect 967 5596 984 5604
rect 1007 5597 1053 5605
rect 576 5580 604 5584
rect 716 5580 744 5584
rect 576 5576 607 5580
rect 716 5576 747 5580
rect 593 5567 607 5576
rect 207 5555 253 5563
rect 733 5567 747 5576
rect 796 5567 804 5593
rect 916 5564 924 5594
rect 956 5564 964 5594
rect 1207 5596 1233 5604
rect 1256 5604 1264 5616
rect 1847 5616 1893 5624
rect 1907 5616 2313 5624
rect 2647 5616 2693 5624
rect 3767 5616 3833 5624
rect 4227 5616 4273 5624
rect 5087 5616 5193 5624
rect 5927 5616 6213 5624
rect 1256 5596 1344 5604
rect 1187 5576 1313 5584
rect 867 5556 924 5564
rect 936 5556 964 5564
rect 1336 5564 1344 5596
rect 1407 5597 1473 5605
rect 1707 5596 1813 5604
rect 1656 5584 1664 5594
rect 1927 5597 2093 5605
rect 2367 5597 2413 5605
rect 2516 5596 2593 5604
rect 1853 5584 1867 5593
rect 1656 5576 1684 5584
rect 1336 5556 1373 5564
rect 936 5547 944 5556
rect 1487 5556 1533 5564
rect 1676 5564 1684 5576
rect 1796 5580 1867 5584
rect 1796 5576 1864 5580
rect 1796 5566 1804 5576
rect 2287 5576 2364 5584
rect 1676 5556 1764 5564
rect 347 5536 553 5544
rect 727 5536 753 5544
rect 927 5536 944 5547
rect 927 5533 940 5536
rect 1047 5536 1173 5544
rect 1587 5536 1733 5544
rect 1756 5544 1764 5556
rect 2047 5555 2213 5563
rect 2356 5564 2364 5576
rect 2356 5556 2373 5564
rect 2516 5566 2524 5596
rect 2727 5597 2773 5605
rect 3127 5597 3173 5605
rect 3287 5597 3313 5605
rect 3367 5596 3493 5604
rect 3516 5596 3593 5604
rect 3276 5584 3284 5594
rect 2896 5576 3284 5584
rect 2896 5566 2904 5576
rect 2427 5556 2473 5564
rect 2627 5555 2733 5563
rect 2947 5555 2973 5563
rect 3067 5556 3112 5564
rect 3147 5556 3193 5564
rect 3516 5566 3524 5596
rect 3856 5596 3893 5604
rect 3636 5567 3644 5593
rect 3696 5567 3704 5594
rect 3307 5556 3333 5564
rect 3687 5556 3704 5567
rect 3736 5567 3744 5594
rect 3736 5556 3753 5567
rect 3687 5553 3700 5556
rect 3740 5553 3753 5556
rect 3856 5566 3864 5596
rect 3947 5597 3973 5605
rect 4167 5597 4193 5605
rect 4427 5596 4513 5604
rect 4567 5597 4633 5605
rect 4827 5596 4873 5604
rect 4056 5564 4064 5593
rect 4256 5584 4264 5594
rect 4987 5597 5033 5605
rect 5127 5596 5173 5604
rect 5296 5596 5313 5604
rect 4256 5576 4384 5584
rect 4376 5566 4384 5576
rect 5296 5584 5304 5596
rect 5627 5596 5773 5604
rect 5147 5576 5304 5584
rect 4056 5556 4133 5564
rect 4407 5556 4533 5564
rect 4667 5556 4773 5564
rect 4887 5555 4913 5563
rect 5067 5555 5113 5563
rect 5347 5555 5393 5563
rect 5507 5555 5553 5563
rect 5727 5555 5753 5563
rect 5947 5555 5993 5563
rect 1756 5536 1953 5544
rect 2707 5536 2793 5544
rect 3007 5536 3033 5544
rect 3667 5536 3713 5544
rect 4167 5536 4333 5544
rect 147 5516 173 5524
rect 427 5516 533 5524
rect 667 5516 872 5524
rect 907 5516 973 5524
rect 1027 5516 1253 5524
rect 1567 5516 1753 5524
rect 1767 5520 1963 5524
rect 1767 5516 1967 5520
rect 656 5504 664 5513
rect 1953 5507 1967 5516
rect 3167 5516 3233 5524
rect 3367 5516 3433 5524
rect 3487 5516 3693 5524
rect 3807 5516 3893 5524
rect 4207 5516 4393 5524
rect 4487 5516 4653 5524
rect 4707 5516 4853 5524
rect 5267 5516 5413 5524
rect 5607 5516 5693 5524
rect 5907 5516 6193 5524
rect 387 5496 664 5504
rect 887 5496 1673 5504
rect 1847 5496 1913 5504
rect 1966 5500 1967 5507
rect 1987 5496 2253 5504
rect 2567 5496 2713 5504
rect 3767 5496 3993 5504
rect 4387 5496 4433 5504
rect 4607 5496 4973 5504
rect 4987 5496 5193 5504
rect 5247 5496 5433 5504
rect 5567 5496 5793 5504
rect 327 5476 393 5484
rect 847 5476 1133 5484
rect 1607 5476 1993 5484
rect 2527 5476 2753 5484
rect 2947 5476 3153 5484
rect 4647 5476 4673 5484
rect 5387 5476 5453 5484
rect 5467 5476 5513 5484
rect 5887 5476 6133 5484
rect 67 5456 473 5464
rect 487 5456 1113 5464
rect 1807 5456 1873 5464
rect 1927 5456 1973 5464
rect 2847 5456 3252 5464
rect 3287 5456 3493 5464
rect 3507 5456 3672 5464
rect 3707 5456 4013 5464
rect 4027 5456 4053 5464
rect 4067 5456 4153 5464
rect 4207 5456 4273 5464
rect 4287 5456 4613 5464
rect 5127 5456 5713 5464
rect 727 5436 933 5444
rect 1296 5436 1373 5444
rect 1296 5427 1304 5436
rect 1867 5436 1893 5444
rect 2047 5436 2493 5444
rect 2987 5436 3393 5444
rect 3827 5436 4173 5444
rect 4807 5436 4893 5444
rect 5027 5436 5233 5444
rect 5327 5436 5653 5444
rect 227 5416 433 5424
rect 947 5416 1293 5424
rect 1467 5416 1493 5424
rect 1516 5416 1593 5424
rect 140 5404 153 5407
rect 136 5394 153 5404
rect 136 5393 160 5394
rect 567 5396 793 5404
rect 116 5344 124 5374
rect 136 5346 144 5393
rect 167 5376 273 5384
rect 407 5376 433 5384
rect 616 5376 653 5384
rect 616 5347 624 5376
rect 87 5336 124 5344
rect 267 5335 332 5343
rect 427 5336 533 5344
rect 676 5346 684 5396
rect 836 5396 913 5404
rect 836 5384 844 5396
rect 1516 5404 1524 5416
rect 1687 5416 1753 5424
rect 1916 5416 2173 5424
rect 1540 5404 1553 5407
rect 1327 5396 1524 5404
rect 1536 5393 1553 5404
rect 1916 5404 1924 5416
rect 2587 5416 2653 5424
rect 3267 5416 3473 5424
rect 3547 5416 3733 5424
rect 4027 5416 4093 5424
rect 4507 5416 4693 5424
rect 5707 5416 6303 5424
rect 1696 5396 1924 5404
rect 816 5376 844 5384
rect 816 5346 824 5376
rect 1007 5377 1053 5385
rect 1107 5377 1233 5385
rect 1387 5384 1400 5387
rect 1387 5373 1404 5384
rect 1536 5384 1544 5393
rect 1427 5376 1544 5384
rect 1696 5384 1704 5396
rect 2027 5396 2093 5404
rect 2867 5396 2893 5404
rect 3587 5396 3613 5404
rect 3927 5396 3973 5404
rect 4427 5396 4453 5404
rect 4867 5396 5053 5404
rect 5527 5396 5612 5404
rect 5987 5396 6033 5404
rect 6087 5396 6153 5404
rect 1607 5376 1704 5384
rect 1396 5364 1404 5373
rect 1596 5364 1604 5374
rect 1396 5356 1584 5364
rect 1596 5356 1644 5364
rect 727 5335 773 5343
rect 927 5336 1033 5344
rect 1087 5335 1153 5343
rect 1576 5346 1584 5356
rect 1267 5336 1293 5344
rect 1367 5335 1393 5343
rect 1636 5344 1644 5356
rect 1636 5336 1693 5344
rect 1616 5324 1624 5332
rect 1507 5316 1624 5324
rect 1636 5316 1673 5324
rect 307 5296 593 5304
rect 647 5296 693 5304
rect 1227 5296 1433 5304
rect 1636 5304 1644 5316
rect 1716 5324 1724 5374
rect 1947 5377 1973 5385
rect 2207 5376 2273 5384
rect 1716 5316 1793 5324
rect 1856 5324 1864 5373
rect 1976 5364 1984 5374
rect 2387 5377 2433 5385
rect 2476 5376 2653 5384
rect 1976 5356 2224 5364
rect 2216 5346 2224 5356
rect 1927 5336 2173 5344
rect 2287 5335 2313 5343
rect 2336 5344 2344 5374
rect 2336 5336 2413 5344
rect 2476 5346 2484 5376
rect 2727 5376 2773 5384
rect 2787 5377 2833 5385
rect 3107 5376 3173 5384
rect 2607 5335 2633 5343
rect 2727 5336 2773 5344
rect 2867 5336 2953 5344
rect 3216 5344 3224 5393
rect 3287 5377 3333 5385
rect 3347 5376 3573 5384
rect 3687 5377 3853 5385
rect 3867 5376 3893 5384
rect 4087 5376 4133 5384
rect 4147 5376 4273 5384
rect 4327 5376 4533 5384
rect 4547 5376 4584 5384
rect 4576 5347 4584 5376
rect 4627 5376 4713 5384
rect 5007 5376 5193 5384
rect 5298 5376 5333 5384
rect 3216 5336 3253 5344
rect 3536 5336 3593 5344
rect 1856 5316 1893 5324
rect 2527 5316 2573 5324
rect 3127 5316 3153 5324
rect 3227 5316 3433 5324
rect 1547 5296 1644 5304
rect 2007 5296 2193 5304
rect 2576 5304 2584 5313
rect 2576 5296 2673 5304
rect 2807 5296 2932 5304
rect 2967 5296 3073 5304
rect 3216 5304 3224 5313
rect 3536 5304 3544 5336
rect 3667 5335 3753 5343
rect 3847 5336 3913 5344
rect 3967 5335 4073 5343
rect 4167 5335 4193 5343
rect 4207 5336 4333 5344
rect 4627 5335 4653 5343
rect 4767 5335 4853 5343
rect 4867 5336 4913 5344
rect 4247 5316 4293 5324
rect 4427 5316 4513 5324
rect 4987 5316 5173 5324
rect 5298 5324 5306 5376
rect 5427 5377 5473 5385
rect 5356 5356 5433 5364
rect 5356 5346 5364 5356
rect 5476 5344 5484 5374
rect 5407 5336 5484 5344
rect 5636 5346 5644 5393
rect 5727 5376 5753 5384
rect 5807 5377 5853 5385
rect 5867 5376 5933 5384
rect 5676 5347 5684 5373
rect 5996 5347 6004 5373
rect 5547 5336 5633 5344
rect 5787 5336 5833 5344
rect 6027 5335 6093 5343
rect 5187 5316 5306 5324
rect 5447 5316 5692 5324
rect 5727 5316 5873 5324
rect 3187 5296 3224 5304
rect 3516 5296 3544 5304
rect 67 5276 193 5284
rect 507 5276 713 5284
rect 1807 5276 1833 5284
rect 1887 5276 2072 5284
rect 2107 5276 2453 5284
rect 2887 5276 2913 5284
rect 2927 5276 2993 5284
rect 3207 5276 3473 5284
rect 1307 5256 1504 5264
rect 767 5236 973 5244
rect 1387 5236 1453 5244
rect 1496 5244 1504 5256
rect 1967 5256 2033 5264
rect 2127 5256 2353 5264
rect 2487 5256 3153 5264
rect 3407 5256 3453 5264
rect 3516 5264 3524 5296
rect 3767 5296 3993 5304
rect 4667 5296 4693 5304
rect 4927 5296 5033 5304
rect 5627 5296 6033 5304
rect 3607 5276 3653 5284
rect 3987 5276 4113 5284
rect 4267 5276 4373 5284
rect 4387 5276 4553 5284
rect 4627 5276 4773 5284
rect 4907 5276 5093 5284
rect 5107 5276 5133 5284
rect 5227 5276 5492 5284
rect 5527 5284 5540 5287
rect 5527 5273 5544 5284
rect 5687 5276 5953 5284
rect 3516 5260 3544 5264
rect 3516 5256 3547 5260
rect 3533 5247 3547 5256
rect 3707 5256 3833 5264
rect 4147 5256 4333 5264
rect 4556 5264 4564 5273
rect 5536 5264 5544 5273
rect 4556 5256 5094 5264
rect 5536 5256 5773 5264
rect 1496 5236 1733 5244
rect 1787 5236 2093 5244
rect 2467 5236 2573 5244
rect 2787 5236 2873 5244
rect 2947 5236 3113 5244
rect 3127 5236 3313 5244
rect 3447 5236 3473 5244
rect 507 5216 873 5224
rect 976 5224 984 5233
rect 3667 5236 3713 5244
rect 3907 5236 4413 5244
rect 4747 5236 4933 5244
rect 976 5216 1672 5224
rect 1707 5216 1953 5224
rect 1967 5216 2433 5224
rect 2507 5216 2793 5224
rect 2847 5216 3333 5224
rect 3347 5216 3733 5224
rect 3807 5216 4133 5224
rect 4527 5216 4713 5224
rect 5086 5224 5094 5256
rect 5167 5236 5393 5244
rect 5467 5236 5813 5244
rect 5827 5236 5913 5244
rect 5086 5216 5433 5224
rect 1007 5196 1073 5204
rect 1147 5196 1533 5204
rect 2067 5196 2172 5204
rect 2207 5196 2473 5204
rect 2527 5196 2653 5204
rect 3507 5196 3713 5204
rect 3947 5196 4433 5204
rect 5067 5196 5453 5204
rect 5607 5196 5733 5204
rect 107 5176 173 5184
rect 187 5176 613 5184
rect 2076 5176 2113 5184
rect 547 5156 573 5164
rect 1047 5156 1293 5164
rect 1447 5156 1513 5164
rect 2076 5164 2084 5176
rect 2547 5176 2873 5184
rect 3076 5176 3173 5184
rect 2007 5156 2084 5164
rect 2167 5156 2493 5164
rect 3076 5164 3084 5176
rect 3227 5176 3353 5184
rect 3367 5176 3433 5184
rect 3527 5176 3553 5184
rect 4187 5176 4213 5184
rect 4647 5176 4753 5184
rect 4807 5176 4993 5184
rect 5327 5176 5513 5184
rect 5847 5176 6113 5184
rect 2587 5156 3084 5164
rect 3467 5156 3533 5164
rect 3967 5156 4253 5164
rect 4407 5156 4513 5164
rect 4967 5156 5113 5164
rect 5287 5156 5573 5164
rect 5947 5156 5993 5164
rect 6007 5156 6093 5164
rect 607 5136 973 5144
rect 1056 5136 1213 5144
rect 547 5116 653 5124
rect 847 5116 953 5124
rect 1056 5124 1064 5136
rect 1467 5136 1693 5144
rect 3007 5136 3133 5144
rect 3207 5136 3393 5144
rect 3447 5136 3593 5144
rect 3747 5136 4193 5144
rect 4307 5136 4544 5144
rect 4536 5127 4544 5136
rect 4847 5136 5152 5144
rect 5187 5136 5413 5144
rect 1027 5116 1064 5124
rect 1247 5116 1424 5124
rect 1416 5104 1424 5116
rect 1596 5116 1753 5124
rect 1416 5096 1444 5104
rect 147 5076 233 5084
rect 327 5077 353 5085
rect 76 5044 84 5073
rect 276 5064 284 5074
rect 196 5060 284 5064
rect 193 5056 284 5060
rect 193 5047 207 5056
rect 76 5036 153 5044
rect 616 5047 624 5074
rect 687 5076 713 5084
rect 467 5036 553 5044
rect 616 5036 633 5047
rect 620 5033 633 5036
rect 735 5027 743 5093
rect 756 5046 764 5093
rect 876 5047 884 5074
rect 767 5036 844 5044
rect 67 5016 133 5024
rect 836 5024 844 5036
rect 867 5036 884 5047
rect 916 5044 924 5074
rect 1147 5076 1173 5084
rect 1227 5076 1333 5084
rect 916 5036 953 5044
rect 867 5033 880 5036
rect 1067 5035 1133 5043
rect 1207 5035 1233 5043
rect 1396 5044 1404 5074
rect 1436 5064 1444 5096
rect 1507 5077 1533 5085
rect 1436 5056 1564 5064
rect 1456 5046 1464 5056
rect 1556 5046 1564 5056
rect 1596 5046 1604 5116
rect 1767 5116 2093 5124
rect 2167 5116 2333 5124
rect 2427 5116 2584 5124
rect 2576 5107 2584 5116
rect 2827 5116 2973 5124
rect 2987 5116 3053 5124
rect 3347 5116 3373 5124
rect 3487 5116 3613 5124
rect 3787 5116 3893 5124
rect 4107 5116 4193 5124
rect 4387 5116 4524 5124
rect 2587 5096 2833 5104
rect 3407 5096 3633 5104
rect 3647 5096 3793 5104
rect 3816 5096 3973 5104
rect 1827 5077 1853 5085
rect 1907 5076 1933 5084
rect 1673 5064 1687 5073
rect 1673 5060 1704 5064
rect 1676 5056 1704 5060
rect 1696 5046 1704 5056
rect 1327 5036 1404 5044
rect 1716 5044 1724 5074
rect 2033 5084 2047 5093
rect 2033 5080 2073 5084
rect 2036 5076 2073 5080
rect 2207 5077 2233 5085
rect 2387 5076 2393 5084
rect 2407 5076 2453 5084
rect 2607 5084 2620 5087
rect 2607 5073 2624 5084
rect 2907 5077 2933 5085
rect 3007 5076 3033 5084
rect 3247 5077 3293 5085
rect 1716 5036 1833 5044
rect 1967 5035 2033 5043
rect 2107 5036 2173 5044
rect 2253 5044 2267 5053
rect 2316 5056 2584 5064
rect 2316 5046 2324 5056
rect 2227 5040 2267 5044
rect 2227 5036 2264 5040
rect 2527 5035 2553 5043
rect 2576 5046 2584 5056
rect 2567 5035 2573 5043
rect 2616 5044 2624 5073
rect 2616 5036 2633 5044
rect 2687 5036 2793 5044
rect 2847 5035 2893 5043
rect 3196 5027 3204 5074
rect 3307 5036 3373 5044
rect 3496 5044 3504 5074
rect 3816 5084 3824 5096
rect 4287 5096 4313 5104
rect 4516 5104 4524 5116
rect 4547 5116 4813 5124
rect 5227 5116 5533 5124
rect 5667 5116 6013 5124
rect 4516 5096 4573 5104
rect 4856 5096 4973 5104
rect 4856 5088 4864 5096
rect 5047 5096 5113 5104
rect 5647 5104 5660 5107
rect 5647 5093 5664 5104
rect 6167 5096 6243 5104
rect 3687 5076 3824 5084
rect 4087 5077 4133 5085
rect 3653 5064 3667 5073
rect 3653 5056 3727 5064
rect 3713 5047 3727 5056
rect 3496 5036 3613 5044
rect 3936 5044 3944 5073
rect 4216 5064 4224 5074
rect 4327 5077 4373 5085
rect 4747 5076 4764 5084
rect 4187 5056 4453 5064
rect 4756 5047 4764 5076
rect 4907 5077 4933 5085
rect 5367 5076 5384 5084
rect 3867 5036 3944 5044
rect 3987 5036 4113 5044
rect 4567 5036 4613 5044
rect 4856 5027 4864 5074
rect 5196 5056 5273 5064
rect 4947 5036 5033 5044
rect 5196 5046 5204 5056
rect 5287 5056 5344 5064
rect 5336 5046 5344 5056
rect 5087 5036 5153 5044
rect 5376 5044 5384 5076
rect 5396 5064 5404 5074
rect 5447 5076 5533 5084
rect 5656 5084 5664 5093
rect 5656 5076 5704 5084
rect 5616 5064 5624 5073
rect 5396 5056 5444 5064
rect 5616 5056 5664 5064
rect 5376 5036 5413 5044
rect 5436 5044 5444 5056
rect 5436 5036 5513 5044
rect 5527 5036 5633 5044
rect 5656 5044 5664 5056
rect 5696 5044 5704 5076
rect 5747 5077 5793 5085
rect 5987 5076 6033 5084
rect 6147 5077 6173 5085
rect 5656 5036 5684 5044
rect 5696 5036 5773 5044
rect 836 5016 913 5024
rect 1387 5016 1413 5024
rect 1767 5016 1793 5024
rect 2887 5016 2953 5024
rect 3327 5016 3433 5024
rect 3827 5016 3953 5024
rect 4007 5016 4032 5024
rect 4067 5016 4393 5024
rect 4516 5016 4633 5024
rect 667 4996 773 5004
rect 827 4996 913 5004
rect 1327 4996 1493 5004
rect 1507 4996 1713 5004
rect 2047 4996 2353 5004
rect 2467 4996 2713 5004
rect 3027 4996 3473 5004
rect 4036 5004 4044 5013
rect 4516 5004 4524 5016
rect 5367 5016 5473 5024
rect 5676 5024 5684 5036
rect 5827 5036 6073 5044
rect 5676 5016 5784 5024
rect 4036 4996 4524 5004
rect 4727 4996 4773 5004
rect 4887 4996 4953 5004
rect 5127 4996 5613 5004
rect 5676 4996 5753 5004
rect 5676 4987 5684 4996
rect 5776 5004 5784 5016
rect 5776 4996 5832 5004
rect 5867 4996 5933 5004
rect 6047 4996 6113 5004
rect 187 4976 253 4984
rect 367 4976 772 4984
rect 807 4976 953 4984
rect 967 4976 1373 4984
rect 1747 4976 1973 4984
rect 3387 4976 3473 4984
rect 3487 4976 3673 4984
rect 3867 4976 3953 4984
rect 4127 4976 4193 4984
rect 4407 4976 4513 4984
rect 4567 4976 5093 4984
rect 5267 4976 5673 4984
rect 447 4956 473 4964
rect 667 4956 733 4964
rect 887 4956 1793 4964
rect 2487 4956 2733 4964
rect 2747 4956 2924 4964
rect 876 4944 884 4953
rect 647 4936 884 4944
rect 927 4936 1013 4944
rect 1787 4936 2072 4944
rect 2107 4936 2193 4944
rect 2216 4936 2513 4944
rect 487 4916 553 4924
rect 927 4916 973 4924
rect 2216 4924 2224 4936
rect 2916 4944 2924 4956
rect 2996 4956 3073 4964
rect 2996 4944 3004 4956
rect 3367 4956 3653 4964
rect 3987 4956 4313 4964
rect 4707 4956 4813 4964
rect 4827 4956 5073 4964
rect 5287 4956 5373 4964
rect 5547 4956 5613 4964
rect 5627 4956 5893 4964
rect 5967 4956 6093 4964
rect 6107 4956 6173 4964
rect 2916 4936 3004 4944
rect 3047 4936 3213 4944
rect 3547 4936 3753 4944
rect 4347 4936 4553 4944
rect 4607 4936 4993 4944
rect 5107 4936 5233 4944
rect 5647 4936 5713 4944
rect 5887 4936 5924 4944
rect 1427 4916 2224 4924
rect 2427 4916 2533 4924
rect 3347 4916 3513 4924
rect 3927 4916 4053 4924
rect 4147 4916 4173 4924
rect 5127 4916 5213 4924
rect 5307 4913 5313 4927
rect 5767 4916 5853 4924
rect 5916 4924 5924 4936
rect 5916 4916 5993 4924
rect 207 4896 413 4904
rect 427 4896 573 4904
rect 787 4896 813 4904
rect 936 4896 993 4904
rect 936 4884 944 4896
rect 1087 4896 1113 4904
rect 1127 4896 1173 4904
rect 1507 4896 1653 4904
rect 1807 4896 2373 4904
rect 2396 4896 2673 4904
rect 567 4876 744 4884
rect 736 4868 744 4876
rect 876 4876 944 4884
rect 956 4876 1053 4884
rect 47 4857 73 4865
rect 147 4856 213 4864
rect 367 4857 393 4865
rect 747 4856 833 4864
rect 536 4824 544 4853
rect 876 4844 884 4876
rect 956 4868 964 4876
rect 1427 4876 1584 4884
rect 1107 4856 1133 4864
rect 1307 4857 1353 4865
rect 1487 4856 1553 4864
rect 796 4840 884 4844
rect 793 4836 884 4840
rect 793 4827 807 4836
rect 467 4816 544 4824
rect 567 4815 613 4823
rect 687 4815 753 4823
rect 896 4824 904 4853
rect 1576 4826 1584 4876
rect 1707 4876 1773 4884
rect 1887 4876 1924 4884
rect 1607 4856 1633 4864
rect 1647 4856 1853 4864
rect 1916 4864 1924 4876
rect 2396 4884 2404 4896
rect 2907 4896 2993 4904
rect 3067 4896 3133 4904
rect 3356 4896 3413 4904
rect 2247 4876 2404 4884
rect 2547 4876 2753 4884
rect 1916 4856 1993 4864
rect 2007 4857 2033 4865
rect 2116 4844 2124 4873
rect 2447 4856 2504 4864
rect 2116 4836 2164 4844
rect 2156 4826 2164 4836
rect 2496 4826 2504 4856
rect 2527 4856 2544 4864
rect 836 4816 904 4824
rect 836 4807 844 4816
rect 1407 4815 1473 4823
rect 1687 4815 1773 4823
rect 2067 4815 2113 4823
rect 2167 4815 2293 4823
rect 2536 4807 2544 4856
rect 2627 4856 2813 4864
rect 2967 4856 3033 4864
rect 3107 4857 3173 4865
rect 3356 4864 3364 4896
rect 3867 4896 4072 4904
rect 4107 4896 4173 4904
rect 4527 4896 4673 4904
rect 4907 4896 5093 4904
rect 4087 4876 4113 4884
rect 4167 4876 4313 4884
rect 4516 4884 4524 4893
rect 5247 4896 5332 4904
rect 5367 4896 5413 4904
rect 5487 4896 5513 4904
rect 5527 4896 5673 4904
rect 5896 4896 6033 4904
rect 4376 4876 4524 4884
rect 3267 4856 3373 4864
rect 3427 4856 3553 4864
rect 3567 4857 3613 4865
rect 3636 4856 3653 4864
rect 2707 4816 2793 4824
rect 2916 4824 2924 4853
rect 3636 4844 3644 4856
rect 3787 4857 3813 4865
rect 4016 4844 4024 4854
rect 3596 4840 3644 4844
rect 2896 4816 2933 4824
rect 87 4796 153 4804
rect 727 4796 773 4804
rect 827 4793 844 4807
rect 1147 4796 1273 4804
rect 1547 4796 1613 4804
rect 1627 4796 1793 4804
rect 2536 4796 2553 4807
rect 2540 4793 2553 4796
rect 2896 4804 2904 4816
rect 2987 4816 3073 4824
rect 3193 4824 3207 4833
rect 3593 4836 3644 4840
rect 3976 4836 4024 4844
rect 3593 4827 3607 4836
rect 3116 4820 3207 4824
rect 3116 4816 3204 4820
rect 2647 4796 2904 4804
rect 3116 4804 3124 4816
rect 3327 4816 3393 4824
rect 3487 4815 3533 4823
rect 3687 4816 3813 4824
rect 3976 4824 3984 4836
rect 4376 4826 4384 4876
rect 4747 4876 4793 4884
rect 5167 4876 5393 4884
rect 5407 4876 5653 4884
rect 4407 4856 4444 4864
rect 4436 4827 4444 4856
rect 4613 4864 4627 4873
rect 4567 4856 4604 4864
rect 4613 4860 4653 4864
rect 4616 4856 4653 4860
rect 4596 4844 4604 4856
rect 4716 4856 4753 4864
rect 4596 4836 4644 4844
rect 3896 4820 3984 4824
rect 3893 4816 3984 4820
rect 2967 4796 3124 4804
rect 3893 4807 3907 4816
rect 4636 4826 4644 4836
rect 4716 4827 4724 4856
rect 4776 4856 4832 4864
rect 4776 4844 4784 4856
rect 5047 4856 5193 4864
rect 5276 4856 5353 4864
rect 4756 4840 4784 4844
rect 4753 4836 4784 4840
rect 4753 4827 4767 4836
rect 4856 4823 4864 4853
rect 5276 4827 5284 4856
rect 5376 4856 5433 4864
rect 5376 4844 5384 4856
rect 5336 4836 5384 4844
rect 4807 4815 4864 4823
rect 5067 4815 5093 4823
rect 5187 4815 5233 4823
rect 5336 4826 5344 4836
rect 5716 4827 5724 4893
rect 5747 4876 5784 4884
rect 5776 4868 5784 4876
rect 5787 4856 5853 4864
rect 5896 4844 5904 4896
rect 5947 4876 5973 4884
rect 5856 4840 5904 4844
rect 5853 4836 5904 4840
rect 5916 4864 5924 4873
rect 5916 4856 6013 4864
rect 5853 4827 5867 4836
rect 5507 4815 5533 4823
rect 5916 4826 5924 4856
rect 6067 4857 6133 4865
rect 4007 4796 4053 4804
rect 4127 4796 4153 4804
rect 4167 4796 4233 4804
rect 5607 4796 5693 4804
rect 5767 4796 5813 4804
rect 5936 4796 6013 4804
rect 1847 4776 2033 4784
rect 2047 4776 2213 4784
rect 2367 4776 2513 4784
rect 2667 4776 2693 4784
rect 2847 4776 2973 4784
rect 3247 4776 3433 4784
rect 3447 4776 3593 4784
rect 3607 4776 3833 4784
rect 4687 4776 4813 4784
rect 4827 4776 4873 4784
rect 5167 4776 5293 4784
rect 5707 4776 5872 4784
rect 5936 4784 5944 4796
rect 6087 4796 6113 4804
rect 5907 4776 5944 4784
rect 1447 4756 1633 4764
rect 1647 4756 1853 4764
rect 2067 4756 2173 4764
rect 2307 4756 2633 4764
rect 2767 4756 2953 4764
rect 3147 4756 3473 4764
rect 3687 4756 3753 4764
rect 3947 4756 3993 4764
rect 4007 4756 4133 4764
rect 4427 4756 4533 4764
rect 4547 4756 4733 4764
rect 4907 4756 5353 4764
rect 5807 4756 5953 4764
rect 6027 4756 6153 4764
rect 407 4736 653 4744
rect 667 4736 733 4744
rect 2207 4736 2273 4744
rect 2287 4736 2613 4744
rect 2807 4736 2913 4744
rect 3067 4736 3153 4744
rect 3327 4736 3613 4744
rect 4267 4736 4313 4744
rect 5827 4736 5933 4744
rect 1187 4716 1793 4724
rect 2127 4716 2833 4724
rect 3047 4716 3173 4724
rect 3287 4716 3853 4724
rect 4367 4716 4453 4724
rect 4887 4716 4953 4724
rect 4967 4716 5133 4724
rect 5887 4716 6133 4724
rect 1167 4696 1413 4704
rect 1787 4696 1933 4704
rect 2107 4696 2953 4704
rect 3007 4696 4224 4704
rect 1107 4676 1753 4684
rect 1807 4676 2113 4684
rect 2167 4676 2313 4684
rect 2567 4676 2813 4684
rect 3587 4676 3793 4684
rect 3847 4676 3893 4684
rect 4216 4684 4224 4696
rect 4327 4696 4633 4704
rect 5327 4696 5373 4704
rect 5387 4696 5753 4704
rect 5987 4696 6013 4704
rect 4216 4676 4373 4684
rect 5107 4676 5724 4684
rect -63 4648 232 4656
rect 1287 4656 1493 4664
rect 2027 4656 2073 4664
rect 2847 4656 2993 4664
rect 3187 4656 3473 4664
rect 3527 4656 4053 4664
rect 4207 4656 4433 4664
rect 5716 4664 5724 4676
rect 5827 4676 6193 4684
rect 6235 4664 6243 5096
rect 5447 4656 5704 4664
rect 5716 4656 6243 4664
rect 1807 4636 2173 4644
rect 2487 4636 2693 4644
rect 3027 4636 3433 4644
rect 3447 4636 4113 4644
rect 4427 4636 4573 4644
rect 4927 4636 5113 4644
rect 5127 4636 5333 4644
rect 5696 4644 5704 4656
rect 5696 4636 5773 4644
rect 5987 4636 6033 4644
rect 67 4616 93 4624
rect 527 4616 633 4624
rect 767 4616 933 4624
rect 1367 4616 1593 4624
rect 2087 4616 2153 4624
rect 2827 4616 3033 4624
rect 3147 4616 3313 4624
rect 3487 4616 3713 4624
rect 4527 4616 4713 4624
rect 5007 4616 5313 4624
rect 5587 4616 5853 4624
rect 27 4596 153 4604
rect 987 4596 1173 4604
rect 1887 4596 2053 4604
rect 2587 4596 2793 4604
rect 2807 4596 3453 4604
rect 3467 4596 3593 4604
rect 4067 4596 4493 4604
rect 4596 4596 4893 4604
rect 387 4576 413 4584
rect 527 4576 573 4584
rect 887 4576 1093 4584
rect 1107 4576 1153 4584
rect 1447 4576 2133 4584
rect 47 4556 93 4564
rect 107 4557 173 4565
rect 316 4544 324 4554
rect 347 4556 493 4564
rect 607 4556 693 4564
rect 736 4556 793 4564
rect 316 4536 473 4544
rect 87 4516 113 4524
rect 367 4516 493 4524
rect 567 4515 593 4523
rect 647 4515 673 4523
rect 736 4524 744 4556
rect 727 4516 744 4524
rect 767 4516 813 4524
rect 836 4524 844 4554
rect 1047 4556 1093 4564
rect 1227 4557 1313 4565
rect 1133 4544 1147 4553
rect 1116 4540 1147 4544
rect 1116 4536 1144 4540
rect 1116 4526 1124 4536
rect 836 4516 993 4524
rect 1136 4516 1193 4524
rect -63 4496 273 4504
rect 1136 4504 1144 4516
rect 1207 4515 1333 4523
rect 1356 4524 1364 4554
rect 1416 4527 1424 4573
rect 1436 4547 1444 4574
rect 2187 4576 2224 4584
rect 1607 4557 1972 4565
rect 1436 4536 1453 4547
rect 1440 4533 1453 4536
rect 1607 4536 1753 4544
rect 1993 4544 2007 4553
rect 1827 4536 1984 4544
rect 1993 4540 2193 4544
rect 1996 4536 2193 4540
rect 1347 4516 1364 4524
rect 1887 4516 1953 4524
rect 1976 4524 1984 4536
rect 1976 4516 2073 4524
rect 2216 4507 2224 4576
rect 2316 4524 2324 4534
rect 2456 4524 2464 4593
rect 2707 4576 3073 4584
rect 4596 4584 4604 4596
rect 5847 4596 5993 4604
rect 6147 4596 6213 4604
rect 3987 4576 4604 4584
rect 4647 4576 4733 4584
rect 4947 4576 4973 4584
rect 5780 4584 5793 4587
rect 5776 4573 5793 4584
rect 2627 4557 2653 4565
rect 2856 4556 3013 4564
rect 2487 4536 2513 4544
rect 2316 4516 2364 4524
rect 2456 4516 2513 4524
rect 1027 4496 1144 4504
rect 1307 4496 1373 4504
rect 1787 4496 1973 4504
rect 2207 4496 2224 4507
rect 2356 4504 2364 4516
rect 2607 4516 2673 4524
rect 2856 4526 2864 4556
rect 3107 4557 3173 4565
rect 3367 4556 3753 4564
rect 3767 4556 3873 4564
rect 2767 4516 2813 4524
rect 3047 4516 3073 4524
rect 3236 4524 3244 4554
rect 4247 4557 4273 4565
rect 4467 4556 4553 4564
rect 3953 4544 3967 4553
rect 3896 4540 3967 4544
rect 3896 4536 3964 4540
rect 3207 4516 3244 4524
rect 3547 4516 3733 4524
rect 3896 4524 3904 4536
rect 3876 4520 3904 4524
rect 3873 4516 3904 4520
rect 3873 4507 3887 4516
rect 4156 4524 4164 4554
rect 4627 4556 4673 4564
rect 4753 4544 4767 4553
rect 4793 4544 4807 4553
rect 4847 4557 4873 4565
rect 5067 4556 5153 4564
rect 5207 4557 5233 4565
rect 5427 4556 5453 4564
rect 5507 4556 5533 4564
rect 4647 4540 4767 4544
rect 4776 4540 4807 4544
rect 4647 4536 4764 4540
rect 4776 4536 4804 4540
rect 4047 4516 4164 4524
rect 4187 4516 4233 4524
rect 4776 4526 4784 4536
rect 4387 4516 4433 4524
rect 4587 4515 4613 4523
rect 4847 4516 4953 4524
rect 4967 4515 5033 4523
rect 5267 4516 5513 4524
rect 5596 4507 5604 4553
rect 5687 4516 5753 4524
rect 5776 4524 5784 4573
rect 5827 4557 5873 4565
rect 6107 4557 6173 4565
rect 5767 4516 5784 4524
rect 2356 4496 2384 4504
rect 2207 4493 2220 4496
rect 487 4476 573 4484
rect 627 4476 693 4484
rect 907 4476 1284 4484
rect 187 4456 393 4464
rect 407 4456 873 4464
rect 1087 4456 1153 4464
rect 1276 4464 1284 4476
rect 1507 4476 1813 4484
rect 1907 4476 1993 4484
rect 2376 4484 2384 4496
rect 2967 4496 3173 4504
rect 3227 4496 3273 4504
rect 3387 4496 3413 4504
rect 3927 4496 3973 4504
rect 5187 4496 5393 4504
rect 5936 4504 5944 4553
rect 5976 4527 5984 4553
rect 6067 4516 6193 4524
rect 5887 4496 6013 4504
rect 2376 4476 2673 4484
rect 2747 4476 2793 4484
rect 2907 4476 2973 4484
rect 2987 4476 3113 4484
rect 3127 4476 3333 4484
rect 3607 4476 3713 4484
rect 4467 4476 4633 4484
rect 4947 4476 5273 4484
rect 5427 4476 5613 4484
rect 5667 4476 5793 4484
rect 6216 4484 6224 4554
rect 6187 4476 6224 4484
rect 1276 4456 1473 4464
rect 2187 4456 2213 4464
rect 2236 4456 2693 4464
rect 787 4436 952 4444
rect 987 4436 1013 4444
rect 1027 4436 1633 4444
rect 1707 4436 1733 4444
rect 1747 4436 1833 4444
rect 2236 4444 2244 4456
rect 2827 4456 3493 4464
rect 3587 4456 3633 4464
rect 3827 4456 4293 4464
rect 5107 4456 5173 4464
rect 5436 4456 5533 4464
rect 2147 4436 2244 4444
rect 2376 4436 2753 4444
rect 387 4416 813 4424
rect 1467 4416 1552 4424
rect 1587 4416 1793 4424
rect 1867 4416 1973 4424
rect 2376 4424 2384 4436
rect 3007 4436 3193 4444
rect 3207 4436 3233 4444
rect 3667 4436 3753 4444
rect 4547 4436 4833 4444
rect 4947 4436 4993 4444
rect 5436 4444 5444 4456
rect 5707 4456 5753 4464
rect 5827 4456 6072 4464
rect 6107 4456 6233 4464
rect 5347 4436 5444 4444
rect 5567 4436 5693 4444
rect 2207 4416 2384 4424
rect 2407 4416 2473 4424
rect 2627 4416 2652 4424
rect 2687 4416 2733 4424
rect 2787 4416 2973 4424
rect 3876 4416 3893 4424
rect 307 4396 333 4404
rect 907 4396 1193 4404
rect 1247 4396 1433 4404
rect 1687 4396 1993 4404
rect 2176 4396 2493 4404
rect 476 4376 613 4384
rect 476 4364 484 4376
rect 1047 4376 1093 4384
rect 1407 4376 1573 4384
rect 2027 4376 2133 4384
rect 2176 4384 2184 4396
rect 2767 4396 2813 4404
rect 3007 4396 3693 4404
rect 3876 4404 3884 4416
rect 3907 4416 3973 4424
rect 4347 4416 4513 4424
rect 5587 4416 5893 4424
rect 3807 4396 3884 4404
rect 4007 4396 4053 4404
rect 4356 4396 4473 4404
rect 4356 4387 4364 4396
rect 2147 4376 2184 4384
rect 2447 4376 2473 4384
rect 3747 4376 4353 4384
rect 5027 4376 5233 4384
rect 5487 4376 5593 4384
rect 5607 4376 5853 4384
rect 6107 4376 6153 4384
rect 247 4356 484 4364
rect 1507 4356 1533 4364
rect 1647 4356 2033 4364
rect 2307 4356 2573 4364
rect 2907 4356 3193 4364
rect 3287 4356 3353 4364
rect 3407 4356 3644 4364
rect 67 4337 93 4345
rect 147 4337 173 4345
rect 387 4336 433 4344
rect 507 4337 533 4345
rect 867 4336 953 4344
rect 576 4304 584 4334
rect 1007 4336 1053 4344
rect 1096 4336 1233 4344
rect 487 4296 653 4304
rect 847 4296 893 4304
rect 947 4295 993 4303
rect 1096 4304 1104 4336
rect 1276 4336 1333 4344
rect 1276 4324 1284 4336
rect 1427 4337 1593 4345
rect 2067 4336 2253 4344
rect 2396 4336 2473 4344
rect 1256 4316 1284 4324
rect 1087 4296 1104 4304
rect 1256 4304 1264 4316
rect 1167 4296 1264 4304
rect 1307 4295 1373 4303
rect 187 4276 393 4284
rect 407 4276 633 4284
rect 936 4284 944 4292
rect 647 4276 944 4284
rect 1676 4287 1684 4333
rect 1733 4324 1747 4333
rect 1733 4320 1813 4324
rect 1736 4316 1813 4320
rect 2236 4316 2293 4324
rect 1693 4304 1707 4313
rect 1693 4300 1724 4304
rect 1696 4296 1724 4300
rect 1676 4276 1693 4287
rect 1680 4273 1693 4276
rect 1147 4256 1293 4264
rect 1347 4256 1393 4264
rect 1716 4264 1724 4296
rect 2236 4306 2244 4316
rect 2396 4306 2404 4336
rect 2607 4336 2673 4344
rect 3636 4347 3644 4356
rect 4307 4356 4353 4364
rect 4427 4356 4533 4364
rect 4767 4356 4973 4364
rect 5427 4356 5453 4364
rect 5647 4356 5673 4364
rect 6087 4356 6113 4364
rect 3147 4336 3173 4344
rect 3196 4336 3524 4344
rect 3636 4336 3653 4347
rect 2047 4295 2193 4303
rect 1827 4276 2033 4284
rect 2516 4284 2524 4333
rect 3196 4324 3204 4336
rect 2827 4316 3204 4324
rect 3367 4316 3493 4324
rect 3516 4324 3524 4336
rect 3640 4333 3653 4336
rect 3676 4336 3773 4344
rect 3676 4324 3684 4336
rect 3847 4336 3913 4344
rect 4027 4336 4193 4344
rect 4207 4337 4253 4345
rect 4496 4336 4513 4344
rect 3516 4316 3684 4324
rect 3727 4316 3904 4324
rect 3896 4307 3904 4316
rect 4276 4316 4344 4324
rect 2687 4295 2713 4303
rect 3227 4295 3293 4303
rect 3896 4296 3913 4307
rect 3900 4293 3913 4296
rect 4276 4306 4284 4316
rect 4336 4306 4344 4316
rect 3967 4295 4053 4303
rect 4347 4295 4433 4303
rect 2427 4276 2524 4284
rect 2547 4276 2573 4284
rect 2587 4276 2653 4284
rect 2847 4276 3013 4284
rect 3147 4275 3333 4283
rect 3347 4276 3493 4284
rect 4307 4276 4353 4284
rect 4456 4284 4464 4333
rect 4496 4307 4504 4336
rect 4567 4336 4673 4344
rect 4727 4336 4773 4344
rect 4796 4336 4813 4344
rect 4796 4324 4804 4336
rect 5107 4337 5133 4345
rect 5187 4336 5293 4344
rect 4656 4316 4933 4324
rect 4656 4306 4664 4316
rect 5176 4324 5184 4334
rect 5627 4337 5653 4345
rect 5767 4336 5833 4344
rect 5967 4336 6053 4344
rect 5116 4320 5184 4324
rect 5113 4316 5184 4320
rect 5416 4324 5424 4333
rect 5416 4316 5513 4324
rect 5113 4307 5127 4316
rect 5876 4307 5884 4333
rect 5976 4307 5984 4336
rect 4587 4296 4653 4304
rect 4847 4295 4913 4303
rect 5007 4295 5073 4303
rect 5487 4296 5573 4304
rect 5587 4295 5753 4303
rect 6116 4306 6124 4353
rect 6147 4336 6193 4344
rect 4427 4276 4464 4284
rect 5047 4276 5373 4284
rect 5387 4276 5453 4284
rect 1716 4256 2073 4264
rect 2627 4256 2753 4264
rect 3867 4256 3993 4264
rect 4227 4256 4553 4264
rect 4667 4256 4893 4264
rect 5327 4256 5373 4264
rect 5907 4256 5953 4264
rect 367 4236 393 4244
rect 767 4236 933 4244
rect 1587 4236 1673 4244
rect 2807 4236 2933 4244
rect 3007 4236 3053 4244
rect 3327 4236 4153 4244
rect 4167 4236 4593 4244
rect 4607 4236 5273 4244
rect 5287 4236 5393 4244
rect 5896 4244 5904 4253
rect 5787 4236 5904 4244
rect 6107 4236 6133 4244
rect 1327 4216 1993 4224
rect 2067 4216 2093 4224
rect 2207 4216 2353 4224
rect 2507 4216 2613 4224
rect 2667 4216 2953 4224
rect 2967 4216 3073 4224
rect 3127 4216 3253 4224
rect 3647 4216 4133 4224
rect 4147 4216 4453 4224
rect 4647 4216 4733 4224
rect 4887 4216 5213 4224
rect 5227 4216 5333 4224
rect 5447 4216 5513 4224
rect 5527 4216 5613 4224
rect 5627 4216 5704 4224
rect 247 4196 1213 4204
rect 1387 4196 1693 4204
rect 2447 4196 2633 4204
rect 2747 4196 3153 4204
rect 3167 4196 3313 4204
rect 3767 4196 3853 4204
rect 4087 4196 4173 4204
rect 5427 4196 5673 4204
rect 5696 4204 5704 4216
rect 5867 4216 5933 4224
rect 5947 4216 5993 4224
rect 5696 4196 5824 4204
rect 1187 4176 1453 4184
rect 1507 4176 2273 4184
rect 3607 4176 3693 4184
rect 4207 4176 4273 4184
rect 4347 4176 4653 4184
rect 5416 4184 5424 4193
rect 5167 4176 5424 4184
rect 5816 4184 5824 4196
rect 5816 4176 5973 4184
rect 6147 4176 6193 4184
rect 447 4156 833 4164
rect 1707 4156 2233 4164
rect 2707 4156 3093 4164
rect 3407 4156 3433 4164
rect 3507 4156 3833 4164
rect 3927 4156 4633 4164
rect 6007 4156 6153 4164
rect 727 4136 953 4144
rect 1627 4136 2453 4144
rect 2476 4136 2813 4144
rect 267 4116 373 4124
rect 607 4116 1193 4124
rect 1207 4116 1353 4124
rect 1527 4116 1873 4124
rect 2476 4124 2484 4136
rect 3516 4136 4673 4144
rect 2007 4116 2484 4124
rect 3516 4124 3524 4136
rect 4787 4136 4833 4144
rect 5107 4136 5213 4144
rect 5967 4136 6113 4144
rect 3107 4116 3524 4124
rect 3827 4116 4333 4124
rect 5847 4116 5884 4124
rect 727 4096 1093 4104
rect 1107 4096 1153 4104
rect 1987 4096 2173 4104
rect 2767 4096 2893 4104
rect 3587 4096 3773 4104
rect 3867 4096 4193 4104
rect 4787 4096 5053 4104
rect 5467 4096 5613 4104
rect 5687 4096 5813 4104
rect 5876 4104 5884 4116
rect 5876 4096 6113 4104
rect 6207 4093 6213 4107
rect 67 4076 193 4084
rect 307 4076 533 4084
rect 547 4076 673 4084
rect 787 4076 973 4084
rect 987 4076 1253 4084
rect 1387 4076 1433 4084
rect 1487 4076 1533 4084
rect 1647 4076 1813 4084
rect 2056 4076 2113 4084
rect 227 4056 273 4064
rect 1847 4056 1893 4064
rect 2056 4064 2064 4076
rect 2667 4076 2733 4084
rect 2780 4084 2793 4087
rect 2776 4073 2793 4084
rect 2867 4076 3053 4084
rect 3807 4076 3973 4084
rect 4487 4076 4533 4084
rect 4667 4076 4753 4084
rect 5376 4076 5733 4084
rect 1956 4056 2064 4064
rect 1956 4048 1964 4056
rect 167 4037 193 4045
rect 327 4037 353 4045
rect 447 4036 573 4044
rect 147 3996 193 4004
rect 396 4004 404 4033
rect 620 4024 633 4027
rect 616 4020 633 4024
rect 613 4013 633 4020
rect 613 4007 627 4013
rect 676 4007 684 4033
rect 956 4007 964 4033
rect 1136 4024 1144 4034
rect 1247 4036 1293 4044
rect 1347 4036 1413 4044
rect 1436 4036 1513 4044
rect 1436 4024 1444 4036
rect 1527 4036 1633 4044
rect 1747 4037 1773 4045
rect 2087 4036 2193 4044
rect 1136 4016 1444 4024
rect 396 3996 413 4004
rect 467 3996 493 4004
rect 1167 3995 1192 4003
rect 1436 4006 1444 4016
rect 1676 4007 1684 4034
rect 1227 3995 1273 4003
rect 1676 3996 1693 4007
rect 1680 3993 1693 3996
rect 1807 3995 1853 4003
rect 1956 4004 1964 4034
rect 1927 3996 1964 4004
rect 1996 4004 2004 4034
rect 2076 4024 2084 4034
rect 2076 4016 2124 4024
rect 1996 3996 2093 4004
rect 2116 4004 2124 4016
rect 2236 4007 2244 4034
rect 2116 3996 2144 4004
rect -63 3976 113 3984
rect 667 3976 693 3984
rect 707 3976 733 3984
rect 947 3976 973 3984
rect 1587 3976 2113 3984
rect 2136 3984 2144 3996
rect 2187 3995 2213 4003
rect 2236 3996 2253 4007
rect 2240 3993 2253 3996
rect 2376 4004 2384 4034
rect 2496 4024 2504 4034
rect 2587 4036 2613 4044
rect 2636 4036 2673 4044
rect 2496 4016 2553 4024
rect 2636 4006 2644 4036
rect 2376 3996 2473 4004
rect 2516 3996 2593 4004
rect 2136 3976 2173 3984
rect 367 3956 433 3964
rect 867 3956 993 3964
rect 1013 3964 1027 3973
rect 2516 3984 2524 3996
rect 2327 3976 2384 3984
rect 1013 3956 1113 3964
rect 1567 3956 1613 3964
rect 1847 3956 1873 3964
rect 1887 3956 1933 3964
rect 1987 3956 2033 3964
rect 2287 3956 2353 3964
rect 2376 3964 2384 3976
rect 2496 3976 2524 3984
rect 2496 3964 2504 3976
rect 2776 3984 2784 4073
rect 5376 4067 5384 4076
rect 2796 4056 2833 4064
rect 2796 4004 2804 4056
rect 3636 4056 3753 4064
rect 2947 4037 2973 4045
rect 2816 4024 2824 4034
rect 3036 4024 3044 4053
rect 3636 4048 3644 4056
rect 4947 4056 4973 4064
rect 5147 4056 5193 4064
rect 5367 4056 5384 4067
rect 5367 4053 5380 4056
rect 5627 4056 5773 4064
rect 6027 4056 6073 4064
rect 3347 4036 3553 4044
rect 3687 4037 3713 4045
rect 3816 4036 3993 4044
rect 2816 4016 2864 4024
rect 3036 4016 3113 4024
rect 2796 3996 2833 4004
rect 2856 4004 2864 4016
rect 3467 4016 3533 4024
rect 3636 4024 3644 4034
rect 3593 4016 3644 4024
rect 3593 4007 3607 4016
rect 3816 4007 3824 4036
rect 4267 4037 4353 4045
rect 4407 4037 4493 4045
rect 4707 4036 4733 4044
rect 4867 4037 4893 4045
rect 5021 4036 5093 4044
rect 3867 4016 3973 4024
rect 5213 4024 5227 4033
rect 5196 4020 5227 4024
rect 5236 4036 5273 4044
rect 5196 4016 5224 4020
rect 2856 3996 2913 4004
rect 3007 3996 3153 4004
rect 3727 3996 3773 4004
rect 4167 3996 4233 4004
rect 4247 3996 4273 4004
rect 4447 3995 4473 4003
rect 4547 3995 4633 4003
rect 4687 3996 4753 4004
rect 4847 3995 5033 4003
rect 5196 4004 5204 4016
rect 5236 4007 5244 4036
rect 5387 4036 5444 4044
rect 5347 4016 5424 4024
rect 5147 3996 5204 4004
rect 5227 3996 5244 4007
rect 5227 3993 5240 3996
rect 2667 3976 2784 3984
rect 3187 3976 3433 3984
rect 3627 3976 3893 3984
rect 4807 3976 4873 3984
rect 4987 3976 5293 3984
rect 5416 3984 5424 4016
rect 5436 4004 5444 4036
rect 5487 4037 5513 4045
rect 5827 4037 5933 4045
rect 5947 4036 5972 4044
rect 5436 3996 5453 4004
rect 5576 4004 5584 4034
rect 5507 3996 5584 4004
rect 5696 4004 5704 4034
rect 6227 4038 6243 4046
rect 5996 4007 6004 4033
rect 5647 3996 5704 4004
rect 6176 4004 6184 4034
rect 6116 3996 6184 4004
rect 5416 3976 5593 3984
rect 5607 3976 5753 3984
rect 6116 3984 6124 3996
rect 6087 3976 6124 3984
rect 2376 3956 2504 3964
rect 2707 3956 2752 3964
rect 2787 3956 2853 3964
rect 2927 3956 3013 3964
rect 3107 3956 3433 3964
rect 3447 3956 3573 3964
rect 3627 3956 3904 3964
rect 107 3936 293 3944
rect 387 3936 533 3944
rect 607 3936 733 3944
rect 827 3936 1093 3944
rect 1167 3936 1193 3944
rect 1707 3936 1872 3944
rect 1907 3936 2213 3944
rect 2347 3936 2513 3944
rect 2887 3936 2973 3944
rect 3107 3936 3453 3944
rect 3567 3936 3653 3944
rect 427 3916 713 3924
rect 736 3916 1204 3924
rect 736 3904 744 3916
rect 447 3896 744 3904
rect 847 3896 913 3904
rect 1196 3904 1204 3916
rect 1287 3916 1373 3924
rect 1416 3916 2613 3924
rect 1416 3904 1424 3916
rect 3147 3916 3213 3924
rect 3307 3916 3833 3924
rect 3896 3924 3904 3956
rect 4307 3956 4513 3964
rect 4927 3956 5093 3964
rect 5347 3956 5433 3964
rect 5727 3956 5753 3964
rect 6147 3956 6213 3964
rect 4987 3936 5553 3944
rect 6235 3944 6243 4038
rect 5987 3936 6243 3944
rect 3896 3916 4033 3924
rect 4367 3916 5784 3924
rect 967 3896 1184 3904
rect 1196 3896 1424 3904
rect 207 3876 393 3884
rect 727 3876 813 3884
rect 1067 3876 1133 3884
rect 1176 3884 1184 3896
rect 1767 3896 1892 3904
rect 1927 3896 1973 3904
rect 2627 3896 2653 3904
rect 2747 3896 2793 3904
rect 3127 3896 3253 3904
rect 3467 3896 3613 3904
rect 3707 3896 3773 3904
rect 4147 3896 4173 3904
rect 5087 3896 5173 3904
rect 5776 3904 5784 3916
rect 6007 3916 6153 3924
rect 5776 3896 5813 3904
rect 5896 3896 6073 3904
rect 5896 3887 5904 3896
rect 1176 3876 1373 3884
rect 2327 3876 2373 3884
rect 2787 3876 3353 3884
rect 3747 3876 3853 3884
rect 4047 3876 4333 3884
rect 5867 3876 5893 3884
rect 867 3856 953 3864
rect 1047 3856 1193 3864
rect 1447 3856 1493 3864
rect 2307 3856 2393 3864
rect 2587 3856 2733 3864
rect 3527 3856 3693 3864
rect 4107 3856 4213 3864
rect 4807 3856 4893 3864
rect 5287 3856 5353 3864
rect 5667 3856 5693 3864
rect 407 3836 444 3844
rect 247 3816 293 3824
rect 116 3804 124 3814
rect 367 3817 413 3825
rect 116 3800 184 3804
rect 116 3796 187 3800
rect 173 3787 187 3796
rect -63 3776 73 3784
rect 436 3784 444 3836
rect 567 3836 593 3844
rect 707 3836 1013 3844
rect 1427 3836 1473 3844
rect 1907 3836 1993 3844
rect 2007 3836 2133 3844
rect 3207 3836 3233 3844
rect 3887 3836 3953 3844
rect 4027 3836 4113 3844
rect 4327 3836 4473 3844
rect 4607 3836 4633 3844
rect 4876 3836 4933 3844
rect 536 3804 544 3814
rect 627 3816 764 3824
rect 536 3800 584 3804
rect 536 3796 587 3800
rect 573 3787 587 3796
rect 436 3776 473 3784
rect 756 3786 764 3816
rect 787 3816 853 3824
rect 947 3816 993 3824
rect 647 3780 684 3784
rect 647 3776 687 3780
rect 673 3767 687 3776
rect 167 3756 213 3764
rect 347 3756 593 3764
rect 896 3764 904 3814
rect 927 3775 953 3783
rect 1056 3784 1064 3814
rect 1307 3816 1333 3824
rect 2087 3816 2204 3824
rect 1096 3787 1104 3813
rect 1007 3776 1064 3784
rect 1167 3776 1393 3784
rect 1407 3775 1453 3783
rect 1476 3767 1484 3813
rect 1887 3796 1953 3804
rect 1573 3784 1587 3793
rect 1527 3780 1587 3784
rect 1527 3776 1584 3780
rect 1727 3776 1853 3784
rect 2196 3786 2204 3816
rect 2267 3816 2353 3824
rect 2467 3816 2513 3824
rect 2667 3816 2684 3824
rect 2027 3776 2053 3784
rect 2427 3775 2453 3783
rect 2567 3776 2593 3784
rect 2676 3784 2684 3816
rect 2707 3817 2753 3825
rect 2676 3776 2733 3784
rect 2776 3786 2784 3833
rect 2796 3767 2804 3814
rect 3327 3817 3373 3825
rect 3487 3816 3553 3824
rect 3633 3824 3647 3833
rect 3633 3820 3673 3824
rect 3636 3816 3673 3820
rect 3756 3816 4133 3824
rect 687 3756 904 3764
rect 1147 3756 1373 3764
rect 1527 3755 1553 3763
rect 2107 3756 2233 3764
rect 2247 3756 2633 3764
rect 2836 3764 2844 3813
rect 2887 3796 3044 3804
rect 3036 3767 3044 3796
rect 3756 3807 3764 3816
rect 4227 3816 4304 3824
rect 3196 3767 3204 3794
rect 3747 3796 3764 3807
rect 3776 3796 3873 3804
rect 3747 3793 3760 3796
rect 3236 3767 3244 3793
rect 3347 3775 3533 3783
rect 3776 3784 3784 3796
rect 3887 3796 4013 3804
rect 3667 3776 3784 3784
rect 3807 3776 3933 3784
rect 4007 3775 4033 3783
rect 4047 3775 4073 3783
rect 4176 3784 4184 3813
rect 4296 3786 4304 3816
rect 4747 3817 4833 3825
rect 4147 3776 4184 3784
rect 2836 3756 2873 3764
rect 3027 3756 3044 3767
rect 3027 3753 3040 3756
rect 3187 3756 3204 3767
rect 3187 3753 3200 3756
rect 4436 3764 4444 3813
rect 4436 3756 4473 3764
rect 4516 3747 4524 3814
rect 4567 3796 4673 3804
rect 4767 3776 4813 3784
rect 4876 3786 4884 3836
rect 5027 3836 5253 3844
rect 5267 3836 5313 3844
rect 5856 3836 5893 3844
rect 4992 3824 5006 3833
rect 4916 3816 5153 3824
rect 4916 3786 4924 3816
rect 5176 3816 5193 3824
rect 5176 3804 5184 3816
rect 5307 3816 5344 3824
rect 5036 3796 5184 3804
rect 5036 3786 5044 3796
rect 5336 3786 5344 3816
rect 5356 3804 5364 3814
rect 5567 3817 5593 3825
rect 5356 3796 5384 3804
rect 5376 3787 5384 3796
rect 5456 3787 5464 3813
rect 5856 3804 5864 3836
rect 5836 3796 5864 3804
rect 5227 3775 5253 3783
rect 5376 3776 5393 3787
rect 5380 3773 5393 3776
rect 5836 3784 5844 3796
rect 5876 3787 5884 3813
rect 6016 3804 6024 3833
rect 6067 3816 6093 3824
rect 6107 3816 6133 3824
rect 5996 3800 6024 3804
rect 6096 3800 6153 3804
rect 5993 3796 6024 3800
rect 6093 3796 6153 3800
rect 5993 3787 6007 3796
rect 5827 3776 5844 3784
rect 6093 3787 6107 3796
rect 5047 3756 5093 3764
rect 6047 3756 6113 3764
rect 267 3736 493 3744
rect 647 3736 753 3744
rect 867 3736 933 3744
rect 1127 3736 1493 3744
rect 2187 3736 2693 3744
rect 2916 3736 2993 3744
rect 607 3716 753 3724
rect 807 3716 833 3724
rect 847 3716 1033 3724
rect 1227 3716 1433 3724
rect 1596 3716 2084 3724
rect 187 3696 453 3704
rect 667 3696 913 3704
rect 1467 3696 1573 3704
rect 1596 3704 1604 3716
rect 1587 3696 1604 3704
rect 2076 3704 2084 3716
rect 2147 3716 2784 3724
rect 2076 3696 2273 3704
rect 2327 3696 2533 3704
rect 2776 3704 2784 3716
rect 2916 3724 2924 3736
rect 3167 3736 3253 3744
rect 3547 3736 3613 3744
rect 3627 3736 3693 3744
rect 4087 3736 4293 3744
rect 4500 3746 4524 3747
rect 4507 3736 4524 3746
rect 4507 3733 4520 3736
rect 5647 3736 5853 3744
rect 2807 3716 2924 3724
rect 3367 3716 3793 3724
rect 3887 3716 3953 3724
rect 4327 3716 4413 3724
rect 4427 3716 4453 3724
rect 4847 3716 5424 3724
rect 2776 3696 2853 3704
rect 3287 3696 3553 3704
rect 3807 3696 4153 3704
rect 4196 3696 4853 3704
rect 4196 3687 4204 3696
rect 5147 3696 5193 3704
rect 5416 3704 5424 3716
rect 5447 3716 5993 3724
rect 6007 3716 6193 3724
rect 5416 3696 5632 3704
rect 5667 3696 5713 3704
rect 5727 3696 5913 3704
rect 487 3676 593 3684
rect 687 3676 993 3684
rect 1387 3676 1553 3684
rect 1707 3676 1973 3684
rect 2067 3676 2453 3684
rect 2747 3676 2813 3684
rect 2907 3676 3293 3684
rect 3827 3676 4133 3684
rect 4187 3676 4204 3687
rect 4187 3673 4200 3676
rect 4647 3676 4773 3684
rect 5007 3676 5173 3684
rect 5387 3676 5513 3684
rect 6087 3676 6233 3684
rect 107 3656 133 3664
rect 727 3656 904 3664
rect 207 3636 292 3644
rect 327 3636 393 3644
rect 447 3636 613 3644
rect 767 3636 873 3644
rect 896 3644 904 3656
rect 967 3656 1133 3664
rect 1407 3656 1433 3664
rect 1487 3656 1593 3664
rect 1847 3656 1913 3664
rect 2027 3656 2372 3664
rect 2407 3656 2433 3664
rect 3007 3656 3233 3664
rect 3407 3656 3733 3664
rect 3787 3656 3844 3664
rect 896 3636 1013 3644
rect 1187 3636 1273 3644
rect 1487 3636 1613 3644
rect 1627 3636 2593 3644
rect 2607 3636 2913 3644
rect 3047 3636 3173 3644
rect 3227 3636 3384 3644
rect 3376 3627 3384 3636
rect 3487 3636 3673 3644
rect 3836 3644 3844 3656
rect 4527 3656 4833 3664
rect 5247 3656 5453 3664
rect 5547 3656 5813 3664
rect 5907 3656 5953 3664
rect 3836 3636 4093 3644
rect 5567 3636 5673 3644
rect 5687 3636 5853 3644
rect 5867 3636 5973 3644
rect 107 3616 653 3624
rect 927 3616 1453 3624
rect 1507 3616 1813 3624
rect 1967 3616 2113 3624
rect 2267 3616 2293 3624
rect 2427 3616 2733 3624
rect 2836 3616 2893 3624
rect 607 3596 853 3604
rect 1107 3596 1333 3604
rect 2836 3604 2844 3616
rect 3156 3616 3313 3624
rect 2467 3596 2844 3604
rect 3156 3604 3164 3616
rect 3387 3616 3413 3624
rect 4207 3616 4633 3624
rect 4687 3616 5573 3624
rect 3027 3596 3164 3604
rect 3187 3596 3393 3604
rect 3567 3596 3773 3604
rect 4147 3596 4393 3604
rect 4707 3596 5013 3604
rect 5127 3596 5493 3604
rect 5787 3596 5893 3604
rect 567 3576 713 3584
rect 807 3576 973 3584
rect 1607 3576 1873 3584
rect 2727 3576 2793 3584
rect 2807 3576 2912 3584
rect 2947 3576 3272 3584
rect 3300 3584 3313 3587
rect 3296 3576 3313 3584
rect 3300 3573 3313 3576
rect 3327 3576 3333 3584
rect 3547 3576 3933 3584
rect 4027 3576 4673 3584
rect 4867 3576 5233 3584
rect 67 3556 324 3564
rect 316 3547 324 3556
rect 867 3556 1253 3564
rect 1267 3556 1453 3564
rect 1616 3556 1793 3564
rect 316 3536 333 3547
rect 16 3507 24 3533
rect 36 3507 44 3534
rect 320 3533 333 3536
rect 707 3536 853 3544
rect 416 3507 424 3533
rect 1067 3536 1193 3544
rect 1616 3544 1624 3556
rect 1867 3556 2413 3564
rect 2747 3556 3993 3564
rect 4207 3556 4313 3564
rect 4387 3556 4793 3564
rect 5667 3556 5693 3564
rect 6007 3556 6153 3564
rect 1496 3536 1624 3544
rect 467 3516 533 3524
rect 587 3516 653 3524
rect 676 3516 733 3524
rect 36 3496 53 3507
rect 40 3493 53 3496
rect 387 3476 433 3484
rect 487 3476 553 3484
rect 676 3484 684 3516
rect 907 3516 953 3524
rect 967 3517 1013 3525
rect 1036 3516 1073 3524
rect 1036 3504 1044 3516
rect 776 3500 1044 3504
rect 607 3476 684 3484
rect 773 3496 1044 3500
rect 773 3487 787 3496
rect 1216 3487 1224 3513
rect 827 3476 993 3484
rect 1107 3475 1153 3483
rect 1276 3486 1284 3533
rect 1496 3524 1504 3536
rect 1647 3536 1753 3544
rect 1987 3537 2092 3545
rect 2127 3536 2233 3544
rect 2687 3536 2813 3544
rect 2827 3536 2933 3544
rect 1407 3516 1504 3524
rect 1296 3487 1304 3513
rect 1356 3487 1364 3513
rect 1296 3476 1313 3487
rect 1300 3473 1313 3476
rect 1476 3484 1484 3516
rect 1527 3516 1544 3524
rect 1536 3504 1544 3516
rect 1567 3516 1713 3524
rect 1827 3516 1893 3524
rect 1907 3516 1953 3524
rect 2076 3520 2653 3524
rect 2073 3516 2653 3520
rect 2073 3507 2087 3516
rect 2967 3517 3113 3525
rect 3247 3517 3293 3525
rect 1536 3500 1564 3504
rect 1536 3496 1567 3500
rect 1553 3487 1567 3496
rect 2147 3496 2233 3504
rect 2707 3496 2824 3504
rect 1476 3476 1493 3484
rect 1787 3476 1933 3484
rect 1947 3476 2053 3484
rect 2816 3484 2824 3496
rect 3376 3487 3384 3534
rect 3847 3536 3893 3544
rect 3916 3536 4173 3544
rect 3547 3516 3673 3524
rect 3696 3520 3813 3524
rect 3693 3516 3813 3520
rect 3693 3507 3707 3516
rect 3916 3524 3924 3536
rect 4367 3536 4613 3544
rect 4907 3536 5053 3544
rect 5127 3536 5273 3544
rect 5287 3536 5353 3544
rect 5400 3544 5413 3547
rect 5396 3534 5413 3544
rect 5736 3536 5812 3544
rect 5396 3533 5420 3534
rect 3867 3516 3924 3524
rect 4227 3517 4273 3525
rect 4447 3516 4533 3524
rect 3427 3496 3513 3504
rect 2816 3476 2933 3484
rect 3236 3476 3313 3484
rect 807 3456 1073 3464
rect 1347 3456 1393 3464
rect 1407 3456 1533 3464
rect 1547 3456 1613 3464
rect 2427 3456 2793 3464
rect 2867 3456 2893 3464
rect 3236 3464 3244 3476
rect 3376 3476 3393 3487
rect 3380 3473 3393 3476
rect 3827 3475 3873 3483
rect 3936 3476 4093 3484
rect 3936 3467 3944 3476
rect 4307 3476 4393 3484
rect 4436 3484 4444 3514
rect 4620 3524 4633 3527
rect 4616 3513 4633 3524
rect 4767 3516 4932 3524
rect 4967 3517 5253 3525
rect 5320 3524 5333 3527
rect 4436 3476 4533 3484
rect 4616 3484 4624 3513
rect 4696 3487 4704 3513
rect 4827 3496 4904 3504
rect 4607 3476 4624 3484
rect 4747 3476 4793 3484
rect 4896 3467 4904 3496
rect 5047 3496 5184 3504
rect 5107 3475 5133 3483
rect 5176 3484 5184 3496
rect 5176 3476 5273 3484
rect 3127 3456 3244 3464
rect 3747 3456 3853 3464
rect 3927 3456 3944 3467
rect 3927 3453 3940 3456
rect 3987 3456 4013 3464
rect 4427 3456 4493 3464
rect 4987 3456 5153 3464
rect 427 3436 473 3444
rect 667 3436 733 3444
rect 847 3436 873 3444
rect 927 3436 1033 3444
rect 1487 3436 1513 3444
rect 1707 3436 1813 3444
rect 1887 3436 2773 3444
rect 3267 3436 3313 3444
rect 736 3424 744 3433
rect 3987 3436 4113 3444
rect 4687 3436 4733 3444
rect 5296 3444 5304 3514
rect 5316 3513 5333 3524
rect 5316 3464 5324 3513
rect 5396 3487 5404 3533
rect 5587 3517 5613 3525
rect 5627 3517 5633 3525
rect 5387 3476 5404 3487
rect 5387 3473 5400 3476
rect 5416 3464 5424 3513
rect 5516 3484 5524 3513
rect 5447 3476 5524 3484
rect 5736 3484 5744 3536
rect 5836 3524 5844 3533
rect 5767 3516 5893 3524
rect 6047 3517 6073 3525
rect 6113 3504 6127 3513
rect 5687 3476 5744 3484
rect 5856 3500 6127 3504
rect 5856 3496 6124 3500
rect 5316 3456 5424 3464
rect 5527 3456 5553 3464
rect 5856 3464 5864 3496
rect 5887 3475 5933 3483
rect 6196 3467 6204 3514
rect 5767 3456 5864 3464
rect 5147 3436 5393 3444
rect 5747 3436 5793 3444
rect 5807 3436 6133 3444
rect 736 3416 1113 3424
rect 1207 3416 1333 3424
rect 1347 3416 1653 3424
rect 2416 3416 2453 3424
rect 107 3396 133 3404
rect 207 3396 393 3404
rect 447 3396 513 3404
rect 607 3396 1373 3404
rect 2416 3404 2424 3416
rect 2507 3416 2593 3424
rect 2767 3416 3173 3424
rect 3807 3416 3873 3424
rect 3887 3416 4053 3424
rect 4136 3416 4173 3424
rect 2347 3396 2424 3404
rect 2807 3396 3033 3404
rect 3247 3396 3573 3404
rect 3587 3396 3733 3404
rect 3867 3396 3953 3404
rect 4136 3404 4144 3416
rect 4527 3416 4553 3424
rect 4707 3416 4773 3424
rect 5447 3416 5524 3424
rect 3967 3396 4144 3404
rect 4167 3396 4213 3404
rect 4236 3396 4372 3404
rect 96 3376 333 3384
rect 96 3367 104 3376
rect 847 3376 932 3384
rect 967 3376 1133 3384
rect 2007 3376 2033 3384
rect 2047 3376 2433 3384
rect 2867 3376 3013 3384
rect 3067 3376 3093 3384
rect 3547 3376 3833 3384
rect 4236 3384 4244 3396
rect 4407 3396 4604 3404
rect 4007 3376 4244 3384
rect 4596 3384 4604 3396
rect 4627 3396 4653 3404
rect 4987 3396 5073 3404
rect 5516 3404 5524 3416
rect 5647 3416 5973 3424
rect 6127 3416 6173 3424
rect 5516 3396 5693 3404
rect 6027 3396 6193 3404
rect 4347 3376 4484 3384
rect 4596 3376 4633 3384
rect 87 3356 104 3367
rect 87 3353 100 3356
rect 647 3356 713 3364
rect 1167 3356 1533 3364
rect 2067 3356 2753 3364
rect 2907 3356 2933 3364
rect 3847 3356 3873 3364
rect 3927 3356 3953 3364
rect 4367 3356 4453 3364
rect 4476 3364 4484 3376
rect 4887 3376 4933 3384
rect 5056 3376 5313 3384
rect 4476 3356 4653 3364
rect 4707 3356 4813 3364
rect 5056 3364 5064 3376
rect 5507 3376 5733 3384
rect 6087 3376 6153 3384
rect 4867 3356 5064 3364
rect 5076 3356 5373 3364
rect 5076 3347 5084 3356
rect 5527 3356 5793 3364
rect 5927 3356 6013 3364
rect 107 3336 493 3344
rect 1187 3336 1213 3344
rect 1576 3336 1853 3344
rect 767 3316 1153 3324
rect 1576 3324 1584 3336
rect 2167 3336 2293 3344
rect 2467 3336 2693 3344
rect 2787 3336 2853 3344
rect 2907 3336 3073 3344
rect 3947 3336 4433 3344
rect 4447 3336 5073 3344
rect 5427 3336 5553 3344
rect 5567 3336 5672 3344
rect 5707 3336 5773 3344
rect 1327 3316 1584 3324
rect 3316 3316 3493 3324
rect 47 3296 133 3304
rect 607 3297 693 3305
rect 760 3304 773 3307
rect 207 3276 312 3284
rect 473 3284 487 3293
rect 347 3280 487 3284
rect 756 3293 773 3304
rect 847 3304 860 3307
rect 847 3293 864 3304
rect 1267 3304 1280 3307
rect 1267 3293 1284 3304
rect 347 3276 484 3280
rect 756 3247 764 3293
rect 856 3284 864 3293
rect 856 3276 933 3284
rect 796 3247 804 3273
rect 1116 3264 1124 3274
rect 1176 3264 1184 3274
rect 847 3256 1124 3264
rect 1156 3260 1184 3264
rect 1153 3256 1184 3260
rect 1153 3247 1167 3256
rect 67 3236 93 3244
rect 107 3236 233 3244
rect 247 3236 553 3244
rect 1276 3247 1284 3293
rect 1513 3284 1527 3293
rect 1476 3280 1527 3284
rect 1576 3296 1633 3304
rect 1476 3276 1524 3280
rect 1476 3264 1484 3276
rect 1576 3267 1584 3296
rect 1656 3296 1753 3304
rect 1327 3256 1484 3264
rect 1507 3255 1533 3263
rect 1656 3266 1664 3296
rect 2447 3297 2513 3305
rect 2567 3296 2693 3304
rect 2767 3296 2833 3304
rect 1736 3276 1953 3284
rect 1736 3266 1744 3276
rect 1907 3256 1973 3264
rect 2387 3256 2413 3264
rect 3053 3264 3067 3273
rect 3316 3284 3324 3316
rect 4207 3316 4233 3324
rect 4247 3316 4573 3324
rect 4847 3316 4913 3324
rect 5027 3316 5053 3324
rect 5227 3316 5293 3324
rect 3476 3296 3653 3304
rect 3227 3276 3324 3284
rect 3347 3276 3464 3284
rect 3036 3260 3067 3264
rect 3036 3256 3064 3260
rect 1276 3236 1293 3247
rect 1280 3233 1293 3236
rect 1347 3236 1373 3244
rect 1387 3236 1453 3244
rect 1736 3244 1744 3252
rect 1627 3236 1744 3244
rect 2007 3236 2033 3244
rect 2127 3236 2253 3244
rect 2307 3236 2473 3244
rect 2487 3236 2733 3244
rect 3036 3244 3044 3256
rect 2847 3236 3044 3244
rect 187 3216 473 3224
rect 556 3224 564 3233
rect 3387 3235 3413 3243
rect 3456 3245 3464 3276
rect 3476 3266 3484 3296
rect 3767 3296 3793 3304
rect 3867 3296 3913 3304
rect 4047 3296 4133 3304
rect 4187 3296 4393 3304
rect 4487 3297 4693 3305
rect 3796 3267 3804 3293
rect 3527 3256 3633 3264
rect 4636 3266 4644 3297
rect 4747 3296 4764 3304
rect 4756 3267 4764 3296
rect 4907 3296 4944 3304
rect 4936 3267 4944 3296
rect 3987 3256 4113 3264
rect 4127 3255 4313 3263
rect 4407 3255 4453 3263
rect 4887 3255 4912 3263
rect 4976 3264 4984 3294
rect 5087 3304 5100 3307
rect 5087 3293 5104 3304
rect 5127 3297 5173 3305
rect 5247 3300 5344 3304
rect 5247 3296 5347 3300
rect 5096 3267 5104 3293
rect 5333 3286 5347 3296
rect 5527 3296 5593 3304
rect 5620 3304 5633 3307
rect 5616 3293 5633 3304
rect 5660 3304 5673 3307
rect 5656 3293 5673 3304
rect 5616 3284 5624 3293
rect 5576 3276 5624 3284
rect 4976 3256 5033 3264
rect 5107 3256 5153 3264
rect 5576 3266 5584 3276
rect 5656 3267 5664 3293
rect 5267 3256 5313 3264
rect 5327 3255 5353 3263
rect 5647 3256 5664 3267
rect 5647 3253 5660 3256
rect 3456 3231 3473 3245
rect 3876 3244 3884 3252
rect 5716 3247 5724 3294
rect 5807 3296 5833 3304
rect 6067 3296 6133 3304
rect 6147 3297 6213 3305
rect 5876 3264 5884 3294
rect 5747 3256 5884 3264
rect 3856 3236 3884 3244
rect 556 3216 773 3224
rect 2276 3216 3313 3224
rect 667 3196 764 3204
rect 507 3176 533 3184
rect 756 3184 764 3196
rect 2276 3204 2284 3216
rect 3327 3216 3613 3224
rect 3856 3224 3864 3236
rect 3927 3236 3953 3244
rect 4547 3236 4693 3244
rect 5507 3236 5564 3244
rect 3687 3216 3864 3224
rect 3947 3216 4093 3224
rect 4107 3216 4153 3224
rect 4567 3216 4673 3224
rect 4687 3216 4833 3224
rect 5107 3216 5173 3224
rect 5556 3224 5564 3236
rect 5556 3216 5613 3224
rect 6047 3216 6213 3224
rect 1787 3196 2284 3204
rect 2667 3196 2773 3204
rect 2787 3196 2913 3204
rect 3667 3196 4353 3204
rect 5227 3196 5473 3204
rect 5747 3196 5973 3204
rect 756 3176 933 3184
rect 1167 3176 1333 3184
rect 2247 3176 2393 3184
rect 2547 3176 2892 3184
rect 2916 3184 2924 3193
rect 2916 3176 3513 3184
rect 3787 3176 4053 3184
rect 4467 3176 4744 3184
rect 967 3156 1133 3164
rect 1227 3156 1253 3164
rect 2647 3156 2673 3164
rect 3027 3156 3433 3164
rect 3596 3156 3853 3164
rect 787 3136 893 3144
rect 1827 3136 1893 3144
rect 3596 3144 3604 3156
rect 4107 3156 4393 3164
rect 4407 3156 4533 3164
rect 4736 3164 4744 3176
rect 4767 3176 4953 3184
rect 4967 3176 5133 3184
rect 5527 3176 5813 3184
rect 5907 3176 6193 3184
rect 4736 3156 5213 3164
rect 5256 3156 5473 3164
rect 2607 3136 3604 3144
rect 4116 3136 4333 3144
rect 267 3116 333 3124
rect 507 3116 833 3124
rect 927 3116 1413 3124
rect 1467 3116 1773 3124
rect 2087 3116 2113 3124
rect 2347 3116 2484 3124
rect 687 3096 713 3104
rect 1227 3096 1293 3104
rect 1567 3096 1593 3104
rect 1707 3096 1733 3104
rect 2476 3104 2484 3116
rect 2827 3116 2953 3124
rect 3207 3116 3553 3124
rect 3596 3116 3813 3124
rect 3596 3107 3604 3116
rect 4116 3124 4124 3136
rect 4516 3136 4593 3144
rect 3867 3116 4124 3124
rect 4516 3124 4524 3136
rect 4607 3136 4633 3144
rect 4787 3136 4973 3144
rect 5256 3144 5264 3156
rect 5667 3156 5793 3164
rect 5127 3136 5264 3144
rect 5427 3136 5893 3144
rect 4147 3116 4524 3124
rect 4547 3116 5052 3124
rect 5087 3116 5633 3124
rect 5927 3116 6093 3124
rect 2476 3096 2753 3104
rect 2847 3096 3593 3104
rect 4227 3096 4453 3104
rect 5407 3096 5553 3104
rect 5727 3096 5773 3104
rect 5787 3096 5853 3104
rect 5867 3096 6073 3104
rect 887 3076 1313 3084
rect 1587 3076 1624 3084
rect 87 3056 193 3064
rect 867 3056 1233 3064
rect 1616 3047 1624 3076
rect 2416 3076 2453 3084
rect 1707 3056 1833 3064
rect 2416 3047 2424 3076
rect 3467 3076 3632 3084
rect 3667 3076 3893 3084
rect 3907 3076 4113 3084
rect 4236 3076 4453 3084
rect 2747 3056 3193 3064
rect 3216 3056 3353 3064
rect 947 3044 960 3047
rect 947 3033 964 3044
rect 1767 3036 1813 3044
rect 1827 3036 2173 3044
rect 2187 3036 2273 3044
rect 3216 3044 3224 3056
rect 3567 3056 3673 3064
rect 4236 3064 4244 3076
rect 4927 3076 5133 3084
rect 5207 3076 5693 3084
rect 3687 3056 4244 3064
rect 4287 3056 4333 3064
rect 4627 3056 4813 3064
rect 5287 3056 5373 3064
rect 5747 3056 5793 3064
rect 5956 3056 5993 3064
rect 2767 3036 3224 3044
rect 3507 3036 3693 3044
rect 4056 3036 4093 3044
rect 956 3024 964 3033
rect 956 3016 1053 3024
rect 1287 3016 1313 3024
rect 2196 3016 2253 3024
rect 47 2997 93 3005
rect 687 2996 753 3004
rect 767 2996 813 3004
rect 407 2976 544 2984
rect 127 2955 153 2963
rect 536 2964 544 2976
rect 876 2967 884 3013
rect 916 2967 924 3013
rect 1216 2987 1224 3013
rect 1607 2996 1724 3004
rect 536 2956 693 2964
rect 796 2960 833 2964
rect 793 2956 833 2960
rect 793 2947 807 2956
rect 907 2956 924 2967
rect 907 2953 920 2956
rect 1036 2944 1044 2973
rect 1367 2975 1453 2983
rect 1716 2964 1724 2996
rect 1736 2987 1744 3013
rect 1796 2987 1804 3013
rect 1887 2976 1973 2984
rect 2196 2984 2204 3016
rect 3267 3017 3373 3025
rect 3836 3016 4013 3024
rect 3427 2996 3653 3004
rect 3836 3004 3844 3016
rect 3727 2996 3844 3004
rect 3867 2996 4004 3004
rect 2147 2976 2204 2984
rect 2433 2984 2447 2993
rect 2307 2976 2593 2984
rect 2687 2975 2893 2983
rect 3227 2976 3313 2984
rect 1716 2956 1833 2964
rect 2227 2956 2273 2964
rect 3436 2956 3513 2964
rect 3436 2947 3444 2956
rect 3647 2955 3693 2963
rect 3827 2956 3953 2964
rect 3996 2947 4004 2996
rect 4036 2967 4044 2993
rect 4056 2947 4064 3036
rect 4267 3036 4513 3044
rect 4667 3036 4713 3044
rect 4947 3036 4993 3044
rect 5087 3036 5173 3044
rect 5227 3036 5293 3044
rect 5956 3044 5964 3056
rect 5707 3036 5964 3044
rect 5987 3036 6144 3044
rect 4436 3016 4553 3024
rect 4147 2996 4213 3004
rect 4227 2997 4313 3005
rect 4436 3007 4444 3016
rect 4647 3016 4853 3024
rect 5067 3016 5153 3024
rect 5267 3016 5433 3024
rect 5707 3016 5893 3024
rect 4096 2984 4104 2994
rect 4507 2996 4593 3004
rect 4747 2997 4773 3005
rect 4796 2996 4973 3004
rect 4096 2980 4164 2984
rect 4096 2976 4167 2980
rect 4153 2967 4167 2976
rect 4187 2976 4613 2984
rect 4327 2956 4413 2964
rect 4467 2960 4564 2964
rect 4467 2956 4567 2960
rect 4553 2947 4567 2956
rect 4627 2955 4673 2963
rect 947 2936 1044 2944
rect 1307 2936 1393 2944
rect 1856 2936 2153 2944
rect 1856 2924 1864 2936
rect 2327 2936 2713 2944
rect 2887 2936 3433 2944
rect 3536 2936 3713 2944
rect 1447 2916 1864 2924
rect 2907 2916 3233 2924
rect 3536 2924 3544 2936
rect 3987 2936 4004 2947
rect 3987 2933 4000 2936
rect 4447 2936 4473 2944
rect 4696 2944 4704 2994
rect 4796 2967 4804 2996
rect 5247 2997 5273 3005
rect 5347 2996 5413 3004
rect 5496 2996 5593 3004
rect 4887 2956 4913 2964
rect 5027 2955 5053 2963
rect 5196 2964 5204 2993
rect 5496 2984 5504 2996
rect 6136 3004 6144 3036
rect 6136 2996 6153 3004
rect 5167 2956 5204 2964
rect 5396 2976 5504 2984
rect 4696 2936 4813 2944
rect 5396 2944 5404 2976
rect 5676 2967 5684 2993
rect 5527 2955 5573 2963
rect 5776 2964 5784 2993
rect 6036 2984 6044 2994
rect 6016 2976 6044 2984
rect 5767 2956 5784 2964
rect 6016 2964 6024 2976
rect 6176 2966 6184 3033
rect 5927 2956 6024 2964
rect 5347 2936 5404 2944
rect 5467 2936 5833 2944
rect 3367 2916 3544 2924
rect 3967 2916 4172 2924
rect 4207 2916 4353 2924
rect 4507 2916 4773 2924
rect 4887 2916 5233 2924
rect 5416 2916 5493 2924
rect 47 2896 653 2904
rect 2036 2900 2293 2904
rect 2033 2896 2293 2900
rect 2033 2887 2047 2896
rect 3347 2896 3573 2904
rect 3807 2896 3993 2904
rect 4307 2896 4333 2904
rect 4407 2896 4453 2904
rect 4647 2896 4713 2904
rect 4787 2896 4833 2904
rect 5116 2896 5313 2904
rect 227 2876 293 2884
rect 307 2876 493 2884
rect 1247 2876 1433 2884
rect 2567 2876 2613 2884
rect 2627 2876 2913 2884
rect 3067 2876 3733 2884
rect 4167 2876 4193 2884
rect 4287 2876 5073 2884
rect 5116 2884 5124 2896
rect 5416 2904 5424 2916
rect 5727 2916 5873 2924
rect 5387 2896 5424 2904
rect 5436 2896 5593 2904
rect 5087 2876 5124 2884
rect 5436 2884 5444 2896
rect 6107 2896 6213 2904
rect 5267 2876 5444 2884
rect 5456 2876 5713 2884
rect 907 2856 1053 2864
rect 1687 2856 1833 2864
rect 2107 2856 2173 2864
rect 2627 2856 2813 2864
rect 3867 2856 4113 2864
rect 4127 2856 4233 2864
rect 4567 2856 4624 2864
rect 67 2836 473 2844
rect 607 2836 833 2844
rect 847 2836 873 2844
rect 1187 2836 1253 2844
rect 1567 2836 1793 2844
rect 2607 2836 2864 2844
rect 2856 2827 2864 2836
rect 3947 2836 3973 2844
rect 3987 2836 4013 2844
rect 4367 2836 4493 2844
rect 4547 2836 4573 2844
rect 4616 2844 4624 2856
rect 4647 2856 4793 2864
rect 5187 2856 5233 2864
rect 5456 2864 5464 2876
rect 5927 2876 6153 2884
rect 5247 2856 5464 2864
rect 5487 2856 5613 2864
rect 5727 2856 5793 2864
rect 6127 2856 6193 2864
rect 4616 2836 4773 2844
rect 4967 2836 5052 2844
rect 5087 2836 5604 2844
rect 5596 2827 5604 2836
rect 6067 2836 6233 2844
rect 547 2816 613 2824
rect 667 2816 753 2824
rect 807 2816 913 2824
rect 1487 2816 1693 2824
rect 1707 2816 1993 2824
rect 2167 2816 2553 2824
rect 2576 2816 2753 2824
rect 67 2796 253 2804
rect 447 2796 513 2804
rect 927 2796 953 2804
rect 1047 2796 1073 2804
rect 1087 2796 1233 2804
rect 1333 2804 1347 2813
rect 1247 2800 1347 2804
rect 1247 2796 1344 2800
rect 1447 2796 1653 2804
rect 1707 2796 1773 2804
rect 1847 2796 1933 2804
rect 2576 2804 2584 2816
rect 2867 2816 2973 2824
rect 2987 2816 3373 2824
rect 3727 2816 3813 2824
rect 4107 2816 4213 2824
rect 4267 2816 4333 2824
rect 4607 2816 4793 2824
rect 4807 2816 4973 2824
rect 5047 2816 5273 2824
rect 5596 2816 5613 2827
rect 5600 2813 5613 2816
rect 5687 2816 5753 2824
rect 2527 2796 2584 2804
rect 3547 2796 3613 2804
rect 3627 2796 3864 2804
rect 27 2777 353 2785
rect 407 2776 424 2784
rect 416 2747 424 2776
rect 787 2776 812 2784
rect 847 2776 973 2784
rect 1147 2777 1193 2785
rect 1287 2776 1344 2784
rect 976 2747 984 2774
rect 1336 2764 1344 2776
rect 1367 2776 1413 2784
rect 1547 2776 1733 2784
rect 1747 2776 1832 2784
rect 1867 2776 1973 2784
rect 2136 2776 2153 2784
rect 1336 2756 1433 2764
rect 2136 2747 2144 2776
rect 2267 2780 2364 2784
rect 2267 2776 2367 2780
rect 2353 2767 2367 2776
rect 2747 2776 2773 2784
rect 3047 2777 3113 2785
rect 3247 2776 3333 2784
rect 3747 2776 3833 2784
rect 3856 2784 3864 2796
rect 3967 2796 4033 2804
rect 4667 2796 4693 2804
rect 5147 2796 5293 2804
rect 5307 2796 5373 2804
rect 5427 2796 5453 2804
rect 5887 2796 5913 2804
rect 3856 2776 4093 2784
rect 4187 2776 4253 2784
rect 4276 2764 4284 2793
rect 4307 2776 4333 2784
rect 4407 2776 4513 2784
rect 4620 2784 4633 2787
rect 4616 2773 4633 2784
rect 4747 2776 4844 2784
rect 4276 2756 4373 2764
rect -63 2736 73 2744
rect 667 2735 713 2743
rect 887 2735 913 2743
rect 967 2736 984 2747
rect 967 2733 980 2736
rect 1087 2735 1113 2743
rect 1136 2736 1533 2744
rect 1136 2724 1144 2736
rect 1807 2735 1853 2743
rect 2387 2736 2573 2744
rect 2727 2736 2833 2744
rect 3027 2736 3093 2744
rect 3107 2736 3193 2744
rect 4047 2736 4193 2744
rect 4207 2736 4273 2744
rect 4327 2735 4353 2743
rect 4556 2744 4564 2773
rect 4616 2746 4624 2773
rect 4836 2747 4844 2776
rect 4876 2764 4884 2774
rect 4927 2776 4964 2784
rect 4876 2756 4944 2764
rect 4556 2736 4573 2744
rect 4767 2735 4793 2743
rect 1027 2716 1144 2724
rect 215 2686 223 2713
rect 1547 2716 1673 2724
rect 2107 2715 2213 2723
rect 3487 2716 3693 2724
rect 3767 2716 4013 2724
rect 4507 2716 4593 2724
rect 4716 2724 4724 2732
rect 4639 2716 4724 2724
rect 4936 2724 4944 2756
rect 4956 2747 4964 2776
rect 5036 2747 5044 2773
rect 5356 2747 5364 2773
rect 5487 2776 5553 2784
rect 5607 2776 5673 2784
rect 5796 2776 5833 2784
rect 5796 2764 5804 2776
rect 6027 2777 6073 2785
rect 5087 2736 5113 2744
rect 5127 2736 5273 2744
rect 5373 2744 5387 2753
rect 5736 2756 5804 2764
rect 5736 2746 5744 2756
rect 5896 2747 5904 2773
rect 5373 2740 5433 2744
rect 5376 2736 5433 2740
rect 5447 2736 5533 2744
rect 5947 2735 5993 2743
rect 4936 2716 5153 2724
rect 527 2696 873 2704
rect 967 2696 993 2704
rect 1007 2696 1253 2704
rect 1307 2696 1473 2704
rect 1707 2696 1813 2704
rect 1927 2696 2113 2704
rect 2827 2696 2953 2704
rect 3607 2696 3664 2704
rect -63 2678 223 2686
rect 347 2676 533 2684
rect 947 2676 1393 2684
rect 1867 2676 2273 2684
rect 2287 2676 2953 2684
rect 3367 2676 3393 2684
rect 3407 2676 3493 2684
rect 3596 2684 3604 2693
rect 3507 2676 3604 2684
rect 3656 2684 3664 2696
rect 3847 2696 4213 2704
rect 4467 2696 4613 2704
rect 3656 2676 3873 2684
rect 3947 2676 4173 2684
rect 4639 2684 4647 2716
rect 5167 2716 5613 2724
rect 5627 2716 5773 2724
rect 5787 2716 5853 2724
rect 5927 2716 6033 2724
rect 5007 2696 5133 2704
rect 5187 2696 5313 2704
rect 5327 2696 5573 2704
rect 5667 2696 5813 2704
rect 4327 2676 4647 2684
rect 4767 2676 4933 2684
rect 5196 2676 5432 2684
rect 5196 2667 5204 2676
rect 5467 2676 5573 2684
rect 147 2656 1513 2664
rect 1767 2656 1913 2664
rect 2167 2656 2813 2664
rect 3647 2656 3993 2664
rect 4087 2656 4153 2664
rect 4176 2656 4653 2664
rect 287 2636 453 2644
rect 467 2636 1013 2644
rect 1247 2636 1493 2644
rect 1987 2636 2033 2644
rect 2187 2636 2513 2644
rect 3687 2636 3973 2644
rect 4176 2644 4184 2656
rect 4807 2656 5193 2664
rect 5247 2656 5593 2664
rect 5667 2656 5893 2664
rect 3987 2636 4184 2644
rect 4527 2636 4773 2644
rect 4847 2636 5113 2644
rect 5356 2636 5373 2644
rect 347 2616 433 2624
rect 767 2616 1073 2624
rect 1527 2616 2073 2624
rect 3787 2616 3833 2624
rect 4067 2616 4313 2624
rect 5356 2624 5364 2636
rect 5387 2636 5452 2644
rect 5487 2636 6073 2644
rect 6087 2636 6133 2644
rect 5207 2616 5364 2624
rect 5676 2616 5893 2624
rect 207 2596 1233 2604
rect 1667 2596 1713 2604
rect 2107 2596 2313 2604
rect 2327 2596 2633 2604
rect 2647 2596 2733 2604
rect 2747 2596 3053 2604
rect 3667 2596 3853 2604
rect 3867 2596 4413 2604
rect 4427 2596 4453 2604
rect 4627 2596 4793 2604
rect 4847 2596 5033 2604
rect 5676 2604 5684 2616
rect 5387 2596 5684 2604
rect 287 2576 373 2584
rect 1067 2576 1093 2584
rect 1447 2576 1473 2584
rect 1487 2576 1813 2584
rect 1827 2576 1973 2584
rect 2607 2576 2773 2584
rect 3387 2576 3753 2584
rect 3887 2576 4173 2584
rect 4267 2576 4413 2584
rect 4667 2576 4773 2584
rect 4827 2576 5153 2584
rect 5447 2576 5693 2584
rect 827 2556 1033 2564
rect 1467 2556 1613 2564
rect 2027 2556 2133 2564
rect 2147 2556 3113 2564
rect 3487 2556 3613 2564
rect 4027 2556 4753 2564
rect 4767 2556 4853 2564
rect 5407 2556 5533 2564
rect 727 2536 1273 2544
rect 1887 2536 2173 2544
rect 2227 2536 2533 2544
rect 3116 2544 3124 2553
rect 3116 2536 3633 2544
rect 3927 2536 4073 2544
rect 4087 2536 4293 2544
rect 4607 2536 4633 2544
rect 4647 2536 4713 2544
rect 1087 2516 1173 2524
rect 1387 2516 1453 2524
rect 1467 2516 1553 2524
rect 1867 2516 2033 2524
rect 2427 2516 2513 2524
rect 2647 2516 2873 2524
rect 3047 2516 3673 2524
rect 3976 2516 4053 2524
rect 247 2496 293 2504
rect 307 2496 513 2504
rect 827 2496 873 2504
rect 1027 2496 1144 2504
rect -63 2476 113 2484
rect 327 2477 353 2485
rect 407 2476 444 2484
rect 436 2447 444 2476
rect 467 2484 480 2487
rect 467 2473 484 2484
rect 476 2466 484 2473
rect 1113 2464 1127 2473
rect 847 2460 1127 2464
rect 847 2456 1124 2460
rect 436 2436 453 2447
rect 440 2433 453 2436
rect 867 2436 973 2444
rect 1016 2436 1112 2444
rect 167 2416 373 2424
rect 387 2416 573 2424
rect 587 2416 833 2424
rect 1016 2424 1024 2436
rect 1136 2446 1144 2496
rect 1407 2496 1583 2504
rect 1575 2488 1583 2496
rect 2067 2496 2273 2504
rect 3976 2504 3984 2516
rect 4227 2516 4493 2524
rect 4847 2516 4893 2524
rect 4907 2516 5293 2524
rect 5307 2516 5413 2524
rect 5587 2516 5673 2524
rect 6007 2516 6093 2524
rect 3767 2496 3984 2504
rect 4167 2496 4204 2504
rect 1167 2476 1233 2484
rect 1387 2476 1413 2484
rect 1496 2476 1533 2484
rect 847 2416 1024 2424
rect 1047 2416 1093 2424
rect 1316 2424 1324 2473
rect 1496 2464 1504 2476
rect 1667 2476 1713 2484
rect 1476 2456 1504 2464
rect 1476 2427 1484 2456
rect 1576 2444 1584 2474
rect 1787 2477 1833 2485
rect 1847 2476 1933 2484
rect 2047 2476 2153 2484
rect 2487 2476 2632 2484
rect 2807 2476 2913 2484
rect 2927 2476 2993 2484
rect 3227 2476 3253 2484
rect 3267 2477 3293 2485
rect 3347 2476 3413 2484
rect 3427 2476 3573 2484
rect 3676 2476 3733 2484
rect 1993 2464 2007 2473
rect 1993 2460 2224 2464
rect 1996 2456 2224 2460
rect 1576 2436 1673 2444
rect 1727 2435 1753 2443
rect 1807 2436 1873 2444
rect 2007 2436 2193 2444
rect 2216 2427 2224 2456
rect 2653 2464 2667 2473
rect 2387 2460 2667 2464
rect 2387 2456 2664 2460
rect 3676 2464 3684 2476
rect 3807 2476 3924 2484
rect 2967 2456 3684 2464
rect 3707 2456 3833 2464
rect 3916 2464 3924 2476
rect 3947 2476 3993 2484
rect 4047 2476 4113 2484
rect 4196 2484 4204 2496
rect 4607 2496 4673 2504
rect 5767 2496 5813 2504
rect 4196 2476 4213 2484
rect 4227 2476 4333 2484
rect 4467 2476 4553 2484
rect 4920 2484 4933 2487
rect 4416 2464 4424 2474
rect 4916 2473 4933 2484
rect 5087 2477 5113 2485
rect 3916 2456 3964 2464
rect 4416 2456 4604 2464
rect 2287 2435 2453 2443
rect 2567 2436 2673 2444
rect 2787 2435 2833 2443
rect 3067 2436 3113 2444
rect 3127 2435 3153 2443
rect 3207 2436 3513 2444
rect 3647 2435 3673 2443
rect 3956 2427 3964 2456
rect 3987 2435 4013 2443
rect 4156 2436 4324 2444
rect 1316 2416 1413 2424
rect 1467 2416 1484 2427
rect 1467 2413 1480 2416
rect 1527 2416 1553 2424
rect 3956 2426 3980 2427
rect 3956 2416 3973 2426
rect 3960 2413 3973 2416
rect 4156 2424 4164 2436
rect 4047 2416 4164 2424
rect 4316 2424 4324 2436
rect 4507 2435 4533 2443
rect 4547 2435 4573 2443
rect 4596 2444 4604 2456
rect 4916 2446 4924 2473
rect 4596 2436 4613 2444
rect 4627 2436 4733 2444
rect 4996 2427 5004 2474
rect 5236 2476 5253 2484
rect 5196 2444 5204 2473
rect 5236 2447 5244 2476
rect 5556 2476 5573 2484
rect 5373 2464 5387 2473
rect 5356 2460 5387 2464
rect 5356 2456 5384 2460
rect 5187 2436 5204 2444
rect 4316 2416 4473 2424
rect 4687 2416 4813 2424
rect 5087 2416 5153 2424
rect 5356 2424 5364 2456
rect 5456 2447 5464 2473
rect 5376 2440 5433 2444
rect 5287 2416 5364 2424
rect 5373 2436 5433 2440
rect 5373 2427 5387 2436
rect 5456 2436 5473 2447
rect 5460 2433 5473 2436
rect 5556 2427 5564 2476
rect 5596 2446 5604 2493
rect 5653 2484 5667 2493
rect 5636 2480 5667 2484
rect 5636 2476 5664 2480
rect 5636 2447 5644 2476
rect 5707 2484 5720 2487
rect 5707 2473 5724 2484
rect 5907 2476 6033 2484
rect 5716 2446 5724 2473
rect 5767 2436 5973 2444
rect 5556 2416 5573 2427
rect 5560 2413 5573 2416
rect 5847 2416 5893 2424
rect 1507 2396 1912 2404
rect 1947 2396 2073 2404
rect 2127 2396 2333 2404
rect 2347 2396 2573 2404
rect 2627 2396 2713 2404
rect 3447 2396 3653 2404
rect 3856 2396 4693 2404
rect 887 2376 1373 2384
rect 1427 2376 1993 2384
rect 2507 2376 2773 2384
rect 3107 2376 3673 2384
rect 3856 2384 3864 2396
rect 5096 2396 5144 2404
rect 3827 2376 3864 2384
rect 3947 2376 4033 2384
rect 5096 2384 5104 2396
rect 5007 2376 5104 2384
rect 5136 2384 5144 2396
rect 6027 2396 6124 2404
rect 5136 2376 5253 2384
rect 5607 2376 5813 2384
rect 6116 2384 6124 2396
rect 6116 2376 6173 2384
rect 207 2356 753 2364
rect 1127 2356 1253 2364
rect 1707 2356 1733 2364
rect 1747 2356 1853 2364
rect 2187 2356 2273 2364
rect 2496 2364 2504 2373
rect 2287 2356 2504 2364
rect 3567 2356 3613 2364
rect 3727 2356 3753 2364
rect 4067 2356 4093 2364
rect 4167 2356 4273 2364
rect 4287 2356 4333 2364
rect 4447 2356 4673 2364
rect 4687 2356 4792 2364
rect 4827 2356 5113 2364
rect 5127 2356 5313 2364
rect 5327 2356 5393 2364
rect 5447 2356 5693 2364
rect 5787 2356 5913 2364
rect 5927 2356 6053 2364
rect 1407 2336 1533 2344
rect 1807 2336 1953 2344
rect 2247 2336 2353 2344
rect 3507 2336 3633 2344
rect 4087 2336 4793 2344
rect 4807 2336 5013 2344
rect 5027 2336 5133 2344
rect 5147 2336 5233 2344
rect 5667 2336 5753 2344
rect 5807 2336 5833 2344
rect 5847 2336 5873 2344
rect 6107 2336 6213 2344
rect 427 2316 853 2324
rect 987 2316 1013 2324
rect 1027 2316 1113 2324
rect 1347 2316 1513 2324
rect 1567 2316 1873 2324
rect 2867 2316 3013 2324
rect 3667 2316 3693 2324
rect 3707 2316 3753 2324
rect 4327 2316 4393 2324
rect 4507 2316 4753 2324
rect 4816 2316 4853 2324
rect 467 2296 513 2304
rect 1027 2296 1073 2304
rect 1287 2296 1453 2304
rect 1847 2296 2013 2304
rect 2247 2296 2632 2304
rect 2667 2296 2833 2304
rect 3047 2296 3153 2304
rect 3267 2296 3312 2304
rect 3347 2296 3453 2304
rect 3527 2296 3593 2304
rect 3847 2296 3933 2304
rect 4007 2296 4112 2304
rect 4147 2296 4233 2304
rect 4327 2296 4373 2304
rect 4816 2304 4824 2316
rect 5267 2316 5473 2324
rect 5627 2316 5653 2324
rect 5667 2316 6073 2324
rect 4776 2296 4824 2304
rect 767 2276 1044 2284
rect 267 2256 473 2264
rect 827 2256 853 2264
rect 1000 2264 1013 2267
rect 996 2253 1013 2264
rect 1036 2264 1044 2276
rect 1187 2276 1673 2284
rect 2907 2276 2953 2284
rect 3007 2276 3513 2284
rect 3627 2276 3893 2284
rect 1036 2256 1073 2264
rect 1127 2257 1193 2265
rect 1247 2256 1313 2264
rect 1367 2256 1453 2264
rect 1587 2256 1613 2264
rect 2007 2256 2053 2264
rect 2096 2256 2133 2264
rect 427 2236 453 2244
rect 527 2235 653 2243
rect 847 2236 944 2244
rect 327 2216 353 2224
rect 936 2224 944 2236
rect 996 2226 1004 2253
rect 2096 2227 2104 2256
rect 2160 2264 2173 2267
rect 2156 2253 2173 2264
rect 2227 2256 2313 2264
rect 2327 2256 2453 2264
rect 936 2216 953 2224
rect 1067 2215 1093 2223
rect 1847 2216 1953 2224
rect 2156 2226 2164 2253
rect 2596 2244 2604 2254
rect 2727 2256 2744 2264
rect 2496 2236 2604 2244
rect 2407 2215 2433 2223
rect 2496 2224 2504 2236
rect 2636 2227 2644 2253
rect 2736 2244 2744 2256
rect 2767 2256 2793 2264
rect 2927 2256 2984 2264
rect 2976 2244 2984 2256
rect 3107 2257 3193 2265
rect 3307 2257 3373 2265
rect 2736 2236 2844 2244
rect 2976 2236 3104 2244
rect 2487 2216 2504 2224
rect 2836 2226 2844 2236
rect 827 2195 853 2203
rect 1227 2196 1333 2204
rect 1427 2196 1693 2204
rect 2007 2196 2044 2204
rect 1007 2176 1033 2184
rect 1387 2176 1573 2184
rect 1587 2176 1973 2184
rect 2036 2184 2044 2196
rect 2467 2196 2513 2204
rect 2567 2196 2593 2204
rect 3096 2204 3104 2236
rect 3127 2216 3313 2224
rect 3393 2224 3407 2233
rect 3367 2220 3407 2224
rect 3367 2216 3404 2220
rect 3556 2207 3564 2254
rect 3576 2226 3584 2273
rect 3716 2268 3724 2276
rect 3987 2276 4273 2284
rect 4347 2276 4713 2284
rect 4776 2284 4784 2296
rect 5687 2296 5733 2304
rect 5893 2306 5907 2316
rect 6007 2296 6053 2304
rect 6147 2296 6213 2304
rect 4756 2276 4784 2284
rect 3687 2264 3700 2267
rect 3687 2253 3704 2264
rect 3767 2256 3884 2264
rect 3696 2226 3704 2253
rect 3716 2224 3724 2254
rect 3716 2216 3793 2224
rect 3876 2226 3884 2256
rect 4116 2256 4153 2264
rect 4116 2227 4124 2256
rect 4256 2227 4264 2253
rect 4456 2224 4464 2254
rect 4567 2256 4613 2264
rect 4636 2256 4693 2264
rect 4636 2226 4644 2256
rect 4756 2227 4764 2276
rect 4847 2276 4913 2284
rect 5187 2276 5213 2284
rect 5327 2276 5353 2284
rect 5467 2276 5493 2284
rect 5516 2276 5613 2284
rect 4807 2264 4820 2267
rect 4807 2253 4824 2264
rect 5033 2264 5047 2273
rect 4967 2260 5047 2264
rect 4967 2256 5044 2260
rect 5287 2256 5344 2264
rect 4816 2244 4824 2253
rect 5336 2244 5344 2256
rect 5516 2264 5524 2276
rect 5676 2276 6113 2284
rect 5387 2256 5524 2264
rect 4816 2236 4844 2244
rect 5336 2236 5364 2244
rect 4347 2216 4464 2224
rect 4547 2215 4593 2223
rect 4836 2226 4844 2236
rect 4927 2215 4973 2223
rect 5027 2216 5093 2224
rect 5107 2216 5153 2224
rect 5167 2216 5213 2224
rect 5356 2224 5364 2236
rect 5536 2244 5544 2254
rect 5487 2236 5544 2244
rect 5356 2216 5633 2224
rect 5676 2226 5684 2276
rect 5747 2256 5804 2264
rect 3096 2196 3173 2204
rect 4407 2196 4473 2204
rect 5796 2204 5804 2256
rect 5816 2256 5893 2264
rect 5816 2226 5824 2256
rect 5936 2227 5944 2253
rect 5976 2207 5984 2254
rect 5996 2226 6004 2276
rect 6127 2276 6164 2284
rect 6016 2244 6024 2254
rect 6016 2240 6044 2244
rect 6016 2236 6047 2240
rect 6033 2227 6047 2236
rect 6156 2226 6164 2276
rect 6087 2215 6113 2223
rect 5796 2196 5853 2204
rect 2036 2176 2113 2184
rect 2127 2176 2193 2184
rect 2427 2176 2513 2184
rect 2707 2176 2873 2184
rect 3907 2176 3953 2184
rect 4107 2176 4193 2184
rect 4327 2176 4353 2184
rect 4407 2176 4433 2184
rect 4607 2176 4633 2184
rect 4787 2176 4873 2184
rect 4887 2176 5253 2184
rect 5647 2176 5773 2184
rect 287 2156 393 2164
rect 1147 2156 1313 2164
rect 1387 2156 1873 2164
rect 2027 2156 2213 2164
rect 2387 2156 2653 2164
rect 2787 2156 3573 2164
rect 3687 2156 3732 2164
rect 3767 2156 3973 2164
rect 3987 2156 4033 2164
rect 4107 2156 4373 2164
rect 4387 2156 4513 2164
rect 4587 2156 4733 2164
rect 5587 2156 6033 2164
rect 1447 2136 1633 2144
rect 1747 2136 1813 2144
rect 1896 2136 1993 2144
rect 1896 2124 1904 2136
rect 2047 2136 2173 2144
rect 2267 2136 4592 2144
rect 4627 2136 4673 2144
rect 4807 2136 5353 2144
rect 5367 2136 5473 2144
rect 1687 2116 1904 2124
rect 2047 2116 2173 2124
rect 2807 2116 3013 2124
rect 3127 2116 3533 2124
rect 3707 2116 3893 2124
rect 3947 2116 4112 2124
rect 4147 2116 4633 2124
rect 4707 2116 5393 2124
rect 767 2096 1073 2104
rect 1207 2096 1473 2104
rect 1987 2096 2113 2104
rect 2207 2096 2353 2104
rect 2367 2096 2453 2104
rect 3667 2096 3753 2104
rect 3927 2096 4093 2104
rect 4207 2096 4533 2104
rect 4716 2096 5033 2104
rect 1267 2076 2013 2084
rect 2487 2076 2793 2084
rect 2967 2076 3413 2084
rect 3547 2076 3833 2084
rect 4207 2076 4273 2084
rect 4716 2084 4724 2096
rect 4687 2076 4724 2084
rect 5187 2076 5453 2084
rect 5607 2076 5833 2084
rect 47 2056 113 2064
rect 347 2056 453 2064
rect 1467 2056 1593 2064
rect 1707 2056 1833 2064
rect 1887 2056 2073 2064
rect 2087 2056 2152 2064
rect 2187 2056 2273 2064
rect 2287 2056 2944 2064
rect 2936 2047 2944 2056
rect 3147 2056 3353 2064
rect 3727 2056 3873 2064
rect 5927 2056 6113 2064
rect 1107 2036 1153 2044
rect 1807 2036 1913 2044
rect 1967 2036 2013 2044
rect 2067 2036 2473 2044
rect 2947 2036 3013 2044
rect 3027 2036 3053 2044
rect 3747 2036 3773 2044
rect 4027 2036 4273 2044
rect 4347 2036 4553 2044
rect 5547 2036 5613 2044
rect 5787 2036 5953 2044
rect 267 2016 313 2024
rect 327 2016 453 2024
rect 1007 2016 1073 2024
rect 1587 2016 1804 2024
rect 147 1996 233 2004
rect 387 1996 933 2004
rect 1547 1996 1773 2004
rect 1796 2004 1804 2016
rect 1907 2016 2172 2024
rect 2207 2016 2373 2024
rect 2447 2016 2533 2024
rect 3467 2016 3753 2024
rect 4167 2016 4353 2024
rect 4707 2016 4853 2024
rect 4867 2016 4893 2024
rect 5147 2016 5473 2024
rect 1796 1996 2033 2004
rect 2647 1996 2733 2004
rect 2967 1996 3213 2004
rect 3227 1996 3233 2004
rect 3327 1996 3373 2004
rect 3567 1996 3793 2004
rect 4847 1996 4993 2004
rect 5247 1996 5313 2004
rect 5567 1996 5653 2004
rect 5916 1996 5933 2004
rect 227 1976 264 1984
rect 107 1956 193 1964
rect 56 1927 64 1953
rect 256 1926 264 1976
rect 667 1976 973 1984
rect 1013 1984 1027 1993
rect 996 1980 1027 1984
rect 996 1976 1024 1980
rect 276 1944 284 1954
rect 996 1964 1004 1976
rect 1976 1976 2093 1984
rect 407 1956 464 1964
rect 836 1960 1004 1964
rect 276 1936 433 1944
rect 456 1944 464 1956
rect 833 1956 1004 1960
rect 833 1947 847 1956
rect 1027 1957 1053 1965
rect 1080 1964 1093 1967
rect 456 1936 493 1944
rect 1076 1953 1093 1964
rect 1156 1956 1193 1964
rect 1076 1944 1084 1953
rect 1016 1936 1084 1944
rect 787 1916 853 1924
rect 1016 1924 1024 1936
rect 1156 1926 1164 1956
rect 1347 1956 1413 1964
rect 1427 1956 1444 1964
rect 1436 1944 1444 1956
rect 1467 1956 1573 1964
rect 1656 1944 1664 1954
rect 1436 1936 1664 1944
rect 1007 1916 1024 1924
rect 1307 1915 1333 1923
rect 1647 1915 1733 1923
rect 1796 1907 1804 1973
rect 1927 1956 1964 1964
rect 1827 1915 1893 1923
rect 1956 1924 1964 1956
rect 1976 1944 1984 1976
rect 2627 1976 3093 1984
rect 3107 1976 3153 1984
rect 3267 1976 3293 1984
rect 3507 1976 3673 1984
rect 3987 1984 4000 1987
rect 3987 1973 4004 1984
rect 2007 1956 2044 1964
rect 1976 1940 2024 1944
rect 1976 1936 2027 1940
rect 2013 1927 2027 1936
rect 1956 1916 1984 1924
rect 847 1896 953 1904
rect 1976 1904 1984 1916
rect 2036 1924 2044 1956
rect 2247 1956 2533 1964
rect 2587 1956 2693 1964
rect 2847 1956 3193 1964
rect 2036 1916 2093 1924
rect 2116 1924 2124 1954
rect 3347 1956 3473 1964
rect 3996 1967 4004 1973
rect 4076 1976 4133 1984
rect 3587 1956 3624 1964
rect 2187 1944 2200 1947
rect 3616 1944 3624 1956
rect 3647 1956 3772 1964
rect 3807 1956 3893 1964
rect 2187 1933 2204 1944
rect 3616 1936 3784 1944
rect 2116 1916 2173 1924
rect 2196 1924 2204 1933
rect 2196 1916 2253 1924
rect 2467 1916 2553 1924
rect 2687 1916 2773 1924
rect 2787 1916 2873 1924
rect 2887 1916 2933 1924
rect 3167 1915 3213 1923
rect 3327 1915 3353 1923
rect 3447 1915 3473 1923
rect 3567 1916 3613 1924
rect 3627 1916 3653 1924
rect 3776 1924 3784 1936
rect 3776 1916 3864 1924
rect 3856 1907 3864 1916
rect 4076 1924 4084 1976
rect 4447 1976 4613 1984
rect 4787 1976 4844 1984
rect 4367 1964 4380 1967
rect 4367 1953 4384 1964
rect 4027 1916 4084 1924
rect 4156 1924 4164 1953
rect 4127 1916 4164 1924
rect 4316 1924 4324 1953
rect 4376 1926 4384 1953
rect 4556 1956 4633 1964
rect 4556 1927 4564 1956
rect 4836 1947 4844 1976
rect 5707 1976 5753 1984
rect 4887 1957 4913 1965
rect 5367 1956 5493 1964
rect 5587 1957 5613 1965
rect 5756 1956 5853 1964
rect 4307 1916 4324 1924
rect 4387 1916 4532 1924
rect 4956 1924 4964 1954
rect 4956 1916 5053 1924
rect 5076 1924 5084 1954
rect 5076 1916 5193 1924
rect 5496 1907 5504 1954
rect 5756 1926 5764 1956
rect 5916 1926 5924 1996
rect 5947 1996 6013 2004
rect 5947 1957 5973 1965
rect 6107 1956 6213 1964
rect 5647 1916 5753 1924
rect 5987 1915 6033 1923
rect 1976 1896 2073 1904
rect 3856 1896 3873 1907
rect 3860 1893 3873 1896
rect 3947 1896 3973 1904
rect 4887 1896 5113 1904
rect 47 1876 393 1884
rect 967 1876 1053 1884
rect 1407 1876 1453 1884
rect 1527 1876 1673 1884
rect 1867 1876 1973 1884
rect 2507 1876 2873 1884
rect 3767 1876 4033 1884
rect 4307 1876 4393 1884
rect 4607 1876 4753 1884
rect 4947 1876 4993 1884
rect 5267 1876 5333 1884
rect 5347 1876 5473 1884
rect 596 1860 753 1864
rect 593 1856 753 1860
rect 593 1847 607 1856
rect 2527 1856 2773 1864
rect 3747 1856 3833 1864
rect 3887 1856 4013 1864
rect 4087 1856 4173 1864
rect 4507 1856 4713 1864
rect 5067 1856 5173 1864
rect 5807 1856 5893 1864
rect 5907 1856 5993 1864
rect 347 1836 373 1844
rect 447 1836 553 1844
rect 687 1836 973 1844
rect 1267 1836 1473 1844
rect 1487 1836 1733 1844
rect 1947 1836 2053 1844
rect 2067 1836 2173 1844
rect 2187 1836 2384 1844
rect 107 1816 313 1824
rect 667 1816 873 1824
rect 1216 1820 1433 1824
rect 1213 1816 1433 1820
rect 1213 1807 1227 1816
rect 1507 1816 1593 1824
rect 2107 1816 2193 1824
rect 2376 1824 2384 1836
rect 2407 1836 2473 1844
rect 3407 1836 3653 1844
rect 3787 1836 4153 1844
rect 4167 1836 4613 1844
rect 5207 1836 5293 1844
rect 2376 1816 2473 1824
rect 2827 1816 3113 1824
rect 4287 1816 4433 1824
rect 5107 1816 5153 1824
rect 5407 1816 5433 1824
rect 5447 1816 5533 1824
rect 5547 1816 5793 1824
rect 727 1796 753 1804
rect 1327 1796 1353 1804
rect 1667 1796 1753 1804
rect 2207 1796 2553 1804
rect 3027 1796 3073 1804
rect 3507 1796 3613 1804
rect 3807 1796 3913 1804
rect 4007 1796 4073 1804
rect 4227 1796 4513 1804
rect 4527 1796 4633 1804
rect 4747 1796 4873 1804
rect 5187 1796 5513 1804
rect 647 1776 773 1784
rect 1167 1776 1353 1784
rect 1847 1776 1873 1784
rect 2487 1776 3193 1784
rect 3207 1776 3524 1784
rect 47 1756 73 1764
rect 687 1744 700 1747
rect 687 1733 704 1744
rect 787 1736 833 1744
rect 1027 1737 1113 1745
rect 1247 1744 1260 1747
rect 1247 1733 1264 1744
rect 1287 1736 1324 1744
rect 147 1715 272 1723
rect 307 1716 413 1724
rect 696 1706 704 1733
rect 487 1695 573 1703
rect 956 1704 964 1733
rect 1256 1724 1264 1733
rect 1036 1716 1264 1724
rect 1316 1724 1324 1736
rect 1347 1744 1360 1747
rect 1513 1744 1527 1753
rect 1947 1756 1993 1764
rect 2096 1756 2153 1764
rect 1347 1733 1364 1744
rect 1513 1740 1564 1744
rect 1516 1736 1564 1740
rect 1356 1724 1364 1733
rect 1316 1720 1344 1724
rect 1316 1716 1347 1720
rect 1356 1716 1424 1724
rect 1036 1706 1044 1716
rect 1256 1706 1264 1716
rect 1333 1707 1347 1716
rect 927 1696 964 1704
rect 1107 1695 1133 1703
rect 1187 1695 1213 1703
rect 1416 1706 1424 1716
rect 1556 1707 1564 1736
rect 1596 1724 1604 1734
rect 1676 1736 1713 1744
rect 1596 1716 1624 1724
rect 447 1675 633 1683
rect 1616 1684 1624 1716
rect 1636 1707 1644 1733
rect 1676 1707 1684 1736
rect 1813 1744 1827 1753
rect 1813 1740 1873 1744
rect 1816 1736 1873 1740
rect 1976 1736 2033 1744
rect 1976 1706 1984 1736
rect 2096 1707 2104 1756
rect 2247 1756 2313 1764
rect 2327 1756 2453 1764
rect 2127 1736 2293 1744
rect 2427 1736 2493 1744
rect 2827 1736 2913 1744
rect 2927 1737 2973 1745
rect 3147 1737 3233 1745
rect 3296 1736 3313 1744
rect 1747 1696 1793 1704
rect 1807 1695 1853 1703
rect 2187 1695 2233 1703
rect 2327 1695 2393 1703
rect 2727 1695 2753 1703
rect 3056 1704 3064 1734
rect 3296 1707 3304 1736
rect 3367 1737 3413 1745
rect 3516 1744 3524 1776
rect 3747 1776 3833 1784
rect 4047 1776 4093 1784
rect 4347 1776 4413 1784
rect 4787 1776 4993 1784
rect 5047 1776 5353 1784
rect 5767 1776 5833 1784
rect 5927 1776 6113 1784
rect 3547 1756 3693 1764
rect 3907 1756 3933 1764
rect 5247 1756 5293 1764
rect 5707 1756 5733 1764
rect 3516 1736 3673 1744
rect 3687 1736 3713 1744
rect 3767 1736 3864 1744
rect 3056 1696 3213 1704
rect 3856 1706 3864 1736
rect 3887 1736 3913 1744
rect 4067 1736 4104 1744
rect 3387 1696 3473 1704
rect 3907 1696 3973 1704
rect 3987 1696 4013 1704
rect 4096 1687 4104 1736
rect 4136 1736 4173 1744
rect 4136 1704 4144 1736
rect 4267 1737 4333 1745
rect 4387 1736 4404 1744
rect 4167 1716 4324 1724
rect 4316 1706 4324 1716
rect 4396 1707 4404 1736
rect 4447 1736 4473 1744
rect 4540 1744 4553 1747
rect 4536 1733 4553 1744
rect 4607 1744 4620 1747
rect 4607 1733 4624 1744
rect 4136 1696 4233 1704
rect 4536 1706 4544 1733
rect 4616 1706 4624 1733
rect 1616 1676 1693 1684
rect 3287 1676 3333 1684
rect 4347 1676 4493 1684
rect 4653 1684 4667 1691
rect 4676 1687 4684 1753
rect 4827 1736 4893 1744
rect 4947 1736 5053 1744
rect 5096 1724 5104 1734
rect 5216 1724 5224 1734
rect 5607 1736 5633 1744
rect 5096 1716 5224 1724
rect 5173 1707 5187 1716
rect 5416 1707 5424 1733
rect 5556 1707 5564 1733
rect 4807 1695 4853 1703
rect 4967 1695 5013 1703
rect 5307 1695 5333 1703
rect 5676 1704 5684 1734
rect 5916 1736 5953 1744
rect 5876 1707 5884 1733
rect 5676 1696 5712 1704
rect 5747 1695 5813 1703
rect 4507 1676 4667 1684
rect 4927 1676 5133 1684
rect 5296 1684 5304 1692
rect 5207 1676 5304 1684
rect 5736 1684 5744 1692
rect 5667 1676 5744 1684
rect 547 1656 653 1664
rect 927 1656 1053 1664
rect 1307 1656 1453 1664
rect 1467 1656 1513 1664
rect 1527 1656 1573 1664
rect 2687 1656 2833 1664
rect 3427 1656 3593 1664
rect 656 1644 664 1653
rect 656 1636 713 1644
rect 767 1636 1093 1644
rect 1576 1644 1584 1653
rect 5707 1656 5853 1664
rect 5916 1664 5924 1736
rect 6087 1737 6113 1745
rect 6167 1736 6193 1744
rect 6027 1695 6173 1703
rect 5896 1656 5924 1664
rect 1576 1636 2053 1644
rect 2987 1636 3093 1644
rect 4047 1636 4353 1644
rect 4367 1636 4973 1644
rect 5896 1644 5904 1656
rect 5947 1656 6193 1664
rect 5867 1636 5904 1644
rect 907 1616 2013 1624
rect 2147 1616 2313 1624
rect 2807 1616 2953 1624
rect 2967 1616 3313 1624
rect 3967 1616 4333 1624
rect 5187 1616 5593 1624
rect 5987 1616 6233 1624
rect 527 1596 653 1604
rect 3007 1596 3753 1604
rect 3947 1596 4073 1604
rect 5387 1596 5513 1604
rect 5527 1596 5673 1604
rect 1087 1576 1853 1584
rect 1907 1576 2133 1584
rect 3747 1576 4113 1584
rect 4127 1576 4193 1584
rect 4307 1576 4893 1584
rect 5247 1576 5333 1584
rect 5347 1576 5933 1584
rect 607 1556 773 1564
rect 2827 1556 3473 1564
rect 3767 1556 4133 1564
rect 4547 1556 4933 1564
rect 5447 1556 5613 1564
rect 5747 1556 5993 1564
rect 567 1536 813 1544
rect 1007 1536 1393 1544
rect 1727 1536 1933 1544
rect 2287 1536 2533 1544
rect 2547 1536 2793 1544
rect 2807 1536 4993 1544
rect 6067 1536 6193 1544
rect 2347 1516 2373 1524
rect 2387 1516 2713 1524
rect 2847 1516 3133 1524
rect 3667 1516 3793 1524
rect 4287 1516 4313 1524
rect 5767 1516 5953 1524
rect 6107 1516 6153 1524
rect 1367 1496 1433 1504
rect 1547 1496 1613 1504
rect 2947 1496 3033 1504
rect 3227 1496 3273 1504
rect 4047 1496 4453 1504
rect 4547 1496 4573 1504
rect 5127 1496 5493 1504
rect 5507 1496 5653 1504
rect 647 1476 1013 1484
rect 1667 1476 1773 1484
rect 1827 1476 1873 1484
rect 2007 1476 2093 1484
rect 2247 1476 2813 1484
rect 2887 1476 3193 1484
rect 3207 1476 3353 1484
rect 3827 1476 3853 1484
rect 3867 1476 3953 1484
rect 4456 1484 4464 1493
rect 4456 1476 4513 1484
rect 4707 1476 5253 1484
rect 5727 1476 5913 1484
rect 147 1456 273 1464
rect 296 1456 653 1464
rect 296 1444 304 1456
rect 1927 1456 1953 1464
rect 2047 1456 2113 1464
rect 3687 1456 4033 1464
rect 116 1436 304 1444
rect 116 1424 124 1436
rect 607 1440 644 1444
rect 607 1436 647 1440
rect 633 1427 647 1436
rect 1567 1437 1613 1445
rect 107 1416 124 1424
rect 307 1416 364 1424
rect 356 1404 364 1416
rect 407 1416 513 1424
rect 987 1416 1253 1424
rect 1616 1407 1624 1434
rect 1867 1436 2313 1444
rect 2427 1436 2533 1444
rect 2707 1437 2733 1445
rect 2987 1437 3013 1445
rect 356 1396 384 1404
rect 376 1387 384 1396
rect 427 1396 493 1404
rect 587 1396 613 1404
rect 1887 1395 1933 1403
rect 2027 1396 2093 1404
rect 2187 1395 2253 1403
rect 2327 1396 2393 1404
rect 2656 1404 2664 1434
rect 3167 1437 3233 1445
rect 3327 1436 3384 1444
rect 3093 1424 3107 1433
rect 3376 1424 3384 1436
rect 3627 1437 3673 1445
rect 3727 1437 3773 1445
rect 3907 1436 3944 1444
rect 3093 1420 3364 1424
rect 3096 1416 3364 1420
rect 3376 1416 3484 1424
rect 2627 1396 2664 1404
rect 2747 1396 2773 1404
rect 2887 1395 2913 1403
rect 3027 1395 3073 1403
rect 3087 1396 3173 1404
rect 3287 1395 3333 1403
rect 3356 1404 3364 1416
rect 3356 1396 3453 1404
rect 3476 1404 3484 1416
rect 3476 1396 3593 1404
rect 376 1376 393 1387
rect 380 1373 393 1376
rect 967 1376 1133 1384
rect 1587 1376 1833 1384
rect 2447 1376 2633 1384
rect 2827 1376 2933 1384
rect 3527 1376 3733 1384
rect 3936 1384 3944 1436
rect 3956 1404 3964 1456
rect 4367 1456 4413 1464
rect 5607 1456 5644 1464
rect 4327 1436 4653 1444
rect 4667 1436 4833 1444
rect 4987 1436 5073 1444
rect 5127 1436 5173 1444
rect 5187 1437 5213 1445
rect 5636 1406 5644 1456
rect 5747 1436 5804 1444
rect 3956 1396 3993 1404
rect 4047 1395 4093 1403
rect 4307 1395 4353 1403
rect 4367 1396 4553 1404
rect 4567 1396 4733 1404
rect 4907 1395 4953 1403
rect 5676 1404 5684 1433
rect 5796 1406 5804 1436
rect 5836 1436 5873 1444
rect 5836 1407 5844 1436
rect 5896 1424 5904 1453
rect 5876 1420 5904 1424
rect 5873 1416 5904 1420
rect 5873 1407 5887 1416
rect 5676 1396 5753 1404
rect 3936 1376 3973 1384
rect 5107 1376 5193 1384
rect 5307 1376 5393 1384
rect 5407 1376 5473 1384
rect 5936 1384 5944 1453
rect 5967 1436 5993 1444
rect 6087 1437 6133 1445
rect 6036 1404 6044 1434
rect 5987 1396 6044 1404
rect 6067 1395 6193 1403
rect 5907 1376 5944 1384
rect 6087 1376 6153 1384
rect 87 1356 113 1364
rect 2047 1356 2093 1364
rect 3127 1356 3213 1364
rect 3227 1356 3373 1364
rect 3507 1356 3633 1364
rect 3647 1356 3873 1364
rect 3896 1356 4393 1364
rect 47 1336 73 1344
rect 1407 1336 1453 1344
rect 1667 1336 1893 1344
rect 2267 1336 2433 1344
rect 2527 1336 2713 1344
rect 3387 1336 3453 1344
rect 3896 1344 3904 1356
rect 5007 1356 5073 1364
rect 5127 1356 5173 1364
rect 6007 1356 6093 1364
rect 3687 1336 3904 1344
rect 3967 1336 4313 1344
rect 4427 1336 5133 1344
rect 5227 1336 5533 1344
rect 5767 1336 5933 1344
rect 347 1316 633 1324
rect 656 1316 893 1324
rect 656 1304 664 1316
rect 1227 1316 1253 1324
rect 1267 1316 1493 1324
rect 3047 1316 3093 1324
rect 3307 1316 4093 1324
rect 4107 1316 4353 1324
rect 4407 1316 5153 1324
rect 5627 1316 5713 1324
rect 5827 1316 5913 1324
rect 487 1296 664 1304
rect 867 1296 1053 1304
rect 2387 1296 2753 1304
rect 2767 1296 3253 1304
rect 3327 1296 3672 1304
rect 3707 1296 3773 1304
rect 3987 1296 4133 1304
rect 5247 1296 5733 1304
rect 5787 1296 5853 1304
rect 5867 1296 5913 1304
rect 567 1276 693 1284
rect 787 1276 1033 1284
rect 1147 1276 1313 1284
rect 2027 1276 2433 1284
rect 2487 1276 2653 1284
rect 2827 1276 2953 1284
rect 3127 1276 3193 1284
rect 3447 1276 3553 1284
rect 3567 1276 3653 1284
rect 3807 1276 3833 1284
rect 4447 1276 5633 1284
rect 5647 1276 5973 1284
rect 227 1256 253 1264
rect 327 1256 373 1264
rect 447 1256 733 1264
rect 1387 1256 1433 1264
rect 1507 1256 1613 1264
rect 1687 1256 1713 1264
rect 1767 1256 1913 1264
rect 1927 1256 1993 1264
rect 2807 1256 2993 1264
rect 3067 1256 3153 1264
rect 3167 1256 3313 1264
rect 3707 1256 3773 1264
rect 4187 1256 4233 1264
rect 4627 1256 4673 1264
rect 4787 1256 5033 1264
rect 5727 1256 5773 1264
rect 296 1236 473 1244
rect 127 1216 253 1224
rect 296 1204 304 1236
rect 807 1236 993 1244
rect 1007 1236 1132 1244
rect 3187 1236 3273 1244
rect 3816 1236 3873 1244
rect 276 1196 304 1204
rect 276 1186 284 1196
rect 107 1176 193 1184
rect 376 1184 384 1214
rect 347 1176 384 1184
rect 516 1204 524 1214
rect 747 1217 933 1225
rect 947 1216 1073 1224
rect 1327 1216 1393 1224
rect 553 1204 567 1213
rect 516 1200 567 1204
rect 516 1196 564 1200
rect 413 1184 427 1193
rect 616 1187 624 1214
rect 1547 1216 1633 1224
rect 1816 1216 1853 1224
rect 1716 1204 1724 1214
rect 1716 1196 1793 1204
rect 413 1180 444 1184
rect 416 1176 447 1180
rect 433 1167 447 1176
rect 507 1175 553 1183
rect 607 1176 624 1187
rect 607 1173 620 1176
rect 767 1176 853 1184
rect 967 1176 1053 1184
rect 1407 1175 1433 1183
rect 1716 1184 1724 1196
rect 1607 1176 1724 1184
rect 1816 1167 1824 1216
rect 1956 1204 1964 1214
rect 2147 1216 2184 1224
rect 1956 1196 2153 1204
rect 1887 1175 1913 1183
rect 2027 1175 2073 1183
rect 2176 1184 2184 1216
rect 2327 1217 2353 1225
rect 2487 1217 2553 1225
rect 2616 1204 2624 1214
rect 2736 1216 2873 1224
rect 2256 1196 2624 1204
rect 2176 1176 2213 1184
rect 2256 1167 2264 1196
rect 2507 1175 2533 1183
rect 2676 1184 2684 1213
rect 2736 1186 2744 1216
rect 3133 1224 3147 1233
rect 3816 1228 3824 1236
rect 3887 1236 3933 1244
rect 4047 1236 4073 1244
rect 4727 1236 4753 1244
rect 5207 1236 5373 1244
rect 5467 1236 5553 1244
rect 5787 1236 5833 1244
rect 6060 1244 6073 1247
rect 6056 1233 6073 1244
rect 2967 1216 3233 1224
rect 3516 1216 3593 1224
rect 3516 1207 3524 1216
rect 3896 1216 3913 1224
rect 3507 1196 3524 1207
rect 3507 1193 3520 1196
rect 3896 1204 3904 1216
rect 3967 1217 4013 1225
rect 4196 1216 4233 1224
rect 3867 1196 3904 1204
rect 4196 1187 4204 1216
rect 4256 1216 4353 1224
rect 2676 1176 2693 1184
rect 3067 1175 3093 1183
rect 3267 1175 3293 1183
rect 3487 1175 3673 1183
rect 4256 1186 4264 1216
rect 4487 1216 4673 1224
rect 4907 1216 4953 1224
rect 5027 1216 5093 1224
rect 5176 1216 5213 1224
rect 4736 1187 4744 1213
rect 5176 1207 5184 1216
rect 5267 1217 5313 1225
rect 4776 1200 4824 1204
rect 4773 1196 4824 1200
rect 4773 1187 4787 1196
rect 4816 1186 4824 1196
rect 5167 1196 5184 1207
rect 5167 1193 5180 1196
rect 5496 1204 5504 1214
rect 5647 1224 5660 1227
rect 5647 1213 5664 1224
rect 6056 1224 6064 1233
rect 5747 1216 5804 1224
rect 5347 1196 5504 1204
rect 5656 1186 5664 1213
rect 5796 1204 5804 1216
rect 5976 1216 6064 1224
rect 6076 1216 6113 1224
rect 5976 1204 5984 1216
rect 6076 1204 6084 1216
rect 5796 1196 5984 1204
rect 6056 1200 6084 1204
rect 6053 1196 6084 1200
rect 5796 1186 5804 1196
rect 6053 1187 6067 1196
rect 4987 1176 5033 1184
rect 5047 1175 5073 1183
rect 5567 1175 5593 1183
rect 6007 1175 6032 1183
rect 6136 1186 6144 1233
rect 367 1156 412 1164
rect 547 1156 653 1164
rect 667 1156 713 1164
rect 1207 1156 1293 1164
rect 1387 1156 1473 1164
rect 1807 1156 1824 1167
rect 1807 1153 1820 1156
rect 2247 1156 2264 1167
rect 2247 1153 2260 1156
rect 2367 1156 2453 1164
rect 2567 1156 2593 1164
rect 3547 1156 3573 1164
rect 3716 1164 3724 1172
rect 3587 1156 3724 1164
rect 4067 1156 4213 1164
rect 4227 1156 4333 1164
rect 4547 1156 4793 1164
rect 4887 1156 4933 1164
rect 5276 1164 5284 1172
rect 5276 1156 5353 1164
rect 5707 1156 5833 1164
rect 687 1136 773 1144
rect 2167 1136 2213 1144
rect 2227 1136 2273 1144
rect 2447 1136 2693 1144
rect 2867 1136 2913 1144
rect 3227 1136 3333 1144
rect 3847 1136 3973 1144
rect 4427 1136 4553 1144
rect 5927 1136 6093 1144
rect 147 1116 233 1124
rect 347 1116 593 1124
rect 647 1116 733 1124
rect 1107 1116 1333 1124
rect 1347 1116 1773 1124
rect 4167 1116 4673 1124
rect 4727 1116 5113 1124
rect 5267 1116 5313 1124
rect 5847 1116 5953 1124
rect 2327 1096 2733 1104
rect 3187 1096 3653 1104
rect 3667 1096 4133 1104
rect 4147 1096 5153 1104
rect 227 1076 333 1084
rect 3247 1076 3413 1084
rect 3627 1076 3873 1084
rect 3947 1076 4473 1084
rect 4627 1076 4713 1084
rect 5367 1076 5693 1084
rect 367 1056 2113 1064
rect 2127 1056 2393 1064
rect 3987 1056 4173 1064
rect 4267 1056 4413 1064
rect 5907 1056 6093 1064
rect 927 1036 1533 1044
rect 2667 1036 2753 1044
rect 3387 1036 3553 1044
rect 3787 1036 3933 1044
rect 4387 1036 4453 1044
rect 4467 1036 4653 1044
rect 4667 1036 4893 1044
rect 5767 1036 5893 1044
rect 5816 1016 6193 1024
rect 307 996 393 1004
rect 1087 996 2193 1004
rect 2687 996 2813 1004
rect 3227 996 3393 1004
rect 3407 996 3853 1004
rect 3867 996 3893 1004
rect 3907 996 4013 1004
rect 4207 996 4733 1004
rect 4747 996 4873 1004
rect 4887 996 4953 1004
rect 5816 1004 5824 1016
rect 5796 996 5824 1004
rect 5796 987 5804 996
rect 1347 976 1393 984
rect 1407 976 1733 984
rect 1907 976 2153 984
rect 2487 976 2513 984
rect 2527 976 2653 984
rect 3727 976 3833 984
rect 4607 976 4633 984
rect 4647 976 4713 984
rect 5596 976 5793 984
rect 5596 967 5604 976
rect 5847 976 5933 984
rect 5947 976 6073 984
rect 1307 956 1793 964
rect 4247 956 4444 964
rect 4436 947 4444 956
rect 5207 956 5313 964
rect 5407 956 5593 964
rect 5647 956 5713 964
rect 5727 956 5813 964
rect 887 936 1844 944
rect 1016 928 1024 936
rect 116 904 124 914
rect 226 913 227 920
rect 407 916 453 924
rect 467 917 513 925
rect 627 917 693 925
rect 787 917 833 925
rect 1227 917 1253 925
rect 1467 916 1573 924
rect 1627 916 1713 924
rect 1836 924 1844 936
rect 2107 936 2273 944
rect 2567 936 2593 944
rect 2707 936 2733 944
rect 2747 936 2793 944
rect 3247 936 3464 944
rect 3456 928 3464 936
rect 4127 936 4224 944
rect 4216 928 4224 936
rect 4447 936 4493 944
rect 5256 936 5365 944
rect 1836 916 1853 924
rect 1947 917 1973 925
rect 2027 917 2073 925
rect 2396 916 2453 924
rect 213 904 227 913
rect 76 900 124 904
rect 73 896 124 900
rect 136 900 227 904
rect 136 896 223 900
rect 73 887 87 896
rect 136 886 144 896
rect 236 887 244 914
rect 276 904 284 914
rect 276 896 304 904
rect 227 876 244 887
rect 296 884 304 896
rect 556 887 564 914
rect 976 904 984 914
rect 936 900 984 904
rect 933 896 984 900
rect 1816 904 1824 914
rect 1936 904 1944 914
rect 1816 896 1944 904
rect 933 887 947 896
rect 2396 887 2404 916
rect 2627 916 2653 924
rect 2827 917 2893 925
rect 3147 917 3393 925
rect 3467 916 3573 924
rect 3587 917 3693 925
rect 3827 916 3933 924
rect 3947 916 4013 924
rect 4227 916 4333 924
rect 4496 916 4633 924
rect 2416 896 2864 904
rect 296 876 493 884
rect 227 873 240 876
rect 556 876 573 887
rect 560 873 573 876
rect 727 876 753 884
rect 1407 875 1433 883
rect 1447 876 1533 884
rect 1607 875 1773 883
rect 1847 876 1993 884
rect 2047 876 2093 884
rect 2416 886 2424 896
rect 2547 876 2833 884
rect 2856 884 2864 896
rect 2927 896 3073 904
rect 4056 904 4064 914
rect 4056 896 4113 904
rect 4496 904 4504 916
rect 4767 916 4933 924
rect 4987 916 5013 924
rect 5256 924 5264 936
rect 5357 928 5365 936
rect 5627 936 5673 944
rect 5167 916 5264 924
rect 4196 896 4264 904
rect 4196 886 4204 896
rect 4256 886 4264 896
rect 4476 896 4504 904
rect 4476 886 4484 896
rect 2856 876 3113 884
rect 3367 876 3433 884
rect 3447 875 3533 883
rect 3547 876 3673 884
rect 3807 875 3853 883
rect 4267 875 4353 883
rect 4567 876 4613 884
rect 5007 875 5033 883
rect 5156 884 5164 914
rect 5367 916 5433 924
rect 5487 916 5533 924
rect 5573 924 5587 933
rect 5573 920 5604 924
rect 5576 916 5604 920
rect 5276 887 5284 913
rect 5596 904 5604 916
rect 5727 917 5753 925
rect 5907 916 5973 924
rect 5596 896 5644 904
rect 5087 876 5164 884
rect 5347 876 5453 884
rect 107 856 153 864
rect 207 856 253 864
rect 387 856 433 864
rect 547 856 613 864
rect 867 856 993 864
rect 1007 856 1073 864
rect 1687 856 1733 864
rect 2767 856 2993 864
rect 3856 864 3864 872
rect 5636 867 5644 896
rect 5707 876 5733 884
rect 6036 867 6044 914
rect 6096 887 6104 913
rect 3167 856 3304 864
rect 3856 856 4033 864
rect 467 836 813 844
rect 1067 836 1173 844
rect 1347 836 1553 844
rect 2127 836 2173 844
rect 2187 836 2233 844
rect 2647 836 2673 844
rect 2687 836 2893 844
rect 3047 836 3273 844
rect 3296 844 3304 856
rect 4747 856 4893 864
rect 4907 856 4973 864
rect 5116 856 5193 864
rect 3296 836 3473 844
rect 5116 844 5124 856
rect 5767 856 5833 864
rect 5887 856 5993 864
rect 4427 836 5124 844
rect 5627 836 5773 844
rect 427 816 733 824
rect 947 816 993 824
rect 1367 816 1673 824
rect 1887 816 2073 824
rect 2087 816 2413 824
rect 2667 816 2913 824
rect 3447 816 3933 824
rect 4327 816 5173 824
rect 5187 816 5333 824
rect 5927 816 6053 824
rect 87 796 353 804
rect 367 796 1153 804
rect 2147 796 2193 804
rect 2607 796 3013 804
rect 3067 796 3233 804
rect 3247 796 3973 804
rect 4087 796 4173 804
rect 4767 796 5004 804
rect 807 776 953 784
rect 1207 776 1453 784
rect 1467 776 2293 784
rect 2807 776 2913 784
rect 3627 776 4193 784
rect 4996 784 5004 796
rect 5207 796 5324 804
rect 4996 776 5173 784
rect 5187 776 5253 784
rect 5316 784 5324 796
rect 5316 776 5373 784
rect 5447 776 5553 784
rect 5567 776 5713 784
rect 5867 776 5953 784
rect 6007 776 6053 784
rect 1587 756 1673 764
rect 2367 756 2653 764
rect 2947 756 3253 764
rect 3727 756 3773 764
rect 4087 756 4113 764
rect 4127 756 4153 764
rect 4287 756 4353 764
rect 4527 756 4973 764
rect 5287 756 5893 764
rect 227 736 253 744
rect 267 736 533 744
rect 547 736 573 744
rect 587 736 953 744
rect 1007 736 1233 744
rect 1307 736 1393 744
rect 1547 736 1633 744
rect 2687 736 2853 744
rect 3927 736 4153 744
rect 4167 736 4373 744
rect 4687 736 4933 744
rect 5787 736 5873 744
rect 5947 736 5973 744
rect 1667 716 1733 724
rect 1907 716 1953 724
rect 2607 716 2704 724
rect 27 697 73 705
rect 307 697 353 705
rect 427 696 444 704
rect 167 655 193 663
rect 436 644 444 696
rect 467 697 493 705
rect 707 696 773 704
rect 787 696 813 704
rect 887 696 913 704
rect 1047 697 1093 705
rect 1136 684 1144 694
rect 1187 696 1353 704
rect 1527 696 1593 704
rect 1700 704 1713 707
rect 1696 693 1713 704
rect 1847 696 2033 704
rect 2087 697 2113 705
rect 2267 697 2293 705
rect 1136 676 1324 684
rect 527 656 633 664
rect 1167 655 1193 663
rect 1267 656 1293 664
rect 1316 664 1324 676
rect 1696 666 1704 693
rect 2487 696 2533 704
rect 2560 704 2573 707
rect 2556 693 2573 704
rect 2627 697 2673 705
rect 2696 704 2704 716
rect 3007 716 3153 724
rect 3167 716 3213 724
rect 3267 724 3280 727
rect 3267 713 3284 724
rect 3647 716 3733 724
rect 3747 716 4213 724
rect 2696 696 2813 704
rect 2827 696 2953 704
rect 3087 696 3113 704
rect 3247 704 3260 707
rect 3247 693 3264 704
rect 1316 656 1413 664
rect 1467 655 1493 663
rect 2067 655 2133 663
rect 2327 656 2373 664
rect 2556 666 2564 693
rect 2747 676 2884 684
rect 2876 666 2884 676
rect 3256 666 3264 693
rect 3276 684 3284 713
rect 3367 697 3393 705
rect 3276 676 3324 684
rect 2427 656 2513 664
rect 3027 655 3053 663
rect 3187 656 3253 664
rect 3316 664 3324 676
rect 3456 667 3464 693
rect 3647 696 3693 704
rect 3767 697 3793 705
rect 3807 697 3833 705
rect 3316 656 3413 664
rect 3587 655 3613 663
rect 436 636 593 644
rect 607 636 793 644
rect 807 636 933 644
rect 947 636 1033 644
rect 1667 636 1773 644
rect 1887 636 1973 644
rect 1987 636 2173 644
rect 2767 636 2973 644
rect 2987 636 3133 644
rect 3687 636 3773 644
rect 407 616 453 624
rect 747 616 1113 624
rect 2147 616 2213 624
rect 2487 616 2793 624
rect 3487 616 3533 624
rect 3547 616 3613 624
rect 3876 624 3884 694
rect 3896 666 3904 716
rect 4327 716 4353 724
rect 5087 716 5113 724
rect 5407 716 5464 724
rect 3927 696 3984 704
rect 3976 666 3984 696
rect 4007 696 4053 704
rect 4387 704 4400 707
rect 4387 693 4404 704
rect 4507 696 4553 704
rect 4607 697 4653 705
rect 4396 666 4404 693
rect 4716 684 4724 694
rect 5027 696 5133 704
rect 5147 696 5273 704
rect 4636 676 4724 684
rect 4027 655 4073 663
rect 4227 655 4293 663
rect 4527 655 4573 663
rect 4636 664 4644 676
rect 4796 667 4804 693
rect 4627 656 4644 664
rect 4876 644 4884 694
rect 5336 667 5344 693
rect 4907 656 4993 664
rect 5047 656 5073 664
rect 5087 655 5113 663
rect 5127 656 5293 664
rect 5456 666 5464 716
rect 5507 716 5533 724
rect 5607 696 5793 704
rect 5920 704 5932 707
rect 5916 693 5932 704
rect 5967 697 6013 705
rect 6033 704 6047 713
rect 6033 696 6084 704
rect 5513 684 5527 693
rect 5513 680 5544 684
rect 5516 676 5544 680
rect 5536 666 5544 676
rect 5916 666 5924 693
rect 6076 666 6084 696
rect 5587 656 5693 664
rect 5807 655 5873 663
rect 4787 636 5153 644
rect 5167 636 5253 644
rect 5267 636 5973 644
rect 6076 644 6084 652
rect 6027 636 6084 644
rect 3876 616 4013 624
rect 4207 616 4493 624
rect 4547 616 4733 624
rect 5647 616 5833 624
rect 5887 616 5953 624
rect 987 596 1013 604
rect 1027 596 1073 604
rect 1827 596 2353 604
rect 3227 596 3293 604
rect 4447 596 4833 604
rect 4847 596 5393 604
rect 5407 596 5413 604
rect 5427 596 5593 604
rect 687 576 1593 584
rect 2327 576 2593 584
rect 3527 576 3853 584
rect 3867 576 4133 584
rect 4507 576 4613 584
rect 5547 576 5733 584
rect 5807 576 6033 584
rect 2227 556 2773 564
rect 2787 556 3073 564
rect 4667 556 4693 564
rect 3947 536 4533 544
rect 5667 536 5713 544
rect 1427 516 1533 524
rect 1547 516 1833 524
rect 2527 516 2673 524
rect 2687 516 2933 524
rect 2947 516 3633 524
rect 4607 516 5313 524
rect 27 496 253 504
rect 267 496 993 504
rect 1007 496 1313 504
rect 3927 496 4053 504
rect 4287 496 4373 504
rect 4387 496 5693 504
rect 5827 496 5853 504
rect 2287 476 2373 484
rect 2387 476 2653 484
rect 4947 476 5013 484
rect 5027 476 5053 484
rect 5187 476 5573 484
rect 5667 476 5833 484
rect 687 456 853 464
rect 1367 456 1504 464
rect 1496 447 1504 456
rect 1927 456 2053 464
rect 2067 456 2253 464
rect 2267 456 2593 464
rect 2867 456 3133 464
rect 3347 456 3553 464
rect 3567 456 3693 464
rect 3707 456 3813 464
rect 4027 456 4053 464
rect 4067 456 4233 464
rect 4276 456 4633 464
rect 67 436 113 444
rect 587 436 873 444
rect 1507 436 1733 444
rect 2647 436 2753 444
rect 2847 436 2893 444
rect 4276 444 4284 456
rect 5907 456 5993 464
rect 6067 456 6113 464
rect 4207 436 4284 444
rect 4796 436 4913 444
rect 107 416 193 424
rect 327 416 433 424
rect 1427 416 1573 424
rect 2327 416 2844 424
rect 227 396 453 404
rect 467 396 513 404
rect 647 396 733 404
rect 747 396 773 404
rect 1187 396 1233 404
rect 27 355 113 363
rect 167 356 193 364
rect 407 355 453 363
rect 507 355 573 363
rect 596 364 604 393
rect 916 384 924 394
rect 876 376 924 384
rect 956 384 964 394
rect 1056 384 1064 394
rect 956 376 1064 384
rect 596 356 613 364
rect 876 364 884 376
rect 1056 367 1064 376
rect 807 356 884 364
rect 1047 356 1064 367
rect 1096 367 1104 394
rect 1576 396 1613 404
rect 1576 387 1584 396
rect 1727 397 1773 405
rect 1827 396 1853 404
rect 1967 397 2013 405
rect 2107 397 2153 405
rect 2627 397 2713 405
rect 2727 396 2784 404
rect 1567 376 1584 387
rect 2236 376 2324 384
rect 1567 373 1580 376
rect 1096 356 1113 367
rect 1047 353 1060 356
rect 1100 353 1113 356
rect 1207 356 1293 364
rect 1347 356 1413 364
rect 1427 355 1473 363
rect 1527 356 1593 364
rect 1707 356 1893 364
rect 1947 356 1992 364
rect 2027 356 2113 364
rect 2236 366 2244 376
rect 2316 366 2324 376
rect 2327 355 2393 363
rect 2556 364 2564 394
rect 2776 367 2784 396
rect 2556 356 2693 364
rect 907 336 1013 344
rect 1647 336 1713 344
rect 2087 340 2144 344
rect 2087 336 2147 340
rect 2133 327 2147 336
rect 2796 344 2804 394
rect 2836 364 2844 416
rect 3207 416 3253 424
rect 3347 416 3393 424
rect 3987 416 4133 424
rect 4147 416 4593 424
rect 4796 424 4804 436
rect 5807 436 6033 444
rect 4727 416 4804 424
rect 5287 416 5333 424
rect 5347 416 5513 424
rect 6107 416 6173 424
rect 2927 397 2973 405
rect 3147 397 3173 405
rect 3307 397 3453 405
rect 3667 396 3853 404
rect 4036 396 4093 404
rect 3796 376 3924 384
rect 2836 356 2873 364
rect 3127 356 3193 364
rect 3796 364 3804 376
rect 3916 367 3924 376
rect 3687 356 3804 364
rect 3856 356 3913 364
rect 3856 347 3864 356
rect 4036 364 4044 396
rect 4367 397 4413 405
rect 4427 396 4553 404
rect 4787 396 4813 404
rect 4887 396 4973 404
rect 5687 397 5753 405
rect 5807 396 5833 404
rect 5976 384 5984 394
rect 5936 376 5984 384
rect 4007 356 4044 364
rect 4067 355 4113 363
rect 4807 355 4853 363
rect 4927 355 4953 363
rect 5067 355 5093 363
rect 5267 356 5313 364
rect 5707 356 5733 364
rect 2727 336 2804 344
rect 2907 336 2993 344
rect 3007 336 3073 344
rect 3847 336 3864 347
rect 3847 333 3860 336
rect 3996 344 4004 352
rect 3887 336 4004 344
rect 367 316 733 324
rect 1047 316 1213 324
rect 1227 316 1793 324
rect 2367 316 2533 324
rect 2547 316 2612 324
rect 2647 316 2673 324
rect 2787 316 2813 324
rect 3187 316 3493 324
rect 3727 316 3813 324
rect 3867 316 3972 324
rect 3996 324 4004 336
rect 4147 336 4433 344
rect 4447 336 4533 344
rect 4796 344 4804 352
rect 5936 347 5944 376
rect 6036 364 6044 393
rect 5967 356 6044 364
rect 6136 364 6144 393
rect 6127 356 6144 364
rect 4707 336 4804 344
rect 5347 336 5373 344
rect 5387 336 5453 344
rect 5507 336 5613 344
rect 5827 336 5873 344
rect 3996 316 4253 324
rect 4607 316 4653 324
rect 4727 316 5053 324
rect 5727 316 5973 324
rect 6087 316 6233 324
rect 1247 296 1393 304
rect 1447 296 1693 304
rect 2607 296 3073 304
rect 3627 296 3653 304
rect 3967 296 4073 304
rect 4327 296 4573 304
rect 4647 296 5693 304
rect 5747 296 5833 304
rect 947 276 1113 284
rect 1127 276 1764 284
rect 1756 267 1764 276
rect 2267 276 3113 284
rect 3367 276 3513 284
rect 3787 276 4193 284
rect 4307 276 4613 284
rect 5187 276 5213 284
rect 5227 276 5293 284
rect 867 256 1073 264
rect 1327 256 1513 264
rect 1767 256 1913 264
rect 1927 256 2073 264
rect 2616 256 2653 264
rect 2616 244 2624 256
rect 2667 256 3273 264
rect 4296 264 4304 273
rect 3967 256 4304 264
rect 4767 256 4853 264
rect 4867 256 5133 264
rect 5427 256 5613 264
rect 5727 256 5793 264
rect 2347 236 2624 244
rect 2687 236 3033 244
rect 3047 236 3333 244
rect 3807 236 3913 244
rect 4027 236 4313 244
rect 4407 236 4473 244
rect 4687 236 4713 244
rect 5616 244 5624 253
rect 5616 236 5673 244
rect 5687 236 5773 244
rect 5847 236 5893 244
rect 5907 236 6153 244
rect 247 216 493 224
rect 667 216 713 224
rect 727 216 764 224
rect 756 204 764 216
rect 807 216 1033 224
rect 1047 216 1093 224
rect 1107 216 1293 224
rect 1307 216 1413 224
rect 1527 216 1553 224
rect 1907 216 2173 224
rect 2227 216 2324 224
rect 756 196 833 204
rect 1887 196 2213 204
rect 47 177 93 185
rect 267 177 293 185
rect 387 177 433 185
rect 507 176 733 184
rect 1187 177 1253 185
rect 736 164 744 174
rect 876 164 884 174
rect 736 156 884 164
rect 427 136 473 144
rect 547 136 713 144
rect 727 135 793 143
rect 1107 135 1153 143
rect 1436 146 1444 193
rect 1467 176 1493 184
rect 1576 146 1584 193
rect 2316 204 2324 216
rect 2447 216 2573 224
rect 2687 216 2733 224
rect 3127 216 3233 224
rect 3247 216 3313 224
rect 3407 216 3753 224
rect 3767 216 4113 224
rect 4447 216 4493 224
rect 4547 216 4573 224
rect 5007 216 5353 224
rect 5367 216 5433 224
rect 5447 216 5573 224
rect 2316 196 2393 204
rect 2416 196 2473 204
rect 1607 176 1713 184
rect 1767 176 1884 184
rect 1876 167 1884 176
rect 1927 184 1940 187
rect 1927 173 1944 184
rect 1967 176 2173 184
rect 1876 156 1893 167
rect 1880 153 1893 156
rect 1936 146 1944 173
rect 2416 146 2424 196
rect 2607 196 2753 204
rect 3467 196 4153 204
rect 2507 176 2553 184
rect 3007 176 3104 184
rect 3096 164 3104 176
rect 3187 176 3233 184
rect 3307 176 3353 184
rect 3567 176 3693 184
rect 3707 177 3793 185
rect 3096 156 3124 164
rect 1267 136 1293 144
rect 1307 136 1393 144
rect 1527 135 1573 143
rect 1707 136 1833 144
rect 1987 136 2053 144
rect 2107 135 2133 143
rect 2187 135 2233 143
rect 2347 135 2373 143
rect 2487 135 2533 143
rect 2627 136 2873 144
rect 2947 135 3033 143
rect 3116 144 3124 156
rect 3816 146 3824 196
rect 4167 196 4393 204
rect 4807 196 4973 204
rect 5087 196 5153 204
rect 5487 196 5653 204
rect 5667 196 5713 204
rect 5787 196 5833 204
rect 5927 196 6193 204
rect 3847 176 3864 184
rect 3116 136 3133 144
rect 3147 136 3213 144
rect 3587 136 3713 144
rect 3727 135 3753 143
rect 3856 127 3864 176
rect 3876 164 3884 174
rect 3967 176 4004 184
rect 3876 156 3933 164
rect 3996 146 4004 176
rect 4516 176 4713 184
rect 4056 147 4064 173
rect 4256 164 4264 174
rect 4516 164 4524 176
rect 5187 176 5233 184
rect 4753 164 4767 173
rect 4176 156 4524 164
rect 4176 146 4184 156
rect 4516 146 4524 156
rect 4736 160 4767 164
rect 4736 156 4764 160
rect 4736 146 4744 156
rect 4287 136 4373 144
rect 4427 135 4473 143
rect 4567 135 4613 143
rect 4807 135 4833 143
rect 5087 135 5113 143
rect 5225 144 5233 176
rect 5736 164 5744 174
rect 5793 164 5807 173
rect 5527 156 5744 164
rect 5756 160 5807 164
rect 5756 156 5804 160
rect 5636 146 5644 156
rect 5756 146 5764 156
rect 5225 136 5273 144
rect 5687 135 5713 143
rect 5847 135 5873 143
rect 5927 135 5993 143
rect 2587 116 2704 124
rect 2696 107 2704 116
rect 3847 116 3864 127
rect 3847 113 3860 116
rect 5276 124 5284 132
rect 3947 116 4044 124
rect 5276 116 5393 124
rect 4036 107 4044 116
rect 5407 116 5553 124
rect 587 96 753 104
rect 867 96 993 104
rect 1207 96 1613 104
rect 1627 96 2493 104
rect 2707 96 2833 104
rect 3107 96 3344 104
rect 1507 76 1593 84
rect 2167 76 2613 84
rect 2887 76 3293 84
rect 3336 84 3344 96
rect 3967 96 3993 104
rect 4047 96 4273 104
rect 4787 96 4873 104
rect 4887 96 4953 104
rect 5607 96 5813 104
rect 6027 96 6213 104
rect 3336 76 3833 84
rect 4147 76 4473 84
rect 3867 56 4073 64
rect 4707 56 4913 64
rect 5987 56 6073 64
rect 767 36 1053 44
rect 3187 36 3373 44
use INVX1  _889_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 1170 0 1 3390
box -12 -8 52 272
use NOR2X1  _890_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 690 0 -1 3390
box -12 -8 74 272
use NAND2X1  _891_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform -1 0 770 0 -1 2870
box -12 -8 72 272
use INVX1  _892_
timestamp 1701862152
transform 1 0 850 0 -1 2870
box -12 -8 52 272
use INVX1  _893_
timestamp 1701862152
transform 1 0 1370 0 1 3390
box -12 -8 52 272
use INVX2  _894_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 1110 0 -1 2870
box -12 -8 52 272
use NOR2X1  _895_
timestamp 1701862152
transform 1 0 1610 0 1 3390
box -12 -8 74 272
use NAND2X1  _896_
timestamp 1702508443
transform -1 0 1810 0 1 3390
box -12 -8 72 272
use INVX1  _897_
timestamp 1701862152
transform -1 0 1010 0 1 3910
box -12 -8 52 272
use NOR2X1  _898_
timestamp 1701862152
transform -1 0 1550 0 1 3390
box -12 -8 74 272
use AOI21X1  _899_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform -1 0 1070 0 1 3390
box -12 -8 92 272
use NOR2X1  _900_
timestamp 1701862152
transform -1 0 470 0 1 3910
box -12 -8 74 272
use OAI21X1  _901_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform -1 0 610 0 1 3910
box -12 -8 92 272
use INVX1  _902_
timestamp 1701862152
transform 1 0 230 0 -1 4430
box -12 -8 52 272
use INVX4  _903_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 650 0 -1 2870
box -12 -8 72 272
use OAI21X1  _904_
timestamp 1702508443
transform -1 0 770 0 1 3390
box -12 -8 92 272
use INVX1  _905_
timestamp 1701862152
transform -1 0 670 0 -1 3910
box -12 -8 52 272
use NOR2X1  _906_
timestamp 1701862152
transform -1 0 1030 0 -1 2870
box -12 -8 74 272
use INVX1  _907_
timestamp 1701862152
transform -1 0 970 0 -1 4430
box -12 -8 52 272
use INVX1  _908_
timestamp 1701862152
transform -1 0 510 0 -1 4430
box -12 -8 52 272
use OAI21X1  _909_
timestamp 1702508443
transform -1 0 930 0 1 3390
box -12 -8 92 272
use OAI21X1  _910_
timestamp 1702508443
transform 1 0 730 0 -1 3910
box -12 -8 92 272
use AOI22X1  _911_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 470 0 -1 3910
box -14 -8 114 272
use NAND2X1  _912_
timestamp 1702508443
transform -1 0 390 0 -1 3910
box -12 -8 72 272
use OAI21X1  _913_
timestamp 1702508443
transform 1 0 250 0 1 4430
box -12 -8 92 272
use OAI21X1  _914_
timestamp 1702508443
transform 1 0 330 0 -1 4430
box -12 -8 92 272
use NAND2X1  _915_
timestamp 1702508443
transform 1 0 1450 0 -1 3390
box -12 -8 72 272
use NOR2X1  _916_
timestamp 1701862152
transform -1 0 630 0 -1 4430
box -12 -8 74 272
use NOR2X1  _917_
timestamp 1701862152
transform 1 0 690 0 1 3910
box -12 -8 74 272
use OAI22X1  _918_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 1170 0 1 3910
box -12 -8 112 272
use OR2X2  _919_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform 1 0 830 0 1 3910
box -12 -8 92 272
use INVX1  _920_
timestamp 1701862152
transform -1 0 1450 0 1 3910
box -12 -8 52 272
use AOI22X1  _921_
timestamp 1701862152
transform -1 0 1350 0 1 3910
box -14 -8 114 272
use NAND3X1  _922_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform 1 0 870 0 -1 3910
box -12 -8 92 272
use AND2X2  _923_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 1250 0 -1 3910
box -12 -8 94 272
use OAI21X1  _924_
timestamp 1702508443
transform 1 0 1010 0 -1 3910
box -12 -8 92 272
use INVX8  _925_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 90 0 1 3910
box -12 -8 114 272
use INVX1  _926_
timestamp 1701862152
transform 1 0 3210 0 1 4430
box -12 -8 52 272
use NAND2X1  _927_
timestamp 1702508443
transform -1 0 3170 0 -1 4430
box -12 -8 72 272
use OAI21X1  _928_
timestamp 1702508443
transform 1 0 3230 0 -1 4430
box -12 -8 92 272
use INVX1  _929_
timestamp 1701862152
transform -1 0 3790 0 -1 4950
box -12 -8 52 272
use NAND2X1  _930_
timestamp 1702508443
transform -1 0 3990 0 -1 3910
box -12 -8 72 272
use OAI21X1  _931_
timestamp 1702508443
transform 1 0 3770 0 -1 3910
box -12 -8 92 272
use INVX1  _932_
timestamp 1701862152
transform 1 0 2210 0 1 3910
box -12 -8 52 272
use NAND2X1  _933_
timestamp 1702508443
transform 1 0 2050 0 -1 3910
box -12 -8 72 272
use OAI21X1  _934_
timestamp 1702508443
transform -1 0 2270 0 -1 3910
box -12 -8 92 272
use INVX1  _935_
timestamp 1701862152
transform 1 0 4410 0 -1 5470
box -12 -8 52 272
use NAND2X1  _936_
timestamp 1702508443
transform -1 0 3690 0 -1 3390
box -12 -8 72 272
use OAI21X1  _937_
timestamp 1702508443
transform -1 0 3550 0 -1 3390
box -12 -8 92 272
use INVX1  _938_
timestamp 1701862152
transform 1 0 2990 0 -1 4430
box -12 -8 52 272
use NAND2X1  _939_
timestamp 1702508443
transform 1 0 2730 0 -1 3390
box -12 -8 72 272
use OAI21X1  _940_
timestamp 1702508443
transform -1 0 2950 0 -1 3390
box -12 -8 92 272
use INVX1  _941_
timestamp 1701862152
transform 1 0 2470 0 -1 4430
box -12 -8 52 272
use NAND2X1  _942_
timestamp 1702508443
transform -1 0 2690 0 -1 3910
box -12 -8 72 272
use OAI21X1  _943_
timestamp 1702508443
transform 1 0 2750 0 -1 3910
box -12 -8 92 272
use INVX1  _944_
timestamp 1701862152
transform 1 0 1470 0 -1 4430
box -12 -8 52 272
use NAND2X1  _945_
timestamp 1702508443
transform -1 0 1690 0 1 3910
box -12 -8 72 272
use OAI21X1  _946_
timestamp 1702508443
transform -1 0 1850 0 1 3910
box -12 -8 92 272
use INVX4  _947_
timestamp 1701862152
transform -1 0 1390 0 -1 4430
box -12 -8 72 272
use NAND2X1  _948_
timestamp 1702508443
transform -1 0 1810 0 -1 2870
box -12 -8 72 272
use OAI21X1  _949_
timestamp 1702508443
transform -1 0 1950 0 -1 2870
box -12 -8 92 272
use INVX1  _950_
timestamp 1701862152
transform -1 0 130 0 1 2870
box -12 -8 52 272
use INVX1  _951_
timestamp 1701862152
transform 1 0 4330 0 1 3910
box -12 -8 52 272
use INVX2  _952_
timestamp 1701862152
transform 1 0 2710 0 -1 2870
box -12 -8 52 272
use NOR2X1  _953_
timestamp 1701862152
transform 1 0 4250 0 -1 4430
box -12 -8 74 272
use AND2X2  _954_
timestamp 1701862152
transform 1 0 4130 0 1 3390
box -12 -8 94 272
use NAND2X1  _955_
timestamp 1702508443
transform 1 0 4390 0 -1 4430
box -12 -8 72 272
use NAND2X1  _956_
timestamp 1702508443
transform 1 0 5030 0 -1 5470
box -12 -8 72 272
use NAND2X1  _957_
timestamp 1702508443
transform 1 0 4690 0 -1 5990
box -12 -8 72 272
use OR2X2  _958_
timestamp 1702508443
transform 1 0 4930 0 1 5990
box -12 -8 92 272
use NAND2X1  _959_
timestamp 1702508443
transform -1 0 5290 0 -1 5990
box -12 -8 72 272
use AND2X2  _960_
timestamp 1701862152
transform -1 0 4870 0 1 5990
box -12 -8 94 272
use OAI21X1  _961_
timestamp 1702508443
transform -1 0 5170 0 1 5990
box -12 -8 92 272
use NAND2X1  _962_
timestamp 1702508443
transform -1 0 5370 0 1 5470
box -12 -8 72 272
use INVX1  _963_
timestamp 1701862152
transform 1 0 6090 0 1 5990
box -12 -8 52 272
use NAND2X1  _964_
timestamp 1702508443
transform 1 0 5730 0 1 4430
box -12 -8 72 272
use NAND2X1  _965_
timestamp 1702508443
transform 1 0 5270 0 -1 4430
box -12 -8 72 272
use OR2X2  _966_
timestamp 1702508443
transform -1 0 6110 0 1 5470
box -12 -8 92 272
use INVX1  _967_
timestamp 1701862152
transform 1 0 4910 0 1 5470
box -12 -8 52 272
use INVX1  _968_
timestamp 1701862152
transform 1 0 3330 0 -1 2870
box -12 -8 52 272
use OAI21X1  _969_
timestamp 1702508443
transform 1 0 5450 0 1 5470
box -12 -8 92 272
use NAND3X1  _970_
timestamp 1702508443
transform -1 0 6030 0 -1 5990
box -12 -8 92 272
use NOR2X1  _971_
timestamp 1701862152
transform -1 0 6130 0 -1 5470
box -12 -8 74 272
use AND2X2  _972_
timestamp 1701862152
transform -1 0 6090 0 -1 270
box -12 -8 94 272
use OAI21X1  _973_
timestamp 1702508443
transform -1 0 5870 0 1 5990
box -12 -8 92 272
use NAND3X1  _974_
timestamp 1702508443
transform 1 0 5490 0 1 5990
box -12 -8 92 272
use INVX1  _975_
timestamp 1701862152
transform 1 0 4770 0 -1 4950
box -12 -8 52 272
use NAND2X1  _976_
timestamp 1702508443
transform -1 0 4510 0 1 3910
box -12 -8 72 272
use INVX2  _977_
timestamp 1701862152
transform 1 0 3090 0 -1 2870
box -12 -8 52 272
use NAND2X1  _978_
timestamp 1702508443
transform -1 0 4510 0 -1 3390
box -12 -8 72 272
use OAI21X1  _979_
timestamp 1702508443
transform 1 0 4570 0 -1 3390
box -12 -8 92 272
use OAI21X1  _980_
timestamp 1702508443
transform 1 0 4830 0 1 4950
box -12 -8 92 272
use AOI21X1  _981_
timestamp 1702508443
transform 1 0 5630 0 1 5990
box -12 -8 92 272
use OAI21X1  _982_
timestamp 1702508443
transform 1 0 5750 0 1 5470
box -12 -8 92 272
use OAI21X1  _983_
timestamp 1702508443
transform 1 0 5890 0 1 5470
box -12 -8 92 272
use AND2X2  _984_
timestamp 1701862152
transform 1 0 4970 0 1 2870
box -12 -8 94 272
use NAND3X1  _985_
timestamp 1702508443
transform 1 0 4950 0 -1 3390
box -12 -8 92 272
use AOI22X1  _986_
timestamp 1701862152
transform 1 0 5390 0 1 3910
box -14 -8 114 272
use INVX1  _987_
timestamp 1701862152
transform -1 0 5970 0 -1 4430
box -12 -8 52 272
use NAND2X1  _988_
timestamp 1702508443
transform -1 0 5370 0 1 4430
box -12 -8 72 272
use INVX1  _989_
timestamp 1701862152
transform 1 0 5550 0 -1 4430
box -12 -8 52 272
use NAND3X1  _990_
timestamp 1702508443
transform 1 0 6030 0 -1 4950
box -12 -8 92 272
use NAND2X1  _991_
timestamp 1702508443
transform -1 0 5150 0 -1 3390
box -12 -8 72 272
use NOR2X1  _992_
timestamp 1701862152
transform -1 0 5190 0 -1 4430
box -12 -8 74 272
use OAI21X1  _993_
timestamp 1702508443
transform 1 0 5650 0 -1 4430
box -12 -8 92 272
use NAND3X1  _994_
timestamp 1702508443
transform -1 0 6150 0 1 4950
box -12 -8 92 272
use AOI21X1  _995_
timestamp 1702508443
transform 1 0 6090 0 -1 5990
box -12 -8 92 272
use OAI21X1  _996_
timestamp 1702508443
transform 1 0 5410 0 -1 4430
box -12 -8 92 272
use NAND3X1  _997_
timestamp 1702508443
transform -1 0 5930 0 1 4430
box -12 -8 92 272
use NAND3X1  _998_
timestamp 1702508443
transform 1 0 5590 0 1 4430
box -12 -8 92 272
use NAND2X1  _999_
timestamp 1702508443
transform 1 0 4070 0 -1 3910
box -12 -8 72 272
use INVX1  _1000_
timestamp 1701862152
transform -1 0 4230 0 -1 3910
box -12 -8 52 272
use AND2X2  _1001_
timestamp 1701862152
transform 1 0 3870 0 -1 3390
box -12 -8 94 272
use NAND2X1  _1002_
timestamp 1702508443
transform -1 0 4330 0 1 3390
box -12 -8 72 272
use INVX1  _1003_
timestamp 1701862152
transform 1 0 4710 0 -1 2350
box -12 -8 52 272
use OAI21X1  _1004_
timestamp 1702508443
transform 1 0 4410 0 1 3390
box -12 -8 92 272
use NAND3X1  _1005_
timestamp 1702508443
transform -1 0 4630 0 1 3390
box -12 -8 92 272
use OAI21X1  _1006_
timestamp 1702508443
transform -1 0 4530 0 -1 3910
box -12 -8 92 272
use INVX1  _1007_
timestamp 1701862152
transform 1 0 3750 0 -1 3390
box -12 -8 52 272
use OAI21X1  _1008_
timestamp 1702508443
transform 1 0 4030 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1009_
timestamp 1702508443
transform 1 0 4290 0 -1 3910
box -12 -8 92 272
use AND2X2  _1010_
timestamp 1701862152
transform -1 0 5950 0 1 3910
box -12 -8 94 272
use NAND3X1  _1011_
timestamp 1702508443
transform -1 0 5810 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1012_
timestamp 1702508443
transform 1 0 5450 0 1 4430
box -12 -8 92 272
use AOI21X1  _1013_
timestamp 1702508443
transform -1 0 5990 0 1 4950
box -12 -8 92 272
use NAND2X1  _1014_
timestamp 1702508443
transform 1 0 6170 0 1 3910
box -12 -8 72 272
use OAI21X1  _1015_
timestamp 1702508443
transform -1 0 5950 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1016_
timestamp 1702508443
transform 1 0 5590 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1017_
timestamp 1702508443
transform -1 0 5510 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1018_
timestamp 1702508443
transform 1 0 4970 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1019_
timestamp 1702508443
transform 1 0 5990 0 1 4430
box -12 -8 92 272
use OAI21X1  _1020_
timestamp 1702508443
transform 1 0 6050 0 -1 4430
box -12 -8 92 272
use AND2X2  _1021_
timestamp 1701862152
transform 1 0 3690 0 -1 2870
box -12 -8 94 272
use NAND2X1  _1022_
timestamp 1702508443
transform -1 0 4910 0 -1 2870
box -12 -8 72 272
use INVX1  _1023_
timestamp 1701862152
transform -1 0 4750 0 -1 3390
box -12 -8 52 272
use INVX2  _1024_
timestamp 1701862152
transform -1 0 2190 0 -1 2870
box -12 -8 52 272
use NAND2X1  _1025_
timestamp 1702508443
transform -1 0 4630 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1026_
timestamp 1702508443
transform 1 0 4690 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1027_
timestamp 1702508443
transform 1 0 5430 0 1 2870
box -12 -8 72 272
use INVX1  _1028_
timestamp 1701862152
transform 1 0 5410 0 -1 2870
box -12 -8 52 272
use NAND3X1  _1029_
timestamp 1702508443
transform 1 0 5110 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1030_
timestamp 1701862152
transform -1 0 5030 0 -1 2870
box -12 -8 74 272
use AOI22X1  _1031_
timestamp 1701862152
transform -1 0 4510 0 -1 2870
box -14 -8 114 272
use OAI21X1  _1032_
timestamp 1702508443
transform 1 0 5670 0 -1 2870
box -12 -8 92 272
use AOI21X1  _1033_
timestamp 1702508443
transform 1 0 5850 0 1 2870
box -12 -8 92 272
use AOI21X1  _1034_
timestamp 1702508443
transform -1 0 5870 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1035_
timestamp 1702508443
transform -1 0 5610 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1036_
timestamp 1702508443
transform 1 0 5810 0 -1 2870
box -12 -8 92 272
use AOI21X1  _1037_
timestamp 1702508443
transform 1 0 6130 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1038_
timestamp 1702508443
transform -1 0 3850 0 1 2870
box -12 -8 72 272
use INVX1  _1039_
timestamp 1701862152
transform -1 0 3970 0 1 2870
box -12 -8 52 272
use AND2X2  _1040_
timestamp 1701862152
transform 1 0 3970 0 -1 2870
box -12 -8 94 272
use AND2X2  _1041_
timestamp 1701862152
transform 1 0 4530 0 1 2870
box -12 -8 94 272
use NAND2X1  _1042_
timestamp 1702508443
transform 1 0 4270 0 -1 2870
box -12 -8 72 272
use INVX2  _1043_
timestamp 1701862152
transform 1 0 4310 0 -1 5990
box -12 -8 52 272
use NAND2X1  _1044_
timestamp 1702508443
transform 1 0 4310 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1045_
timestamp 1702508443
transform 1 0 4370 0 1 2870
box -12 -8 92 272
use NAND3X1  _1046_
timestamp 1702508443
transform 1 0 4210 0 1 2870
box -12 -8 92 272
use OAI21X1  _1047_
timestamp 1702508443
transform 1 0 4130 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1048_
timestamp 1702508443
transform 1 0 4670 0 1 2870
box -12 -8 92 272
use NAND3X1  _1049_
timestamp 1702508443
transform 1 0 4810 0 1 2870
box -12 -8 92 272
use AND2X2  _1050_
timestamp 1701862152
transform 1 0 5270 0 1 2870
box -12 -8 94 272
use OAI21X1  _1051_
timestamp 1702508443
transform 1 0 6130 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1052_
timestamp 1702508443
transform -1 0 6050 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1053_
timestamp 1702508443
transform 1 0 5690 0 1 2870
box -12 -8 92 272
use NAND2X1  _1054_
timestamp 1702508443
transform -1 0 5190 0 1 2870
box -12 -8 72 272
use NAND3X1  _1055_
timestamp 1702508443
transform 1 0 5690 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1056_
timestamp 1702508443
transform -1 0 6230 0 1 4430
box -12 -8 92 272
use OAI21X1  _1057_
timestamp 1702508443
transform 1 0 6010 0 1 3910
box -12 -8 92 272
use NAND3X1  _1058_
timestamp 1702508443
transform 1 0 5850 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1059_
timestamp 1702508443
transform -1 0 6070 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1060_
timestamp 1702508443
transform -1 0 6210 0 1 3390
box -12 -8 92 272
use INVX4  _1061_
timestamp 1701862152
transform 1 0 1370 0 -1 2870
box -12 -8 72 272
use NOR2X1  _1062_
timestamp 1701862152
transform 1 0 4190 0 -1 3390
box -12 -8 74 272
use OAI21X1  _1063_
timestamp 1702508443
transform 1 0 4810 0 -1 3390
box -12 -8 92 272
use XNOR2X1  _1064_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform 1 0 5350 0 -1 3390
box -12 -8 132 272
use INVX1  _1065_
timestamp 1701862152
transform 1 0 5890 0 -1 3910
box -12 -8 52 272
use NAND3X1  _1066_
timestamp 1702508443
transform -1 0 5770 0 1 3390
box -12 -8 92 272
use AOI21X1  _1067_
timestamp 1702508443
transform -1 0 6050 0 1 3390
box -12 -8 92 272
use AOI21X1  _1068_
timestamp 1702508443
transform -1 0 6090 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1069_
timestamp 1702508443
transform -1 0 5610 0 1 3390
box -12 -8 92 272
use NAND3X1  _1070_
timestamp 1702508443
transform -1 0 5390 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1071_
timestamp 1702508443
transform 1 0 5210 0 -1 3390
box -12 -8 72 272
use INVX1  _1072_
timestamp 1701862152
transform 1 0 5470 0 1 1310
box -12 -8 52 272
use OAI21X1  _1073_
timestamp 1702508443
transform 1 0 5550 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1074_
timestamp 1702508443
transform 1 0 6150 0 1 2870
box -12 -8 92 272
use OAI21X1  _1075_
timestamp 1702508443
transform 1 0 5710 0 1 2350
box -12 -8 92 272
use NAND3X1  _1076_
timestamp 1702508443
transform 1 0 4710 0 1 2350
box -12 -8 92 272
use AOI22X1  _1077_
timestamp 1701862152
transform -1 0 4650 0 1 2350
box -14 -8 114 272
use INVX1  _1078_
timestamp 1701862152
transform -1 0 5130 0 -1 2350
box -12 -8 52 272
use NAND2X1  _1079_
timestamp 1702508443
transform -1 0 4110 0 -1 2350
box -12 -8 72 272
use INVX1  _1080_
timestamp 1701862152
transform -1 0 5030 0 1 2350
box -12 -8 52 272
use NAND3X1  _1081_
timestamp 1702508443
transform 1 0 5210 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1082_
timestamp 1702508443
transform -1 0 4470 0 1 2350
box -12 -8 72 272
use NOR2X1  _1083_
timestamp 1701862152
transform -1 0 4930 0 1 2350
box -12 -8 74 272
use OAI21X1  _1084_
timestamp 1702508443
transform -1 0 5330 0 1 2350
box -12 -8 92 272
use AOI21X1  _1085_
timestamp 1702508443
transform 1 0 6030 0 1 2350
box -12 -8 92 272
use OAI21X1  _1086_
timestamp 1702508443
transform 1 0 5390 0 1 2350
box -12 -8 92 272
use NAND3X1  _1087_
timestamp 1702508443
transform 1 0 5110 0 1 2350
box -12 -8 92 272
use AOI22X1  _1088_
timestamp 1701862152
transform -1 0 5630 0 1 2350
box -14 -8 114 272
use NAND2X1  _1089_
timestamp 1702508443
transform -1 0 4150 0 1 1830
box -12 -8 72 272
use INVX1  _1090_
timestamp 1701862152
transform 1 0 4370 0 1 1830
box -12 -8 52 272
use AND2X2  _1091_
timestamp 1701862152
transform 1 0 3650 0 1 2870
box -12 -8 94 272
use AND2X2  _1092_
timestamp 1701862152
transform 1 0 3850 0 1 2350
box -12 -8 94 272
use NAND2X1  _1093_
timestamp 1702508443
transform -1 0 4350 0 1 2350
box -12 -8 72 272
use AOI22X1  _1094_
timestamp 1701862152
transform 1 0 3870 0 -1 2350
box -14 -8 114 272
use INVX1  _1095_
timestamp 1701862152
transform 1 0 4310 0 -1 2350
box -12 -8 52 272
use NAND3X1  _1096_
timestamp 1702508443
transform 1 0 4430 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1097_
timestamp 1702508443
transform 1 0 4150 0 1 2350
box -12 -8 92 272
use OAI21X1  _1098_
timestamp 1702508443
transform 1 0 4010 0 1 2350
box -12 -8 92 272
use NAND3X1  _1099_
timestamp 1702508443
transform 1 0 4170 0 -1 2350
box -12 -8 92 272
use AND2X2  _1100_
timestamp 1701862152
transform 1 0 5490 0 -1 2350
box -12 -8 94 272
use OAI21X1  _1101_
timestamp 1702508443
transform -1 0 6030 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1102_
timestamp 1702508443
transform 1 0 5270 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1103_
timestamp 1702508443
transform 1 0 5550 0 1 2870
box -12 -8 92 272
use NAND3X1  _1104_
timestamp 1702508443
transform -1 0 5950 0 1 2350
box -12 -8 92 272
use NAND2X1  _1105_
timestamp 1702508443
transform 1 0 5350 0 -1 2350
box -12 -8 72 272
use NAND3X1  _1106_
timestamp 1702508443
transform 1 0 5810 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1107_
timestamp 1702508443
transform 1 0 6010 0 1 1830
box -12 -8 92 272
use OAI21X1  _1108_
timestamp 1702508443
transform 1 0 6010 0 1 2870
box -12 -8 92 272
use NAND3X1  _1109_
timestamp 1702508443
transform 1 0 5730 0 1 1830
box -12 -8 92 272
use OAI21X1  _1110_
timestamp 1702508443
transform -1 0 6190 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1111_
timestamp 1702508443
transform 1 0 6050 0 1 270
box -12 -8 92 272
use NAND2X1  _1112_
timestamp 1702508443
transform -1 0 3790 0 1 2350
box -12 -8 72 272
use INVX1  _1113_
timestamp 1701862152
transform 1 0 4610 0 1 1830
box -12 -8 52 272
use AOI22X1  _1114_
timestamp 1701862152
transform 1 0 4050 0 1 2870
box -14 -8 114 272
use INVX1  _1115_
timestamp 1701862152
transform -1 0 4010 0 -1 1830
box -12 -8 52 272
use OAI21X1  _1116_
timestamp 1702508443
transform 1 0 3830 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1117_
timestamp 1701862152
transform 1 0 3710 0 -1 1830
box -12 -8 74 272
use NAND2X1  _1118_
timestamp 1702508443
transform 1 0 4190 0 -1 1830
box -12 -8 72 272
use NAND3X1  _1119_
timestamp 1702508443
transform -1 0 4550 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1120_
timestamp 1702508443
transform -1 0 4130 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1121_
timestamp 1702508443
transform -1 0 4310 0 1 1830
box -12 -8 92 272
use NAND3X1  _1122_
timestamp 1702508443
transform 1 0 4310 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1123_
timestamp 1702508443
transform 1 0 4410 0 1 1310
box -12 -8 72 272
use NAND3X1  _1124_
timestamp 1702508443
transform 1 0 6030 0 1 1310
box -12 -8 92 272
use AOI21X1  _1125_
timestamp 1702508443
transform -1 0 6030 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1126_
timestamp 1702508443
transform -1 0 5950 0 1 1830
box -12 -8 92 272
use NAND3X1  _1127_
timestamp 1702508443
transform 1 0 4930 0 1 1310
box -12 -8 92 272
use NAND3X1  _1128_
timestamp 1702508443
transform 1 0 4610 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1129_
timestamp 1702508443
transform 1 0 5210 0 1 1310
box -12 -8 72 272
use OAI21X1  _1130_
timestamp 1702508443
transform -1 0 5870 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1131_
timestamp 1702508443
transform -1 0 5830 0 1 1310
box -12 -8 92 272
use AOI21X1  _1132_
timestamp 1702508443
transform -1 0 5910 0 1 3390
box -12 -8 92 272
use OAI21X1  _1133_
timestamp 1702508443
transform -1 0 5730 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1134_
timestamp 1702508443
transform 1 0 6090 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1135_
timestamp 1702508443
transform -1 0 5870 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1136_
timestamp 1702508443
transform -1 0 5550 0 -1 1830
box -12 -8 92 272
use NAND3X1  _1137_
timestamp 1702508443
transform -1 0 5710 0 -1 1830
box -12 -8 92 272
use NAND3X1  _1138_
timestamp 1702508443
transform -1 0 5970 0 1 1310
box -12 -8 92 272
use NAND3X1  _1139_
timestamp 1702508443
transform 1 0 5190 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1140_
timestamp 1702508443
transform -1 0 5370 0 1 1830
box -12 -8 92 272
use INVX1  _1141_
timestamp 1701862152
transform -1 0 5210 0 1 1830
box -12 -8 52 272
use INVX1  _1142_
timestamp 1701862152
transform 1 0 5030 0 1 4430
box -12 -8 52 272
use NOR2X1  _1143_
timestamp 1701862152
transform -1 0 5010 0 -1 5990
box -12 -8 74 272
use INVX1  _1144_
timestamp 1701862152
transform -1 0 5430 0 1 5990
box -12 -8 52 272
use OAI21X1  _1145_
timestamp 1702508443
transform 1 0 4810 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1146_
timestamp 1702508443
transform 1 0 5370 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1147_
timestamp 1702508443
transform 1 0 5930 0 1 5990
box -12 -8 92 272
use NAND3X1  _1148_
timestamp 1702508443
transform -1 0 5890 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1149_
timestamp 1702508443
transform -1 0 5590 0 -1 5990
box -12 -8 92 272
use AND2X2  _1150_
timestamp 1701862152
transform 1 0 4990 0 1 4950
box -12 -8 94 272
use NAND3X1  _1151_
timestamp 1702508443
transform 1 0 5650 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1152_
timestamp 1702508443
transform 1 0 5910 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1153_
timestamp 1702508443
transform -1 0 5690 0 1 4950
box -12 -8 92 272
use NAND3X1  _1154_
timestamp 1702508443
transform -1 0 5850 0 1 4950
box -12 -8 92 272
use NAND3X1  _1155_
timestamp 1702508443
transform -1 0 5550 0 1 4950
box -12 -8 92 272
use NAND3X1  _1156_
timestamp 1702508443
transform 1 0 5150 0 1 4430
box -12 -8 92 272
use OAI21X1  _1157_
timestamp 1702508443
transform 1 0 5590 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1158_
timestamp 1702508443
transform -1 0 5830 0 -1 3910
box -12 -8 92 272
use AOI22X1  _1159_
timestamp 1701862152
transform -1 0 5790 0 1 3910
box -14 -8 114 272
use NAND3X1  _1160_
timestamp 1702508443
transform -1 0 5130 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1161_
timestamp 1702508443
transform -1 0 5410 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1162_
timestamp 1702508443
transform -1 0 4970 0 -1 1830
box -12 -8 92 272
use NAND3X1  _1163_
timestamp 1702508443
transform -1 0 5830 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1164_
timestamp 1702508443
transform -1 0 5310 0 1 5990
box -12 -8 92 272
use NAND2X1  _1165_
timestamp 1702508443
transform -1 0 4170 0 -1 4430
box -12 -8 72 272
use OR2X2  _1166_
timestamp 1702508443
transform 1 0 4210 0 1 4950
box -12 -8 92 272
use NAND2X1  _1167_
timestamp 1702508443
transform -1 0 4430 0 1 4950
box -12 -8 72 272
use AOI22X1  _1168_
timestamp 1701862152
transform 1 0 4770 0 -1 5470
box -14 -8 114 272
use OAI21X1  _1169_
timestamp 1702508443
transform 1 0 4510 0 1 4950
box -12 -8 92 272
use OAI21X1  _1170_
timestamp 1702508443
transform 1 0 5070 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1171_
timestamp 1702508443
transform 1 0 5170 0 1 5470
box -12 -8 92 272
use AOI21X1  _1172_
timestamp 1702508443
transform -1 0 5090 0 1 5470
box -12 -8 92 272
use OAI21X1  _1173_
timestamp 1702508443
transform 1 0 5330 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1174_
timestamp 1702508443
transform 1 0 5590 0 1 5470
box -12 -8 92 272
use NAND3X1  _1175_
timestamp 1702508443
transform 1 0 5590 0 -1 5470
box -12 -8 92 272
use INVX1  _1176_
timestamp 1701862152
transform -1 0 4910 0 -1 4950
box -12 -8 52 272
use AOI22X1  _1177_
timestamp 1701862152
transform 1 0 5310 0 1 4950
box -14 -8 114 272
use OAI21X1  _1178_
timestamp 1702508443
transform -1 0 4950 0 1 4430
box -12 -8 92 272
use NAND3X1  _1179_
timestamp 1702508443
transform -1 0 4890 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1180_
timestamp 1702508443
transform -1 0 5470 0 1 3390
box -12 -8 92 272
use NOR3X1  _1181_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 5190 0 1 3390
box -12 -8 172 272
use INVX1  _1182_
timestamp 1701862152
transform -1 0 4970 0 -1 5470
box -12 -8 52 272
use NAND3X1  _1183_
timestamp 1702508443
transform -1 0 4750 0 1 4950
box -12 -8 92 272
use INVX1  _1184_
timestamp 1701862152
transform -1 0 4310 0 -1 4950
box -12 -8 52 272
use OAI21X1  _1185_
timestamp 1702508443
transform 1 0 4130 0 -1 4950
box -12 -8 92 272
use OR2X2  _1186_
timestamp 1702508443
transform -1 0 3950 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1187_
timestamp 1702508443
transform 1 0 3090 0 1 4430
box -12 -8 72 272
use NOR2X1  _1188_
timestamp 1701862152
transform -1 0 3390 0 1 4430
box -12 -8 74 272
use INVX1  _1189_
timestamp 1701862152
transform 1 0 3830 0 -1 4430
box -12 -8 52 272
use OAI21X1  _1190_
timestamp 1702508443
transform -1 0 4030 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1191_
timestamp 1702508443
transform 1 0 3870 0 1 4430
box -12 -8 92 272
use INVX1  _1192_
timestamp 1701862152
transform 1 0 4030 0 1 4430
box -12 -8 52 272
use INVX1  _1193_
timestamp 1701862152
transform 1 0 5470 0 -1 5470
box -12 -8 52 272
use OAI21X1  _1194_
timestamp 1702508443
transform -1 0 5250 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1195_
timestamp 1702508443
transform 1 0 4490 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1196_
timestamp 1702508443
transform -1 0 5230 0 1 4950
box -12 -8 92 272
use NOR3X1  _1197_
timestamp 1701862152
transform -1 0 4810 0 1 4430
box -12 -8 172 272
use OAI21X1  _1198_
timestamp 1702508443
transform -1 0 5370 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1199_
timestamp 1702508443
transform 1 0 5130 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1200_
timestamp 1702508443
transform -1 0 5070 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1201_
timestamp 1702508443
transform 1 0 4650 0 -1 4430
box -12 -8 92 272
use INVX1  _1202_
timestamp 1701862152
transform 1 0 4730 0 -1 3910
box -12 -8 52 272
use OAI21X1  _1203_
timestamp 1702508443
transform -1 0 5330 0 1 3390
box -12 -8 92 272
use AOI21X1  _1204_
timestamp 1702508443
transform -1 0 4950 0 1 3390
box -12 -8 92 272
use OAI21X1  _1205_
timestamp 1702508443
transform -1 0 4830 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1206_
timestamp 1702508443
transform -1 0 5670 0 1 1310
box -12 -8 92 272
use NAND2X1  _1207_
timestamp 1702508443
transform 1 0 5070 0 1 1310
box -12 -8 72 272
use OAI21X1  _1208_
timestamp 1702508443
transform 1 0 6070 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1209_
timestamp 1702508443
transform 1 0 4130 0 1 1310
box -12 -8 72 272
use INVX1  _1210_
timestamp 1701862152
transform 1 0 5090 0 1 270
box -12 -8 52 272
use NOR2X1  _1211_
timestamp 1701862152
transform -1 0 4570 0 -1 1310
box -12 -8 74 272
use OAI21X1  _1212_
timestamp 1702508443
transform -1 0 4550 0 1 1830
box -12 -8 92 272
use NAND2X1  _1213_
timestamp 1702508443
transform 1 0 4830 0 -1 270
box -12 -8 72 272
use OR2X2  _1214_
timestamp 1702508443
transform 1 0 4950 0 -1 270
box -12 -8 92 272
use NAND3X1  _1215_
timestamp 1702508443
transform 1 0 5110 0 -1 270
box -12 -8 92 272
use AND2X2  _1216_
timestamp 1701862152
transform 1 0 4810 0 1 270
box -12 -8 94 272
use NOR2X1  _1217_
timestamp 1701862152
transform 1 0 4690 0 1 270
box -12 -8 74 272
use OAI21X1  _1218_
timestamp 1702508443
transform 1 0 4950 0 1 270
box -12 -8 92 272
use NAND2X1  _1219_
timestamp 1702508443
transform -1 0 5330 0 -1 270
box -12 -8 72 272
use AOI21X1  _1220_
timestamp 1702508443
transform -1 0 5670 0 1 1830
box -12 -8 92 272
use NAND2X1  _1221_
timestamp 1702508443
transform -1 0 3590 0 1 1830
box -12 -8 72 272
use AND2X2  _1222_
timestamp 1701862152
transform 1 0 3190 0 -1 2870
box -12 -8 94 272
use OAI21X1  _1223_
timestamp 1702508443
transform 1 0 3150 0 1 2350
box -12 -8 92 272
use AND2X2  _1224_
timestamp 1701862152
transform -1 0 3490 0 1 2350
box -12 -8 94 272
use OAI21X1  _1225_
timestamp 1702508443
transform -1 0 3650 0 1 2350
box -12 -8 92 272
use NAND3X1  _1226_
timestamp 1702508443
transform -1 0 3630 0 -1 2350
box -12 -8 92 272
use INVX1  _1227_
timestamp 1701862152
transform -1 0 3510 0 -1 1830
box -12 -8 52 272
use NAND2X1  _1228_
timestamp 1702508443
transform 1 0 3290 0 1 2350
box -12 -8 72 272
use AOI22X1  _1229_
timestamp 1701862152
transform -1 0 3790 0 -1 2350
box -14 -8 114 272
use INVX1  _1230_
timestamp 1701862152
transform -1 0 3630 0 -1 1830
box -12 -8 52 272
use NAND3X1  _1231_
timestamp 1702508443
transform -1 0 3390 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1232_
timestamp 1702508443
transform -1 0 4270 0 -1 1310
box -12 -8 72 272
use AOI21X1  _1233_
timestamp 1702508443
transform -1 0 5030 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1234_
timestamp 1702508443
transform -1 0 4650 0 -1 2350
box -12 -8 72 272
use XOR2X1  _1235_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform -1 0 4850 0 1 1310
box -12 -8 132 272
use NAND2X1  _1236_
timestamp 1702508443
transform 1 0 5070 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1237_
timestamp 1702508443
transform 1 0 4810 0 -1 2350
box -12 -8 92 272
use XNOR2X1  _1238_
timestamp 1702508443
transform -1 0 4670 0 1 1310
box -12 -8 132 272
use NAND2X1  _1239_
timestamp 1702508443
transform -1 0 4770 0 1 790
box -12 -8 72 272
use NAND3X1  _1240_
timestamp 1702508443
transform 1 0 5010 0 1 790
box -12 -8 92 272
use AND2X2  _1241_
timestamp 1701862152
transform 1 0 4050 0 -1 1310
box -12 -8 94 272
use NAND2X1  _1242_
timestamp 1702508443
transform 1 0 4930 0 -1 1310
box -12 -8 72 272
use NAND2X1  _1243_
timestamp 1702508443
transform -1 0 4650 0 1 790
box -12 -8 72 272
use NAND3X1  _1244_
timestamp 1702508443
transform -1 0 4390 0 1 790
box -12 -8 92 272
use NAND3X1  _1245_
timestamp 1702508443
transform 1 0 5430 0 1 790
box -12 -8 92 272
use OAI21X1  _1246_
timestamp 1702508443
transform 1 0 5650 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1247_
timestamp 1701862152
transform 1 0 4330 0 -1 1310
box -14 -8 114 272
use AOI21X1  _1248_
timestamp 1702508443
transform -1 0 4930 0 1 790
box -12 -8 92 272
use OAI21X1  _1249_
timestamp 1702508443
transform 1 0 5390 0 -1 790
box -12 -8 92 272
use NAND3X1  _1250_
timestamp 1702508443
transform 1 0 5690 0 -1 790
box -12 -8 92 272
use AND2X2  _1251_
timestamp 1701862152
transform 1 0 5390 0 -1 270
box -12 -8 94 272
use NAND3X1  _1252_
timestamp 1702508443
transform -1 0 5370 0 1 790
box -12 -8 92 272
use OAI21X1  _1253_
timestamp 1702508443
transform 1 0 5370 0 1 270
box -12 -8 92 272
use NAND3X1  _1254_
timestamp 1702508443
transform 1 0 5710 0 -1 270
box -12 -8 92 272
use NAND3X1  _1255_
timestamp 1702508443
transform 1 0 5870 0 -1 270
box -12 -8 92 272
use AOI21X1  _1256_
timestamp 1702508443
transform -1 0 6010 0 -1 1310
box -12 -8 92 272
use AOI22X1  _1257_
timestamp 1701862152
transform 1 0 5550 0 -1 270
box -14 -8 114 272
use AOI21X1  _1258_
timestamp 1702508443
transform 1 0 5530 0 -1 790
box -12 -8 92 272
use OAI21X1  _1259_
timestamp 1702508443
transform 1 0 5850 0 -1 790
box -12 -8 92 272
use AOI21X1  _1260_
timestamp 1702508443
transform 1 0 5250 0 -1 790
box -12 -8 92 272
use INVX1  _1261_
timestamp 1701862152
transform 1 0 5370 0 -1 1310
box -12 -8 52 272
use NAND3X1  _1262_
timestamp 1702508443
transform -1 0 5950 0 1 790
box -12 -8 92 272
use OAI21X1  _1263_
timestamp 1702508443
transform 1 0 6010 0 -1 790
box -12 -8 92 272
use AOI21X1  _1264_
timestamp 1702508443
transform -1 0 5650 0 1 790
box -12 -8 92 272
use OAI21X1  _1265_
timestamp 1702508443
transform 1 0 5490 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1266_
timestamp 1702508443
transform -1 0 5410 0 1 1310
box -12 -8 92 272
use NAND3X1  _1267_
timestamp 1702508443
transform -1 0 5810 0 1 790
box -12 -8 92 272
use NAND3X1  _1268_
timestamp 1702508443
transform 1 0 5110 0 -1 790
box -12 -8 92 272
use NAND3X1  _1269_
timestamp 1702508443
transform -1 0 5290 0 -1 1310
box -12 -8 92 272
use AND2X2  _1270_
timestamp 1701862152
transform -1 0 3490 0 -1 1310
box -12 -8 94 272
use XOR2X1  _1271_
timestamp 1702508443
transform 1 0 2550 0 -1 1830
box -12 -8 132 272
use NOR2X1  _1272_
timestamp 1701862152
transform 1 0 1130 0 -1 4950
box -12 -8 74 272
use NOR2X1  _1273_
timestamp 1701862152
transform 1 0 1590 0 -1 4430
box -12 -8 74 272
use OAI21X1  _1274_
timestamp 1702508443
transform -1 0 2530 0 1 3910
box -12 -8 92 272
use AOI21X1  _1275_
timestamp 1702508443
transform -1 0 2670 0 1 3910
box -12 -8 92 272
use OAI21X1  _1276_
timestamp 1702508443
transform -1 0 2270 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1277_
timestamp 1702508443
transform 1 0 2310 0 1 3910
box -12 -8 92 272
use NAND2X1  _1278_
timestamp 1702508443
transform 1 0 810 0 1 2870
box -12 -8 72 272
use OAI21X1  _1279_
timestamp 1702508443
transform 1 0 650 0 1 2870
box -12 -8 92 272
use INVX1  _1280_
timestamp 1701862152
transform 1 0 1130 0 1 2350
box -12 -8 52 272
use INVX1  _1281_
timestamp 1701862152
transform -1 0 1690 0 1 2350
box -12 -8 52 272
use OAI21X1  _1282_
timestamp 1702508443
transform 1 0 1230 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1283_
timestamp 1702508443
transform 1 0 1750 0 1 2350
box -12 -8 92 272
use NAND3X1  _1284_
timestamp 1702508443
transform 1 0 5450 0 1 1830
box -12 -8 92 272
use INVX1  _1285_
timestamp 1701862152
transform -1 0 5310 0 1 3910
box -12 -8 52 272
use NAND2X1  _1286_
timestamp 1702508443
transform -1 0 5530 0 -1 3910
box -12 -8 72 272
use NAND3X1  _1287_
timestamp 1702508443
transform -1 0 5630 0 1 3910
box -12 -8 92 272
use NAND3X1  _1288_
timestamp 1702508443
transform -1 0 5230 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1289_
timestamp 1702508443
transform 1 0 4990 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1290_
timestamp 1702508443
transform 1 0 4850 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1291_
timestamp 1702508443
transform 1 0 5030 0 1 1830
box -12 -8 92 272
use NAND2X1  _1292_
timestamp 1702508443
transform -1 0 3910 0 1 1310
box -12 -8 72 272
use OAI21X1  _1293_
timestamp 1702508443
transform -1 0 3650 0 1 1310
box -12 -8 92 272
use INVX1  _1294_
timestamp 1701862152
transform 1 0 4870 0 -1 790
box -12 -8 52 272
use AOI21X1  _1295_
timestamp 1702508443
transform -1 0 5050 0 -1 790
box -12 -8 92 272
use OAI21X1  _1296_
timestamp 1702508443
transform 1 0 4670 0 -1 270
box -12 -8 92 272
use INVX1  _1297_
timestamp 1701862152
transform 1 0 4250 0 -1 270
box -12 -8 52 272
use AOI21X1  _1298_
timestamp 1702508443
transform 1 0 5150 0 1 790
box -12 -8 92 272
use OAI21X1  _1299_
timestamp 1702508443
transform 1 0 5210 0 1 270
box -12 -8 92 272
use NAND2X1  _1300_
timestamp 1702508443
transform 1 0 3710 0 1 1310
box -12 -8 72 272
use NOR2X1  _1301_
timestamp 1701862152
transform -1 0 4050 0 1 1310
box -12 -8 74 272
use NAND2X1  _1302_
timestamp 1702508443
transform -1 0 3870 0 1 1830
box -12 -8 72 272
use NAND2X1  _1303_
timestamp 1702508443
transform -1 0 4010 0 1 1830
box -12 -8 72 272
use OAI22X1  _1304_
timestamp 1701862152
transform -1 0 3750 0 1 1830
box -12 -8 112 272
use XNOR2X1  _1305_
timestamp 1702508443
transform 1 0 3710 0 -1 1310
box -12 -8 132 272
use XNOR2X1  _1306_
timestamp 1702508443
transform 1 0 3570 0 1 790
box -12 -8 132 272
use NOR2X1  _1307_
timestamp 1701862152
transform 1 0 4470 0 1 790
box -12 -8 74 272
use AOI21X1  _1308_
timestamp 1702508443
transform -1 0 4230 0 1 790
box -12 -8 92 272
use NAND2X1  _1309_
timestamp 1702508443
transform -1 0 3490 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1310_
timestamp 1702508443
transform 1 0 2650 0 1 1830
box -12 -8 72 272
use INVX1  _1311_
timestamp 1701862152
transform 1 0 2930 0 1 1830
box -12 -8 52 272
use AND2X2  _1312_
timestamp 1701862152
transform 1 0 2410 0 1 2350
box -12 -8 94 272
use AND2X2  _1313_
timestamp 1701862152
transform 1 0 2730 0 1 2350
box -12 -8 94 272
use NAND2X1  _1314_
timestamp 1702508443
transform 1 0 2870 0 1 2350
box -12 -8 72 272
use AOI22X1  _1315_
timestamp 1701862152
transform -1 0 2530 0 -1 2350
box -14 -8 114 272
use INVX1  _1316_
timestamp 1701862152
transform 1 0 2590 0 -1 2350
box -12 -8 52 272
use AOI21X1  _1317_
timestamp 1702508443
transform 1 0 3190 0 1 1830
box -12 -8 92 272
use INVX2  _1318_
timestamp 1701862152
transform 1 0 2310 0 1 2350
box -12 -8 52 272
use OAI21X1  _1319_
timestamp 1702508443
transform 1 0 2570 0 1 2350
box -12 -8 92 272
use OAI21X1  _1320_
timestamp 1702508443
transform -1 0 3070 0 1 2350
box -12 -8 92 272
use AOI21X1  _1321_
timestamp 1702508443
transform 1 0 2830 0 -1 2350
box -12 -8 92 272
use OAI22X1  _1322_
timestamp 1701862152
transform 1 0 3350 0 1 1830
box -12 -8 112 272
use NAND3X1  _1323_
timestamp 1702508443
transform 1 0 2690 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1324_
timestamp 1702508443
transform -1 0 3230 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1325_
timestamp 1701862152
transform -1 0 3350 0 -1 2350
box -12 -8 74 272
use NAND3X1  _1326_
timestamp 1702508443
transform -1 0 3070 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1327_
timestamp 1702508443
transform 1 0 3890 0 1 790
box -12 -8 72 272
use NOR2X1  _1328_
timestamp 1701862152
transform -1 0 4170 0 -1 790
box -12 -8 74 272
use NOR2X1  _1329_
timestamp 1701862152
transform -1 0 4850 0 -1 1310
box -12 -8 74 272
use OAI21X1  _1330_
timestamp 1702508443
transform -1 0 4730 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1331_
timestamp 1702508443
transform -1 0 3830 0 1 790
box -12 -8 92 272
use OAI21X1  _1332_
timestamp 1702508443
transform 1 0 3830 0 -1 790
box -12 -8 92 272
use XOR2X1  _1333_
timestamp 1702508443
transform 1 0 3250 0 1 790
box -12 -8 132 272
use NAND3X1  _1334_
timestamp 1702508443
transform -1 0 3990 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1335_
timestamp 1702508443
transform 1 0 3970 0 -1 790
box -12 -8 72 272
use NAND3X1  _1336_
timestamp 1702508443
transform 1 0 3810 0 1 270
box -12 -8 92 272
use NAND3X1  _1337_
timestamp 1702508443
transform 1 0 4090 0 1 270
box -12 -8 92 272
use NOR3X1  _1338_
timestamp 1701862152
transform 1 0 5530 0 1 270
box -12 -8 172 272
use AOI21X1  _1339_
timestamp 1702508443
transform 1 0 5750 0 1 270
box -12 -8 92 272
use AOI21X1  _1340_
timestamp 1702508443
transform 1 0 3650 0 1 270
box -12 -8 92 272
use NAND3X1  _1341_
timestamp 1702508443
transform 1 0 4010 0 1 790
box -12 -8 92 272
use OAI21X1  _1342_
timestamp 1702508443
transform -1 0 4470 0 -1 790
box -12 -8 92 272
use AOI21X1  _1343_
timestamp 1702508443
transform 1 0 4250 0 -1 790
box -12 -8 92 272
use OAI21X1  _1344_
timestamp 1702508443
transform -1 0 4450 0 1 270
box -12 -8 92 272
use NAND3X1  _1345_
timestamp 1702508443
transform 1 0 4370 0 -1 270
box -12 -8 92 272
use NAND3X1  _1346_
timestamp 1702508443
transform 1 0 4230 0 1 270
box -12 -8 92 272
use OAI21X1  _1347_
timestamp 1702508443
transform 1 0 4530 0 1 270
box -12 -8 92 272
use NAND3X1  _1348_
timestamp 1702508443
transform 1 0 4510 0 -1 270
box -12 -8 92 272
use NAND3X1  _1349_
timestamp 1702508443
transform -1 0 4630 0 -1 790
box -12 -8 92 272
use AOI21X1  _1350_
timestamp 1702508443
transform -1 0 6090 0 1 790
box -12 -8 92 272
use OAI21X1  _1351_
timestamp 1702508443
transform 1 0 5910 0 1 270
box -12 -8 92 272
use NAND3X1  _1352_
timestamp 1702508443
transform -1 0 4190 0 -1 270
box -12 -8 92 272
use NAND3X1  _1353_
timestamp 1702508443
transform -1 0 4050 0 -1 270
box -12 -8 92 272
use NAND3X1  _1354_
timestamp 1702508443
transform -1 0 3730 0 -1 270
box -12 -8 92 272
use NAND2X1  _1355_
timestamp 1702508443
transform 1 0 3530 0 -1 790
box -12 -8 72 272
use AND2X2  _1356_
timestamp 1701862152
transform -1 0 2970 0 -1 1830
box -12 -8 94 272
use OAI21X1  _1357_
timestamp 1702508443
transform -1 0 2830 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1358_
timestamp 1702508443
transform -1 0 2250 0 1 2350
box -12 -8 92 272
use AND2X2  _1359_
timestamp 1701862152
transform -1 0 3030 0 1 4430
box -12 -8 94 272
use NAND2X1  _1360_
timestamp 1702508443
transform 1 0 1930 0 1 4430
box -12 -8 72 272
use OAI21X1  _1361_
timestamp 1702508443
transform -1 0 2870 0 1 4430
box -12 -8 92 272
use OAI21X1  _1362_
timestamp 1702508443
transform -1 0 2130 0 1 4430
box -12 -8 92 272
use AOI21X1  _1363_
timestamp 1702508443
transform -1 0 1370 0 -1 3390
box -12 -8 92 272
use AOI22X1  _1364_
timestamp 1701862152
transform 1 0 1230 0 1 2350
box -14 -8 114 272
use OAI21X1  _1365_
timestamp 1702508443
transform -1 0 610 0 1 3390
box -12 -8 92 272
use AOI21X1  _1366_
timestamp 1702508443
transform -1 0 3590 0 -1 270
box -12 -8 92 272
use AOI22X1  _1367_
timestamp 1701862152
transform -1 0 4790 0 -1 790
box -14 -8 114 272
use NOR2X1  _1368_
timestamp 1701862152
transform -1 0 3450 0 -1 790
box -12 -8 74 272
use NAND3X1  _1369_
timestamp 1702508443
transform -1 0 2850 0 1 1310
box -12 -8 92 272
use AOI21X1  _1370_
timestamp 1702508443
transform -1 0 3190 0 1 790
box -12 -8 92 272
use INVX1  _1371_
timestamp 1701862152
transform 1 0 2410 0 1 790
box -12 -8 52 272
use NAND2X1  _1372_
timestamp 1702508443
transform -1 0 3630 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1373_
timestamp 1702508443
transform 1 0 3430 0 1 790
box -12 -8 92 272
use INVX1  _1374_
timestamp 1701862152
transform -1 0 3430 0 1 270
box -12 -8 52 272
use AOI21X1  _1375_
timestamp 1702508443
transform -1 0 3570 0 1 270
box -12 -8 92 272
use NAND2X1  _1376_
timestamp 1702508443
transform -1 0 3110 0 1 1830
box -12 -8 72 272
use INVX1  _1377_
timestamp 1701862152
transform -1 0 3090 0 1 1310
box -12 -8 52 272
use NOR2X1  _1378_
timestamp 1701862152
transform -1 0 3250 0 -1 1830
box -12 -8 74 272
use OAI21X1  _1379_
timestamp 1702508443
transform 1 0 2770 0 1 1830
box -12 -8 92 272
use NAND2X1  _1380_
timestamp 1702508443
transform 1 0 3290 0 -1 1310
box -12 -8 72 272
use OR2X2  _1381_
timestamp 1702508443
transform -1 0 3210 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1382_
timestamp 1702508443
transform -1 0 3070 0 -1 1310
box -12 -8 92 272
use AND2X2  _1383_
timestamp 1701862152
transform -1 0 3110 0 -1 1830
box -12 -8 94 272
use NOR2X1  _1384_
timestamp 1701862152
transform 1 0 3330 0 1 1310
box -12 -8 74 272
use OAI21X1  _1385_
timestamp 1702508443
transform 1 0 2910 0 1 1310
box -12 -8 92 272
use NAND2X1  _1386_
timestamp 1702508443
transform 1 0 2650 0 1 790
box -12 -8 72 272
use OR2X2  _1387_
timestamp 1702508443
transform -1 0 4330 0 1 1310
box -12 -8 92 272
use NAND2X1  _1388_
timestamp 1702508443
transform 1 0 2530 0 1 1830
box -12 -8 72 272
use NAND2X1  _1389_
timestamp 1702508443
transform 1 0 2110 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1390_
timestamp 1702508443
transform 1 0 1970 0 -1 2350
box -12 -8 72 272
use AOI22X1  _1391_
timestamp 1701862152
transform 1 0 2250 0 -1 2350
box -14 -8 114 272
use INVX1  _1392_
timestamp 1701862152
transform -1 0 2470 0 -1 1830
box -12 -8 52 272
use OAI21X1  _1393_
timestamp 1702508443
transform 1 0 2290 0 -1 1830
box -12 -8 92 272
use XNOR2X1  _1394_
timestamp 1702508443
transform 1 0 2350 0 1 1830
box -12 -8 132 272
use AOI21X1  _1395_
timestamp 1702508443
transform -1 0 3190 0 -1 790
box -12 -8 92 272
use NAND3X1  _1396_
timestamp 1702508443
transform -1 0 3030 0 -1 790
box -12 -8 92 272
use INVX1  _1397_
timestamp 1701862152
transform -1 0 2870 0 -1 270
box -12 -8 52 272
use OAI21X1  _1398_
timestamp 1702508443
transform 1 0 2670 0 -1 270
box -12 -8 92 272
use AND2X2  _1399_
timestamp 1701862152
transform -1 0 2730 0 -1 790
box -12 -8 94 272
use NAND2X1  _1400_
timestamp 1702508443
transform 1 0 3250 0 -1 790
box -12 -8 72 272
use INVX1  _1401_
timestamp 1701862152
transform -1 0 2450 0 -1 790
box -12 -8 52 272
use NAND2X1  _1402_
timestamp 1702508443
transform -1 0 2570 0 -1 790
box -12 -8 72 272
use NAND3X1  _1403_
timestamp 1702508443
transform -1 0 2430 0 1 270
box -12 -8 92 272
use NAND3X1  _1404_
timestamp 1702508443
transform 1 0 2790 0 1 270
box -12 -8 92 272
use OAI21X1  _1405_
timestamp 1702508443
transform -1 0 3750 0 -1 790
box -12 -8 92 272
use AOI22X1  _1406_
timestamp 1701862152
transform -1 0 2890 0 -1 790
box -14 -8 114 272
use OR2X2  _1407_
timestamp 1702508443
transform -1 0 3030 0 1 790
box -12 -8 92 272
use NAND2X1  _1408_
timestamp 1702508443
transform 1 0 2510 0 1 790
box -12 -8 72 272
use AOI21X1  _1409_
timestamp 1702508443
transform -1 0 2870 0 1 790
box -12 -8 92 272
use OAI21X1  _1410_
timestamp 1702508443
transform -1 0 3010 0 1 270
box -12 -8 92 272
use NAND3X1  _1411_
timestamp 1702508443
transform 1 0 2930 0 -1 270
box -12 -8 92 272
use NAND3X1  _1412_
timestamp 1702508443
transform -1 0 2730 0 1 270
box -12 -8 92 272
use OAI21X1  _1413_
timestamp 1702508443
transform 1 0 3070 0 1 270
box -12 -8 92 272
use NAND3X1  _1414_
timestamp 1702508443
transform -1 0 3310 0 1 270
box -12 -8 92 272
use NAND2X1  _1415_
timestamp 1702508443
transform -1 0 3270 0 -1 270
box -12 -8 72 272
use NAND3X1  _1416_
timestamp 1702508443
transform -1 0 3430 0 -1 270
box -12 -8 92 272
use AOI21X1  _1417_
timestamp 1702508443
transform -1 0 4030 0 1 270
box -12 -8 92 272
use OAI21X1  _1418_
timestamp 1702508443
transform -1 0 3890 0 -1 270
box -12 -8 92 272
use NAND3X1  _1419_
timestamp 1702508443
transform -1 0 3150 0 -1 270
box -12 -8 92 272
use NAND2X1  _1420_
timestamp 1702508443
transform 1 0 2050 0 1 270
box -12 -8 72 272
use AOI21X1  _1421_
timestamp 1702508443
transform -1 0 2710 0 1 1310
box -12 -8 92 272
use NAND2X1  _1422_
timestamp 1702508443
transform -1 0 2910 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1423_
timestamp 1702508443
transform -1 0 2770 0 -1 1310
box -12 -8 92 272
use INVX1  _1424_
timestamp 1701862152
transform -1 0 2630 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1425_
timestamp 1701862152
transform -1 0 2570 0 1 1310
box -12 -8 74 272
use OAI21X1  _1426_
timestamp 1702508443
transform -1 0 2450 0 1 1310
box -12 -8 92 272
use NOR2X1  _1427_
timestamp 1701862152
transform 1 0 390 0 1 4430
box -12 -8 74 272
use NOR2X1  _1428_
timestamp 1701862152
transform 1 0 810 0 -1 4430
box -12 -8 74 272
use AOI21X1  _1429_
timestamp 1702508443
transform -1 0 3810 0 1 4430
box -12 -8 92 272
use OAI21X1  _1430_
timestamp 1702508443
transform -1 0 3550 0 1 4430
box -12 -8 92 272
use NOR2X1  _1431_
timestamp 1701862152
transform 1 0 1070 0 1 4430
box -12 -8 74 272
use NOR2X1  _1432_
timestamp 1701862152
transform -1 0 1110 0 -1 4430
box -12 -8 74 272
use AOI22X1  _1433_
timestamp 1701862152
transform -1 0 1270 0 -1 4430
box -14 -8 114 272
use OAI21X1  _1434_
timestamp 1702508443
transform 1 0 190 0 -1 3910
box -12 -8 92 272
use INVX1  _1435_
timestamp 1701862152
transform -1 0 590 0 1 1310
box -12 -8 52 272
use INVX1  _1436_
timestamp 1701862152
transform -1 0 230 0 -1 4950
box -12 -8 52 272
use OAI21X1  _1437_
timestamp 1702508443
transform 1 0 1910 0 1 2350
box -12 -8 92 272
use INVX1  _1438_
timestamp 1701862152
transform 1 0 2290 0 -1 790
box -12 -8 52 272
use OAI21X1  _1439_
timestamp 1702508443
transform 1 0 3170 0 1 1310
box -12 -8 92 272
use INVX1  _1440_
timestamp 1701862152
transform -1 0 1870 0 -1 270
box -12 -8 52 272
use AOI21X1  _1441_
timestamp 1702508443
transform -1 0 2270 0 1 270
box -12 -8 92 272
use NAND2X1  _1442_
timestamp 1702508443
transform -1 0 2030 0 -1 1830
box -12 -8 72 272
use INVX1  _1443_
timestamp 1701862152
transform -1 0 1750 0 1 790
box -12 -8 52 272
use NOR2X1  _1444_
timestamp 1701862152
transform -1 0 1630 0 -1 1310
box -12 -8 74 272
use OAI22X1  _1445_
timestamp 1701862152
transform 1 0 2110 0 -1 1830
box -12 -8 112 272
use NAND2X1  _1446_
timestamp 1702508443
transform 1 0 1830 0 -1 1310
box -12 -8 72 272
use NOR2X1  _1447_
timestamp 1701862152
transform 1 0 1710 0 -1 1310
box -12 -8 74 272
use INVX1  _1448_
timestamp 1701862152
transform 1 0 1430 0 1 790
box -12 -8 52 272
use NAND3X1  _1449_
timestamp 1702508443
transform -1 0 1630 0 1 790
box -12 -8 92 272
use INVX1  _1450_
timestamp 1701862152
transform -1 0 1810 0 -1 790
box -12 -8 52 272
use OAI21X1  _1451_
timestamp 1702508443
transform 1 0 1630 0 -1 790
box -12 -8 92 272
use NAND2X1  _1452_
timestamp 1702508443
transform -1 0 2110 0 1 2350
box -12 -8 72 272
use NAND2X1  _1453_
timestamp 1702508443
transform 1 0 1370 0 -1 2350
box -12 -8 72 272
use OR2X2  _1454_
timestamp 1702508443
transform -1 0 1910 0 -1 2350
box -12 -8 92 272
use INVX1  _1455_
timestamp 1701862152
transform 1 0 1730 0 -1 2350
box -12 -8 52 272
use OAI21X1  _1456_
timestamp 1702508443
transform 1 0 1830 0 -1 1830
box -12 -8 92 272
use AND2X2  _1457_
timestamp 1701862152
transform -1 0 1990 0 1 1310
box -12 -8 94 272
use AOI21X1  _1458_
timestamp 1702508443
transform 1 0 1450 0 1 270
box -12 -8 92 272
use INVX1  _1459_
timestamp 1701862152
transform -1 0 1330 0 -1 270
box -12 -8 52 272
use NAND3X1  _1460_
timestamp 1702508443
transform -1 0 1370 0 1 270
box -12 -8 92 272
use NAND3X1  _1461_
timestamp 1702508443
transform 1 0 1390 0 -1 270
box -12 -8 92 272
use OAI21X1  _1462_
timestamp 1702508443
transform -1 0 2610 0 -1 270
box -12 -8 92 272
use INVX1  _1463_
timestamp 1701862152
transform -1 0 1210 0 1 270
box -12 -8 52 272
use OAI21X1  _1464_
timestamp 1702508443
transform 1 0 1550 0 -1 270
box -12 -8 92 272
use NAND3X1  _1465_
timestamp 1702508443
transform 1 0 1690 0 -1 270
box -12 -8 92 272
use NAND3X1  _1466_
timestamp 1702508443
transform 1 0 1150 0 -1 270
box -12 -8 92 272
use OAI21X1  _1467_
timestamp 1702508443
transform 1 0 1590 0 1 270
box -12 -8 92 272
use NAND3X1  _1468_
timestamp 1702508443
transform -1 0 1830 0 1 270
box -12 -8 92 272
use NAND2X1  _1469_
timestamp 1702508443
transform 1 0 1930 0 -1 270
box -12 -8 72 272
use NAND3X1  _1470_
timestamp 1702508443
transform -1 0 2290 0 -1 270
box -12 -8 92 272
use AOI21X1  _1471_
timestamp 1702508443
transform -1 0 2570 0 1 270
box -12 -8 92 272
use OAI21X1  _1472_
timestamp 1702508443
transform -1 0 2450 0 -1 270
box -12 -8 92 272
use NAND3X1  _1473_
timestamp 1702508443
transform 1 0 2050 0 -1 270
box -12 -8 92 272
use NAND2X1  _1474_
timestamp 1702508443
transform -1 0 2230 0 -1 790
box -12 -8 72 272
use NOR3X1  _1475_
timestamp 1701862152
transform -1 0 2350 0 -1 1310
box -12 -8 172 272
use AOI21X1  _1476_
timestamp 1702508443
transform -1 0 2510 0 -1 1310
box -12 -8 92 272
use INVX1  _1477_
timestamp 1701862152
transform 1 0 1950 0 -1 1310
box -12 -8 52 272
use OAI21X1  _1478_
timestamp 1702508443
transform 1 0 2050 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1479_
timestamp 1702508443
transform -1 0 2150 0 1 1310
box -12 -8 92 272
use NAND2X1  _1480_
timestamp 1702508443
transform 1 0 4370 0 -1 4950
box -12 -8 72 272
use NAND2X1  _1481_
timestamp 1702508443
transform 1 0 4150 0 1 4430
box -12 -8 72 272
use NAND2X1  _1482_
timestamp 1702508443
transform -1 0 4330 0 1 4430
box -12 -8 72 272
use NAND2X1  _1483_
timestamp 1702508443
transform -1 0 1410 0 1 4430
box -12 -8 72 272
use OAI21X1  _1484_
timestamp 1702508443
transform 1 0 1190 0 1 4430
box -12 -8 92 272
use AOI21X1  _1485_
timestamp 1702508443
transform -1 0 1010 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1486_
timestamp 1701862152
transform 1 0 810 0 -1 1830
box -14 -8 114 272
use INVX1  _1487_
timestamp 1701862152
transform -1 0 390 0 -1 2350
box -12 -8 52 272
use OAI21X1  _1488_
timestamp 1702508443
transform -1 0 1370 0 1 790
box -12 -8 92 272
use INVX1  _1489_
timestamp 1701862152
transform -1 0 130 0 1 270
box -12 -8 52 272
use INVX1  _1490_
timestamp 1701862152
transform 1 0 1610 0 -1 2350
box -12 -8 52 272
use NAND2X1  _1491_
timestamp 1702508443
transform 1 0 2230 0 1 1830
box -12 -8 72 272
use OAI21X1  _1492_
timestamp 1702508443
transform -1 0 2150 0 1 1830
box -12 -8 92 272
use OAI21X1  _1493_
timestamp 1702508443
transform 1 0 1930 0 1 1830
box -12 -8 92 272
use OR2X2  _1494_
timestamp 1702508443
transform -1 0 1850 0 1 1830
box -12 -8 92 272
use INVX1  _1495_
timestamp 1701862152
transform 1 0 1390 0 1 1830
box -12 -8 52 272
use OAI21X1  _1496_
timestamp 1702508443
transform 1 0 1630 0 1 1830
box -12 -8 92 272
use NAND2X1  _1497_
timestamp 1702508443
transform 1 0 1570 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1498_
timestamp 1702508443
transform -1 0 1770 0 -1 1830
box -12 -8 92 272
use INVX1  _1499_
timestamp 1701862152
transform -1 0 1550 0 -1 2350
box -12 -8 52 272
use NAND3X1  _1500_
timestamp 1702508443
transform 1 0 1490 0 1 1830
box -12 -8 92 272
use NAND2X1  _1501_
timestamp 1702508443
transform 1 0 1630 0 1 1310
box -12 -8 72 272
use NOR2X1  _1502_
timestamp 1701862152
transform -1 0 550 0 1 270
box -12 -8 74 272
use NAND2X1  _1503_
timestamp 1702508443
transform 1 0 710 0 -1 270
box -12 -8 72 272
use INVX1  _1504_
timestamp 1701862152
transform -1 0 510 0 -1 270
box -12 -8 52 272
use OAI21X1  _1505_
timestamp 1702508443
transform -1 0 410 0 1 270
box -12 -8 92 272
use OR2X2  _1506_
timestamp 1702508443
transform -1 0 1070 0 -1 270
box -12 -8 92 272
use NAND3X1  _1507_
timestamp 1702508443
transform -1 0 910 0 -1 270
box -12 -8 92 272
use NAND2X1  _1508_
timestamp 1702508443
transform -1 0 830 0 1 270
box -12 -8 72 272
use NAND3X1  _1509_
timestamp 1702508443
transform -1 0 970 0 1 270
box -12 -8 92 272
use NAND2X1  _1510_
timestamp 1702508443
transform 1 0 1050 0 1 270
box -12 -8 72 272
use NAND3X1  _1511_
timestamp 1702508443
transform -1 0 690 0 1 270
box -12 -8 92 272
use NAND2X1  _1512_
timestamp 1702508443
transform 1 0 790 0 -1 790
box -12 -8 72 272
use NOR2X1  _1513_
timestamp 1701862152
transform -1 0 3510 0 1 1310
box -12 -8 74 272
use NOR2X1  _1514_
timestamp 1701862152
transform 1 0 2130 0 1 790
box -12 -8 74 272
use NAND3X1  _1515_
timestamp 1702508443
transform -1 0 2290 0 1 1310
box -12 -8 92 272
use NAND2X1  _1516_
timestamp 1702508443
transform -1 0 1970 0 1 270
box -12 -8 72 272
use AOI22X1  _1517_
timestamp 1701862152
transform 1 0 1810 0 1 790
box -14 -8 114 272
use AOI21X1  _1518_
timestamp 1702508443
transform -1 0 890 0 1 790
box -12 -8 92 272
use NAND2X1  _1519_
timestamp 1702508443
transform 1 0 1870 0 -1 790
box -12 -8 72 272
use OAI21X1  _1520_
timestamp 1702508443
transform -1 0 2090 0 -1 790
box -12 -8 92 272
use AOI21X1  _1521_
timestamp 1702508443
transform 1 0 1970 0 1 790
box -12 -8 92 272
use OAI21X1  _1522_
timestamp 1702508443
transform -1 0 2350 0 1 790
box -12 -8 92 272
use AOI22X1  _1523_
timestamp 1701862152
transform 1 0 1070 0 -1 790
box -14 -8 114 272
use OAI21X1  _1524_
timestamp 1702508443
transform -1 0 430 0 1 790
box -12 -8 92 272
use OR2X2  _1525_
timestamp 1702508443
transform 1 0 90 0 1 4430
box -12 -8 92 272
use NAND3X1  _1526_
timestamp 1702508443
transform 1 0 330 0 -1 2870
box -12 -8 92 272
use INVX1  _1527_
timestamp 1701862152
transform -1 0 4590 0 1 4430
box -12 -8 52 272
use OAI21X1  _1528_
timestamp 1702508443
transform -1 0 4710 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1529_
timestamp 1702508443
transform 1 0 4410 0 1 4430
box -12 -8 72 272
use NAND2X1  _1530_
timestamp 1702508443
transform 1 0 790 0 1 4430
box -12 -8 72 272
use OAI21X1  _1531_
timestamp 1702508443
transform -1 0 1010 0 1 4430
box -12 -8 92 272
use AOI21X1  _1532_
timestamp 1702508443
transform -1 0 1050 0 1 2350
box -12 -8 92 272
use AOI22X1  _1533_
timestamp 1701862152
transform 1 0 350 0 1 2350
box -14 -8 114 272
use INVX1  _1534_
timestamp 1701862152
transform 1 0 350 0 1 1830
box -12 -8 52 272
use INVX1  _1535_
timestamp 1701862152
transform -1 0 1450 0 1 2350
box -12 -8 52 272
use NAND2X1  _1536_
timestamp 1702508443
transform -1 0 1550 0 -1 790
box -12 -8 72 272
use INVX1  _1537_
timestamp 1701862152
transform -1 0 430 0 -1 790
box -12 -8 52 272
use AOI21X1  _1538_
timestamp 1702508443
transform -1 0 270 0 1 270
box -12 -8 92 272
use OAI21X1  _1539_
timestamp 1702508443
transform -1 0 1850 0 1 1310
box -12 -8 92 272
use NOR2X1  _1540_
timestamp 1701862152
transform 1 0 1250 0 1 1830
box -12 -8 74 272
use NAND3X1  _1541_
timestamp 1702508443
transform -1 0 1190 0 1 1830
box -12 -8 92 272
use OAI22X1  _1542_
timestamp 1701862152
transform -1 0 1490 0 -1 1830
box -12 -8 112 272
use NAND2X1  _1543_
timestamp 1702508443
transform -1 0 1190 0 -1 1830
box -12 -8 72 272
use XNOR2X1  _1544_
timestamp 1702508443
transform -1 0 1570 0 1 1310
box -12 -8 132 272
use XOR2X1  _1545_
timestamp 1702508443
transform -1 0 1230 0 1 790
box -12 -8 132 272
use XOR2X1  _1546_
timestamp 1702508443
transform 1 0 190 0 -1 790
box -12 -8 132 272
use NOR2X1  _1547_
timestamp 1701862152
transform 1 0 490 0 -1 790
box -12 -8 74 272
use OAI21X1  _1548_
timestamp 1702508443
transform -1 0 710 0 -1 790
box -12 -8 92 272
use OAI21X1  _1549_
timestamp 1702508443
transform 1 0 490 0 1 790
box -12 -8 92 272
use NAND3X1  _1550_
timestamp 1702508443
transform 1 0 650 0 1 790
box -12 -8 92 272
use AOI21X1  _1551_
timestamp 1702508443
transform -1 0 4590 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1552_
timestamp 1702508443
transform -1 0 4790 0 1 3390
box -12 -8 92 272
use INVX1  _1553_
timestamp 1701862152
transform 1 0 690 0 -1 4430
box -12 -8 52 272
use AOI21X1  _1554_
timestamp 1702508443
transform -1 0 1410 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1555_
timestamp 1702508443
transform -1 0 1310 0 1 3390
box -12 -8 92 272
use AOI22X1  _1556_
timestamp 1701862152
transform 1 0 930 0 1 1830
box -14 -8 114 272
use INVX1  _1557_
timestamp 1701862152
transform 1 0 70 0 -1 1310
box -12 -8 52 272
use NAND3X1  _1558_
timestamp 1702508443
transform 1 0 930 0 -1 790
box -12 -8 92 272
use INVX1  _1559_
timestamp 1701862152
transform 1 0 1230 0 -1 790
box -12 -8 52 272
use NAND3X1  _1560_
timestamp 1702508443
transform -1 0 1430 0 -1 790
box -12 -8 92 272
use NAND2X1  _1561_
timestamp 1702508443
transform -1 0 290 0 1 790
box -12 -8 72 272
use OAI21X1  _1562_
timestamp 1702508443
transform 1 0 90 0 1 790
box -12 -8 92 272
use INVX1  _1563_
timestamp 1701862152
transform -1 0 390 0 -1 1310
box -12 -8 52 272
use INVX1  _1564_
timestamp 1701862152
transform -1 0 1230 0 -1 1310
box -12 -8 52 272
use NAND2X1  _1565_
timestamp 1702508443
transform -1 0 1350 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1566_
timestamp 1702508443
transform -1 0 1510 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1567_
timestamp 1702508443
transform -1 0 1330 0 -1 1830
box -12 -8 92 272
use XOR2X1  _1568_
timestamp 1702508443
transform -1 0 1390 0 1 1310
box -12 -8 132 272
use NAND3X1  _1569_
timestamp 1702508443
transform -1 0 1110 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1570_
timestamp 1702508443
transform -1 0 1030 0 1 790
box -12 -8 92 272
use INVX1  _1571_
timestamp 1701862152
transform -1 0 810 0 -1 1310
box -12 -8 52 272
use OAI21X1  _1572_
timestamp 1702508443
transform 1 0 610 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1573_
timestamp 1702508443
transform -1 0 550 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1574_
timestamp 1702508443
transform -1 0 5210 0 1 3910
box -12 -8 72 272
use NOR2X1  _1575_
timestamp 1701862152
transform 1 0 5030 0 1 3910
box -12 -8 74 272
use AOI21X1  _1576_
timestamp 1702508443
transform -1 0 4950 0 1 3910
box -12 -8 92 272
use OAI21X1  _1577_
timestamp 1702508443
transform -1 0 4810 0 1 3910
box -12 -8 92 272
use NOR2X1  _1578_
timestamp 1701862152
transform 1 0 70 0 -1 4950
box -12 -8 74 272
use NOR2X1  _1579_
timestamp 1701862152
transform 1 0 90 0 -1 4430
box -12 -8 74 272
use AOI21X1  _1580_
timestamp 1702508443
transform -1 0 330 0 1 3910
box -12 -8 92 272
use AOI22X1  _1581_
timestamp 1701862152
transform 1 0 190 0 -1 1310
box -14 -8 114 272
use INVX1  _1582_
timestamp 1701862152
transform 1 0 70 0 1 1830
box -12 -8 52 272
use AOI21X1  _1583_
timestamp 1702508443
transform -1 0 970 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1584_
timestamp 1702508443
transform -1 0 1050 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1585_
timestamp 1702508443
transform -1 0 750 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1586_
timestamp 1702508443
transform -1 0 610 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1587_
timestamp 1702508443
transform -1 0 4970 0 1 1830
box -12 -8 72 272
use XNOR2X1  _1588_
timestamp 1702508443
transform -1 0 4830 0 1 1830
box -12 -8 132 272
use NAND2X1  _1589_
timestamp 1702508443
transform -1 0 1590 0 1 2350
box -12 -8 72 272
use OAI21X1  _1590_
timestamp 1702508443
transform -1 0 1290 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1591_
timestamp 1702508443
transform -1 0 1150 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1592_
timestamp 1701862152
transform 1 0 190 0 1 1830
box -14 -8 114 272
use NAND2X1  _1593_
timestamp 1702508443
transform 1 0 2570 0 -1 4430
box -12 -8 72 272
use OAI21X1  _1594_
timestamp 1702508443
transform -1 0 2790 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1595_
timestamp 1702508443
transform 1 0 3650 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1596_
timestamp 1702508443
transform 1 0 3510 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1597_
timestamp 1702508443
transform -1 0 2550 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1598_
timestamp 1702508443
transform 1 0 2350 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1599_
timestamp 1702508443
transform -1 0 3810 0 1 3910
box -12 -8 72 272
use OAI21X1  _1600_
timestamp 1702508443
transform 1 0 3610 0 1 3910
box -12 -8 92 272
use NAND2X1  _1601_
timestamp 1702508443
transform 1 0 3290 0 1 3390
box -12 -8 72 272
use OAI21X1  _1602_
timestamp 1702508443
transform 1 0 2890 0 1 3390
box -12 -8 92 272
use NAND2X1  _1603_
timestamp 1702508443
transform -1 0 2950 0 1 3910
box -12 -8 72 272
use OAI21X1  _1604_
timestamp 1702508443
transform 1 0 2750 0 1 3910
box -12 -8 92 272
use NAND2X1  _1605_
timestamp 1702508443
transform 1 0 2070 0 1 3910
box -12 -8 72 272
use OAI21X1  _1606_
timestamp 1702508443
transform 1 0 1930 0 1 3910
box -12 -8 92 272
use NAND2X1  _1607_
timestamp 1702508443
transform -1 0 1790 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1608_
timestamp 1702508443
transform 1 0 1590 0 -1 3390
box -12 -8 92 272
use DFFSR  _1609_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 3310 0 -1 4430
box -12 -8 474 272
use DFFSR  _1610_
timestamp 1701862152
transform 1 0 3810 0 1 3910
box -12 -8 474 272
use DFFSR  _1611_
timestamp 1701862152
transform 1 0 1650 0 -1 4430
box -12 -8 474 272
use DFFSR  _1612_
timestamp 1701862152
transform -1 0 3410 0 -1 3390
box -12 -8 474 272
use DFFSR  _1613_
timestamp 1701862152
transform -1 0 3290 0 1 2870
box -12 -8 474 272
use DFFSR  _1614_
timestamp 1701862152
transform 1 0 2830 0 -1 3910
box -12 -8 474 272
use DFFSR  _1615_
timestamp 1701862152
transform 1 0 1530 0 -1 3910
box -12 -8 474 272
use DFFSR  _1616_
timestamp 1701862152
transform 1 0 1790 0 1 2870
box -12 -8 474 272
use DFFSR  _1617_
timestamp 1701862152
transform -1 0 590 0 1 2870
box -12 -8 474 272
use DFFSR  _1618_
timestamp 1701862152
transform -1 0 910 0 1 2350
box -12 -8 474 272
use DFFSR  _1619_
timestamp 1701862152
transform 1 0 10 0 1 3390
box -12 -8 474 272
use DFFSR  _1620_
timestamp 1701862152
transform -1 0 1050 0 1 1310
box -12 -8 474 272
use DFFSR  _1621_
timestamp 1701862152
transform -1 0 850 0 -1 2350
box -12 -8 474 272
use DFFSR  _1622_
timestamp 1701862152
transform -1 0 850 0 1 1830
box -12 -8 474 272
use DFFSR  _1623_
timestamp 1701862152
transform -1 0 470 0 1 1310
box -12 -8 474 272
use DFFSR  _1624_
timestamp 1701862152
transform -1 0 470 0 -1 1830
box -12 -8 474 272
use DFFSR  _1625_
timestamp 1701862152
transform 1 0 2130 0 1 4430
box -12 -8 474 272
use DFFSR  _1626_
timestamp 1701862152
transform 1 0 3350 0 1 3390
box -12 -8 474 272
use DFFSR  _1627_
timestamp 1701862152
transform 1 0 2070 0 1 3390
box -12 -8 474 272
use DFFSR  _1628_
timestamp 1701862152
transform -1 0 3530 0 1 3910
box -12 -8 474 272
use DFFSR  _1629_
timestamp 1701862152
transform 1 0 2250 0 1 2870
box -12 -8 474 272
use DFFSR  _1630_
timestamp 1701862152
transform 1 0 2190 0 -1 2870
box -12 -8 474 272
use DFFSR  _1631_
timestamp 1701862152
transform 1 0 1410 0 1 4430
box -12 -8 474 272
use DFFSR  _1632_
timestamp 1701862152
transform -1 0 1790 0 1 2870
box -12 -8 474 272
use DFFSR  _1633_
timestamp 1701862152
transform 1 0 150 0 -1 3390
box -12 -8 474 272
use DFFSR  _1634_
timestamp 1701862152
transform 1 0 750 0 -1 3390
box -12 -8 474 272
use DFFSR  _1635_
timestamp 1701862152
transform 1 0 870 0 1 2870
box -12 -8 474 272
use INVX1  _1636_
timestamp 1701862152
transform -1 0 4290 0 1 5990
box -12 -8 52 272
use INVX4  _1637_
timestamp 1701862152
transform -1 0 4430 0 1 5990
box -12 -8 72 272
use OAI21X1  _1638_
timestamp 1702508443
transform -1 0 4190 0 1 5990
box -12 -8 92 272
use NOR2X1  _1639_
timestamp 1701862152
transform 1 0 3990 0 1 5990
box -12 -8 74 272
use INVX1  _1640_
timestamp 1701862152
transform -1 0 3750 0 1 5990
box -12 -8 52 272
use INVX2  _1641_
timestamp 1701862152
transform -1 0 3690 0 -1 4950
box -12 -8 52 272
use NAND2X1  _1642_
timestamp 1702508443
transform -1 0 3290 0 -1 4950
box -12 -8 72 272
use INVX2  _1643_
timestamp 1701862152
transform -1 0 4150 0 1 4950
box -12 -8 52 272
use NAND2X1  _1644_
timestamp 1702508443
transform -1 0 4170 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1645_
timestamp 1702508443
transform 1 0 4510 0 -1 5470
box -12 -8 72 272
use AOI22X1  _1646_
timestamp 1701862152
transform -1 0 4350 0 -1 5470
box -14 -8 114 272
use INVX2  _1647_
timestamp 1701862152
transform 1 0 3330 0 1 4950
box -12 -8 52 272
use INVX1  _1648_
timestamp 1701862152
transform -1 0 4290 0 1 5470
box -12 -8 52 272
use INVX1  _1649_
timestamp 1701862152
transform -1 0 3870 0 -1 5470
box -12 -8 52 272
use OAI21X1  _1650_
timestamp 1702508443
transform -1 0 4050 0 1 5470
box -12 -8 92 272
use NAND2X1  _1651_
timestamp 1702508443
transform 1 0 3690 0 1 5470
box -12 -8 72 272
use NAND2X1  _1652_
timestamp 1702508443
transform 1 0 3710 0 -1 5990
box -12 -8 72 272
use OAI21X1  _1653_
timestamp 1702508443
transform 1 0 3810 0 1 5470
box -12 -8 92 272
use OAI21X1  _1654_
timestamp 1702508443
transform -1 0 4730 0 1 5990
box -12 -8 92 272
use AOI21X1  _1655_
timestamp 1702508443
transform -1 0 4570 0 1 5990
box -12 -8 92 272
use NOR2X1  _1656_
timestamp 1701862152
transform 1 0 1510 0 1 5990
box -12 -8 74 272
use OAI21X1  _1657_
timestamp 1702508443
transform 1 0 3130 0 1 5990
box -12 -8 92 272
use OAI21X1  _1658_
timestamp 1702508443
transform 1 0 3290 0 1 5990
box -12 -8 92 272
use XOR2X1  _1659_
timestamp 1702508443
transform -1 0 3330 0 -1 5990
box -12 -8 132 272
use NOR2X1  _1660_
timestamp 1701862152
transform 1 0 3590 0 1 5990
box -12 -8 74 272
use OAI21X1  _1661_
timestamp 1702508443
transform -1 0 3510 0 1 5990
box -12 -8 92 272
use NAND2X1  _1662_
timestamp 1702508443
transform 1 0 3590 0 1 4950
box -12 -8 72 272
use NAND3X1  _1663_
timestamp 1702508443
transform -1 0 3590 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1664_
timestamp 1701862152
transform -1 0 3450 0 -1 4950
box -14 -8 114 272
use INVX1  _1665_
timestamp 1701862152
transform -1 0 4050 0 1 4950
box -12 -8 52 272
use NOR2X1  _1666_
timestamp 1701862152
transform 1 0 3870 0 1 4950
box -12 -8 74 272
use OAI21X1  _1667_
timestamp 1702508443
transform -1 0 3810 0 1 4950
box -12 -8 92 272
use OAI21X1  _1668_
timestamp 1702508443
transform 1 0 3430 0 1 4950
box -12 -8 92 272
use OAI21X1  _1669_
timestamp 1702508443
transform -1 0 3630 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1670_
timestamp 1702508443
transform -1 0 3470 0 -1 5990
box -12 -8 92 272
use INVX1  _1671_
timestamp 1701862152
transform -1 0 3150 0 -1 5990
box -12 -8 52 272
use OAI21X1  _1672_
timestamp 1702508443
transform 1 0 2770 0 -1 5990
box -12 -8 92 272
use MUX2X1  _1673_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform -1 0 3030 0 -1 5990
box -12 -8 114 272
use NAND2X1  _1674_
timestamp 1702508443
transform 1 0 3010 0 1 5990
box -12 -8 72 272
use INVX1  _1675_
timestamp 1701862152
transform -1 0 4470 0 -1 5990
box -12 -8 52 272
use OAI21X1  _1676_
timestamp 1702508443
transform 1 0 4150 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1677_
timestamp 1702508443
transform 1 0 3850 0 -1 5990
box -12 -8 92 272
use MUX2X1  _1678_
timestamp 1701862152
transform 1 0 4350 0 1 5470
box -12 -8 114 272
use NAND2X1  _1679_
timestamp 1702508443
transform 1 0 4650 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1680_
timestamp 1702508443
transform -1 0 4570 0 1 5470
box -12 -8 72 272
use AOI21X1  _1681_
timestamp 1702508443
transform 1 0 3950 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1682_
timestamp 1702508443
transform 1 0 4110 0 1 5470
box -12 -8 72 272
use NAND3X1  _1683_
timestamp 1702508443
transform 1 0 4010 0 -1 5990
box -12 -8 92 272
use AOI22X1  _1684_
timestamp 1701862152
transform 1 0 3810 0 1 5990
box -14 -8 114 272
use OAI21X1  _1685_
timestamp 1702508443
transform -1 0 2950 0 1 5990
box -12 -8 92 272
use OAI21X1  _1686_
timestamp 1702508443
transform -1 0 2650 0 1 5990
box -12 -8 92 272
use NAND2X1  _1687_
timestamp 1702508443
transform 1 0 2450 0 1 5990
box -12 -8 72 272
use NAND2X1  _1688_
timestamp 1702508443
transform -1 0 2250 0 1 5990
box -12 -8 72 272
use INVX1  _1689_
timestamp 1701862152
transform -1 0 1710 0 -1 4950
box -12 -8 52 272
use NOR2X1  _1690_
timestamp 1701862152
transform 1 0 2730 0 1 5990
box -12 -8 74 272
use OAI21X1  _1691_
timestamp 1702508443
transform -1 0 2390 0 1 5990
box -12 -8 92 272
use NAND2X1  _1692_
timestamp 1702508443
transform -1 0 3090 0 1 5470
box -12 -8 72 272
use NAND3X1  _1693_
timestamp 1702508443
transform 1 0 3190 0 1 4950
box -12 -8 92 272
use AOI22X1  _1694_
timestamp 1701862152
transform 1 0 3210 0 -1 5470
box -14 -8 114 272
use INVX1  _1695_
timestamp 1701862152
transform -1 0 3630 0 1 5470
box -12 -8 52 272
use NOR2X1  _1696_
timestamp 1701862152
transform 1 0 3470 0 1 5470
box -12 -8 74 272
use OAI21X1  _1697_
timestamp 1702508443
transform -1 0 3390 0 1 5470
box -12 -8 92 272
use OAI21X1  _1698_
timestamp 1702508443
transform -1 0 3250 0 1 5470
box -12 -8 92 272
use OAI21X1  _1699_
timestamp 1702508443
transform -1 0 2530 0 1 5470
box -12 -8 92 272
use AOI21X1  _1700_
timestamp 1702508443
transform 1 0 2310 0 1 5470
box -12 -8 92 272
use OAI21X1  _1701_
timestamp 1702508443
transform -1 0 2310 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1702_
timestamp 1702508443
transform 1 0 2090 0 -1 5990
box -12 -8 92 272
use XOR2X1  _1703_
timestamp 1702508443
transform 1 0 1310 0 1 5990
box -12 -8 132 272
use INVX1  _1704_
timestamp 1701862152
transform -1 0 1310 0 -1 4950
box -12 -8 52 272
use INVX1  _1705_
timestamp 1701862152
transform 1 0 2370 0 -1 5990
box -12 -8 52 272
use OAI21X1  _1706_
timestamp 1702508443
transform -1 0 2570 0 -1 5990
box -12 -8 92 272
use INVX1  _1707_
timestamp 1701862152
transform 1 0 1930 0 1 5990
box -12 -8 52 272
use AOI22X1  _1708_
timestamp 1701862152
transform -1 0 2010 0 -1 5990
box -14 -8 114 272
use NAND2X1  _1709_
timestamp 1702508443
transform -1 0 2710 0 1 4430
box -12 -8 72 272
use AND2X2  _1710_
timestamp 1701862152
transform -1 0 3130 0 1 4950
box -12 -8 94 272
use NAND2X1  _1711_
timestamp 1702508443
transform 1 0 2930 0 1 4950
box -12 -8 72 272
use AOI22X1  _1712_
timestamp 1701862152
transform 1 0 2450 0 1 4950
box -14 -8 114 272
use OAI21X1  _1713_
timestamp 1702508443
transform -1 0 2850 0 1 4950
box -12 -8 92 272
use OAI21X1  _1714_
timestamp 1702508443
transform -1 0 2690 0 1 4950
box -12 -8 92 272
use OAI21X1  _1715_
timestamp 1702508443
transform 1 0 2750 0 1 5470
box -12 -8 92 272
use AOI21X1  _1716_
timestamp 1702508443
transform 1 0 2590 0 1 5470
box -12 -8 92 272
use OAI21X1  _1717_
timestamp 1702508443
transform -1 0 2710 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1718_
timestamp 1702508443
transform -1 0 2550 0 -1 5470
box -12 -8 92 272
use XOR2X1  _1719_
timestamp 1702508443
transform 1 0 2110 0 1 5470
box -12 -8 132 272
use XNOR2X1  _1720_
timestamp 1702508443
transform 1 0 1910 0 1 5470
box -12 -8 132 272
use NAND2X1  _1721_
timestamp 1702508443
transform 1 0 1650 0 1 5990
box -12 -8 72 272
use NAND3X1  _1722_
timestamp 1702508443
transform -1 0 2110 0 1 5990
box -12 -8 92 272
use NAND3X1  _1723_
timestamp 1702508443
transform 1 0 1790 0 1 5990
box -12 -8 92 272
use NAND2X1  _1724_
timestamp 1702508443
transform 1 0 1230 0 1 5470
box -12 -8 72 272
use OAI21X1  _1725_
timestamp 1702508443
transform 1 0 2030 0 -1 5470
box -12 -8 92 272
use INVX1  _1726_
timestamp 1701862152
transform -1 0 950 0 -1 5470
box -12 -8 52 272
use OAI21X1  _1727_
timestamp 1702508443
transform -1 0 1110 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1728_
timestamp 1702508443
transform 1 0 2650 0 -1 4950
box -12 -8 72 272
use AND2X2  _1729_
timestamp 1701862152
transform 1 0 1950 0 -1 4950
box -12 -8 94 272
use NAND2X1  _1730_
timestamp 1702508443
transform -1 0 2290 0 -1 4950
box -12 -8 72 272
use AOI22X1  _1731_
timestamp 1701862152
transform -1 0 2390 0 1 4950
box -14 -8 114 272
use OAI21X1  _1732_
timestamp 1702508443
transform 1 0 2090 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1733_
timestamp 1702508443
transform 1 0 2130 0 1 4950
box -12 -8 92 272
use OAI21X1  _1734_
timestamp 1702508443
transform -1 0 1870 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1735_
timestamp 1702508443
transform -1 0 1910 0 1 4950
box -12 -8 92 272
use OAI21X1  _1736_
timestamp 1702508443
transform 1 0 1690 0 1 4950
box -12 -8 92 272
use OAI21X1  _1737_
timestamp 1702508443
transform -1 0 1610 0 1 4950
box -12 -8 92 272
use INVX1  _1738_
timestamp 1701862152
transform -1 0 1210 0 1 4950
box -12 -8 52 272
use XOR2X1  _1739_
timestamp 1702508443
transform -1 0 1070 0 -1 4950
box -12 -8 132 272
use INVX1  _1740_
timestamp 1701862152
transform -1 0 1330 0 1 4950
box -12 -8 52 272
use AOI21X1  _1741_
timestamp 1702508443
transform -1 0 1090 0 1 4950
box -12 -8 92 272
use NAND2X1  _1742_
timestamp 1702508443
transform -1 0 2410 0 -1 4430
box -12 -8 72 272
use AND2X2  _1743_
timestamp 1701862152
transform -1 0 3150 0 -1 4950
box -12 -8 94 272
use NAND2X1  _1744_
timestamp 1702508443
transform 1 0 2790 0 -1 4950
box -12 -8 72 272
use AOI22X1  _1745_
timestamp 1701862152
transform 1 0 2490 0 -1 4950
box -14 -8 114 272
use OAI21X1  _1746_
timestamp 1702508443
transform -1 0 3010 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1747_
timestamp 1702508443
transform -1 0 2430 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1748_
timestamp 1702508443
transform -1 0 1610 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1749_
timestamp 1702508443
transform -1 0 1450 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1750_
timestamp 1702508443
transform -1 0 950 0 1 4950
box -12 -8 92 272
use OAI21X1  _1751_
timestamp 1702508443
transform -1 0 890 0 -1 4950
box -12 -8 92 272
use INVX1  _1752_
timestamp 1701862152
transform -1 0 490 0 -1 4950
box -12 -8 52 272
use XOR2X1  _1753_
timestamp 1702508443
transform 1 0 350 0 1 4950
box -12 -8 132 272
use INVX1  _1754_
timestamp 1701862152
transform -1 0 590 0 -1 4950
box -12 -8 52 272
use OAI21X1  _1755_
timestamp 1702508443
transform -1 0 750 0 -1 4950
box -12 -8 92 272
use INVX1  _1756_
timestamp 1701862152
transform -1 0 1330 0 -1 5470
box -12 -8 52 272
use AND2X2  _1757_
timestamp 1701862152
transform 1 0 1990 0 1 4950
box -12 -8 94 272
use NAND2X1  _1758_
timestamp 1702508443
transform -1 0 2230 0 -1 5470
box -12 -8 72 272
use AOI22X1  _1759_
timestamp 1701862152
transform -1 0 2410 0 -1 5470
box -14 -8 114 272
use OAI21X1  _1760_
timestamp 1702508443
transform -1 0 1950 0 -1 5470
box -12 -8 92 272
use OAI22X1  _1761_
timestamp 1701862152
transform 1 0 1710 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1762_
timestamp 1702508443
transform -1 0 1590 0 1 5470
box -12 -8 92 272
use AOI21X1  _1763_
timestamp 1702508443
transform -1 0 1450 0 1 5470
box -12 -8 92 272
use OAI21X1  _1764_
timestamp 1702508443
transform -1 0 990 0 1 5470
box -12 -8 92 272
use OAI21X1  _1765_
timestamp 1702508443
transform -1 0 850 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1766_
timestamp 1702508443
transform -1 0 690 0 -1 5470
box -12 -8 72 272
use INVX1  _1767_
timestamp 1701862152
transform 1 0 1190 0 -1 5470
box -12 -8 52 272
use AOI21X1  _1768_
timestamp 1702508443
transform 1 0 1390 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1769_
timestamp 1702508443
transform -1 0 1630 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1770_
timestamp 1702508443
transform -1 0 1470 0 1 4950
box -12 -8 92 272
use OR2X2  _1771_
timestamp 1702508443
transform -1 0 790 0 1 4950
box -12 -8 92 272
use AOI22X1  _1772_
timestamp 1701862152
transform -1 0 630 0 1 4950
box -14 -8 114 272
use INVX1  _1773_
timestamp 1701862152
transform 1 0 810 0 1 5470
box -12 -8 52 272
use NAND2X1  _1774_
timestamp 1702508443
transform 1 0 370 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1775_
timestamp 1702508443
transform 1 0 90 0 1 4950
box -12 -8 72 272
use OAI21X1  _1776_
timestamp 1702508443
transform -1 0 570 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1777_
timestamp 1702508443
transform -1 0 3770 0 -1 5470
box -12 -8 72 272
use AND2X2  _1778_
timestamp 1701862152
transform 1 0 2790 0 -1 5470
box -12 -8 94 272
use NAND2X1  _1779_
timestamp 1702508443
transform -1 0 3130 0 -1 5470
box -12 -8 72 272
use AOI22X1  _1780_
timestamp 1701862152
transform -1 0 3650 0 -1 5470
box -14 -8 114 272
use OAI21X1  _1781_
timestamp 1702508443
transform 1 0 2930 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1782_
timestamp 1702508443
transform 1 0 3390 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1783_
timestamp 1702508443
transform -1 0 1590 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1784_
timestamp 1702508443
transform -1 0 1450 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1785_
timestamp 1702508443
transform -1 0 1250 0 1 5990
box -12 -8 92 272
use OAI21X1  _1786_
timestamp 1702508443
transform -1 0 1110 0 1 5990
box -12 -8 92 272
use NAND2X1  _1787_
timestamp 1702508443
transform -1 0 630 0 1 5990
box -12 -8 72 272
use NAND2X1  _1788_
timestamp 1702508443
transform 1 0 670 0 1 5470
box -12 -8 72 272
use INVX1  _1789_
timestamp 1701862152
transform -1 0 670 0 -1 5990
box -12 -8 52 272
use NAND3X1  _1790_
timestamp 1702508443
transform -1 0 570 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1791_
timestamp 1702508443
transform -1 0 410 0 -1 5990
box -12 -8 72 272
use NOR2X1  _1792_
timestamp 1701862152
transform -1 0 1850 0 1 5470
box -12 -8 74 272
use NAND2X1  _1793_
timestamp 1702508443
transform 1 0 1650 0 1 5470
box -12 -8 72 272
use NOR2X1  _1794_
timestamp 1701862152
transform 1 0 670 0 1 4430
box -12 -8 74 272
use NAND3X1  _1795_
timestamp 1702508443
transform -1 0 290 0 1 4950
box -12 -8 92 272
use NOR2X1  _1796_
timestamp 1701862152
transform 1 0 310 0 -1 4950
box -12 -8 74 272
use AND2X2  _1797_
timestamp 1701862152
transform 1 0 510 0 1 4430
box -12 -8 94 272
use NAND3X1  _1798_
timestamp 1702508443
transform -1 0 790 0 1 5990
box -12 -8 92 272
use NAND2X1  _1799_
timestamp 1702508443
transform 1 0 450 0 1 5990
box -12 -8 72 272
use NAND2X1  _1800_
timestamp 1702508443
transform 1 0 230 0 1 5990
box -12 -8 72 272
use NAND2X1  _1801_
timestamp 1702508443
transform -1 0 310 0 -1 5470
box -12 -8 72 272
use NOR2X1  _1802_
timestamp 1701862152
transform -1 0 2950 0 1 5470
box -12 -8 74 272
use OAI21X1  _1803_
timestamp 1702508443
transform 1 0 870 0 1 5990
box -12 -8 92 272
use NOR2X1  _1804_
timestamp 1701862152
transform -1 0 790 0 -1 5990
box -12 -8 74 272
use AOI21X1  _1805_
timestamp 1702508443
transform 1 0 870 0 -1 5990
box -12 -8 92 272
use XOR2X1  _1806_
timestamp 1702508443
transform 1 0 1050 0 1 5470
box -12 -8 132 272
use OAI21X1  _1807_
timestamp 1702508443
transform -1 0 170 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1808_
timestamp 1702508443
transform -1 0 590 0 1 5470
box -12 -8 92 272
use AOI21X1  _1809_
timestamp 1702508443
transform -1 0 1290 0 -1 5990
box -12 -8 92 272
use XOR2X1  _1810_
timestamp 1702508443
transform -1 0 1130 0 -1 5990
box -12 -8 132 272
use NAND3X1  _1811_
timestamp 1702508443
transform -1 0 290 0 -1 5990
box -12 -8 92 272
use INVX1  _1812_
timestamp 1701862152
transform -1 0 390 0 1 5990
box -12 -8 52 272
use NAND3X1  _1813_
timestamp 1702508443
transform -1 0 170 0 1 5990
box -12 -8 92 272
use NAND2X1  _1814_
timestamp 1702508443
transform -1 0 130 0 -1 5990
box -12 -8 72 272
use NAND3X1  _1815_
timestamp 1702508443
transform -1 0 450 0 1 5470
box -12 -8 92 272
use NAND3X1  _1816_
timestamp 1702508443
transform 1 0 70 0 1 5470
box -12 -8 92 272
use NAND2X1  _1817_
timestamp 1702508443
transform -1 0 290 0 1 5470
box -12 -8 72 272
use BUFX2  _1818_ ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1702508443
transform -1 0 130 0 -1 2870
box -12 -8 72 272
use BUFX2  _1819_
timestamp 1702508443
transform -1 0 270 0 -1 2870
box -12 -8 72 272
use BUFX2  _1820_
timestamp 1702508443
transform -1 0 130 0 -1 3910
box -12 -8 72 272
use BUFX2  _1821_
timestamp 1702508443
transform 1 0 590 0 -1 270
box -12 -8 72 272
use BUFX2  _1822_
timestamp 1702508443
transform -1 0 390 0 -1 270
box -12 -8 72 272
use BUFX2  _1823_
timestamp 1702508443
transform -1 0 270 0 -1 270
box -12 -8 72 272
use BUFX2  _1824_
timestamp 1702508443
transform 1 0 90 0 -1 270
box -12 -8 72 272
use BUFX2  _1825_
timestamp 1702508443
transform 1 0 70 0 -1 790
box -12 -8 72 272
use BUFX2  _1826_
timestamp 1702508443
transform 1 0 1130 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert0
timestamp 1702508443
transform -1 0 2890 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert1
timestamp 1702508443
transform 1 0 3430 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert2
timestamp 1702508443
transform 1 0 3510 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert3
timestamp 1702508443
transform -1 0 2910 0 -1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert4
timestamp 1702508443
transform -1 0 4650 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert5
timestamp 1702508443
transform 1 0 4590 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert6
timestamp 1702508443
transform 1 0 4650 0 1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert7
timestamp 1702508443
transform 1 0 4770 0 1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert13
timestamp 1702508443
transform 1 0 3170 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert14
timestamp 1702508443
transform 1 0 2750 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert15
timestamp 1702508443
transform -1 0 2070 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert16
timestamp 1702508443
transform -1 0 1950 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert17
timestamp 1702508443
transform 1 0 470 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert18
timestamp 1702508443
transform 1 0 3370 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert19
timestamp 1702508443
transform 1 0 1850 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert20
timestamp 1702508443
transform 1 0 1470 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert21
timestamp 1702508443
transform -1 0 150 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert22
timestamp 1702508443
transform -1 0 2830 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert23
timestamp 1702508443
transform 1 0 3570 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert24
timestamp 1702508443
transform 1 0 3870 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert25
timestamp 1702508443
transform -1 0 3110 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert26
timestamp 1702508443
transform 1 0 3010 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert27
timestamp 1702508443
transform 1 0 2610 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert28
timestamp 1702508443
transform -1 0 1570 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert29
timestamp 1702508443
transform 1 0 2610 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert30
timestamp 1702508443
transform -1 0 2530 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert31
timestamp 1702508443
transform 1 0 2970 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert32
timestamp 1702508443
transform 1 0 2010 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert33
timestamp 1702508443
transform 1 0 3370 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert34
timestamp 1702508443
transform -1 0 3670 0 1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert35
timestamp 1702508443
transform -1 0 4070 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert36
timestamp 1702508443
transform 1 0 4010 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert37
timestamp 1702508443
transform -1 0 3910 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert38
timestamp 1702508443
transform 1 0 1770 0 -1 5990
box -12 -8 72 272
use BUFX2  BUFX2_insert39
timestamp 1702508443
transform -1 0 4610 0 -1 5990
box -12 -8 72 272
use BUFX2  BUFX2_insert40
timestamp 1702508443
transform -1 0 1710 0 -1 5990
box -12 -8 72 272
use BUFX2  BUFX2_insert41
timestamp 1702508443
transform -1 0 2710 0 -1 5990
box -12 -8 72 272
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701862152
transform 1 0 2230 0 -1 3390
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1701862152
transform 1 0 1490 0 -1 2870
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1701862152
transform 1 0 90 0 1 2350
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1701862152
transform -1 0 2150 0 -1 3390
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1701862152
transform 1 0 90 0 -1 2350
box -12 -8 192 272
use FILL  FILL91350x150 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/layout/digital_ETRI
timestamp 1701859473
transform -1 0 6110 0 -1 270
box -12 -8 32 272
use FILL  FILL91350x7950
timestamp 1701859473
transform -1 0 6110 0 -1 790
box -12 -8 32 272
use FILL  FILL91350x11850
timestamp 1701859473
transform 1 0 6090 0 1 790
box -12 -8 32 272
use FILL  FILL91350x27450
timestamp 1701859473
transform 1 0 6090 0 1 1830
box -12 -8 32 272
use FILL  FILL91350x54750
timestamp 1701859473
transform -1 0 6110 0 -1 3910
box -12 -8 32 272
use FILL  FILL91650x150
timestamp 1701859473
transform -1 0 6130 0 -1 270
box -12 -8 32 272
use FILL  FILL91650x7950
timestamp 1701859473
transform -1 0 6130 0 -1 790
box -12 -8 32 272
use FILL  FILL91650x11850
timestamp 1701859473
transform 1 0 6110 0 1 790
box -12 -8 32 272
use FILL  FILL91650x19650
timestamp 1701859473
transform 1 0 6110 0 1 1310
box -12 -8 32 272
use FILL  FILL91650x27450
timestamp 1701859473
transform 1 0 6110 0 1 1830
box -12 -8 32 272
use FILL  FILL91650x35250
timestamp 1701859473
transform 1 0 6110 0 1 2350
box -12 -8 32 272
use FILL  FILL91650x54750
timestamp 1701859473
transform -1 0 6130 0 -1 3910
box -12 -8 32 272
use FILL  FILL91650x70350
timestamp 1701859473
transform -1 0 6130 0 -1 4950
box -12 -8 32 272
use FILL  FILL91650x82050
timestamp 1701859473
transform 1 0 6110 0 1 5470
box -12 -8 32 272
use FILL  FILL91950x150
timestamp 1701859473
transform -1 0 6150 0 -1 270
box -12 -8 32 272
use FILL  FILL91950x4050
timestamp 1701859473
transform 1 0 6130 0 1 270
box -12 -8 32 272
use FILL  FILL91950x7950
timestamp 1701859473
transform -1 0 6150 0 -1 790
box -12 -8 32 272
use FILL  FILL91950x11850
timestamp 1701859473
transform 1 0 6130 0 1 790
box -12 -8 32 272
use FILL  FILL91950x19650
timestamp 1701859473
transform 1 0 6130 0 1 1310
box -12 -8 32 272
use FILL  FILL91950x27450
timestamp 1701859473
transform 1 0 6130 0 1 1830
box -12 -8 32 272
use FILL  FILL91950x35250
timestamp 1701859473
transform 1 0 6130 0 1 2350
box -12 -8 32 272
use FILL  FILL91950x54750
timestamp 1701859473
transform -1 0 6150 0 -1 3910
box -12 -8 32 272
use FILL  FILL91950x62550
timestamp 1701859473
transform -1 0 6150 0 -1 4430
box -12 -8 32 272
use FILL  FILL91950x70350
timestamp 1701859473
transform -1 0 6150 0 -1 4950
box -12 -8 32 272
use FILL  FILL91950x78150
timestamp 1701859473
transform -1 0 6150 0 -1 5470
box -12 -8 32 272
use FILL  FILL91950x82050
timestamp 1701859473
transform 1 0 6130 0 1 5470
box -12 -8 32 272
use FILL  FILL91950x89850
timestamp 1701859473
transform 1 0 6130 0 1 5990
box -12 -8 32 272
use FILL  FILL92250x150
timestamp 1701859473
transform -1 0 6170 0 -1 270
box -12 -8 32 272
use FILL  FILL92250x4050
timestamp 1701859473
transform 1 0 6150 0 1 270
box -12 -8 32 272
use FILL  FILL92250x7950
timestamp 1701859473
transform -1 0 6170 0 -1 790
box -12 -8 32 272
use FILL  FILL92250x11850
timestamp 1701859473
transform 1 0 6150 0 1 790
box -12 -8 32 272
use FILL  FILL92250x15750
timestamp 1701859473
transform -1 0 6170 0 -1 1310
box -12 -8 32 272
use FILL  FILL92250x19650
timestamp 1701859473
transform 1 0 6150 0 1 1310
box -12 -8 32 272
use FILL  FILL92250x27450
timestamp 1701859473
transform 1 0 6150 0 1 1830
box -12 -8 32 272
use FILL  FILL92250x35250
timestamp 1701859473
transform 1 0 6150 0 1 2350
box -12 -8 32 272
use FILL  FILL92250x54750
timestamp 1701859473
transform -1 0 6170 0 -1 3910
box -12 -8 32 272
use FILL  FILL92250x62550
timestamp 1701859473
transform -1 0 6170 0 -1 4430
box -12 -8 32 272
use FILL  FILL92250x70350
timestamp 1701859473
transform -1 0 6170 0 -1 4950
box -12 -8 32 272
use FILL  FILL92250x74250
timestamp 1701859473
transform 1 0 6150 0 1 4950
box -12 -8 32 272
use FILL  FILL92250x78150
timestamp 1701859473
transform -1 0 6170 0 -1 5470
box -12 -8 32 272
use FILL  FILL92250x82050
timestamp 1701859473
transform 1 0 6150 0 1 5470
box -12 -8 32 272
use FILL  FILL92250x89850
timestamp 1701859473
transform 1 0 6150 0 1 5990
box -12 -8 32 272
use FILL  FILL92550x150
timestamp 1701859473
transform -1 0 6190 0 -1 270
box -12 -8 32 272
use FILL  FILL92550x4050
timestamp 1701859473
transform 1 0 6170 0 1 270
box -12 -8 32 272
use FILL  FILL92550x7950
timestamp 1701859473
transform -1 0 6190 0 -1 790
box -12 -8 32 272
use FILL  FILL92550x11850
timestamp 1701859473
transform 1 0 6170 0 1 790
box -12 -8 32 272
use FILL  FILL92550x15750
timestamp 1701859473
transform -1 0 6190 0 -1 1310
box -12 -8 32 272
use FILL  FILL92550x19650
timestamp 1701859473
transform 1 0 6170 0 1 1310
box -12 -8 32 272
use FILL  FILL92550x23550
timestamp 1701859473
transform -1 0 6190 0 -1 1830
box -12 -8 32 272
use FILL  FILL92550x27450
timestamp 1701859473
transform 1 0 6170 0 1 1830
box -12 -8 32 272
use FILL  FILL92550x35250
timestamp 1701859473
transform 1 0 6170 0 1 2350
box -12 -8 32 272
use FILL  FILL92550x54750
timestamp 1701859473
transform -1 0 6190 0 -1 3910
box -12 -8 32 272
use FILL  FILL92550x62550
timestamp 1701859473
transform -1 0 6190 0 -1 4430
box -12 -8 32 272
use FILL  FILL92550x70350
timestamp 1701859473
transform -1 0 6190 0 -1 4950
box -12 -8 32 272
use FILL  FILL92550x74250
timestamp 1701859473
transform 1 0 6170 0 1 4950
box -12 -8 32 272
use FILL  FILL92550x78150
timestamp 1701859473
transform -1 0 6190 0 -1 5470
box -12 -8 32 272
use FILL  FILL92550x82050
timestamp 1701859473
transform 1 0 6170 0 1 5470
box -12 -8 32 272
use FILL  FILL92550x85950
timestamp 1701859473
transform -1 0 6190 0 -1 5990
box -12 -8 32 272
use FILL  FILL92550x89850
timestamp 1701859473
transform 1 0 6170 0 1 5990
box -12 -8 32 272
use FILL  FILL92850x150
timestamp 1701859473
transform -1 0 6210 0 -1 270
box -12 -8 32 272
use FILL  FILL92850x4050
timestamp 1701859473
transform 1 0 6190 0 1 270
box -12 -8 32 272
use FILL  FILL92850x7950
timestamp 1701859473
transform -1 0 6210 0 -1 790
box -12 -8 32 272
use FILL  FILL92850x11850
timestamp 1701859473
transform 1 0 6190 0 1 790
box -12 -8 32 272
use FILL  FILL92850x15750
timestamp 1701859473
transform -1 0 6210 0 -1 1310
box -12 -8 32 272
use FILL  FILL92850x19650
timestamp 1701859473
transform 1 0 6190 0 1 1310
box -12 -8 32 272
use FILL  FILL92850x23550
timestamp 1701859473
transform -1 0 6210 0 -1 1830
box -12 -8 32 272
use FILL  FILL92850x27450
timestamp 1701859473
transform 1 0 6190 0 1 1830
box -12 -8 32 272
use FILL  FILL92850x31350
timestamp 1701859473
transform -1 0 6210 0 -1 2350
box -12 -8 32 272
use FILL  FILL92850x35250
timestamp 1701859473
transform 1 0 6190 0 1 2350
box -12 -8 32 272
use FILL  FILL92850x54750
timestamp 1701859473
transform -1 0 6210 0 -1 3910
box -12 -8 32 272
use FILL  FILL92850x62550
timestamp 1701859473
transform -1 0 6210 0 -1 4430
box -12 -8 32 272
use FILL  FILL92850x70350
timestamp 1701859473
transform -1 0 6210 0 -1 4950
box -12 -8 32 272
use FILL  FILL92850x74250
timestamp 1701859473
transform 1 0 6190 0 1 4950
box -12 -8 32 272
use FILL  FILL92850x78150
timestamp 1701859473
transform -1 0 6210 0 -1 5470
box -12 -8 32 272
use FILL  FILL92850x82050
timestamp 1701859473
transform 1 0 6190 0 1 5470
box -12 -8 32 272
use FILL  FILL92850x85950
timestamp 1701859473
transform -1 0 6210 0 -1 5990
box -12 -8 32 272
use FILL  FILL92850x89850
timestamp 1701859473
transform 1 0 6190 0 1 5990
box -12 -8 32 272
use FILL  FILL93150x150
timestamp 1701859473
transform -1 0 6230 0 -1 270
box -12 -8 32 272
use FILL  FILL93150x4050
timestamp 1701859473
transform 1 0 6210 0 1 270
box -12 -8 32 272
use FILL  FILL93150x7950
timestamp 1701859473
transform -1 0 6230 0 -1 790
box -12 -8 32 272
use FILL  FILL93150x11850
timestamp 1701859473
transform 1 0 6210 0 1 790
box -12 -8 32 272
use FILL  FILL93150x15750
timestamp 1701859473
transform -1 0 6230 0 -1 1310
box -12 -8 32 272
use FILL  FILL93150x19650
timestamp 1701859473
transform 1 0 6210 0 1 1310
box -12 -8 32 272
use FILL  FILL93150x23550
timestamp 1701859473
transform -1 0 6230 0 -1 1830
box -12 -8 32 272
use FILL  FILL93150x27450
timestamp 1701859473
transform 1 0 6210 0 1 1830
box -12 -8 32 272
use FILL  FILL93150x31350
timestamp 1701859473
transform -1 0 6230 0 -1 2350
box -12 -8 32 272
use FILL  FILL93150x35250
timestamp 1701859473
transform 1 0 6210 0 1 2350
box -12 -8 32 272
use FILL  FILL93150x39150
timestamp 1701859473
transform -1 0 6230 0 -1 2870
box -12 -8 32 272
use FILL  FILL93150x46950
timestamp 1701859473
transform -1 0 6230 0 -1 3390
box -12 -8 32 272
use FILL  FILL93150x50850
timestamp 1701859473
transform 1 0 6210 0 1 3390
box -12 -8 32 272
use FILL  FILL93150x54750
timestamp 1701859473
transform -1 0 6230 0 -1 3910
box -12 -8 32 272
use FILL  FILL93150x62550
timestamp 1701859473
transform -1 0 6230 0 -1 4430
box -12 -8 32 272
use FILL  FILL93150x70350
timestamp 1701859473
transform -1 0 6230 0 -1 4950
box -12 -8 32 272
use FILL  FILL93150x74250
timestamp 1701859473
transform 1 0 6210 0 1 4950
box -12 -8 32 272
use FILL  FILL93150x78150
timestamp 1701859473
transform -1 0 6230 0 -1 5470
box -12 -8 32 272
use FILL  FILL93150x82050
timestamp 1701859473
transform 1 0 6210 0 1 5470
box -12 -8 32 272
use FILL  FILL93150x85950
timestamp 1701859473
transform -1 0 6230 0 -1 5990
box -12 -8 32 272
use FILL  FILL93150x89850
timestamp 1701859473
transform 1 0 6210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__889_
timestamp 1701859473
transform -1 0 1090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__890_
timestamp 1701859473
transform 1 0 610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__891_
timestamp 1701859473
transform -1 0 670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__892_
timestamp 1701859473
transform 1 0 770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__893_
timestamp 1701859473
transform 1 0 1310 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__894_
timestamp 1701859473
transform 1 0 1030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__895_
timestamp 1701859473
transform 1 0 1550 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__896_
timestamp 1701859473
transform -1 0 1690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__897_
timestamp 1701859473
transform -1 0 930 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__898_
timestamp 1701859473
transform -1 0 1430 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__899_
timestamp 1701859473
transform -1 0 950 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__900_
timestamp 1701859473
transform -1 0 350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__901_
timestamp 1701859473
transform -1 0 490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__902_
timestamp 1701859473
transform 1 0 150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__903_
timestamp 1701859473
transform -1 0 550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__904_
timestamp 1701859473
transform -1 0 630 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__905_
timestamp 1701859473
transform -1 0 590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__906_
timestamp 1701859473
transform -1 0 910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__907_
timestamp 1701859473
transform -1 0 890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__908_
timestamp 1701859473
transform -1 0 430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__909_
timestamp 1701859473
transform -1 0 790 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__910_
timestamp 1701859473
transform 1 0 670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__911_
timestamp 1701859473
transform 1 0 390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__912_
timestamp 1701859473
transform -1 0 290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__913_
timestamp 1701859473
transform 1 0 170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__914_
timestamp 1701859473
transform 1 0 270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__915_
timestamp 1701859473
transform 1 0 1370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__916_
timestamp 1701859473
transform -1 0 530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__917_
timestamp 1701859473
transform 1 0 610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__918_
timestamp 1701859473
transform -1 0 1030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__919_
timestamp 1701859473
transform 1 0 750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__920_
timestamp 1701859473
transform -1 0 1370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__921_
timestamp 1701859473
transform -1 0 1190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1701859473
transform 1 0 810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1701859473
transform -1 0 1110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1701859473
transform 1 0 950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1701859473
transform 1 0 10 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1701859473
transform 1 0 3150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1701859473
transform -1 0 3050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1701859473
transform 1 0 3170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1701859473
transform -1 0 3710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1701859473
transform -1 0 3870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1701859473
transform 1 0 3710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1701859473
transform 1 0 2130 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1701859473
transform 1 0 1990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1701859473
transform -1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1701859473
transform 1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1701859473
transform -1 0 3570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1701859473
transform -1 0 3430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1701859473
transform 1 0 2910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1701859473
transform 1 0 2670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1701859473
transform -1 0 2810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1701859473
transform 1 0 2410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1701859473
transform -1 0 2570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1701859473
transform 1 0 2690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1701859473
transform 1 0 1390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1701859473
transform -1 0 1590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1701859473
transform -1 0 1710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1701859473
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1701859473
transform -1 0 1690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1701859473
transform -1 0 1830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1701859473
transform -1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1701859473
transform 1 0 4270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1701859473
transform 1 0 2650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1701859473
transform 1 0 4170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1701859473
transform 1 0 4070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1701859473
transform 1 0 4310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1701859473
transform 1 0 4970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1701859473
transform 1 0 4610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1701859473
transform 1 0 4870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1701859473
transform -1 0 5170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1701859473
transform -1 0 4750 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1701859473
transform -1 0 5030 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1701859473
transform -1 0 5270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1701859473
transform 1 0 6010 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1701859473
transform 1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1701859473
transform 1 0 5190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1701859473
transform -1 0 5990 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1701859473
transform 1 0 4830 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1701859473
transform 1 0 3270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1701859473
transform 1 0 5370 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1701859473
transform -1 0 5910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1701859473
transform -1 0 6010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1701859473
transform -1 0 5970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1701859473
transform -1 0 5730 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1701859473
transform 1 0 5430 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1701859473
transform 1 0 4710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1701859473
transform -1 0 4390 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1701859473
transform 1 0 3030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1701859473
transform -1 0 4390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1701859473
transform 1 0 4510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1701859473
transform 1 0 4750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1701859473
transform 1 0 5570 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1701859473
transform 1 0 5670 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1701859473
transform 1 0 5830 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1701859473
transform 1 0 4890 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1701859473
transform 1 0 4890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1701859473
transform 1 0 5310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1701859473
transform -1 0 5890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1701859473
transform -1 0 5250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1701859473
transform 1 0 5490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1701859473
transform 1 0 5950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1701859473
transform -1 0 5050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1701859473
transform -1 0 5070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1701859473
transform 1 0 5590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1701859473
transform -1 0 6010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1701859473
transform 1 0 6030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1701859473
transform 1 0 5330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1701859473
transform -1 0 5810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1701859473
transform 1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1701859473
transform 1 0 3990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1701859473
transform -1 0 4150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1701859473
transform 1 0 3790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1701859473
transform -1 0 4230 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1701859473
transform 1 0 4650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1701859473
transform 1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1701859473
transform -1 0 4510 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1701859473
transform -1 0 4390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1701859473
transform 1 0 3690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1701859473
transform 1 0 3950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1701859473
transform 1 0 4230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1701859473
transform -1 0 5810 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1701859473
transform -1 0 5690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1701859473
transform 1 0 5370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1701859473
transform -1 0 5870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1701859473
transform 1 0 6090 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1701859473
transform -1 0 5830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1701859473
transform 1 0 5510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1701859473
transform -1 0 5390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1701859473
transform 1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1701859473
transform 1 0 5930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1701859473
transform 1 0 5970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1701859473
transform 1 0 3630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1701859473
transform -1 0 4790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1701859473
transform -1 0 4670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1701859473
transform -1 0 2090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1701859473
transform -1 0 4530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1701859473
transform 1 0 4630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1701859473
transform 1 0 5350 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1701859473
transform 1 0 5350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1701859473
transform 1 0 5030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1701859473
transform -1 0 4930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1701859473
transform -1 0 4350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1701859473
transform 1 0 5610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1701859473
transform 1 0 5770 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1701859473
transform -1 0 5750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1701859473
transform -1 0 5470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1701859473
transform 1 0 5750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1701859473
transform 1 0 6050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1701859473
transform -1 0 3750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1701859473
transform -1 0 3870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1701859473
transform 1 0 3910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1701859473
transform 1 0 4450 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1701859473
transform 1 0 4210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1701859473
transform 1 0 4230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1701859473
transform 1 0 4250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1701859473
transform 1 0 4290 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1701859473
transform 1 0 4150 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1701859473
transform 1 0 4050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1701859473
transform 1 0 4610 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1701859473
transform 1 0 4750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1701859473
transform 1 0 5190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1701859473
transform 1 0 6070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1701859473
transform -1 0 5910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1701859473
transform 1 0 5630 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1701859473
transform -1 0 5070 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1701859473
transform 1 0 5630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1701859473
transform -1 0 6090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1701859473
transform 1 0 5950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1701859473
transform 1 0 5770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1701859473
transform -1 0 5950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1701859473
transform -1 0 6070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1701859473
transform 1 0 1310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1701859473
transform 1 0 4110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1701859473
transform 1 0 4750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1701859473
transform 1 0 5270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1701859473
transform 1 0 5830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1701859473
transform -1 0 5630 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1701859473
transform -1 0 5930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1701859473
transform -1 0 5950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1701859473
transform -1 0 5490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1701859473
transform -1 0 5250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1701859473
transform 1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1701859473
transform 1 0 5410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1701859473
transform 1 0 5470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1701859473
transform 1 0 6090 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1701859473
transform 1 0 5630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1701859473
transform 1 0 4650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1701859473
transform -1 0 4490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1701859473
transform -1 0 5050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1701859473
transform -1 0 3990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1701859473
transform -1 0 4950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1701859473
transform 1 0 5130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1701859473
transform -1 0 4370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1701859473
transform -1 0 4810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1701859473
transform -1 0 5210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1701859473
transform 1 0 5950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1701859473
transform 1 0 5330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1701859473
transform 1 0 5030 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1701859473
transform -1 0 5490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1701859473
transform -1 0 4030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1701859473
transform 1 0 4310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1701859473
transform 1 0 3570 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1701859473
transform 1 0 3790 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1701859473
transform -1 0 4250 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1701859473
transform 1 0 3790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1701859473
transform 1 0 4250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1701859473
transform 1 0 4350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1701859473
transform 1 0 4090 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1701859473
transform 1 0 3930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1701859473
transform 1 0 4110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1701859473
transform 1 0 5410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1701859473
transform -1 0 5910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1701859473
transform 1 0 5190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1701859473
transform 1 0 5490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1701859473
transform -1 0 5810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1701859473
transform 1 0 5290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1701859473
transform 1 0 5730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1701859473
transform 1 0 5950 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1701859473
transform 1 0 5930 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1701859473
transform 1 0 5670 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1701859473
transform -1 0 6050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1701859473
transform 1 0 5990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1701859473
transform -1 0 3670 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1701859473
transform 1 0 4550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1701859473
transform 1 0 3970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1701859473
transform -1 0 3930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1701859473
transform 1 0 3770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1701859473
transform 1 0 3630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1701859473
transform 1 0 4130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1701859473
transform -1 0 4410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1701859473
transform -1 0 4030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1701859473
transform -1 0 4170 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1701859473
transform 1 0 4250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1701859473
transform 1 0 4330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1701859473
transform 1 0 5970 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1701859473
transform -1 0 5890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1701859473
transform -1 0 5830 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1701859473
transform 1 0 4850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1701859473
transform 1 0 4550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1701859473
transform 1 0 5130 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1701859473
transform -1 0 5750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1701859473
transform -1 0 5690 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1701859473
transform -1 0 5790 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1701859473
transform -1 0 5590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1701859473
transform 1 0 6030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1701859473
transform -1 0 5730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1701859473
transform -1 0 5430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1701859473
transform -1 0 5570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1701859473
transform -1 0 5850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1701859473
transform 1 0 5130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1701859473
transform -1 0 5230 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1701859473
transform -1 0 5130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1701859473
transform 1 0 4950 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1701859473
transform -1 0 4910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1701859473
transform -1 0 5330 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1701859473
transform 1 0 4750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1701859473
transform 1 0 5290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1701859473
transform 1 0 5870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1701859473
transform -1 0 5750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1701859473
transform -1 0 5470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1701859473
transform 1 0 4910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1701859473
transform 1 0 5590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1701859473
transform 1 0 5830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1701859473
transform -1 0 5570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1701859473
transform -1 0 5710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1701859473
transform -1 0 5430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1701859473
transform 1 0 5070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1701859473
transform 1 0 5530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1701859473
transform -1 0 5690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1701859473
transform -1 0 5650 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1701859473
transform -1 0 4990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1701859473
transform -1 0 5290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1701859473
transform -1 0 4850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1701859473
transform -1 0 5690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1701859473
transform -1 0 5190 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1701859473
transform -1 0 4050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1701859473
transform 1 0 4150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1701859473
transform -1 0 4310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1701859473
transform 1 0 4710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1701859473
transform 1 0 4430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1701859473
transform 1 0 5010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1701859473
transform 1 0 5090 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1701859473
transform -1 0 4970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1701859473
transform 1 0 5250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1701859473
transform 1 0 5530 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1701859473
transform 1 0 5510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1701859473
transform -1 0 4830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1701859473
transform 1 0 5230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1701859473
transform -1 0 4830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1701859473
transform -1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1701859473
transform -1 0 5350 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1701859473
transform -1 0 4970 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1701859473
transform -1 0 4890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1701859473
transform -1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1701859473
transform -1 0 4230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1701859473
transform 1 0 4070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1701859473
transform -1 0 3810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1701859473
transform 1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1701859473
transform -1 0 3270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1701859473
transform 1 0 3770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1701859473
transform -1 0 3890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1701859473
transform 1 0 3810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1701859473
transform 1 0 3950 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1701859473
transform 1 0 5410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1701859473
transform -1 0 5110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1701859473
transform 1 0 4430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1701859473
transform -1 0 5090 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1701859473
transform -1 0 4610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1701859473
transform -1 0 5230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1701859473
transform 1 0 5070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1701859473
transform -1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1701859473
transform 1 0 4590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1701859473
transform 1 0 4650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1701859473
transform -1 0 5210 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1701859473
transform -1 0 4810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1701859473
transform -1 0 4710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1701859473
transform -1 0 5530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1701859473
transform 1 0 5010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1701859473
transform 1 0 6010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1701859473
transform 1 0 4050 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1701859473
transform 1 0 5030 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1701859473
transform -1 0 4450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1701859473
transform -1 0 4430 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1701859473
transform 1 0 4750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1701859473
transform 1 0 4890 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1701859473
transform 1 0 5030 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1701859473
transform 1 0 4750 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1701859473
transform 1 0 4610 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1701859473
transform 1 0 4890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1701859473
transform -1 0 5210 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1701859473
transform -1 0 5550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1701859473
transform -1 0 3470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1701859473
transform 1 0 3130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1701859473
transform 1 0 3070 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1701859473
transform -1 0 3370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1701859473
transform -1 0 3510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1701859473
transform -1 0 3510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1701859473
transform -1 0 3410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1701859473
transform 1 0 3230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1701859473
transform -1 0 3650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1701859473
transform -1 0 3530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1701859473
transform -1 0 3270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1701859473
transform -1 0 4150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1701859473
transform -1 0 4910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1701859473
transform -1 0 4530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1701859473
transform -1 0 4690 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1701859473
transform 1 0 4990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1701859473
transform 1 0 4750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1701859473
transform -1 0 4490 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1701859473
transform -1 0 4670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1701859473
transform 1 0 4930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1701859473
transform 1 0 3990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1701859473
transform 1 0 4850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1701859473
transform -1 0 4550 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1701859473
transform -1 0 4250 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1701859473
transform 1 0 5370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1701859473
transform 1 0 5570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1701859473
transform 1 0 4270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1701859473
transform -1 0 4790 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1701859473
transform 1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1701859473
transform 1 0 5610 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1701859473
transform 1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1701859473
transform -1 0 5250 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1701859473
transform 1 0 5290 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1701859473
transform 1 0 5650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1701859473
transform 1 0 5790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1701859473
transform -1 0 5890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1701859473
transform 1 0 5470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1701859473
transform 1 0 5470 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1701859473
transform 1 0 5770 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1701859473
transform 1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1701859473
transform 1 0 5290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1701859473
transform -1 0 5830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1701859473
transform 1 0 5930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1701859473
transform -1 0 5530 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1701859473
transform 1 0 5410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1701859473
transform -1 0 5290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1701859473
transform -1 0 5670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1701859473
transform 1 0 5050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1701859473
transform -1 0 5150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1701859473
transform -1 0 3370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1701859473
transform 1 0 2470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1701859473
transform 1 0 1070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1701859473
transform 1 0 1510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1701859473
transform -1 0 2410 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1701859473
transform -1 0 2550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1701859473
transform -1 0 2130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1701859473
transform 1 0 2250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1701859473
transform 1 0 730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1701859473
transform 1 0 590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1701859473
transform 1 0 1050 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1701859473
transform -1 0 1610 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1701859473
transform 1 0 1150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1701859473
transform 1 0 1690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1701859473
transform 1 0 5370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1701859473
transform -1 0 5230 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1701859473
transform -1 0 5410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1701859473
transform -1 0 5510 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1701859473
transform -1 0 5090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1701859473
transform 1 0 4930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1701859473
transform 1 0 4770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1701859473
transform 1 0 4970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1701859473
transform -1 0 3790 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1701859473
transform -1 0 3530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1701859473
transform 1 0 4790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1701859473
transform -1 0 4930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1701859473
transform 1 0 4590 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1701859473
transform 1 0 4190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1701859473
transform 1 0 5090 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1701859473
transform 1 0 5130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1701859473
transform 1 0 3650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1701859473
transform -1 0 3930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1701859473
transform -1 0 3770 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1701859473
transform -1 0 3890 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1701859473
transform -1 0 3610 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1701859473
transform 1 0 3630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1701859473
transform 1 0 3510 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1701859473
transform 1 0 4390 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1701859473
transform -1 0 4110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1701859473
transform -1 0 3370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1701859473
transform 1 0 2590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1701859473
transform 1 0 2850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1701859473
transform 1 0 2350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1701859473
transform 1 0 2650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1701859473
transform 1 0 2810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1701859473
transform -1 0 2370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1701859473
transform 1 0 2530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1701859473
transform 1 0 3110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1701859473
transform 1 0 2250 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1701859473
transform 1 0 2490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1701859473
transform -1 0 2950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1701859473
transform 1 0 2770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1701859473
transform 1 0 3270 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1701859473
transform 1 0 2630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1701859473
transform -1 0 3090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1701859473
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1701859473
transform -1 0 2930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1701859473
transform 1 0 3830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1701859473
transform -1 0 4050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1701859473
transform -1 0 4750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1701859473
transform -1 0 4590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1701859473
transform -1 0 3710 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1701859473
transform 1 0 3750 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1701859473
transform 1 0 3190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1701859473
transform -1 0 3850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1701859473
transform 1 0 3910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1701859473
transform 1 0 3730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1701859473
transform 1 0 4030 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1701859473
transform 1 0 5450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1701859473
transform 1 0 5690 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1701859473
transform 1 0 3570 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1701859473
transform 1 0 3950 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1701859473
transform -1 0 4350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1701859473
transform 1 0 4170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1701859473
transform -1 0 4330 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1701859473
transform 1 0 4290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1701859473
transform 1 0 4170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1701859473
transform 1 0 4450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1701859473
transform 1 0 4450 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1701859473
transform -1 0 4490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1701859473
transform -1 0 5970 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1701859473
transform 1 0 5830 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1701859473
transform -1 0 4070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1701859473
transform -1 0 3910 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1701859473
transform -1 0 3610 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1701859473
transform 1 0 3450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1701859473
transform -1 0 2850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1701859473
transform -1 0 2690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1701859473
transform -1 0 2130 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1701859473
transform -1 0 2890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1701859473
transform 1 0 1870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1701859473
transform -1 0 2730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1701859473
transform -1 0 2010 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1701859473
transform -1 0 1230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1701859473
transform 1 0 1170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1701859473
transform -1 0 490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1701859473
transform -1 0 3450 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1701859473
transform -1 0 4650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1701859473
transform -1 0 3330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1701859473
transform -1 0 2730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1701859473
transform -1 0 3050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1701859473
transform 1 0 2350 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1701859473
transform -1 0 3510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1701859473
transform 1 0 3370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1701859473
transform -1 0 3330 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1701859473
transform -1 0 3450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1701859473
transform -1 0 2990 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1701859473
transform -1 0 3010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1701859473
transform -1 0 3130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1701859473
transform 1 0 2710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1701859473
transform 1 0 3210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1701859473
transform -1 0 3090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1701859473
transform -1 0 2930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1701859473
transform -1 0 2990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1701859473
transform 1 0 3250 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1701859473
transform 1 0 2850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1701859473
transform 1 0 2570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1701859473
transform -1 0 4210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1701859473
transform 1 0 2470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1701859473
transform 1 0 2030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1701859473
transform 1 0 1910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1701859473
transform 1 0 2170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1701859473
transform -1 0 2390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1701859473
transform 1 0 2210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1701859473
transform 1 0 2290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1701859473
transform -1 0 3050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1701859473
transform -1 0 2910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1701859473
transform -1 0 2770 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1701859473
transform 1 0 2610 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1701859473
transform -1 0 2590 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1701859473
transform 1 0 3190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1701859473
transform -1 0 2350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1701859473
transform -1 0 2470 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1701859473
transform -1 0 2290 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1701859473
transform 1 0 2730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1701859473
transform -1 0 3610 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1701859473
transform -1 0 2750 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1701859473
transform -1 0 2890 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1701859473
transform 1 0 2450 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1701859473
transform -1 0 2730 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1701859473
transform -1 0 2890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1701859473
transform 1 0 2870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1701859473
transform -1 0 2590 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1701859473
transform 1 0 3010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1701859473
transform -1 0 3170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1701859473
transform -1 0 3170 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1701859473
transform -1 0 3290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1701859473
transform -1 0 3910 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1701859473
transform -1 0 3750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1701859473
transform -1 0 3030 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1701859473
transform 1 0 1970 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1701859473
transform -1 0 2590 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1701859473
transform -1 0 2790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1701859473
transform -1 0 2650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1701859473
transform -1 0 2530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1701859473
transform -1 0 2470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1701859473
transform -1 0 2310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1701859473
transform 1 0 330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1701859473
transform 1 0 730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1701859473
transform -1 0 3690 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1701859473
transform -1 0 3410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1701859473
transform 1 0 1010 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1701859473
transform -1 0 990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1701859473
transform -1 0 1130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1701859473
transform 1 0 130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1701859473
transform -1 0 490 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1701859473
transform -1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1701859473
transform 1 0 1830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1701859473
transform 1 0 2230 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1701859473
transform 1 0 3090 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1701859473
transform -1 0 1790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1701859473
transform -1 0 2130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1701859473
transform -1 0 1930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1701859473
transform -1 0 1650 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1701859473
transform -1 0 1530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1701859473
transform 1 0 2030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1701859473
transform 1 0 1770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1701859473
transform 1 0 1630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1701859473
transform 1 0 1370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1701859473
transform -1 0 1490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1701859473
transform -1 0 1730 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1701859473
transform 1 0 1550 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1452_
timestamp 1701859473
transform -1 0 2010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1453_
timestamp 1701859473
transform 1 0 1290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1454_
timestamp 1701859473
transform -1 0 1790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1455_
timestamp 1701859473
transform 1 0 1650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1456_
timestamp 1701859473
transform 1 0 1770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1457_
timestamp 1701859473
transform -1 0 1870 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1458_
timestamp 1701859473
transform 1 0 1370 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1459_
timestamp 1701859473
transform -1 0 1250 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1460_
timestamp 1701859473
transform -1 0 1230 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1461_
timestamp 1701859473
transform 1 0 1330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1462_
timestamp 1701859473
transform -1 0 2470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1463_
timestamp 1701859473
transform -1 0 1130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1464_
timestamp 1701859473
transform 1 0 1470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1465_
timestamp 1701859473
transform 1 0 1630 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1466_
timestamp 1701859473
transform 1 0 1070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1467_
timestamp 1701859473
transform 1 0 1530 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1468_
timestamp 1701859473
transform -1 0 1690 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1469_
timestamp 1701859473
transform 1 0 1870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1470_
timestamp 1701859473
transform -1 0 2150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1471_
timestamp 1701859473
transform -1 0 2450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1472_
timestamp 1701859473
transform -1 0 2310 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1473_
timestamp 1701859473
transform 1 0 1990 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1474_
timestamp 1701859473
transform -1 0 2110 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1475_
timestamp 1701859473
transform -1 0 2150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1476_
timestamp 1701859473
transform -1 0 2370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1477_
timestamp 1701859473
transform 1 0 1890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1478_
timestamp 1701859473
transform 1 0 1990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1479_
timestamp 1701859473
transform -1 0 2010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1480_
timestamp 1701859473
transform 1 0 4310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1481_
timestamp 1701859473
transform 1 0 4070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1482_
timestamp 1701859473
transform -1 0 4230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1483_
timestamp 1701859473
transform -1 0 1290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1484_
timestamp 1701859473
transform 1 0 1130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1485_
timestamp 1701859473
transform -1 0 870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1486_
timestamp 1701859473
transform 1 0 750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1487_
timestamp 1701859473
transform -1 0 290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1488_
timestamp 1701859473
transform -1 0 1250 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1489_
timestamp 1701859473
transform -1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1490_
timestamp 1701859473
transform 1 0 1550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1491_
timestamp 1701859473
transform 1 0 2150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1492_
timestamp 1701859473
transform -1 0 2030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1493_
timestamp 1701859473
transform 1 0 1850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1494_
timestamp 1701859473
transform -1 0 1730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1495_
timestamp 1701859473
transform 1 0 1310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1496_
timestamp 1701859473
transform 1 0 1570 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1497_
timestamp 1701859473
transform 1 0 1490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1498_
timestamp 1701859473
transform -1 0 1650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1499_
timestamp 1701859473
transform -1 0 1450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1500_
timestamp 1701859473
transform 1 0 1430 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1501_
timestamp 1701859473
transform 1 0 1570 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1502_
timestamp 1701859473
transform -1 0 430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1503_
timestamp 1701859473
transform 1 0 650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1504_
timestamp 1701859473
transform -1 0 410 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1505_
timestamp 1701859473
transform -1 0 290 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1506_
timestamp 1701859473
transform -1 0 930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1507_
timestamp 1701859473
transform -1 0 790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1508_
timestamp 1701859473
transform -1 0 710 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1509_
timestamp 1701859473
transform -1 0 850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1510_
timestamp 1701859473
transform 1 0 970 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1511_
timestamp 1701859473
transform -1 0 570 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1512_
timestamp 1701859473
transform 1 0 710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1513_
timestamp 1701859473
transform -1 0 3410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1514_
timestamp 1701859473
transform 1 0 2050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1515_
timestamp 1701859473
transform -1 0 2170 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1516_
timestamp 1701859473
transform -1 0 1850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1517_
timestamp 1701859473
transform 1 0 1750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1518_
timestamp 1701859473
transform -1 0 750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1519_
timestamp 1701859473
transform 1 0 1810 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1520_
timestamp 1701859473
transform -1 0 1950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1521_
timestamp 1701859473
transform 1 0 1910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1522_
timestamp 1701859473
transform -1 0 2210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1523_
timestamp 1701859473
transform 1 0 1010 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1524_
timestamp 1701859473
transform -1 0 310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1525_
timestamp 1701859473
transform 1 0 10 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1526_
timestamp 1701859473
transform 1 0 270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1527_
timestamp 1701859473
transform -1 0 4490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1528_
timestamp 1701859473
transform -1 0 4590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1529_
timestamp 1701859473
transform 1 0 4330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1530_
timestamp 1701859473
transform 1 0 730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1531_
timestamp 1701859473
transform -1 0 870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1532_
timestamp 1701859473
transform -1 0 930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1533_
timestamp 1701859473
transform 1 0 270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1534_
timestamp 1701859473
transform 1 0 290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1535_
timestamp 1701859473
transform -1 0 1350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1536_
timestamp 1701859473
transform -1 0 1450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1537_
timestamp 1701859473
transform -1 0 330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1538_
timestamp 1701859473
transform -1 0 150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1539_
timestamp 1701859473
transform -1 0 1710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1540_
timestamp 1701859473
transform 1 0 1190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1541_
timestamp 1701859473
transform -1 0 1050 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1542_
timestamp 1701859473
transform -1 0 1350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1543_
timestamp 1701859473
transform -1 0 1070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1544_
timestamp 1701859473
transform -1 0 1410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1545_
timestamp 1701859473
transform -1 0 1050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1546_
timestamp 1701859473
transform 1 0 130 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1547_
timestamp 1701859473
transform 1 0 430 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1548_
timestamp 1701859473
transform -1 0 570 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1549_
timestamp 1701859473
transform 1 0 430 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1550_
timestamp 1701859473
transform 1 0 570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1551_
timestamp 1701859473
transform -1 0 4470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1552_
timestamp 1701859473
transform -1 0 4650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1553_
timestamp 1701859473
transform 1 0 630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1554_
timestamp 1701859473
transform -1 0 1270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1555_
timestamp 1701859473
transform -1 0 1190 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1556_
timestamp 1701859473
transform 1 0 850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1557_
timestamp 1701859473
transform 1 0 10 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1558_
timestamp 1701859473
transform 1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1559_
timestamp 1701859473
transform 1 0 1170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1560_
timestamp 1701859473
transform -1 0 1290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1561_
timestamp 1701859473
transform -1 0 190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1562_
timestamp 1701859473
transform 1 0 10 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1563_
timestamp 1701859473
transform -1 0 310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1564_
timestamp 1701859473
transform -1 0 1130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1565_
timestamp 1701859473
transform -1 0 1250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1566_
timestamp 1701859473
transform -1 0 1370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1567_
timestamp 1701859473
transform -1 0 1210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1568_
timestamp 1701859473
transform -1 0 1210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1569_
timestamp 1701859473
transform -1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1570_
timestamp 1701859473
transform -1 0 910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1571_
timestamp 1701859473
transform -1 0 710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1572_
timestamp 1701859473
transform 1 0 550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1573_
timestamp 1701859473
transform -1 0 410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1574_
timestamp 1701859473
transform -1 0 5110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1575_
timestamp 1701859473
transform 1 0 4950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1576_
timestamp 1701859473
transform -1 0 4830 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1577_
timestamp 1701859473
transform -1 0 4670 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1578_
timestamp 1701859473
transform 1 0 10 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1579_
timestamp 1701859473
transform 1 0 10 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1580_
timestamp 1701859473
transform -1 0 210 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1581_
timestamp 1701859473
transform 1 0 110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1582_
timestamp 1701859473
transform 1 0 10 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1583_
timestamp 1701859473
transform -1 0 830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1584_
timestamp 1701859473
transform -1 0 930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1585_
timestamp 1701859473
transform -1 0 630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1586_
timestamp 1701859473
transform -1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1587_
timestamp 1701859473
transform -1 0 4850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1588_
timestamp 1701859473
transform -1 0 4670 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1589_
timestamp 1701859473
transform -1 0 1470 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1590_
timestamp 1701859473
transform -1 0 1170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1591_
timestamp 1701859473
transform -1 0 1030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1592_
timestamp 1701859473
transform 1 0 110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1593_
timestamp 1701859473
transform 1 0 2510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1594_
timestamp 1701859473
transform -1 0 2650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1595_
timestamp 1701859473
transform 1 0 3590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1596_
timestamp 1701859473
transform 1 0 3430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1597_
timestamp 1701859473
transform -1 0 2450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1598_
timestamp 1701859473
transform 1 0 2270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1599_
timestamp 1701859473
transform -1 0 3710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1600_
timestamp 1701859473
transform 1 0 3530 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1601_
timestamp 1701859473
transform 1 0 3230 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1602_
timestamp 1701859473
transform 1 0 2810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1603_
timestamp 1701859473
transform -1 0 2850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1604_
timestamp 1701859473
transform 1 0 2670 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1605_
timestamp 1701859473
transform 1 0 2010 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1606_
timestamp 1701859473
transform 1 0 1850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1607_
timestamp 1701859473
transform -1 0 1690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1608_
timestamp 1701859473
transform 1 0 1510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1636_
timestamp 1701859473
transform -1 0 4210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1637_
timestamp 1701859473
transform -1 0 4310 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1638_
timestamp 1701859473
transform -1 0 4070 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1639_
timestamp 1701859473
transform 1 0 3910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1640_
timestamp 1701859473
transform -1 0 3670 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1641_
timestamp 1701859473
transform -1 0 3610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1642_
timestamp 1701859473
transform -1 0 3170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1643_
timestamp 1701859473
transform -1 0 4070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1644_
timestamp 1701859473
transform -1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1645_
timestamp 1701859473
transform 1 0 4450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1646_
timestamp 1701859473
transform -1 0 4190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1647_
timestamp 1701859473
transform 1 0 3270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1648_
timestamp 1701859473
transform -1 0 4190 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1649_
timestamp 1701859473
transform -1 0 3790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1650_
timestamp 1701859473
transform -1 0 3910 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1651_
timestamp 1701859473
transform 1 0 3630 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1652_
timestamp 1701859473
transform 1 0 3630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1653_
timestamp 1701859473
transform 1 0 3750 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1654_
timestamp 1701859473
transform -1 0 4590 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1655_
timestamp 1701859473
transform -1 0 4450 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1656_
timestamp 1701859473
transform 1 0 1430 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1657_
timestamp 1701859473
transform 1 0 3070 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1658_
timestamp 1701859473
transform 1 0 3210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1659_
timestamp 1701859473
transform -1 0 3170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1660_
timestamp 1701859473
transform 1 0 3510 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1661_
timestamp 1701859473
transform -1 0 3390 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1662_
timestamp 1701859473
transform 1 0 3510 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1663_
timestamp 1701859473
transform -1 0 3470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1664_
timestamp 1701859473
transform -1 0 3310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1665_
timestamp 1701859473
transform -1 0 3950 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1666_
timestamp 1701859473
transform 1 0 3810 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1667_
timestamp 1701859473
transform -1 0 3670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1668_
timestamp 1701859473
transform 1 0 3370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1669_
timestamp 1701859473
transform -1 0 3490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1670_
timestamp 1701859473
transform -1 0 3350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1671_
timestamp 1701859473
transform -1 0 3050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1672_
timestamp 1701859473
transform 1 0 2710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1673_
timestamp 1701859473
transform -1 0 2870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1674_
timestamp 1701859473
transform 1 0 2950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1675_
timestamp 1701859473
transform -1 0 4370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1676_
timestamp 1701859473
transform 1 0 4090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1677_
timestamp 1701859473
transform 1 0 3770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1678_
timestamp 1701859473
transform 1 0 4290 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1679_
timestamp 1701859473
transform 1 0 4570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1680_
timestamp 1701859473
transform -1 0 4470 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1681_
timestamp 1701859473
transform 1 0 3870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1682_
timestamp 1701859473
transform 1 0 4050 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1683_
timestamp 1701859473
transform 1 0 3930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1684_
timestamp 1701859473
transform 1 0 3750 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1685_
timestamp 1701859473
transform -1 0 2810 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1686_
timestamp 1701859473
transform -1 0 2530 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1687_
timestamp 1701859473
transform 1 0 2390 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1688_
timestamp 1701859473
transform -1 0 2130 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1689_
timestamp 1701859473
transform -1 0 1630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1690_
timestamp 1701859473
transform 1 0 2650 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1691_
timestamp 1701859473
transform -1 0 2270 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1692_
timestamp 1701859473
transform -1 0 2970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1693_
timestamp 1701859473
transform 1 0 3130 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1694_
timestamp 1701859473
transform 1 0 3130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1695_
timestamp 1701859473
transform -1 0 3550 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1696_
timestamp 1701859473
transform 1 0 3390 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1697_
timestamp 1701859473
transform -1 0 3270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1698_
timestamp 1701859473
transform -1 0 3110 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1699_
timestamp 1701859473
transform -1 0 2410 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1700_
timestamp 1701859473
transform 1 0 2230 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1701_
timestamp 1701859473
transform -1 0 2190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1702_
timestamp 1701859473
transform 1 0 2010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1703_
timestamp 1701859473
transform 1 0 1250 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1704_
timestamp 1701859473
transform -1 0 1210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1705_
timestamp 1701859473
transform 1 0 2310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1706_
timestamp 1701859473
transform -1 0 2430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1707_
timestamp 1701859473
transform 1 0 1870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1708_
timestamp 1701859473
transform -1 0 1850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1709_
timestamp 1701859473
transform -1 0 2610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1710_
timestamp 1701859473
transform -1 0 3010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1711_
timestamp 1701859473
transform 1 0 2850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1712_
timestamp 1701859473
transform 1 0 2390 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1713_
timestamp 1701859473
transform -1 0 2710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1714_
timestamp 1701859473
transform -1 0 2570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1715_
timestamp 1701859473
transform 1 0 2670 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1716_
timestamp 1701859473
transform 1 0 2530 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1717_
timestamp 1701859473
transform -1 0 2570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1718_
timestamp 1701859473
transform -1 0 2430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1719_
timestamp 1701859473
transform 1 0 2030 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1720_
timestamp 1701859473
transform 1 0 1850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1721_
timestamp 1701859473
transform 1 0 1570 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1722_
timestamp 1701859473
transform -1 0 1990 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1723_
timestamp 1701859473
transform 1 0 1710 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1724_
timestamp 1701859473
transform 1 0 1170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1725_
timestamp 1701859473
transform 1 0 1950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1726_
timestamp 1701859473
transform -1 0 870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1727_
timestamp 1701859473
transform -1 0 970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1728_
timestamp 1701859473
transform 1 0 2590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1729_
timestamp 1701859473
transform 1 0 1870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1730_
timestamp 1701859473
transform -1 0 2190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1731_
timestamp 1701859473
transform -1 0 2230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1732_
timestamp 1701859473
transform 1 0 2030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1733_
timestamp 1701859473
transform 1 0 2070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1734_
timestamp 1701859473
transform -1 0 1730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1735_
timestamp 1701859473
transform -1 0 1790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1736_
timestamp 1701859473
transform 1 0 1610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1737_
timestamp 1701859473
transform -1 0 1490 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1738_
timestamp 1701859473
transform -1 0 1110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1739_
timestamp 1701859473
transform -1 0 910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1740_
timestamp 1701859473
transform -1 0 1230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1741_
timestamp 1701859473
transform -1 0 970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1742_
timestamp 1701859473
transform -1 0 2290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1743_
timestamp 1701859473
transform -1 0 3030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1744_
timestamp 1701859473
transform 1 0 2710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1745_
timestamp 1701859473
transform 1 0 2430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1746_
timestamp 1701859473
transform -1 0 2870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1747_
timestamp 1701859473
transform -1 0 2310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1748_
timestamp 1701859473
transform -1 0 1470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1749_
timestamp 1701859473
transform -1 0 1330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1750_
timestamp 1701859473
transform -1 0 810 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1751_
timestamp 1701859473
transform -1 0 770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1752_
timestamp 1701859473
transform -1 0 390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1753_
timestamp 1701859473
transform 1 0 290 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1754_
timestamp 1701859473
transform -1 0 510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1755_
timestamp 1701859473
transform -1 0 610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1756_
timestamp 1701859473
transform -1 0 1250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1757_
timestamp 1701859473
transform 1 0 1910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1758_
timestamp 1701859473
transform -1 0 2130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1759_
timestamp 1701859473
transform -1 0 2250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1760_
timestamp 1701859473
transform -1 0 1830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1761_
timestamp 1701859473
transform 1 0 1630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1762_
timestamp 1701859473
transform -1 0 1470 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1763_
timestamp 1701859473
transform -1 0 1310 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1764_
timestamp 1701859473
transform -1 0 870 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1765_
timestamp 1701859473
transform -1 0 710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1766_
timestamp 1701859473
transform -1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1767_
timestamp 1701859473
transform 1 0 1110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1768_
timestamp 1701859473
transform 1 0 1330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1769_
timestamp 1701859473
transform -1 0 1490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1770_
timestamp 1701859473
transform -1 0 1350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1771_
timestamp 1701859473
transform -1 0 650 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1772_
timestamp 1701859473
transform -1 0 490 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1773_
timestamp 1701859473
transform 1 0 730 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1774_
timestamp 1701859473
transform 1 0 310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1775_
timestamp 1701859473
transform 1 0 10 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1776_
timestamp 1701859473
transform -1 0 450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1777_
timestamp 1701859473
transform -1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1778_
timestamp 1701859473
transform 1 0 2710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1779_
timestamp 1701859473
transform -1 0 3030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1780_
timestamp 1701859473
transform -1 0 3490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1781_
timestamp 1701859473
transform 1 0 2870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1782_
timestamp 1701859473
transform 1 0 3310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1783_
timestamp 1701859473
transform -1 0 1470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1784_
timestamp 1701859473
transform -1 0 1310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1785_
timestamp 1701859473
transform -1 0 1130 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1786_
timestamp 1701859473
transform -1 0 970 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1787_
timestamp 1701859473
transform -1 0 530 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1788_
timestamp 1701859473
transform 1 0 590 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1789_
timestamp 1701859473
transform -1 0 590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1790_
timestamp 1701859473
transform -1 0 430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1791_
timestamp 1701859473
transform -1 0 310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1792_
timestamp 1701859473
transform -1 0 1730 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1793_
timestamp 1701859473
transform 1 0 1590 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1794_
timestamp 1701859473
transform 1 0 590 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1795_
timestamp 1701859473
transform -1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1796_
timestamp 1701859473
transform 1 0 230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1797_
timestamp 1701859473
transform 1 0 450 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1798_
timestamp 1701859473
transform -1 0 650 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1799_
timestamp 1701859473
transform 1 0 390 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1800_
timestamp 1701859473
transform 1 0 170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1801_
timestamp 1701859473
transform -1 0 190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1802_
timestamp 1701859473
transform -1 0 2850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1803_
timestamp 1701859473
transform 1 0 790 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1804_
timestamp 1701859473
transform -1 0 690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1805_
timestamp 1701859473
transform 1 0 790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1806_
timestamp 1701859473
transform 1 0 990 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1807_
timestamp 1701859473
transform -1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1808_
timestamp 1701859473
transform -1 0 470 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1809_
timestamp 1701859473
transform -1 0 1150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1810_
timestamp 1701859473
transform -1 0 970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1811_
timestamp 1701859473
transform -1 0 150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1812_
timestamp 1701859473
transform -1 0 310 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1813_
timestamp 1701859473
transform -1 0 30 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1814_
timestamp 1701859473
transform -1 0 30 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1815_
timestamp 1701859473
transform -1 0 310 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1816_
timestamp 1701859473
transform 1 0 10 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1817_
timestamp 1701859473
transform -1 0 170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1818_
timestamp 1701859473
transform -1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1819_
timestamp 1701859473
transform -1 0 150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1820_
timestamp 1701859473
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1821_
timestamp 1701859473
transform 1 0 510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1822_
timestamp 1701859473
transform -1 0 290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1823_
timestamp 1701859473
transform -1 0 170 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1824_
timestamp 1701859473
transform 1 0 10 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1825_
timestamp 1701859473
transform 1 0 10 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1826_
timestamp 1701859473
transform 1 0 1050 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1701859473
transform -1 0 2770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1701859473
transform 1 0 3370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1701859473
transform 1 0 3430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1701859473
transform -1 0 2810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1701859473
transform -1 0 4530 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1701859473
transform 1 0 4530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1701859473
transform 1 0 4570 0 1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1701859473
transform 1 0 4710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert13
timestamp 1701859473
transform 1 0 3110 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert14
timestamp 1701859473
transform 1 0 2670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1701859473
transform -1 0 1970 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1701859473
transform -1 0 1830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1701859473
transform 1 0 410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1701859473
transform 1 0 3290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1701859473
transform 1 0 1790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1701859473
transform 1 0 1410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1701859473
transform -1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1701859473
transform -1 0 2730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1701859473
transform 1 0 3490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1701859473
transform 1 0 3810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1701859473
transform -1 0 2990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1701859473
transform 1 0 2950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1701859473
transform 1 0 2530 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1701859473
transform -1 0 1470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1701859473
transform 1 0 2530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1701859473
transform -1 0 2430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1701859473
transform 1 0 2890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1701859473
transform 1 0 1950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1701859473
transform 1 0 3290 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert34
timestamp 1701859473
transform -1 0 3570 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert35
timestamp 1701859473
transform -1 0 3950 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert36
timestamp 1701859473
transform 1 0 3950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert37
timestamp 1701859473
transform -1 0 3790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert38
timestamp 1701859473
transform 1 0 1710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert39
timestamp 1701859473
transform -1 0 4490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert40
timestamp 1701859473
transform -1 0 1610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert41
timestamp 1701859473
transform -1 0 2590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1701859473
transform 1 0 2150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1701859473
transform 1 0 1430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 10 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 1930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1701859473
transform 1 0 10 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__889_
timestamp 1701859473
transform -1 0 1110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__890_
timestamp 1701859473
transform 1 0 630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__891_
timestamp 1701859473
transform -1 0 690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__892_
timestamp 1701859473
transform 1 0 790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__893_
timestamp 1701859473
transform 1 0 1330 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__894_
timestamp 1701859473
transform 1 0 1050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__895_
timestamp 1701859473
transform 1 0 1570 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__896_
timestamp 1701859473
transform -1 0 1710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__897_
timestamp 1701859473
transform -1 0 950 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__898_
timestamp 1701859473
transform -1 0 1450 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__899_
timestamp 1701859473
transform -1 0 970 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__900_
timestamp 1701859473
transform -1 0 370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__901_
timestamp 1701859473
transform -1 0 510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__902_
timestamp 1701859473
transform 1 0 170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__903_
timestamp 1701859473
transform -1 0 570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__904_
timestamp 1701859473
transform -1 0 650 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__905_
timestamp 1701859473
transform -1 0 610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__906_
timestamp 1701859473
transform -1 0 930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__907_
timestamp 1701859473
transform -1 0 910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__908_
timestamp 1701859473
transform -1 0 450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__909_
timestamp 1701859473
transform -1 0 810 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__910_
timestamp 1701859473
transform 1 0 690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__911_
timestamp 1701859473
transform 1 0 410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__912_
timestamp 1701859473
transform -1 0 310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__913_
timestamp 1701859473
transform 1 0 190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__914_
timestamp 1701859473
transform 1 0 290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__915_
timestamp 1701859473
transform 1 0 1390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__916_
timestamp 1701859473
transform -1 0 550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__917_
timestamp 1701859473
transform 1 0 630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__918_
timestamp 1701859473
transform -1 0 1050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__919_
timestamp 1701859473
transform 1 0 770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__920_
timestamp 1701859473
transform -1 0 1390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__921_
timestamp 1701859473
transform -1 0 1210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__922_
timestamp 1701859473
transform 1 0 830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1701859473
transform -1 0 1130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1701859473
transform 1 0 970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__925_
timestamp 1701859473
transform 1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1701859473
transform 1 0 3170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__927_
timestamp 1701859473
transform -1 0 3070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1701859473
transform 1 0 3190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__929_
timestamp 1701859473
transform -1 0 3730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1701859473
transform -1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1701859473
transform 1 0 3730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__932_
timestamp 1701859473
transform 1 0 2150 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1701859473
transform 1 0 2010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__934_
timestamp 1701859473
transform -1 0 2150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1701859473
transform 1 0 4370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__936_
timestamp 1701859473
transform -1 0 3590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1701859473
transform -1 0 3450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1701859473
transform 1 0 2930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__939_
timestamp 1701859473
transform 1 0 2690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1701859473
transform -1 0 2830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__941_
timestamp 1701859473
transform 1 0 2430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1701859473
transform -1 0 2590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__943_
timestamp 1701859473
transform 1 0 2710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1701859473
transform 1 0 1410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__945_
timestamp 1701859473
transform -1 0 1610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1701859473
transform -1 0 1730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1701859473
transform -1 0 1310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__948_
timestamp 1701859473
transform -1 0 1710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1701859473
transform -1 0 1850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__950_
timestamp 1701859473
transform -1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1701859473
transform 1 0 4290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__952_
timestamp 1701859473
transform 1 0 2670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1701859473
transform 1 0 4190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1701859473
transform 1 0 4090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__955_
timestamp 1701859473
transform 1 0 4330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1701859473
transform 1 0 4990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__957_
timestamp 1701859473
transform 1 0 4630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1701859473
transform 1 0 4890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__959_
timestamp 1701859473
transform -1 0 5190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1701859473
transform -1 0 4770 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1701859473
transform -1 0 5050 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__962_
timestamp 1701859473
transform -1 0 5290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1701859473
transform 1 0 6030 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__964_
timestamp 1701859473
transform 1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1701859473
transform 1 0 5210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__966_
timestamp 1701859473
transform -1 0 6010 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1701859473
transform 1 0 4850 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1701859473
transform 1 0 3290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__969_
timestamp 1701859473
transform 1 0 5390 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1701859473
transform -1 0 5930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__971_
timestamp 1701859473
transform -1 0 6030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1701859473
transform -1 0 5990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__973_
timestamp 1701859473
transform -1 0 5750 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1701859473
transform 1 0 5450 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1701859473
transform 1 0 4730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__976_
timestamp 1701859473
transform -1 0 4410 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1701859473
transform 1 0 3050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__978_
timestamp 1701859473
transform -1 0 4410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1701859473
transform 1 0 4530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__980_
timestamp 1701859473
transform 1 0 4770 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1701859473
transform 1 0 5590 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1701859473
transform 1 0 5690 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__983_
timestamp 1701859473
transform 1 0 5850 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1701859473
transform 1 0 4910 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__985_
timestamp 1701859473
transform 1 0 4910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1701859473
transform 1 0 5330 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__987_
timestamp 1701859473
transform -1 0 5910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1701859473
transform -1 0 5270 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__989_
timestamp 1701859473
transform 1 0 5510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1701859473
transform 1 0 5970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1701859473
transform -1 0 5070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__992_
timestamp 1701859473
transform -1 0 5090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1701859473
transform 1 0 5610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__994_
timestamp 1701859473
transform -1 0 6030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1701859473
transform 1 0 6050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__996_
timestamp 1701859473
transform 1 0 5350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1701859473
transform -1 0 5830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1701859473
transform 1 0 5550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__999_
timestamp 1701859473
transform 1 0 4010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1000_
timestamp 1701859473
transform -1 0 4170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1701859473
transform 1 0 3810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1701859473
transform -1 0 4250 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1003_
timestamp 1701859473
transform 1 0 4670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1701859473
transform 1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1005_
timestamp 1701859473
transform -1 0 4530 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1701859473
transform -1 0 4410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1007_
timestamp 1701859473
transform 1 0 3710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1701859473
transform 1 0 3970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1701859473
transform 1 0 4250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1010_
timestamp 1701859473
transform -1 0 5830 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1701859473
transform -1 0 5710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1012_
timestamp 1701859473
transform 1 0 5390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1701859473
transform -1 0 5890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1014_
timestamp 1701859473
transform 1 0 6110 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1701859473
transform -1 0 5850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1016_
timestamp 1701859473
transform 1 0 5530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1701859473
transform -1 0 5410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1701859473
transform 1 0 4910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1019_
timestamp 1701859473
transform 1 0 5950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1701859473
transform 1 0 5990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1021_
timestamp 1701859473
transform 1 0 3650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1701859473
transform -1 0 4810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1023_
timestamp 1701859473
transform -1 0 4690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1701859473
transform -1 0 2110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1701859473
transform -1 0 4550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1026_
timestamp 1701859473
transform 1 0 4650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1701859473
transform 1 0 5370 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1028_
timestamp 1701859473
transform 1 0 5370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1701859473
transform 1 0 5050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1030_
timestamp 1701859473
transform -1 0 4950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1701859473
transform -1 0 4370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1701859473
transform 1 0 5630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1033_
timestamp 1701859473
transform 1 0 5790 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1701859473
transform -1 0 5770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1035_
timestamp 1701859473
transform -1 0 5490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1701859473
transform 1 0 5770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1037_
timestamp 1701859473
transform 1 0 6070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1701859473
transform -1 0 3770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1701859473
transform -1 0 3890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1040_
timestamp 1701859473
transform 1 0 3930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1701859473
transform 1 0 4470 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1042_
timestamp 1701859473
transform 1 0 4230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1701859473
transform 1 0 4250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1044_
timestamp 1701859473
transform 1 0 4270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1701859473
transform 1 0 4310 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1701859473
transform 1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1047_
timestamp 1701859473
transform 1 0 4070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1701859473
transform 1 0 4630 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1049_
timestamp 1701859473
transform 1 0 4770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1701859473
transform 1 0 5210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1051_
timestamp 1701859473
transform 1 0 6090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1701859473
transform -1 0 5930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1701859473
transform 1 0 5650 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1054_
timestamp 1701859473
transform -1 0 5090 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1701859473
transform 1 0 5650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1056_
timestamp 1701859473
transform -1 0 6110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1701859473
transform 1 0 5970 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1058_
timestamp 1701859473
transform 1 0 5790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1701859473
transform -1 0 5970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1060_
timestamp 1701859473
transform -1 0 6090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1701859473
transform 1 0 1330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1701859473
transform 1 0 4130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1063_
timestamp 1701859473
transform 1 0 4770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1701859473
transform 1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1065_
timestamp 1701859473
transform 1 0 5850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1701859473
transform -1 0 5650 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1067_
timestamp 1701859473
transform -1 0 5950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1701859473
transform -1 0 5970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1701859473
transform -1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1070_
timestamp 1701859473
transform -1 0 5270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1701859473
transform 1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1072_
timestamp 1701859473
transform 1 0 5430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1701859473
transform 1 0 5490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1074_
timestamp 1701859473
transform 1 0 6110 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1701859473
transform 1 0 5650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1701859473
transform 1 0 4670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1077_
timestamp 1701859473
transform -1 0 4510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1701859473
transform -1 0 5070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1079_
timestamp 1701859473
transform -1 0 4010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1701859473
transform -1 0 4970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1081_
timestamp 1701859473
transform 1 0 5150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1701859473
transform -1 0 4390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1701859473
transform -1 0 4830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1084_
timestamp 1701859473
transform -1 0 5230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1701859473
transform 1 0 5970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1086_
timestamp 1701859473
transform 1 0 5350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1701859473
transform 1 0 5050 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1088_
timestamp 1701859473
transform -1 0 5510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1701859473
transform -1 0 4050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1701859473
transform 1 0 4330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1091_
timestamp 1701859473
transform 1 0 3590 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1701859473
transform 1 0 3810 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1093_
timestamp 1701859473
transform -1 0 4270 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1701859473
transform 1 0 3810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1095_
timestamp 1701859473
transform 1 0 4270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1701859473
transform 1 0 4370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1701859473
transform 1 0 4110 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1098_
timestamp 1701859473
transform 1 0 3950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1701859473
transform 1 0 4130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1100_
timestamp 1701859473
transform 1 0 5430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1701859473
transform -1 0 5930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1102_
timestamp 1701859473
transform 1 0 5210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1701859473
transform 1 0 5510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1104_
timestamp 1701859473
transform -1 0 5830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1701859473
transform 1 0 5310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1701859473
transform 1 0 5750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1107_
timestamp 1701859473
transform 1 0 5970 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1701859473
transform 1 0 5950 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1109_
timestamp 1701859473
transform 1 0 5690 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1701859473
transform -1 0 6070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1111_
timestamp 1701859473
transform 1 0 6010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1701859473
transform -1 0 3690 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1701859473
transform 1 0 4570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1114_
timestamp 1701859473
transform 1 0 3990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1701859473
transform -1 0 3950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1116_
timestamp 1701859473
transform 1 0 3790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1701859473
transform 1 0 3650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1118_
timestamp 1701859473
transform 1 0 4150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1701859473
transform -1 0 4430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1701859473
transform -1 0 4050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1121_
timestamp 1701859473
transform -1 0 4190 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1701859473
transform 1 0 4270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1123_
timestamp 1701859473
transform 1 0 4350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1701859473
transform 1 0 5990 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1125_
timestamp 1701859473
transform -1 0 5910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1701859473
transform -1 0 5850 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1701859473
transform 1 0 4870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1128_
timestamp 1701859473
transform 1 0 4570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1701859473
transform 1 0 5150 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1130_
timestamp 1701859473
transform -1 0 5770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1701859473
transform -1 0 5710 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1132_
timestamp 1701859473
transform -1 0 5810 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1701859473
transform -1 0 5610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1701859473
transform 1 0 6050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1135_
timestamp 1701859473
transform -1 0 5750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1701859473
transform -1 0 5450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1137_
timestamp 1701859473
transform -1 0 5590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1701859473
transform -1 0 5870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1139_
timestamp 1701859473
transform 1 0 5150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1701859473
transform -1 0 5250 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1701859473
transform -1 0 5150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1142_
timestamp 1701859473
transform 1 0 4970 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1701859473
transform -1 0 4930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1144_
timestamp 1701859473
transform -1 0 5350 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1701859473
transform 1 0 4770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1146_
timestamp 1701859473
transform 1 0 5310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1701859473
transform 1 0 5890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1148_
timestamp 1701859473
transform -1 0 5770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1701859473
transform -1 0 5490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1701859473
transform 1 0 4930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1151_
timestamp 1701859473
transform 1 0 5610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1701859473
transform 1 0 5850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1153_
timestamp 1701859473
transform -1 0 5590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1701859473
transform -1 0 5730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1155_
timestamp 1701859473
transform -1 0 5450 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1701859473
transform 1 0 5090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1701859473
transform 1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1158_
timestamp 1701859473
transform -1 0 5710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1701859473
transform -1 0 5670 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1160_
timestamp 1701859473
transform -1 0 5010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1701859473
transform -1 0 5310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1162_
timestamp 1701859473
transform -1 0 4870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1701859473
transform -1 0 5710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1701859473
transform -1 0 5210 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1165_
timestamp 1701859473
transform -1 0 4070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1701859473
transform 1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1167_
timestamp 1701859473
transform -1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1701859473
transform 1 0 4730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1169_
timestamp 1701859473
transform 1 0 4450 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1701859473
transform 1 0 5030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1701859473
transform 1 0 5110 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1172_
timestamp 1701859473
transform -1 0 4990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1701859473
transform 1 0 5270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1174_
timestamp 1701859473
transform 1 0 5550 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1701859473
transform 1 0 5530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1176_
timestamp 1701859473
transform -1 0 4850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1701859473
transform 1 0 5250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1701859473
transform -1 0 4850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1179_
timestamp 1701859473
transform -1 0 4770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1701859473
transform -1 0 5370 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1181_
timestamp 1701859473
transform -1 0 4990 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1701859473
transform -1 0 4910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1183_
timestamp 1701859473
transform -1 0 4630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1701859473
transform -1 0 4250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1701859473
transform 1 0 4090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1186_
timestamp 1701859473
transform -1 0 3830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1701859473
transform 1 0 3050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1188_
timestamp 1701859473
transform -1 0 3290 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1701859473
transform 1 0 3790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1190_
timestamp 1701859473
transform -1 0 3910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1701859473
transform 1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1192_
timestamp 1701859473
transform 1 0 3970 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1701859473
transform 1 0 5430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1701859473
transform -1 0 5130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1195_
timestamp 1701859473
transform 1 0 4450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1701859473
transform -1 0 5110 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1197_
timestamp 1701859473
transform -1 0 4630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1701859473
transform -1 0 5250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1199_
timestamp 1701859473
transform 1 0 5090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1701859473
transform -1 0 4950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1701859473
transform 1 0 4610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1202_
timestamp 1701859473
transform 1 0 4670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1701859473
transform -1 0 5230 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1204_
timestamp 1701859473
transform -1 0 4830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1701859473
transform -1 0 4730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1206_
timestamp 1701859473
transform -1 0 5550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1701859473
transform 1 0 5030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1701859473
transform 1 0 6030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1209_
timestamp 1701859473
transform 1 0 4070 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1701859473
transform 1 0 5050 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1211_
timestamp 1701859473
transform -1 0 4470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1701859473
transform -1 0 4450 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1213_
timestamp 1701859473
transform 1 0 4770 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1701859473
transform 1 0 4910 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1701859473
transform 1 0 5050 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1216_
timestamp 1701859473
transform 1 0 4770 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1701859473
transform 1 0 4630 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1218_
timestamp 1701859473
transform 1 0 4910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1701859473
transform -1 0 5230 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1220_
timestamp 1701859473
transform -1 0 5570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1701859473
transform -1 0 3490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1701859473
transform 1 0 3150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1223_
timestamp 1701859473
transform 1 0 3090 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1701859473
transform -1 0 3390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1225_
timestamp 1701859473
transform -1 0 3530 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1701859473
transform -1 0 3530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1227_
timestamp 1701859473
transform -1 0 3430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1701859473
transform 1 0 3250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1701859473
transform -1 0 3670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1230_
timestamp 1701859473
transform -1 0 3550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1701859473
transform -1 0 3290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1232_
timestamp 1701859473
transform -1 0 4170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1701859473
transform -1 0 4930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1234_
timestamp 1701859473
transform -1 0 4550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1701859473
transform -1 0 4710 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1236_
timestamp 1701859473
transform 1 0 5010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1701859473
transform 1 0 4770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1701859473
transform -1 0 4510 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1239_
timestamp 1701859473
transform -1 0 4690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1701859473
transform 1 0 4950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1241_
timestamp 1701859473
transform 1 0 4010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1701859473
transform 1 0 4870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1243_
timestamp 1701859473
transform -1 0 4570 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1701859473
transform -1 0 4270 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1701859473
transform 1 0 5390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1246_
timestamp 1701859473
transform 1 0 5590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1701859473
transform 1 0 4290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1248_
timestamp 1701859473
transform -1 0 4810 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1701859473
transform 1 0 5350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1250_
timestamp 1701859473
transform 1 0 5630 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1701859473
transform 1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1701859473
transform -1 0 5270 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1253_
timestamp 1701859473
transform 1 0 5310 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1701859473
transform 1 0 5670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1255_
timestamp 1701859473
transform 1 0 5810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1701859473
transform -1 0 5910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1257_
timestamp 1701859473
transform 1 0 5490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1701859473
transform 1 0 5490 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1701859473
transform 1 0 5790 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1260_
timestamp 1701859473
transform 1 0 5210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1701859473
transform 1 0 5310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1262_
timestamp 1701859473
transform -1 0 5850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1701859473
transform 1 0 5950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1264_
timestamp 1701859473
transform -1 0 5550 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1701859473
transform 1 0 5430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1701859473
transform -1 0 5310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1267_
timestamp 1701859473
transform -1 0 5690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1701859473
transform 1 0 5070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1269_
timestamp 1701859473
transform -1 0 5170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1701859473
transform -1 0 3390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1271_
timestamp 1701859473
transform 1 0 2490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1701859473
transform 1 0 1090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1701859473
transform 1 0 1530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1274_
timestamp 1701859473
transform -1 0 2430 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1701859473
transform -1 0 2570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1276_
timestamp 1701859473
transform -1 0 2150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1701859473
transform 1 0 2270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1278_
timestamp 1701859473
transform 1 0 750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1701859473
transform 1 0 610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1280_
timestamp 1701859473
transform 1 0 1070 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1701859473
transform -1 0 1630 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1701859473
transform 1 0 1170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1283_
timestamp 1701859473
transform 1 0 1710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1701859473
transform 1 0 5390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1285_
timestamp 1701859473
transform -1 0 5250 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1701859473
transform -1 0 5430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1287_
timestamp 1701859473
transform -1 0 5530 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1701859473
transform -1 0 5110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1701859473
transform 1 0 4950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1290_
timestamp 1701859473
transform 1 0 4790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1701859473
transform 1 0 4990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1292_
timestamp 1701859473
transform -1 0 3810 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1701859473
transform -1 0 3550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1294_
timestamp 1701859473
transform 1 0 4810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1701859473
transform -1 0 4950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1701859473
transform 1 0 4610 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1297_
timestamp 1701859473
transform 1 0 4210 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1701859473
transform 1 0 5110 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1299_
timestamp 1701859473
transform 1 0 5150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1701859473
transform 1 0 3670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1301_
timestamp 1701859473
transform -1 0 3950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1701859473
transform -1 0 3790 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1701859473
transform -1 0 3910 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1304_
timestamp 1701859473
transform -1 0 3630 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1701859473
transform 1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1306_
timestamp 1701859473
transform 1 0 3530 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1701859473
transform 1 0 4410 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1308_
timestamp 1701859473
transform -1 0 4130 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1701859473
transform -1 0 3390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1701859473
transform 1 0 2610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1311_
timestamp 1701859473
transform 1 0 2870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1701859473
transform 1 0 2370 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1313_
timestamp 1701859473
transform 1 0 2670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1701859473
transform 1 0 2830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1315_
timestamp 1701859473
transform -1 0 2390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1701859473
transform 1 0 2550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1701859473
transform 1 0 3130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1318_
timestamp 1701859473
transform 1 0 2270 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1701859473
transform 1 0 2510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1320_
timestamp 1701859473
transform -1 0 2970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1701859473
transform 1 0 2790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1322_
timestamp 1701859473
transform 1 0 3290 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1701859473
transform 1 0 2650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1324_
timestamp 1701859473
transform -1 0 3110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1701859473
transform -1 0 3270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1701859473
transform -1 0 2950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1327_
timestamp 1701859473
transform 1 0 3850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1701859473
transform -1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1329_
timestamp 1701859473
transform -1 0 4770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1701859473
transform -1 0 4610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1331_
timestamp 1701859473
transform -1 0 3730 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1701859473
transform 1 0 3770 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1701859473
transform 1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1334_
timestamp 1701859473
transform -1 0 3870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1701859473
transform 1 0 3930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1336_
timestamp 1701859473
transform 1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1701859473
transform 1 0 4050 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1338_
timestamp 1701859473
transform 1 0 5470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1701859473
transform 1 0 5710 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1701859473
transform 1 0 3590 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1341_
timestamp 1701859473
transform 1 0 3970 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1701859473
transform -1 0 4370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1343_
timestamp 1701859473
transform 1 0 4190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1701859473
transform -1 0 4350 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1345_
timestamp 1701859473
transform 1 0 4310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1701859473
transform 1 0 4190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1701859473
transform 1 0 4470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1348_
timestamp 1701859473
transform 1 0 4470 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1701859473
transform -1 0 4510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1350_
timestamp 1701859473
transform -1 0 5990 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1701859473
transform 1 0 5850 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1352_
timestamp 1701859473
transform -1 0 4090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1701859473
transform -1 0 3930 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1701859473
transform -1 0 3630 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1355_
timestamp 1701859473
transform 1 0 3470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1701859473
transform -1 0 2870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1357_
timestamp 1701859473
transform -1 0 2710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1701859473
transform -1 0 2150 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1359_
timestamp 1701859473
transform -1 0 2910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1701859473
transform 1 0 1890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1701859473
transform -1 0 2750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1362_
timestamp 1701859473
transform -1 0 2030 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1701859473
transform -1 0 1250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1364_
timestamp 1701859473
transform 1 0 1190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1701859473
transform -1 0 510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1366_
timestamp 1701859473
transform -1 0 3470 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1701859473
transform -1 0 4670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1368_
timestamp 1701859473
transform -1 0 3350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1701859473
transform -1 0 2750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1701859473
transform -1 0 3070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1371_
timestamp 1701859473
transform 1 0 2370 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1701859473
transform -1 0 3530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1373_
timestamp 1701859473
transform 1 0 3390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1701859473
transform -1 0 3350 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1375_
timestamp 1701859473
transform -1 0 3470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1701859473
transform -1 0 3010 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1701859473
transform -1 0 3030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1378_
timestamp 1701859473
transform -1 0 3150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1701859473
transform 1 0 2730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1380_
timestamp 1701859473
transform 1 0 3230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1701859473
transform -1 0 3110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1382_
timestamp 1701859473
transform -1 0 2950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1701859473
transform -1 0 3010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1701859473
transform 1 0 3270 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1385_
timestamp 1701859473
transform 1 0 2870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1701859473
transform 1 0 2590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1387_
timestamp 1701859473
transform -1 0 4230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1701859473
transform 1 0 2490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1389_
timestamp 1701859473
transform 1 0 2050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1701859473
transform 1 0 1930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1701859473
transform 1 0 2190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1392_
timestamp 1701859473
transform -1 0 2410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1701859473
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1394_
timestamp 1701859473
transform 1 0 2310 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1701859473
transform -1 0 3070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1396_
timestamp 1701859473
transform -1 0 2930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1701859473
transform -1 0 2790 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1701859473
transform 1 0 2630 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1399_
timestamp 1701859473
transform -1 0 2610 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1701859473
transform 1 0 3210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1401_
timestamp 1701859473
transform -1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1701859473
transform -1 0 2490 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1403_
timestamp 1701859473
transform -1 0 2310 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1701859473
transform 1 0 2750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1701859473
transform -1 0 3630 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1406_
timestamp 1701859473
transform -1 0 2770 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1701859473
transform -1 0 2910 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1408_
timestamp 1701859473
transform 1 0 2470 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1701859473
transform -1 0 2750 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1410_
timestamp 1701859473
transform -1 0 2910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1701859473
transform 1 0 2890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1412_
timestamp 1701859473
transform -1 0 2610 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1701859473
transform 1 0 3030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1701859473
transform -1 0 3190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1415_
timestamp 1701859473
transform -1 0 3190 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1701859473
transform -1 0 3310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1417_
timestamp 1701859473
transform -1 0 3930 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1701859473
transform -1 0 3770 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1419_
timestamp 1701859473
transform -1 0 3050 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1701859473
transform 1 0 1990 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1701859473
transform -1 0 2610 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1422_
timestamp 1701859473
transform -1 0 2810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1701859473
transform -1 0 2670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1424_
timestamp 1701859473
transform -1 0 2550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1701859473
transform -1 0 2490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1426_
timestamp 1701859473
transform -1 0 2330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1701859473
transform 1 0 350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1701859473
transform 1 0 750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1429_
timestamp 1701859473
transform -1 0 3710 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1701859473
transform -1 0 3430 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1431_
timestamp 1701859473
transform 1 0 1030 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1701859473
transform -1 0 1010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1433_
timestamp 1701859473
transform -1 0 1150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1701859473
transform 1 0 150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1701859473
transform -1 0 510 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1436_
timestamp 1701859473
transform -1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1701859473
transform 1 0 1850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1438_
timestamp 1701859473
transform 1 0 2250 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1701859473
transform 1 0 3110 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1440_
timestamp 1701859473
transform -1 0 1810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1701859473
transform -1 0 2150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1701859473
transform -1 0 1950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1443_
timestamp 1701859473
transform -1 0 1670 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1701859473
transform -1 0 1550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1445_
timestamp 1701859473
transform 1 0 2050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1701859473
transform 1 0 1790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1447_
timestamp 1701859473
transform 1 0 1650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1701859473
transform 1 0 1390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1701859473
transform -1 0 1510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1450_
timestamp 1701859473
transform -1 0 1750 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1701859473
transform 1 0 1570 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1452_
timestamp 1701859473
transform -1 0 2030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1453_
timestamp 1701859473
transform 1 0 1310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1454_
timestamp 1701859473
transform -1 0 1810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1455_
timestamp 1701859473
transform 1 0 1670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1456_
timestamp 1701859473
transform 1 0 1790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1457_
timestamp 1701859473
transform -1 0 1890 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1458_
timestamp 1701859473
transform 1 0 1390 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1459_
timestamp 1701859473
transform -1 0 1270 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1460_
timestamp 1701859473
transform -1 0 1250 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1461_
timestamp 1701859473
transform 1 0 1350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1462_
timestamp 1701859473
transform -1 0 2490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1463_
timestamp 1701859473
transform -1 0 1150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1464_
timestamp 1701859473
transform 1 0 1490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1465_
timestamp 1701859473
transform 1 0 1650 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1466_
timestamp 1701859473
transform 1 0 1090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1467_
timestamp 1701859473
transform 1 0 1550 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1468_
timestamp 1701859473
transform -1 0 1710 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1469_
timestamp 1701859473
transform 1 0 1890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1470_
timestamp 1701859473
transform -1 0 2170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1471_
timestamp 1701859473
transform -1 0 2470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1472_
timestamp 1701859473
transform -1 0 2330 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1473_
timestamp 1701859473
transform 1 0 2010 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1474_
timestamp 1701859473
transform -1 0 2130 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1475_
timestamp 1701859473
transform -1 0 2170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1476_
timestamp 1701859473
transform -1 0 2390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1477_
timestamp 1701859473
transform 1 0 1910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1478_
timestamp 1701859473
transform 1 0 2010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1479_
timestamp 1701859473
transform -1 0 2030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1480_
timestamp 1701859473
transform 1 0 4330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1481_
timestamp 1701859473
transform 1 0 4090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1482_
timestamp 1701859473
transform -1 0 4250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1483_
timestamp 1701859473
transform -1 0 1310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1484_
timestamp 1701859473
transform 1 0 1150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1485_
timestamp 1701859473
transform -1 0 890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1486_
timestamp 1701859473
transform 1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1487_
timestamp 1701859473
transform -1 0 310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1488_
timestamp 1701859473
transform -1 0 1270 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1489_
timestamp 1701859473
transform -1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1490_
timestamp 1701859473
transform 1 0 1570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1491_
timestamp 1701859473
transform 1 0 2170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1492_
timestamp 1701859473
transform -1 0 2050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1493_
timestamp 1701859473
transform 1 0 1870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1494_
timestamp 1701859473
transform -1 0 1750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1495_
timestamp 1701859473
transform 1 0 1330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1496_
timestamp 1701859473
transform 1 0 1590 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1497_
timestamp 1701859473
transform 1 0 1510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1498_
timestamp 1701859473
transform -1 0 1670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1499_
timestamp 1701859473
transform -1 0 1470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1500_
timestamp 1701859473
transform 1 0 1450 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1501_
timestamp 1701859473
transform 1 0 1590 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1502_
timestamp 1701859473
transform -1 0 450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1503_
timestamp 1701859473
transform 1 0 670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1504_
timestamp 1701859473
transform -1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1505_
timestamp 1701859473
transform -1 0 310 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1506_
timestamp 1701859473
transform -1 0 950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1507_
timestamp 1701859473
transform -1 0 810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1508_
timestamp 1701859473
transform -1 0 730 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1509_
timestamp 1701859473
transform -1 0 870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1510_
timestamp 1701859473
transform 1 0 990 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1511_
timestamp 1701859473
transform -1 0 590 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1512_
timestamp 1701859473
transform 1 0 730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1513_
timestamp 1701859473
transform -1 0 3430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1514_
timestamp 1701859473
transform 1 0 2070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1515_
timestamp 1701859473
transform -1 0 2190 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1516_
timestamp 1701859473
transform -1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1517_
timestamp 1701859473
transform 1 0 1770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1518_
timestamp 1701859473
transform -1 0 770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1519_
timestamp 1701859473
transform 1 0 1830 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1520_
timestamp 1701859473
transform -1 0 1970 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1521_
timestamp 1701859473
transform 1 0 1930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1522_
timestamp 1701859473
transform -1 0 2230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1523_
timestamp 1701859473
transform 1 0 1030 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1524_
timestamp 1701859473
transform -1 0 330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1525_
timestamp 1701859473
transform 1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1526_
timestamp 1701859473
transform 1 0 290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1527_
timestamp 1701859473
transform -1 0 4510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1528_
timestamp 1701859473
transform -1 0 4610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1529_
timestamp 1701859473
transform 1 0 4350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1530_
timestamp 1701859473
transform 1 0 750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1531_
timestamp 1701859473
transform -1 0 890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1532_
timestamp 1701859473
transform -1 0 950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1533_
timestamp 1701859473
transform 1 0 290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1534_
timestamp 1701859473
transform 1 0 310 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1535_
timestamp 1701859473
transform -1 0 1370 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1536_
timestamp 1701859473
transform -1 0 1470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1537_
timestamp 1701859473
transform -1 0 350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1538_
timestamp 1701859473
transform -1 0 170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1539_
timestamp 1701859473
transform -1 0 1730 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1540_
timestamp 1701859473
transform 1 0 1210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1541_
timestamp 1701859473
transform -1 0 1070 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1542_
timestamp 1701859473
transform -1 0 1370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1543_
timestamp 1701859473
transform -1 0 1090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1544_
timestamp 1701859473
transform -1 0 1430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1545_
timestamp 1701859473
transform -1 0 1070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1546_
timestamp 1701859473
transform 1 0 150 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1547_
timestamp 1701859473
transform 1 0 450 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1548_
timestamp 1701859473
transform -1 0 590 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1549_
timestamp 1701859473
transform 1 0 450 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1550_
timestamp 1701859473
transform 1 0 590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1551_
timestamp 1701859473
transform -1 0 4490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1552_
timestamp 1701859473
transform -1 0 4670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1553_
timestamp 1701859473
transform 1 0 650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1554_
timestamp 1701859473
transform -1 0 1290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1555_
timestamp 1701859473
transform -1 0 1210 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1556_
timestamp 1701859473
transform 1 0 870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1557_
timestamp 1701859473
transform 1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1558_
timestamp 1701859473
transform 1 0 870 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1559_
timestamp 1701859473
transform 1 0 1190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1560_
timestamp 1701859473
transform -1 0 1310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1561_
timestamp 1701859473
transform -1 0 210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1562_
timestamp 1701859473
transform 1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1563_
timestamp 1701859473
transform -1 0 330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1564_
timestamp 1701859473
transform -1 0 1150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1565_
timestamp 1701859473
transform -1 0 1270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1566_
timestamp 1701859473
transform -1 0 1390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1567_
timestamp 1701859473
transform -1 0 1230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1568_
timestamp 1701859473
transform -1 0 1230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1569_
timestamp 1701859473
transform -1 0 1010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1570_
timestamp 1701859473
transform -1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1571_
timestamp 1701859473
transform -1 0 730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1572_
timestamp 1701859473
transform 1 0 570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1573_
timestamp 1701859473
transform -1 0 430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1574_
timestamp 1701859473
transform -1 0 5130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1575_
timestamp 1701859473
transform 1 0 4970 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1576_
timestamp 1701859473
transform -1 0 4850 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1577_
timestamp 1701859473
transform -1 0 4690 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1578_
timestamp 1701859473
transform 1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1579_
timestamp 1701859473
transform 1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1580_
timestamp 1701859473
transform -1 0 230 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1581_
timestamp 1701859473
transform 1 0 130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1582_
timestamp 1701859473
transform 1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1583_
timestamp 1701859473
transform -1 0 850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1584_
timestamp 1701859473
transform -1 0 950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1585_
timestamp 1701859473
transform -1 0 650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1586_
timestamp 1701859473
transform -1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1587_
timestamp 1701859473
transform -1 0 4870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1588_
timestamp 1701859473
transform -1 0 4690 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1589_
timestamp 1701859473
transform -1 0 1490 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1590_
timestamp 1701859473
transform -1 0 1190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1591_
timestamp 1701859473
transform -1 0 1050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1592_
timestamp 1701859473
transform 1 0 130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1593_
timestamp 1701859473
transform 1 0 2530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1594_
timestamp 1701859473
transform -1 0 2670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1595_
timestamp 1701859473
transform 1 0 3610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1596_
timestamp 1701859473
transform 1 0 3450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1597_
timestamp 1701859473
transform -1 0 2470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1598_
timestamp 1701859473
transform 1 0 2290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1599_
timestamp 1701859473
transform -1 0 3730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1600_
timestamp 1701859473
transform 1 0 3550 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1601_
timestamp 1701859473
transform 1 0 3250 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1602_
timestamp 1701859473
transform 1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1603_
timestamp 1701859473
transform -1 0 2870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1604_
timestamp 1701859473
transform 1 0 2690 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1605_
timestamp 1701859473
transform 1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1606_
timestamp 1701859473
transform 1 0 1870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1607_
timestamp 1701859473
transform -1 0 1710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1608_
timestamp 1701859473
transform 1 0 1530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1636_
timestamp 1701859473
transform -1 0 4230 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1637_
timestamp 1701859473
transform -1 0 4330 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1638_
timestamp 1701859473
transform -1 0 4090 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1639_
timestamp 1701859473
transform 1 0 3930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1640_
timestamp 1701859473
transform -1 0 3690 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1641_
timestamp 1701859473
transform -1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1642_
timestamp 1701859473
transform -1 0 3190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1643_
timestamp 1701859473
transform -1 0 4090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1644_
timestamp 1701859473
transform -1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1645_
timestamp 1701859473
transform 1 0 4470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1646_
timestamp 1701859473
transform -1 0 4210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1647_
timestamp 1701859473
transform 1 0 3290 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1648_
timestamp 1701859473
transform -1 0 4210 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1649_
timestamp 1701859473
transform -1 0 3810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1650_
timestamp 1701859473
transform -1 0 3930 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1651_
timestamp 1701859473
transform 1 0 3650 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1652_
timestamp 1701859473
transform 1 0 3650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1653_
timestamp 1701859473
transform 1 0 3770 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1654_
timestamp 1701859473
transform -1 0 4610 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1655_
timestamp 1701859473
transform -1 0 4470 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1656_
timestamp 1701859473
transform 1 0 1450 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1657_
timestamp 1701859473
transform 1 0 3090 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1658_
timestamp 1701859473
transform 1 0 3230 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1659_
timestamp 1701859473
transform -1 0 3190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1660_
timestamp 1701859473
transform 1 0 3530 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1661_
timestamp 1701859473
transform -1 0 3410 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1662_
timestamp 1701859473
transform 1 0 3530 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1663_
timestamp 1701859473
transform -1 0 3490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1664_
timestamp 1701859473
transform -1 0 3330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1665_
timestamp 1701859473
transform -1 0 3970 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1666_
timestamp 1701859473
transform 1 0 3830 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1667_
timestamp 1701859473
transform -1 0 3690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1668_
timestamp 1701859473
transform 1 0 3390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1669_
timestamp 1701859473
transform -1 0 3510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1670_
timestamp 1701859473
transform -1 0 3370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1671_
timestamp 1701859473
transform -1 0 3070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1672_
timestamp 1701859473
transform 1 0 2730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1673_
timestamp 1701859473
transform -1 0 2890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1674_
timestamp 1701859473
transform 1 0 2970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1675_
timestamp 1701859473
transform -1 0 4390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1676_
timestamp 1701859473
transform 1 0 4110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1677_
timestamp 1701859473
transform 1 0 3790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1678_
timestamp 1701859473
transform 1 0 4310 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1679_
timestamp 1701859473
transform 1 0 4590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1680_
timestamp 1701859473
transform -1 0 4490 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1681_
timestamp 1701859473
transform 1 0 3890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1682_
timestamp 1701859473
transform 1 0 4070 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1683_
timestamp 1701859473
transform 1 0 3950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1684_
timestamp 1701859473
transform 1 0 3770 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1685_
timestamp 1701859473
transform -1 0 2830 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1686_
timestamp 1701859473
transform -1 0 2550 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1687_
timestamp 1701859473
transform 1 0 2410 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1688_
timestamp 1701859473
transform -1 0 2150 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1689_
timestamp 1701859473
transform -1 0 1650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1690_
timestamp 1701859473
transform 1 0 2670 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1691_
timestamp 1701859473
transform -1 0 2290 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1692_
timestamp 1701859473
transform -1 0 2990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1693_
timestamp 1701859473
transform 1 0 3150 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1694_
timestamp 1701859473
transform 1 0 3150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1695_
timestamp 1701859473
transform -1 0 3570 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1696_
timestamp 1701859473
transform 1 0 3410 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1697_
timestamp 1701859473
transform -1 0 3290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1698_
timestamp 1701859473
transform -1 0 3130 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1699_
timestamp 1701859473
transform -1 0 2430 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1700_
timestamp 1701859473
transform 1 0 2250 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1701_
timestamp 1701859473
transform -1 0 2210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1702_
timestamp 1701859473
transform 1 0 2030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1703_
timestamp 1701859473
transform 1 0 1270 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1704_
timestamp 1701859473
transform -1 0 1230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1705_
timestamp 1701859473
transform 1 0 2330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1706_
timestamp 1701859473
transform -1 0 2450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1707_
timestamp 1701859473
transform 1 0 1890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1708_
timestamp 1701859473
transform -1 0 1870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1709_
timestamp 1701859473
transform -1 0 2630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1710_
timestamp 1701859473
transform -1 0 3030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1711_
timestamp 1701859473
transform 1 0 2870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1712_
timestamp 1701859473
transform 1 0 2410 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1713_
timestamp 1701859473
transform -1 0 2730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1714_
timestamp 1701859473
transform -1 0 2590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1715_
timestamp 1701859473
transform 1 0 2690 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1716_
timestamp 1701859473
transform 1 0 2550 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1717_
timestamp 1701859473
transform -1 0 2590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1718_
timestamp 1701859473
transform -1 0 2450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1719_
timestamp 1701859473
transform 1 0 2050 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1720_
timestamp 1701859473
transform 1 0 1870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1721_
timestamp 1701859473
transform 1 0 1590 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1722_
timestamp 1701859473
transform -1 0 2010 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1723_
timestamp 1701859473
transform 1 0 1730 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1724_
timestamp 1701859473
transform 1 0 1190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1725_
timestamp 1701859473
transform 1 0 1970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1726_
timestamp 1701859473
transform -1 0 890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1727_
timestamp 1701859473
transform -1 0 990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1728_
timestamp 1701859473
transform 1 0 2610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1729_
timestamp 1701859473
transform 1 0 1890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1730_
timestamp 1701859473
transform -1 0 2210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1731_
timestamp 1701859473
transform -1 0 2250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1732_
timestamp 1701859473
transform 1 0 2050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1733_
timestamp 1701859473
transform 1 0 2090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1734_
timestamp 1701859473
transform -1 0 1750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1735_
timestamp 1701859473
transform -1 0 1810 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1736_
timestamp 1701859473
transform 1 0 1630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1737_
timestamp 1701859473
transform -1 0 1510 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1738_
timestamp 1701859473
transform -1 0 1130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1739_
timestamp 1701859473
transform -1 0 930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1740_
timestamp 1701859473
transform -1 0 1250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1741_
timestamp 1701859473
transform -1 0 990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1742_
timestamp 1701859473
transform -1 0 2310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1743_
timestamp 1701859473
transform -1 0 3050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1744_
timestamp 1701859473
transform 1 0 2730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1745_
timestamp 1701859473
transform 1 0 2450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1746_
timestamp 1701859473
transform -1 0 2890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1747_
timestamp 1701859473
transform -1 0 2330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1748_
timestamp 1701859473
transform -1 0 1490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1749_
timestamp 1701859473
transform -1 0 1350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1750_
timestamp 1701859473
transform -1 0 830 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1751_
timestamp 1701859473
transform -1 0 790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1752_
timestamp 1701859473
transform -1 0 410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1753_
timestamp 1701859473
transform 1 0 310 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1754_
timestamp 1701859473
transform -1 0 530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1755_
timestamp 1701859473
transform -1 0 630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1756_
timestamp 1701859473
transform -1 0 1270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1757_
timestamp 1701859473
transform 1 0 1930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1758_
timestamp 1701859473
transform -1 0 2150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1759_
timestamp 1701859473
transform -1 0 2270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1760_
timestamp 1701859473
transform -1 0 1850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1761_
timestamp 1701859473
transform 1 0 1650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1762_
timestamp 1701859473
transform -1 0 1490 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1763_
timestamp 1701859473
transform -1 0 1330 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1764_
timestamp 1701859473
transform -1 0 890 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1765_
timestamp 1701859473
transform -1 0 730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1766_
timestamp 1701859473
transform -1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1767_
timestamp 1701859473
transform 1 0 1130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1768_
timestamp 1701859473
transform 1 0 1350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1769_
timestamp 1701859473
transform -1 0 1510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1770_
timestamp 1701859473
transform -1 0 1370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1771_
timestamp 1701859473
transform -1 0 670 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1772_
timestamp 1701859473
transform -1 0 510 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1773_
timestamp 1701859473
transform 1 0 750 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1774_
timestamp 1701859473
transform 1 0 330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1775_
timestamp 1701859473
transform 1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1776_
timestamp 1701859473
transform -1 0 470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1777_
timestamp 1701859473
transform -1 0 3690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1778_
timestamp 1701859473
transform 1 0 2730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1779_
timestamp 1701859473
transform -1 0 3050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1780_
timestamp 1701859473
transform -1 0 3510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1781_
timestamp 1701859473
transform 1 0 2890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1782_
timestamp 1701859473
transform 1 0 3330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1783_
timestamp 1701859473
transform -1 0 1490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1784_
timestamp 1701859473
transform -1 0 1330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1785_
timestamp 1701859473
transform -1 0 1150 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1786_
timestamp 1701859473
transform -1 0 990 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1787_
timestamp 1701859473
transform -1 0 550 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1788_
timestamp 1701859473
transform 1 0 610 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1789_
timestamp 1701859473
transform -1 0 610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1790_
timestamp 1701859473
transform -1 0 450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1791_
timestamp 1701859473
transform -1 0 330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1792_
timestamp 1701859473
transform -1 0 1750 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1793_
timestamp 1701859473
transform 1 0 1610 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1794_
timestamp 1701859473
transform 1 0 610 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1795_
timestamp 1701859473
transform -1 0 190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1796_
timestamp 1701859473
transform 1 0 250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1797_
timestamp 1701859473
transform 1 0 470 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1798_
timestamp 1701859473
transform -1 0 670 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1799_
timestamp 1701859473
transform 1 0 410 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1800_
timestamp 1701859473
transform 1 0 190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1801_
timestamp 1701859473
transform -1 0 210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1802_
timestamp 1701859473
transform -1 0 2870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1803_
timestamp 1701859473
transform 1 0 810 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1804_
timestamp 1701859473
transform -1 0 710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1805_
timestamp 1701859473
transform 1 0 810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1806_
timestamp 1701859473
transform 1 0 1010 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1807_
timestamp 1701859473
transform -1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1808_
timestamp 1701859473
transform -1 0 490 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1809_
timestamp 1701859473
transform -1 0 1170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1810_
timestamp 1701859473
transform -1 0 990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1811_
timestamp 1701859473
transform -1 0 170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1812_
timestamp 1701859473
transform -1 0 330 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1813_
timestamp 1701859473
transform -1 0 50 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1814_
timestamp 1701859473
transform -1 0 50 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1815_
timestamp 1701859473
transform -1 0 330 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1816_
timestamp 1701859473
transform 1 0 30 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1817_
timestamp 1701859473
transform -1 0 190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1818_
timestamp 1701859473
transform -1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1819_
timestamp 1701859473
transform -1 0 170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1820_
timestamp 1701859473
transform -1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1821_
timestamp 1701859473
transform 1 0 530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1822_
timestamp 1701859473
transform -1 0 310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1823_
timestamp 1701859473
transform -1 0 190 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1824_
timestamp 1701859473
transform 1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1825_
timestamp 1701859473
transform 1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1826_
timestamp 1701859473
transform 1 0 1070 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1701859473
transform -1 0 2790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1701859473
transform 1 0 3390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1701859473
transform 1 0 3450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1701859473
transform -1 0 2830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1701859473
transform -1 0 4550 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1701859473
transform 1 0 4550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1701859473
transform 1 0 4590 0 1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1701859473
transform 1 0 4730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert13
timestamp 1701859473
transform 1 0 3130 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert14
timestamp 1701859473
transform 1 0 2690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1701859473
transform -1 0 1990 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1701859473
transform -1 0 1850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1701859473
transform 1 0 430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1701859473
transform 1 0 3310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1701859473
transform 1 0 1810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1701859473
transform 1 0 1430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1701859473
transform -1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1701859473
transform -1 0 2750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1701859473
transform 1 0 3510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1701859473
transform 1 0 3830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1701859473
transform -1 0 3010 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1701859473
transform 1 0 2970 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1701859473
transform 1 0 2550 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1701859473
transform -1 0 1490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1701859473
transform 1 0 2550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1701859473
transform -1 0 2450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1701859473
transform 1 0 2910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1701859473
transform 1 0 1970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1701859473
transform 1 0 3310 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert34
timestamp 1701859473
transform -1 0 3590 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert35
timestamp 1701859473
transform -1 0 3970 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert36
timestamp 1701859473
transform 1 0 3970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert37
timestamp 1701859473
transform -1 0 3810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert38
timestamp 1701859473
transform 1 0 1730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert39
timestamp 1701859473
transform -1 0 4510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert40
timestamp 1701859473
transform -1 0 1630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert41
timestamp 1701859473
transform -1 0 2610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1701859473
transform 1 0 2170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1701859473
transform 1 0 1450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 1950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1701859473
transform 1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__889_
timestamp 1701859473
transform -1 0 1130 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__890_
timestamp 1701859473
transform 1 0 650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__891_
timestamp 1701859473
transform -1 0 710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__892_
timestamp 1701859473
transform 1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__893_
timestamp 1701859473
transform 1 0 1350 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__894_
timestamp 1701859473
transform 1 0 1070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__895_
timestamp 1701859473
transform 1 0 1590 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__896_
timestamp 1701859473
transform -1 0 1730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__897_
timestamp 1701859473
transform -1 0 970 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__898_
timestamp 1701859473
transform -1 0 1470 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__899_
timestamp 1701859473
transform -1 0 990 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__900_
timestamp 1701859473
transform -1 0 390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__901_
timestamp 1701859473
transform -1 0 530 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__902_
timestamp 1701859473
transform 1 0 190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__903_
timestamp 1701859473
transform -1 0 590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__904_
timestamp 1701859473
transform -1 0 670 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__905_
timestamp 1701859473
transform -1 0 630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__906_
timestamp 1701859473
transform -1 0 950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__907_
timestamp 1701859473
transform -1 0 930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__908_
timestamp 1701859473
transform -1 0 470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__909_
timestamp 1701859473
transform -1 0 830 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__910_
timestamp 1701859473
transform 1 0 710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__911_
timestamp 1701859473
transform 1 0 430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__912_
timestamp 1701859473
transform -1 0 330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__913_
timestamp 1701859473
transform 1 0 210 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__914_
timestamp 1701859473
transform 1 0 310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__915_
timestamp 1701859473
transform 1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__916_
timestamp 1701859473
transform -1 0 570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__917_
timestamp 1701859473
transform 1 0 650 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__918_
timestamp 1701859473
transform -1 0 1070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__919_
timestamp 1701859473
transform 1 0 790 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__920_
timestamp 1701859473
transform -1 0 1410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__921_
timestamp 1701859473
transform -1 0 1230 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__922_
timestamp 1701859473
transform 1 0 850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__923_
timestamp 1701859473
transform -1 0 1150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__924_
timestamp 1701859473
transform 1 0 990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__925_
timestamp 1701859473
transform 1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__926_
timestamp 1701859473
transform 1 0 3190 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__927_
timestamp 1701859473
transform -1 0 3090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__928_
timestamp 1701859473
transform 1 0 3210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__929_
timestamp 1701859473
transform -1 0 3750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__930_
timestamp 1701859473
transform -1 0 3910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__931_
timestamp 1701859473
transform 1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__932_
timestamp 1701859473
transform 1 0 2170 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__933_
timestamp 1701859473
transform 1 0 2030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__934_
timestamp 1701859473
transform -1 0 2170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__935_
timestamp 1701859473
transform 1 0 4390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__936_
timestamp 1701859473
transform -1 0 3610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__937_
timestamp 1701859473
transform -1 0 3470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__938_
timestamp 1701859473
transform 1 0 2950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__939_
timestamp 1701859473
transform 1 0 2710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__940_
timestamp 1701859473
transform -1 0 2850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__941_
timestamp 1701859473
transform 1 0 2450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__942_
timestamp 1701859473
transform -1 0 2610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__943_
timestamp 1701859473
transform 1 0 2730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__944_
timestamp 1701859473
transform 1 0 1430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__945_
timestamp 1701859473
transform -1 0 1630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__946_
timestamp 1701859473
transform -1 0 1750 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__947_
timestamp 1701859473
transform -1 0 1330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__948_
timestamp 1701859473
transform -1 0 1730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__949_
timestamp 1701859473
transform -1 0 1870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__950_
timestamp 1701859473
transform -1 0 70 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__951_
timestamp 1701859473
transform 1 0 4310 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__952_
timestamp 1701859473
transform 1 0 2690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__953_
timestamp 1701859473
transform 1 0 4210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__954_
timestamp 1701859473
transform 1 0 4110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__955_
timestamp 1701859473
transform 1 0 4350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__956_
timestamp 1701859473
transform 1 0 5010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__957_
timestamp 1701859473
transform 1 0 4650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__958_
timestamp 1701859473
transform 1 0 4910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__959_
timestamp 1701859473
transform -1 0 5210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__960_
timestamp 1701859473
transform -1 0 4790 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__961_
timestamp 1701859473
transform -1 0 5070 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__962_
timestamp 1701859473
transform -1 0 5310 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__963_
timestamp 1701859473
transform 1 0 6050 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__964_
timestamp 1701859473
transform 1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__965_
timestamp 1701859473
transform 1 0 5230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__966_
timestamp 1701859473
transform -1 0 6030 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__967_
timestamp 1701859473
transform 1 0 4870 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__968_
timestamp 1701859473
transform 1 0 3310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__969_
timestamp 1701859473
transform 1 0 5410 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__970_
timestamp 1701859473
transform -1 0 5950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__971_
timestamp 1701859473
transform -1 0 6050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__972_
timestamp 1701859473
transform -1 0 6010 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__973_
timestamp 1701859473
transform -1 0 5770 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__974_
timestamp 1701859473
transform 1 0 5470 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__975_
timestamp 1701859473
transform 1 0 4750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__976_
timestamp 1701859473
transform -1 0 4430 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__977_
timestamp 1701859473
transform 1 0 3070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__978_
timestamp 1701859473
transform -1 0 4430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__979_
timestamp 1701859473
transform 1 0 4550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__980_
timestamp 1701859473
transform 1 0 4790 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__981_
timestamp 1701859473
transform 1 0 5610 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__982_
timestamp 1701859473
transform 1 0 5710 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__983_
timestamp 1701859473
transform 1 0 5870 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__984_
timestamp 1701859473
transform 1 0 4930 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__985_
timestamp 1701859473
transform 1 0 4930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__986_
timestamp 1701859473
transform 1 0 5350 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__987_
timestamp 1701859473
transform -1 0 5930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__988_
timestamp 1701859473
transform -1 0 5290 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__989_
timestamp 1701859473
transform 1 0 5530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__990_
timestamp 1701859473
transform 1 0 5990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__991_
timestamp 1701859473
transform -1 0 5090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__992_
timestamp 1701859473
transform -1 0 5110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__993_
timestamp 1701859473
transform 1 0 5630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__994_
timestamp 1701859473
transform -1 0 6050 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__995_
timestamp 1701859473
transform 1 0 6070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__996_
timestamp 1701859473
transform 1 0 5370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__997_
timestamp 1701859473
transform -1 0 5850 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__998_
timestamp 1701859473
transform 1 0 5570 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__999_
timestamp 1701859473
transform 1 0 4030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1000_
timestamp 1701859473
transform -1 0 4190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1001_
timestamp 1701859473
transform 1 0 3830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1002_
timestamp 1701859473
transform -1 0 4270 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1003_
timestamp 1701859473
transform 1 0 4690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1004_
timestamp 1701859473
transform 1 0 4370 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1005_
timestamp 1701859473
transform -1 0 4550 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1006_
timestamp 1701859473
transform -1 0 4430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1007_
timestamp 1701859473
transform 1 0 3730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1008_
timestamp 1701859473
transform 1 0 3990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1009_
timestamp 1701859473
transform 1 0 4270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1010_
timestamp 1701859473
transform -1 0 5850 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1011_
timestamp 1701859473
transform -1 0 5730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1012_
timestamp 1701859473
transform 1 0 5410 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1013_
timestamp 1701859473
transform -1 0 5910 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1014_
timestamp 1701859473
transform 1 0 6130 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1015_
timestamp 1701859473
transform -1 0 5870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1016_
timestamp 1701859473
transform 1 0 5550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1017_
timestamp 1701859473
transform -1 0 5430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1018_
timestamp 1701859473
transform 1 0 4930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1019_
timestamp 1701859473
transform 1 0 5970 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1020_
timestamp 1701859473
transform 1 0 6010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1021_
timestamp 1701859473
transform 1 0 3670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1022_
timestamp 1701859473
transform -1 0 4830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1023_
timestamp 1701859473
transform -1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1024_
timestamp 1701859473
transform -1 0 2130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1025_
timestamp 1701859473
transform -1 0 4570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1026_
timestamp 1701859473
transform 1 0 4670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1027_
timestamp 1701859473
transform 1 0 5390 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1028_
timestamp 1701859473
transform 1 0 5390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1029_
timestamp 1701859473
transform 1 0 5070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1030_
timestamp 1701859473
transform -1 0 4970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1031_
timestamp 1701859473
transform -1 0 4390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1032_
timestamp 1701859473
transform 1 0 5650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1033_
timestamp 1701859473
transform 1 0 5810 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1034_
timestamp 1701859473
transform -1 0 5790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1035_
timestamp 1701859473
transform -1 0 5510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1036_
timestamp 1701859473
transform 1 0 5790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1037_
timestamp 1701859473
transform 1 0 6090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1038_
timestamp 1701859473
transform -1 0 3790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1039_
timestamp 1701859473
transform -1 0 3910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1040_
timestamp 1701859473
transform 1 0 3950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1041_
timestamp 1701859473
transform 1 0 4490 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1042_
timestamp 1701859473
transform 1 0 4250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1043_
timestamp 1701859473
transform 1 0 4270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1044_
timestamp 1701859473
transform 1 0 4290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1045_
timestamp 1701859473
transform 1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1046_
timestamp 1701859473
transform 1 0 4190 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1047_
timestamp 1701859473
transform 1 0 4090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1048_
timestamp 1701859473
transform 1 0 4650 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1049_
timestamp 1701859473
transform 1 0 4790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1050_
timestamp 1701859473
transform 1 0 5230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1051_
timestamp 1701859473
transform 1 0 6110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1052_
timestamp 1701859473
transform -1 0 5950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1053_
timestamp 1701859473
transform 1 0 5670 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1054_
timestamp 1701859473
transform -1 0 5110 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1055_
timestamp 1701859473
transform 1 0 5670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1056_
timestamp 1701859473
transform -1 0 6130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1057_
timestamp 1701859473
transform 1 0 5990 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1058_
timestamp 1701859473
transform 1 0 5810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1059_
timestamp 1701859473
transform -1 0 5990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1060_
timestamp 1701859473
transform -1 0 6110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1061_
timestamp 1701859473
transform 1 0 1350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1062_
timestamp 1701859473
transform 1 0 4150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1063_
timestamp 1701859473
transform 1 0 4790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1064_
timestamp 1701859473
transform 1 0 5310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1065_
timestamp 1701859473
transform 1 0 5870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1066_
timestamp 1701859473
transform -1 0 5670 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1067_
timestamp 1701859473
transform -1 0 5970 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1068_
timestamp 1701859473
transform -1 0 5990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1069_
timestamp 1701859473
transform -1 0 5530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1070_
timestamp 1701859473
transform -1 0 5290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1071_
timestamp 1701859473
transform 1 0 5190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1072_
timestamp 1701859473
transform 1 0 5450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1073_
timestamp 1701859473
transform 1 0 5510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1074_
timestamp 1701859473
transform 1 0 6130 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1075_
timestamp 1701859473
transform 1 0 5670 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1076_
timestamp 1701859473
transform 1 0 4690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1077_
timestamp 1701859473
transform -1 0 4530 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1078_
timestamp 1701859473
transform -1 0 5090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1079_
timestamp 1701859473
transform -1 0 4030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1080_
timestamp 1701859473
transform -1 0 4990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1081_
timestamp 1701859473
transform 1 0 5170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1082_
timestamp 1701859473
transform -1 0 4410 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1083_
timestamp 1701859473
transform -1 0 4850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1084_
timestamp 1701859473
transform -1 0 5250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1085_
timestamp 1701859473
transform 1 0 5990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1086_
timestamp 1701859473
transform 1 0 5370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1087_
timestamp 1701859473
transform 1 0 5070 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1088_
timestamp 1701859473
transform -1 0 5530 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1089_
timestamp 1701859473
transform -1 0 4070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1090_
timestamp 1701859473
transform 1 0 4350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1091_
timestamp 1701859473
transform 1 0 3610 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1092_
timestamp 1701859473
transform 1 0 3830 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1093_
timestamp 1701859473
transform -1 0 4290 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1094_
timestamp 1701859473
transform 1 0 3830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1095_
timestamp 1701859473
transform 1 0 4290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1096_
timestamp 1701859473
transform 1 0 4390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1097_
timestamp 1701859473
transform 1 0 4130 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1098_
timestamp 1701859473
transform 1 0 3970 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1099_
timestamp 1701859473
transform 1 0 4150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1100_
timestamp 1701859473
transform 1 0 5450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1101_
timestamp 1701859473
transform -1 0 5950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1102_
timestamp 1701859473
transform 1 0 5230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1103_
timestamp 1701859473
transform 1 0 5530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1104_
timestamp 1701859473
transform -1 0 5850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1105_
timestamp 1701859473
transform 1 0 5330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1106_
timestamp 1701859473
transform 1 0 5770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1107_
timestamp 1701859473
transform 1 0 5990 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1108_
timestamp 1701859473
transform 1 0 5970 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1109_
timestamp 1701859473
transform 1 0 5710 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1110_
timestamp 1701859473
transform -1 0 6090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1111_
timestamp 1701859473
transform 1 0 6030 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1112_
timestamp 1701859473
transform -1 0 3710 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1113_
timestamp 1701859473
transform 1 0 4590 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1114_
timestamp 1701859473
transform 1 0 4010 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1115_
timestamp 1701859473
transform -1 0 3970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1116_
timestamp 1701859473
transform 1 0 3810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1117_
timestamp 1701859473
transform 1 0 3670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1118_
timestamp 1701859473
transform 1 0 4170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1119_
timestamp 1701859473
transform -1 0 4450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1120_
timestamp 1701859473
transform -1 0 4070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1121_
timestamp 1701859473
transform -1 0 4210 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1122_
timestamp 1701859473
transform 1 0 4290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1123_
timestamp 1701859473
transform 1 0 4370 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1124_
timestamp 1701859473
transform 1 0 6010 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1125_
timestamp 1701859473
transform -1 0 5930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1126_
timestamp 1701859473
transform -1 0 5870 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1127_
timestamp 1701859473
transform 1 0 4890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1128_
timestamp 1701859473
transform 1 0 4590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1129_
timestamp 1701859473
transform 1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1130_
timestamp 1701859473
transform -1 0 5790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1131_
timestamp 1701859473
transform -1 0 5730 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1132_
timestamp 1701859473
transform -1 0 5830 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1133_
timestamp 1701859473
transform -1 0 5630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1134_
timestamp 1701859473
transform 1 0 6070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1135_
timestamp 1701859473
transform -1 0 5770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1136_
timestamp 1701859473
transform -1 0 5470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1137_
timestamp 1701859473
transform -1 0 5610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1138_
timestamp 1701859473
transform -1 0 5890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1139_
timestamp 1701859473
transform 1 0 5170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1140_
timestamp 1701859473
transform -1 0 5270 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1141_
timestamp 1701859473
transform -1 0 5170 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1142_
timestamp 1701859473
transform 1 0 4990 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1143_
timestamp 1701859473
transform -1 0 4950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1144_
timestamp 1701859473
transform -1 0 5370 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1145_
timestamp 1701859473
transform 1 0 4790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1146_
timestamp 1701859473
transform 1 0 5330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1147_
timestamp 1701859473
transform 1 0 5910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1148_
timestamp 1701859473
transform -1 0 5790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1149_
timestamp 1701859473
transform -1 0 5510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1150_
timestamp 1701859473
transform 1 0 4950 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1151_
timestamp 1701859473
transform 1 0 5630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1152_
timestamp 1701859473
transform 1 0 5870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1153_
timestamp 1701859473
transform -1 0 5610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1154_
timestamp 1701859473
transform -1 0 5750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1155_
timestamp 1701859473
transform -1 0 5470 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1156_
timestamp 1701859473
transform 1 0 5110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1157_
timestamp 1701859473
transform 1 0 5570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1158_
timestamp 1701859473
transform -1 0 5730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1159_
timestamp 1701859473
transform -1 0 5690 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1160_
timestamp 1701859473
transform -1 0 5030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1161_
timestamp 1701859473
transform -1 0 5330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1162_
timestamp 1701859473
transform -1 0 4890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1163_
timestamp 1701859473
transform -1 0 5730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1164_
timestamp 1701859473
transform -1 0 5230 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1165_
timestamp 1701859473
transform -1 0 4090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1166_
timestamp 1701859473
transform 1 0 4190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1167_
timestamp 1701859473
transform -1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1168_
timestamp 1701859473
transform 1 0 4750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1169_
timestamp 1701859473
transform 1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1170_
timestamp 1701859473
transform 1 0 5050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1171_
timestamp 1701859473
transform 1 0 5130 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1172_
timestamp 1701859473
transform -1 0 5010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1173_
timestamp 1701859473
transform 1 0 5290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1174_
timestamp 1701859473
transform 1 0 5570 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1175_
timestamp 1701859473
transform 1 0 5550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1176_
timestamp 1701859473
transform -1 0 4870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1177_
timestamp 1701859473
transform 1 0 5270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1178_
timestamp 1701859473
transform -1 0 4870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1179_
timestamp 1701859473
transform -1 0 4790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1180_
timestamp 1701859473
transform -1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1181_
timestamp 1701859473
transform -1 0 5010 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1182_
timestamp 1701859473
transform -1 0 4930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1183_
timestamp 1701859473
transform -1 0 4650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1184_
timestamp 1701859473
transform -1 0 4270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1185_
timestamp 1701859473
transform 1 0 4110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1186_
timestamp 1701859473
transform -1 0 3850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1187_
timestamp 1701859473
transform 1 0 3070 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1188_
timestamp 1701859473
transform -1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1189_
timestamp 1701859473
transform 1 0 3810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1190_
timestamp 1701859473
transform -1 0 3930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1191_
timestamp 1701859473
transform 1 0 3850 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1192_
timestamp 1701859473
transform 1 0 3990 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1193_
timestamp 1701859473
transform 1 0 5450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1194_
timestamp 1701859473
transform -1 0 5150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1195_
timestamp 1701859473
transform 1 0 4470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1196_
timestamp 1701859473
transform -1 0 5130 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1197_
timestamp 1701859473
transform -1 0 4650 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1198_
timestamp 1701859473
transform -1 0 5270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1199_
timestamp 1701859473
transform 1 0 5110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1200_
timestamp 1701859473
transform -1 0 4970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1201_
timestamp 1701859473
transform 1 0 4630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1202_
timestamp 1701859473
transform 1 0 4690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1203_
timestamp 1701859473
transform -1 0 5250 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1204_
timestamp 1701859473
transform -1 0 4850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1205_
timestamp 1701859473
transform -1 0 4750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1206_
timestamp 1701859473
transform -1 0 5570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1207_
timestamp 1701859473
transform 1 0 5050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1208_
timestamp 1701859473
transform 1 0 6050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1209_
timestamp 1701859473
transform 1 0 4090 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1210_
timestamp 1701859473
transform 1 0 5070 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1211_
timestamp 1701859473
transform -1 0 4490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1212_
timestamp 1701859473
transform -1 0 4470 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1213_
timestamp 1701859473
transform 1 0 4790 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1214_
timestamp 1701859473
transform 1 0 4930 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1215_
timestamp 1701859473
transform 1 0 5070 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1216_
timestamp 1701859473
transform 1 0 4790 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1217_
timestamp 1701859473
transform 1 0 4650 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1218_
timestamp 1701859473
transform 1 0 4930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1219_
timestamp 1701859473
transform -1 0 5250 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1220_
timestamp 1701859473
transform -1 0 5590 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1221_
timestamp 1701859473
transform -1 0 3510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1222_
timestamp 1701859473
transform 1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1223_
timestamp 1701859473
transform 1 0 3110 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1224_
timestamp 1701859473
transform -1 0 3410 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1225_
timestamp 1701859473
transform -1 0 3550 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1226_
timestamp 1701859473
transform -1 0 3550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1227_
timestamp 1701859473
transform -1 0 3450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1228_
timestamp 1701859473
transform 1 0 3270 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1229_
timestamp 1701859473
transform -1 0 3690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1230_
timestamp 1701859473
transform -1 0 3570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1231_
timestamp 1701859473
transform -1 0 3310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1232_
timestamp 1701859473
transform -1 0 4190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1233_
timestamp 1701859473
transform -1 0 4950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1234_
timestamp 1701859473
transform -1 0 4570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1235_
timestamp 1701859473
transform -1 0 4730 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1236_
timestamp 1701859473
transform 1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1237_
timestamp 1701859473
transform 1 0 4790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1238_
timestamp 1701859473
transform -1 0 4530 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1239_
timestamp 1701859473
transform -1 0 4710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1240_
timestamp 1701859473
transform 1 0 4970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1241_
timestamp 1701859473
transform 1 0 4030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1242_
timestamp 1701859473
transform 1 0 4890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1243_
timestamp 1701859473
transform -1 0 4590 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1244_
timestamp 1701859473
transform -1 0 4290 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1245_
timestamp 1701859473
transform 1 0 5410 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1246_
timestamp 1701859473
transform 1 0 5610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1247_
timestamp 1701859473
transform 1 0 4310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1248_
timestamp 1701859473
transform -1 0 4830 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1249_
timestamp 1701859473
transform 1 0 5370 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1250_
timestamp 1701859473
transform 1 0 5650 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1251_
timestamp 1701859473
transform 1 0 5370 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1252_
timestamp 1701859473
transform -1 0 5290 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1253_
timestamp 1701859473
transform 1 0 5330 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1254_
timestamp 1701859473
transform 1 0 5690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1255_
timestamp 1701859473
transform 1 0 5830 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1256_
timestamp 1701859473
transform -1 0 5930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1257_
timestamp 1701859473
transform 1 0 5510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1258_
timestamp 1701859473
transform 1 0 5510 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1259_
timestamp 1701859473
transform 1 0 5810 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1260_
timestamp 1701859473
transform 1 0 5230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1261_
timestamp 1701859473
transform 1 0 5330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1262_
timestamp 1701859473
transform -1 0 5870 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1263_
timestamp 1701859473
transform 1 0 5970 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1264_
timestamp 1701859473
transform -1 0 5570 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1265_
timestamp 1701859473
transform 1 0 5450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1266_
timestamp 1701859473
transform -1 0 5330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1267_
timestamp 1701859473
transform -1 0 5710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1268_
timestamp 1701859473
transform 1 0 5090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1269_
timestamp 1701859473
transform -1 0 5190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1270_
timestamp 1701859473
transform -1 0 3410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1271_
timestamp 1701859473
transform 1 0 2510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1272_
timestamp 1701859473
transform 1 0 1110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1273_
timestamp 1701859473
transform 1 0 1550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1274_
timestamp 1701859473
transform -1 0 2450 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1275_
timestamp 1701859473
transform -1 0 2590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1276_
timestamp 1701859473
transform -1 0 2170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1277_
timestamp 1701859473
transform 1 0 2290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1278_
timestamp 1701859473
transform 1 0 770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1279_
timestamp 1701859473
transform 1 0 630 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1280_
timestamp 1701859473
transform 1 0 1090 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1281_
timestamp 1701859473
transform -1 0 1650 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1282_
timestamp 1701859473
transform 1 0 1190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1283_
timestamp 1701859473
transform 1 0 1730 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1284_
timestamp 1701859473
transform 1 0 5410 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1285_
timestamp 1701859473
transform -1 0 5270 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1286_
timestamp 1701859473
transform -1 0 5450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1287_
timestamp 1701859473
transform -1 0 5550 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1288_
timestamp 1701859473
transform -1 0 5130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1289_
timestamp 1701859473
transform 1 0 4970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1290_
timestamp 1701859473
transform 1 0 4810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1291_
timestamp 1701859473
transform 1 0 5010 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1292_
timestamp 1701859473
transform -1 0 3830 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1293_
timestamp 1701859473
transform -1 0 3570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1294_
timestamp 1701859473
transform 1 0 4830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1295_
timestamp 1701859473
transform -1 0 4970 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1296_
timestamp 1701859473
transform 1 0 4630 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1297_
timestamp 1701859473
transform 1 0 4230 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1298_
timestamp 1701859473
transform 1 0 5130 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1299_
timestamp 1701859473
transform 1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1300_
timestamp 1701859473
transform 1 0 3690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1301_
timestamp 1701859473
transform -1 0 3970 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1302_
timestamp 1701859473
transform -1 0 3810 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1303_
timestamp 1701859473
transform -1 0 3930 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1304_
timestamp 1701859473
transform -1 0 3650 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1305_
timestamp 1701859473
transform 1 0 3670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1306_
timestamp 1701859473
transform 1 0 3550 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1307_
timestamp 1701859473
transform 1 0 4430 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1308_
timestamp 1701859473
transform -1 0 4150 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1309_
timestamp 1701859473
transform -1 0 3410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1310_
timestamp 1701859473
transform 1 0 2630 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1311_
timestamp 1701859473
transform 1 0 2890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1312_
timestamp 1701859473
transform 1 0 2390 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1313_
timestamp 1701859473
transform 1 0 2690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1314_
timestamp 1701859473
transform 1 0 2850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1315_
timestamp 1701859473
transform -1 0 2410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1316_
timestamp 1701859473
transform 1 0 2570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1317_
timestamp 1701859473
transform 1 0 3150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1318_
timestamp 1701859473
transform 1 0 2290 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1319_
timestamp 1701859473
transform 1 0 2530 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1320_
timestamp 1701859473
transform -1 0 2990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1321_
timestamp 1701859473
transform 1 0 2810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1322_
timestamp 1701859473
transform 1 0 3310 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1323_
timestamp 1701859473
transform 1 0 2670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1324_
timestamp 1701859473
transform -1 0 3130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1325_
timestamp 1701859473
transform -1 0 3290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1326_
timestamp 1701859473
transform -1 0 2970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1327_
timestamp 1701859473
transform 1 0 3870 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1328_
timestamp 1701859473
transform -1 0 4090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1329_
timestamp 1701859473
transform -1 0 4790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1330_
timestamp 1701859473
transform -1 0 4630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1331_
timestamp 1701859473
transform -1 0 3750 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1332_
timestamp 1701859473
transform 1 0 3790 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1333_
timestamp 1701859473
transform 1 0 3230 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1334_
timestamp 1701859473
transform -1 0 3890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1335_
timestamp 1701859473
transform 1 0 3950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1336_
timestamp 1701859473
transform 1 0 3770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1337_
timestamp 1701859473
transform 1 0 4070 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1338_
timestamp 1701859473
transform 1 0 5490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1339_
timestamp 1701859473
transform 1 0 5730 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1340_
timestamp 1701859473
transform 1 0 3610 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1341_
timestamp 1701859473
transform 1 0 3990 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1342_
timestamp 1701859473
transform -1 0 4390 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1343_
timestamp 1701859473
transform 1 0 4210 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1344_
timestamp 1701859473
transform -1 0 4370 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1345_
timestamp 1701859473
transform 1 0 4330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1346_
timestamp 1701859473
transform 1 0 4210 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1347_
timestamp 1701859473
transform 1 0 4490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1348_
timestamp 1701859473
transform 1 0 4490 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1349_
timestamp 1701859473
transform -1 0 4530 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1350_
timestamp 1701859473
transform -1 0 6010 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1351_
timestamp 1701859473
transform 1 0 5870 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1352_
timestamp 1701859473
transform -1 0 4110 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1353_
timestamp 1701859473
transform -1 0 3950 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1354_
timestamp 1701859473
transform -1 0 3650 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1355_
timestamp 1701859473
transform 1 0 3490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1356_
timestamp 1701859473
transform -1 0 2890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1357_
timestamp 1701859473
transform -1 0 2730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1358_
timestamp 1701859473
transform -1 0 2170 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1359_
timestamp 1701859473
transform -1 0 2930 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1360_
timestamp 1701859473
transform 1 0 1910 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1361_
timestamp 1701859473
transform -1 0 2770 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1362_
timestamp 1701859473
transform -1 0 2050 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1363_
timestamp 1701859473
transform -1 0 1270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1364_
timestamp 1701859473
transform 1 0 1210 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1365_
timestamp 1701859473
transform -1 0 530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1366_
timestamp 1701859473
transform -1 0 3490 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1367_
timestamp 1701859473
transform -1 0 4690 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1368_
timestamp 1701859473
transform -1 0 3370 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1369_
timestamp 1701859473
transform -1 0 2770 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1370_
timestamp 1701859473
transform -1 0 3090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1371_
timestamp 1701859473
transform 1 0 2390 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1372_
timestamp 1701859473
transform -1 0 3550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1373_
timestamp 1701859473
transform 1 0 3410 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1374_
timestamp 1701859473
transform -1 0 3370 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1375_
timestamp 1701859473
transform -1 0 3490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1376_
timestamp 1701859473
transform -1 0 3030 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1377_
timestamp 1701859473
transform -1 0 3050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1378_
timestamp 1701859473
transform -1 0 3170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1379_
timestamp 1701859473
transform 1 0 2750 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1380_
timestamp 1701859473
transform 1 0 3250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1381_
timestamp 1701859473
transform -1 0 3130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1382_
timestamp 1701859473
transform -1 0 2970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1383_
timestamp 1701859473
transform -1 0 3030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1384_
timestamp 1701859473
transform 1 0 3290 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1385_
timestamp 1701859473
transform 1 0 2890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1386_
timestamp 1701859473
transform 1 0 2610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1387_
timestamp 1701859473
transform -1 0 4250 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1388_
timestamp 1701859473
transform 1 0 2510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1389_
timestamp 1701859473
transform 1 0 2070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1390_
timestamp 1701859473
transform 1 0 1950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1391_
timestamp 1701859473
transform 1 0 2210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1392_
timestamp 1701859473
transform -1 0 2430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1393_
timestamp 1701859473
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1394_
timestamp 1701859473
transform 1 0 2330 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1395_
timestamp 1701859473
transform -1 0 3090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1396_
timestamp 1701859473
transform -1 0 2950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1397_
timestamp 1701859473
transform -1 0 2810 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1398_
timestamp 1701859473
transform 1 0 2650 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1399_
timestamp 1701859473
transform -1 0 2630 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1400_
timestamp 1701859473
transform 1 0 3230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1401_
timestamp 1701859473
transform -1 0 2390 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1402_
timestamp 1701859473
transform -1 0 2510 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1403_
timestamp 1701859473
transform -1 0 2330 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1404_
timestamp 1701859473
transform 1 0 2770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1405_
timestamp 1701859473
transform -1 0 3650 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1406_
timestamp 1701859473
transform -1 0 2790 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1407_
timestamp 1701859473
transform -1 0 2930 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1408_
timestamp 1701859473
transform 1 0 2490 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1409_
timestamp 1701859473
transform -1 0 2770 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1410_
timestamp 1701859473
transform -1 0 2930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1411_
timestamp 1701859473
transform 1 0 2910 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1412_
timestamp 1701859473
transform -1 0 2630 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1413_
timestamp 1701859473
transform 1 0 3050 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1414_
timestamp 1701859473
transform -1 0 3210 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1415_
timestamp 1701859473
transform -1 0 3210 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1416_
timestamp 1701859473
transform -1 0 3330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1417_
timestamp 1701859473
transform -1 0 3950 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1418_
timestamp 1701859473
transform -1 0 3790 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1419_
timestamp 1701859473
transform -1 0 3070 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1420_
timestamp 1701859473
transform 1 0 2010 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1421_
timestamp 1701859473
transform -1 0 2630 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1422_
timestamp 1701859473
transform -1 0 2830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1423_
timestamp 1701859473
transform -1 0 2690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1424_
timestamp 1701859473
transform -1 0 2570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1425_
timestamp 1701859473
transform -1 0 2510 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1426_
timestamp 1701859473
transform -1 0 2350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1427_
timestamp 1701859473
transform 1 0 370 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1428_
timestamp 1701859473
transform 1 0 770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1429_
timestamp 1701859473
transform -1 0 3730 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1430_
timestamp 1701859473
transform -1 0 3450 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1431_
timestamp 1701859473
transform 1 0 1050 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1432_
timestamp 1701859473
transform -1 0 1030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1433_
timestamp 1701859473
transform -1 0 1170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1434_
timestamp 1701859473
transform 1 0 170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1435_
timestamp 1701859473
transform -1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1436_
timestamp 1701859473
transform -1 0 190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1437_
timestamp 1701859473
transform 1 0 1870 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1438_
timestamp 1701859473
transform 1 0 2270 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1439_
timestamp 1701859473
transform 1 0 3130 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1440_
timestamp 1701859473
transform -1 0 1830 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1441_
timestamp 1701859473
transform -1 0 2170 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1442_
timestamp 1701859473
transform -1 0 1970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1443_
timestamp 1701859473
transform -1 0 1690 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1444_
timestamp 1701859473
transform -1 0 1570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1445_
timestamp 1701859473
transform 1 0 2070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1446_
timestamp 1701859473
transform 1 0 1810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1447_
timestamp 1701859473
transform 1 0 1670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1448_
timestamp 1701859473
transform 1 0 1410 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1449_
timestamp 1701859473
transform -1 0 1530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1450_
timestamp 1701859473
transform -1 0 1770 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1451_
timestamp 1701859473
transform 1 0 1590 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1452_
timestamp 1701859473
transform -1 0 2050 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1453_
timestamp 1701859473
transform 1 0 1330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1454_
timestamp 1701859473
transform -1 0 1830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1455_
timestamp 1701859473
transform 1 0 1690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1456_
timestamp 1701859473
transform 1 0 1810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1457_
timestamp 1701859473
transform -1 0 1910 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1458_
timestamp 1701859473
transform 1 0 1410 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1459_
timestamp 1701859473
transform -1 0 1290 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1460_
timestamp 1701859473
transform -1 0 1270 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1461_
timestamp 1701859473
transform 1 0 1370 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1462_
timestamp 1701859473
transform -1 0 2510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1463_
timestamp 1701859473
transform -1 0 1170 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1464_
timestamp 1701859473
transform 1 0 1510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1465_
timestamp 1701859473
transform 1 0 1670 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1466_
timestamp 1701859473
transform 1 0 1110 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1467_
timestamp 1701859473
transform 1 0 1570 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1468_
timestamp 1701859473
transform -1 0 1730 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1469_
timestamp 1701859473
transform 1 0 1910 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1470_
timestamp 1701859473
transform -1 0 2190 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1471_
timestamp 1701859473
transform -1 0 2490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1472_
timestamp 1701859473
transform -1 0 2350 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1473_
timestamp 1701859473
transform 1 0 2030 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1474_
timestamp 1701859473
transform -1 0 2150 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1475_
timestamp 1701859473
transform -1 0 2190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1476_
timestamp 1701859473
transform -1 0 2410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1477_
timestamp 1701859473
transform 1 0 1930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1478_
timestamp 1701859473
transform 1 0 2030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1479_
timestamp 1701859473
transform -1 0 2050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1480_
timestamp 1701859473
transform 1 0 4350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1481_
timestamp 1701859473
transform 1 0 4110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1482_
timestamp 1701859473
transform -1 0 4270 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1483_
timestamp 1701859473
transform -1 0 1330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1484_
timestamp 1701859473
transform 1 0 1170 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1485_
timestamp 1701859473
transform -1 0 910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1486_
timestamp 1701859473
transform 1 0 790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1487_
timestamp 1701859473
transform -1 0 330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1488_
timestamp 1701859473
transform -1 0 1290 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1489_
timestamp 1701859473
transform -1 0 70 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1490_
timestamp 1701859473
transform 1 0 1590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1491_
timestamp 1701859473
transform 1 0 2190 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1492_
timestamp 1701859473
transform -1 0 2070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1493_
timestamp 1701859473
transform 1 0 1890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1494_
timestamp 1701859473
transform -1 0 1770 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1495_
timestamp 1701859473
transform 1 0 1350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1496_
timestamp 1701859473
transform 1 0 1610 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1497_
timestamp 1701859473
transform 1 0 1530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1498_
timestamp 1701859473
transform -1 0 1690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1499_
timestamp 1701859473
transform -1 0 1490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1500_
timestamp 1701859473
transform 1 0 1470 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1501_
timestamp 1701859473
transform 1 0 1610 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1502_
timestamp 1701859473
transform -1 0 470 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1503_
timestamp 1701859473
transform 1 0 690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1504_
timestamp 1701859473
transform -1 0 450 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1505_
timestamp 1701859473
transform -1 0 330 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1506_
timestamp 1701859473
transform -1 0 970 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1507_
timestamp 1701859473
transform -1 0 830 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1508_
timestamp 1701859473
transform -1 0 750 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1509_
timestamp 1701859473
transform -1 0 890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1510_
timestamp 1701859473
transform 1 0 1010 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1511_
timestamp 1701859473
transform -1 0 610 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1512_
timestamp 1701859473
transform 1 0 750 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1513_
timestamp 1701859473
transform -1 0 3450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1514_
timestamp 1701859473
transform 1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1515_
timestamp 1701859473
transform -1 0 2210 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1516_
timestamp 1701859473
transform -1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1517_
timestamp 1701859473
transform 1 0 1790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1518_
timestamp 1701859473
transform -1 0 790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1519_
timestamp 1701859473
transform 1 0 1850 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1520_
timestamp 1701859473
transform -1 0 1990 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1521_
timestamp 1701859473
transform 1 0 1950 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1522_
timestamp 1701859473
transform -1 0 2250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1523_
timestamp 1701859473
transform 1 0 1050 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1524_
timestamp 1701859473
transform -1 0 350 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1525_
timestamp 1701859473
transform 1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1526_
timestamp 1701859473
transform 1 0 310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1527_
timestamp 1701859473
transform -1 0 4530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1528_
timestamp 1701859473
transform -1 0 4630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1529_
timestamp 1701859473
transform 1 0 4370 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1530_
timestamp 1701859473
transform 1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1531_
timestamp 1701859473
transform -1 0 910 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1532_
timestamp 1701859473
transform -1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1533_
timestamp 1701859473
transform 1 0 310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1534_
timestamp 1701859473
transform 1 0 330 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1535_
timestamp 1701859473
transform -1 0 1390 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1536_
timestamp 1701859473
transform -1 0 1490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1537_
timestamp 1701859473
transform -1 0 370 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1538_
timestamp 1701859473
transform -1 0 190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1539_
timestamp 1701859473
transform -1 0 1750 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1540_
timestamp 1701859473
transform 1 0 1230 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1541_
timestamp 1701859473
transform -1 0 1090 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1542_
timestamp 1701859473
transform -1 0 1390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1543_
timestamp 1701859473
transform -1 0 1110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1544_
timestamp 1701859473
transform -1 0 1450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1545_
timestamp 1701859473
transform -1 0 1090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1546_
timestamp 1701859473
transform 1 0 170 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1547_
timestamp 1701859473
transform 1 0 470 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1548_
timestamp 1701859473
transform -1 0 610 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1549_
timestamp 1701859473
transform 1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1550_
timestamp 1701859473
transform 1 0 610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1551_
timestamp 1701859473
transform -1 0 4510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1552_
timestamp 1701859473
transform -1 0 4690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1553_
timestamp 1701859473
transform 1 0 670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1554_
timestamp 1701859473
transform -1 0 1310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1555_
timestamp 1701859473
transform -1 0 1230 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1556_
timestamp 1701859473
transform 1 0 890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1557_
timestamp 1701859473
transform 1 0 50 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1558_
timestamp 1701859473
transform 1 0 890 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1559_
timestamp 1701859473
transform 1 0 1210 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1560_
timestamp 1701859473
transform -1 0 1330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1561_
timestamp 1701859473
transform -1 0 230 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1562_
timestamp 1701859473
transform 1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1563_
timestamp 1701859473
transform -1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1564_
timestamp 1701859473
transform -1 0 1170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1565_
timestamp 1701859473
transform -1 0 1290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1566_
timestamp 1701859473
transform -1 0 1410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1567_
timestamp 1701859473
transform -1 0 1250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1568_
timestamp 1701859473
transform -1 0 1250 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1569_
timestamp 1701859473
transform -1 0 1030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1570_
timestamp 1701859473
transform -1 0 950 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1571_
timestamp 1701859473
transform -1 0 750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1572_
timestamp 1701859473
transform 1 0 590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1573_
timestamp 1701859473
transform -1 0 450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1574_
timestamp 1701859473
transform -1 0 5150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1575_
timestamp 1701859473
transform 1 0 4990 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1576_
timestamp 1701859473
transform -1 0 4870 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1577_
timestamp 1701859473
transform -1 0 4710 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1578_
timestamp 1701859473
transform 1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1579_
timestamp 1701859473
transform 1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1580_
timestamp 1701859473
transform -1 0 250 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1581_
timestamp 1701859473
transform 1 0 150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1582_
timestamp 1701859473
transform 1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1583_
timestamp 1701859473
transform -1 0 870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1584_
timestamp 1701859473
transform -1 0 970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1585_
timestamp 1701859473
transform -1 0 670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1586_
timestamp 1701859473
transform -1 0 530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1587_
timestamp 1701859473
transform -1 0 4890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1588_
timestamp 1701859473
transform -1 0 4710 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1589_
timestamp 1701859473
transform -1 0 1510 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1590_
timestamp 1701859473
transform -1 0 1210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1591_
timestamp 1701859473
transform -1 0 1070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1592_
timestamp 1701859473
transform 1 0 150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1593_
timestamp 1701859473
transform 1 0 2550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1594_
timestamp 1701859473
transform -1 0 2690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1595_
timestamp 1701859473
transform 1 0 3630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1596_
timestamp 1701859473
transform 1 0 3470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1597_
timestamp 1701859473
transform -1 0 2490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1598_
timestamp 1701859473
transform 1 0 2310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1599_
timestamp 1701859473
transform -1 0 3750 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1600_
timestamp 1701859473
transform 1 0 3570 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1601_
timestamp 1701859473
transform 1 0 3270 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1602_
timestamp 1701859473
transform 1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1603_
timestamp 1701859473
transform -1 0 2890 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1604_
timestamp 1701859473
transform 1 0 2710 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1605_
timestamp 1701859473
transform 1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1606_
timestamp 1701859473
transform 1 0 1890 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1607_
timestamp 1701859473
transform -1 0 1730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1608_
timestamp 1701859473
transform 1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1636_
timestamp 1701859473
transform -1 0 4250 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1637_
timestamp 1701859473
transform -1 0 4350 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1638_
timestamp 1701859473
transform -1 0 4110 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1639_
timestamp 1701859473
transform 1 0 3950 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1640_
timestamp 1701859473
transform -1 0 3710 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1641_
timestamp 1701859473
transform -1 0 3650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1642_
timestamp 1701859473
transform -1 0 3210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1643_
timestamp 1701859473
transform -1 0 4110 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1644_
timestamp 1701859473
transform -1 0 4090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1645_
timestamp 1701859473
transform 1 0 4490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1646_
timestamp 1701859473
transform -1 0 4230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1647_
timestamp 1701859473
transform 1 0 3310 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1648_
timestamp 1701859473
transform -1 0 4230 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1649_
timestamp 1701859473
transform -1 0 3830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1650_
timestamp 1701859473
transform -1 0 3950 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1651_
timestamp 1701859473
transform 1 0 3670 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1652_
timestamp 1701859473
transform 1 0 3670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1653_
timestamp 1701859473
transform 1 0 3790 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1654_
timestamp 1701859473
transform -1 0 4630 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1655_
timestamp 1701859473
transform -1 0 4490 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1656_
timestamp 1701859473
transform 1 0 1470 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1657_
timestamp 1701859473
transform 1 0 3110 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1658_
timestamp 1701859473
transform 1 0 3250 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1659_
timestamp 1701859473
transform -1 0 3210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1660_
timestamp 1701859473
transform 1 0 3550 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1661_
timestamp 1701859473
transform -1 0 3430 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1662_
timestamp 1701859473
transform 1 0 3550 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1663_
timestamp 1701859473
transform -1 0 3510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1664_
timestamp 1701859473
transform -1 0 3350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1665_
timestamp 1701859473
transform -1 0 3990 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1666_
timestamp 1701859473
transform 1 0 3850 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1667_
timestamp 1701859473
transform -1 0 3710 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1668_
timestamp 1701859473
transform 1 0 3410 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1669_
timestamp 1701859473
transform -1 0 3530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1670_
timestamp 1701859473
transform -1 0 3390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1671_
timestamp 1701859473
transform -1 0 3090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1672_
timestamp 1701859473
transform 1 0 2750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1673_
timestamp 1701859473
transform -1 0 2910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1674_
timestamp 1701859473
transform 1 0 2990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1675_
timestamp 1701859473
transform -1 0 4410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1676_
timestamp 1701859473
transform 1 0 4130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1677_
timestamp 1701859473
transform 1 0 3810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1678_
timestamp 1701859473
transform 1 0 4330 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1679_
timestamp 1701859473
transform 1 0 4610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1680_
timestamp 1701859473
transform -1 0 4510 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1681_
timestamp 1701859473
transform 1 0 3910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1682_
timestamp 1701859473
transform 1 0 4090 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1683_
timestamp 1701859473
transform 1 0 3970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1684_
timestamp 1701859473
transform 1 0 3790 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1685_
timestamp 1701859473
transform -1 0 2850 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1686_
timestamp 1701859473
transform -1 0 2570 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1687_
timestamp 1701859473
transform 1 0 2430 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1688_
timestamp 1701859473
transform -1 0 2170 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1689_
timestamp 1701859473
transform -1 0 1670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1690_
timestamp 1701859473
transform 1 0 2690 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1691_
timestamp 1701859473
transform -1 0 2310 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1692_
timestamp 1701859473
transform -1 0 3010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1693_
timestamp 1701859473
transform 1 0 3170 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1694_
timestamp 1701859473
transform 1 0 3170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1695_
timestamp 1701859473
transform -1 0 3590 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1696_
timestamp 1701859473
transform 1 0 3430 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1697_
timestamp 1701859473
transform -1 0 3310 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1698_
timestamp 1701859473
transform -1 0 3150 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1699_
timestamp 1701859473
transform -1 0 2450 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1700_
timestamp 1701859473
transform 1 0 2270 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1701_
timestamp 1701859473
transform -1 0 2230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1702_
timestamp 1701859473
transform 1 0 2050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1703_
timestamp 1701859473
transform 1 0 1290 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1704_
timestamp 1701859473
transform -1 0 1250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1705_
timestamp 1701859473
transform 1 0 2350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1706_
timestamp 1701859473
transform -1 0 2470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1707_
timestamp 1701859473
transform 1 0 1910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1708_
timestamp 1701859473
transform -1 0 1890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1709_
timestamp 1701859473
transform -1 0 2650 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1710_
timestamp 1701859473
transform -1 0 3050 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1711_
timestamp 1701859473
transform 1 0 2890 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1712_
timestamp 1701859473
transform 1 0 2430 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1713_
timestamp 1701859473
transform -1 0 2750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1714_
timestamp 1701859473
transform -1 0 2610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1715_
timestamp 1701859473
transform 1 0 2710 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1716_
timestamp 1701859473
transform 1 0 2570 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1717_
timestamp 1701859473
transform -1 0 2610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1718_
timestamp 1701859473
transform -1 0 2470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1719_
timestamp 1701859473
transform 1 0 2070 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1720_
timestamp 1701859473
transform 1 0 1890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1721_
timestamp 1701859473
transform 1 0 1610 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1722_
timestamp 1701859473
transform -1 0 2030 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1723_
timestamp 1701859473
transform 1 0 1750 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1724_
timestamp 1701859473
transform 1 0 1210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1725_
timestamp 1701859473
transform 1 0 1990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1726_
timestamp 1701859473
transform -1 0 910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1727_
timestamp 1701859473
transform -1 0 1010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1728_
timestamp 1701859473
transform 1 0 2630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1729_
timestamp 1701859473
transform 1 0 1910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1730_
timestamp 1701859473
transform -1 0 2230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1731_
timestamp 1701859473
transform -1 0 2270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1732_
timestamp 1701859473
transform 1 0 2070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1733_
timestamp 1701859473
transform 1 0 2110 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1734_
timestamp 1701859473
transform -1 0 1770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1735_
timestamp 1701859473
transform -1 0 1830 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1736_
timestamp 1701859473
transform 1 0 1650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1737_
timestamp 1701859473
transform -1 0 1530 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1738_
timestamp 1701859473
transform -1 0 1150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1739_
timestamp 1701859473
transform -1 0 950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1740_
timestamp 1701859473
transform -1 0 1270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1741_
timestamp 1701859473
transform -1 0 1010 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1742_
timestamp 1701859473
transform -1 0 2330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1743_
timestamp 1701859473
transform -1 0 3070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1744_
timestamp 1701859473
transform 1 0 2750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1745_
timestamp 1701859473
transform 1 0 2470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1746_
timestamp 1701859473
transform -1 0 2910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1747_
timestamp 1701859473
transform -1 0 2350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1748_
timestamp 1701859473
transform -1 0 1510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1749_
timestamp 1701859473
transform -1 0 1370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1750_
timestamp 1701859473
transform -1 0 850 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1751_
timestamp 1701859473
transform -1 0 810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1752_
timestamp 1701859473
transform -1 0 430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1753_
timestamp 1701859473
transform 1 0 330 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1754_
timestamp 1701859473
transform -1 0 550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1755_
timestamp 1701859473
transform -1 0 650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1756_
timestamp 1701859473
transform -1 0 1290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1757_
timestamp 1701859473
transform 1 0 1950 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1758_
timestamp 1701859473
transform -1 0 2170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1759_
timestamp 1701859473
transform -1 0 2290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1760_
timestamp 1701859473
transform -1 0 1870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1761_
timestamp 1701859473
transform 1 0 1670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1762_
timestamp 1701859473
transform -1 0 1510 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1763_
timestamp 1701859473
transform -1 0 1350 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1764_
timestamp 1701859473
transform -1 0 910 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1765_
timestamp 1701859473
transform -1 0 750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1766_
timestamp 1701859473
transform -1 0 630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1767_
timestamp 1701859473
transform 1 0 1150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1768_
timestamp 1701859473
transform 1 0 1370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1769_
timestamp 1701859473
transform -1 0 1530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1770_
timestamp 1701859473
transform -1 0 1390 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1771_
timestamp 1701859473
transform -1 0 690 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1772_
timestamp 1701859473
transform -1 0 530 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1773_
timestamp 1701859473
transform 1 0 770 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1774_
timestamp 1701859473
transform 1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1775_
timestamp 1701859473
transform 1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1776_
timestamp 1701859473
transform -1 0 490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1777_
timestamp 1701859473
transform -1 0 3710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1778_
timestamp 1701859473
transform 1 0 2750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1779_
timestamp 1701859473
transform -1 0 3070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1780_
timestamp 1701859473
transform -1 0 3530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1781_
timestamp 1701859473
transform 1 0 2910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1782_
timestamp 1701859473
transform 1 0 3350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1783_
timestamp 1701859473
transform -1 0 1510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1784_
timestamp 1701859473
transform -1 0 1350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1785_
timestamp 1701859473
transform -1 0 1170 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1786_
timestamp 1701859473
transform -1 0 1010 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1787_
timestamp 1701859473
transform -1 0 570 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1788_
timestamp 1701859473
transform 1 0 630 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1789_
timestamp 1701859473
transform -1 0 630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1790_
timestamp 1701859473
transform -1 0 470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1791_
timestamp 1701859473
transform -1 0 350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1792_
timestamp 1701859473
transform -1 0 1770 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1793_
timestamp 1701859473
transform 1 0 1630 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1794_
timestamp 1701859473
transform 1 0 630 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1795_
timestamp 1701859473
transform -1 0 210 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1796_
timestamp 1701859473
transform 1 0 270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1797_
timestamp 1701859473
transform 1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1798_
timestamp 1701859473
transform -1 0 690 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1799_
timestamp 1701859473
transform 1 0 430 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1800_
timestamp 1701859473
transform 1 0 210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1801_
timestamp 1701859473
transform -1 0 230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1802_
timestamp 1701859473
transform -1 0 2890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1803_
timestamp 1701859473
transform 1 0 830 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1804_
timestamp 1701859473
transform -1 0 730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1805_
timestamp 1701859473
transform 1 0 830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1806_
timestamp 1701859473
transform 1 0 1030 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1807_
timestamp 1701859473
transform -1 0 70 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1808_
timestamp 1701859473
transform -1 0 510 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1809_
timestamp 1701859473
transform -1 0 1190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1810_
timestamp 1701859473
transform -1 0 1010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1811_
timestamp 1701859473
transform -1 0 190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1812_
timestamp 1701859473
transform -1 0 350 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1813_
timestamp 1701859473
transform -1 0 70 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1814_
timestamp 1701859473
transform -1 0 70 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1815_
timestamp 1701859473
transform -1 0 350 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1816_
timestamp 1701859473
transform 1 0 50 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1817_
timestamp 1701859473
transform -1 0 210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1818_
timestamp 1701859473
transform -1 0 70 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1819_
timestamp 1701859473
transform -1 0 190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1820_
timestamp 1701859473
transform -1 0 70 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1821_
timestamp 1701859473
transform 1 0 550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1822_
timestamp 1701859473
transform -1 0 330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1823_
timestamp 1701859473
transform -1 0 210 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1824_
timestamp 1701859473
transform 1 0 50 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1825_
timestamp 1701859473
transform 1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1826_
timestamp 1701859473
transform 1 0 1090 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1701859473
transform -1 0 2810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1701859473
transform 1 0 3410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1701859473
transform 1 0 3470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1701859473
transform -1 0 2850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1701859473
transform -1 0 4570 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert5
timestamp 1701859473
transform 1 0 4570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1701859473
transform 1 0 4610 0 1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert7
timestamp 1701859473
transform 1 0 4750 0 1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert13
timestamp 1701859473
transform 1 0 3150 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert14
timestamp 1701859473
transform 1 0 2710 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert15
timestamp 1701859473
transform -1 0 2010 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1701859473
transform -1 0 1870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1701859473
transform 1 0 450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1701859473
transform 1 0 3330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1701859473
transform 1 0 1830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1701859473
transform 1 0 1450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1701859473
transform -1 0 70 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1701859473
transform -1 0 2770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1701859473
transform 1 0 3530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1701859473
transform 1 0 3850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1701859473
transform -1 0 3030 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1701859473
transform 1 0 2990 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert27
timestamp 1701859473
transform 1 0 2570 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1701859473
transform -1 0 1510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1701859473
transform 1 0 2570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert30
timestamp 1701859473
transform -1 0 2470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1701859473
transform 1 0 2930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1701859473
transform 1 0 1990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert33
timestamp 1701859473
transform 1 0 3330 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert34
timestamp 1701859473
transform -1 0 3610 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert35
timestamp 1701859473
transform -1 0 3990 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert36
timestamp 1701859473
transform 1 0 3990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert37
timestamp 1701859473
transform -1 0 3830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert38
timestamp 1701859473
transform 1 0 1750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert39
timestamp 1701859473
transform -1 0 4530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert40
timestamp 1701859473
transform -1 0 1650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert41
timestamp 1701859473
transform -1 0 2630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert8
timestamp 1701859473
transform 1 0 2190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1701859473
transform 1 0 1470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 1970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1701859473
transform 1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__890_
timestamp 1701859473
transform 1 0 670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__892_
timestamp 1701859473
transform 1 0 830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__894_
timestamp 1701859473
transform 1 0 1090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__896_
timestamp 1701859473
transform -1 0 1750 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__898_
timestamp 1701859473
transform -1 0 1490 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__900_
timestamp 1701859473
transform -1 0 410 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__902_
timestamp 1701859473
transform 1 0 210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__904_
timestamp 1701859473
transform -1 0 690 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__906_
timestamp 1701859473
transform -1 0 970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__909_
timestamp 1701859473
transform -1 0 850 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__911_
timestamp 1701859473
transform 1 0 450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__913_
timestamp 1701859473
transform 1 0 230 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__915_
timestamp 1701859473
transform 1 0 1430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__917_
timestamp 1701859473
transform 1 0 670 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__919_
timestamp 1701859473
transform 1 0 810 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__921_
timestamp 1701859473
transform -1 0 1250 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__923_
timestamp 1701859473
transform -1 0 1170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__925_
timestamp 1701859473
transform 1 0 70 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__927_
timestamp 1701859473
transform -1 0 3110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__930_
timestamp 1701859473
transform -1 0 3930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__932_
timestamp 1701859473
transform 1 0 2190 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__934_
timestamp 1701859473
transform -1 0 2190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__936_
timestamp 1701859473
transform -1 0 3630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__938_
timestamp 1701859473
transform 1 0 2970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__940_
timestamp 1701859473
transform -1 0 2870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__942_
timestamp 1701859473
transform -1 0 2630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__944_
timestamp 1701859473
transform 1 0 1450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__946_
timestamp 1701859473
transform -1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__948_
timestamp 1701859473
transform -1 0 1750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__950_
timestamp 1701859473
transform -1 0 90 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__953_
timestamp 1701859473
transform 1 0 4230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__955_
timestamp 1701859473
transform 1 0 4370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__957_
timestamp 1701859473
transform 1 0 4670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__959_
timestamp 1701859473
transform -1 0 5230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__961_
timestamp 1701859473
transform -1 0 5090 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__963_
timestamp 1701859473
transform 1 0 6070 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__965_
timestamp 1701859473
transform 1 0 5250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__967_
timestamp 1701859473
transform 1 0 4890 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__969_
timestamp 1701859473
transform 1 0 5430 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__971_
timestamp 1701859473
transform -1 0 6070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__973_
timestamp 1701859473
transform -1 0 5790 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__976_
timestamp 1701859473
transform -1 0 4450 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__978_
timestamp 1701859473
transform -1 0 4450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__980_
timestamp 1701859473
transform 1 0 4810 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__982_
timestamp 1701859473
transform 1 0 5730 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__984_
timestamp 1701859473
transform 1 0 4950 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__986_
timestamp 1701859473
transform 1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__988_
timestamp 1701859473
transform -1 0 5310 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__990_
timestamp 1701859473
transform 1 0 6010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__992_
timestamp 1701859473
transform -1 0 5130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__994_
timestamp 1701859473
transform -1 0 6070 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__996_
timestamp 1701859473
transform 1 0 5390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__999_
timestamp 1701859473
transform 1 0 4050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1001_
timestamp 1701859473
transform 1 0 3850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1004_
timestamp 1701859473
transform 1 0 4390 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1006_
timestamp 1701859473
transform -1 0 4450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1008_
timestamp 1701859473
transform 1 0 4010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1010_
timestamp 1701859473
transform -1 0 5870 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1012_
timestamp 1701859473
transform 1 0 5430 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1014_
timestamp 1701859473
transform 1 0 6150 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1016_
timestamp 1701859473
transform 1 0 5570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1018_
timestamp 1701859473
transform 1 0 4950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1020_
timestamp 1701859473
transform 1 0 6030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1022_
timestamp 1701859473
transform -1 0 4850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1024_
timestamp 1701859473
transform -1 0 2150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1027_
timestamp 1701859473
transform 1 0 5410 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1029_
timestamp 1701859473
transform 1 0 5090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1031_
timestamp 1701859473
transform -1 0 4410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1033_
timestamp 1701859473
transform 1 0 5830 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1035_
timestamp 1701859473
transform -1 0 5530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1037_
timestamp 1701859473
transform 1 0 6110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1039_
timestamp 1701859473
transform -1 0 3930 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1041_
timestamp 1701859473
transform 1 0 4510 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1043_
timestamp 1701859473
transform 1 0 4290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1045_
timestamp 1701859473
transform 1 0 4350 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1047_
timestamp 1701859473
transform 1 0 4110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1050_
timestamp 1701859473
transform 1 0 5250 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1052_
timestamp 1701859473
transform -1 0 5970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1054_
timestamp 1701859473
transform -1 0 5130 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1056_
timestamp 1701859473
transform -1 0 6150 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1058_
timestamp 1701859473
transform 1 0 5830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1060_
timestamp 1701859473
transform -1 0 6130 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1062_
timestamp 1701859473
transform 1 0 4170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1064_
timestamp 1701859473
transform 1 0 5330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1066_
timestamp 1701859473
transform -1 0 5690 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1068_
timestamp 1701859473
transform -1 0 6010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1070_
timestamp 1701859473
transform -1 0 5310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1073_
timestamp 1701859473
transform 1 0 5530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1075_
timestamp 1701859473
transform 1 0 5690 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1077_
timestamp 1701859473
transform -1 0 4550 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1079_
timestamp 1701859473
transform -1 0 4050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1081_
timestamp 1701859473
transform 1 0 5190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1083_
timestamp 1701859473
transform -1 0 4870 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1085_
timestamp 1701859473
transform 1 0 6010 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1087_
timestamp 1701859473
transform 1 0 5090 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1089_
timestamp 1701859473
transform -1 0 4090 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1091_
timestamp 1701859473
transform 1 0 3630 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1094_
timestamp 1701859473
transform 1 0 3850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1096_
timestamp 1701859473
transform 1 0 4410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1098_
timestamp 1701859473
transform 1 0 3990 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1100_
timestamp 1701859473
transform 1 0 5470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1102_
timestamp 1701859473
transform 1 0 5250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1104_
timestamp 1701859473
transform -1 0 5870 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1106_
timestamp 1701859473
transform 1 0 5790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1108_
timestamp 1701859473
transform 1 0 5990 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1110_
timestamp 1701859473
transform -1 0 6110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1112_
timestamp 1701859473
transform -1 0 3730 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1114_
timestamp 1701859473
transform 1 0 4030 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1117_
timestamp 1701859473
transform 1 0 3690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1119_
timestamp 1701859473
transform -1 0 4470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1121_
timestamp 1701859473
transform -1 0 4230 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1123_
timestamp 1701859473
transform 1 0 4390 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1125_
timestamp 1701859473
transform -1 0 5950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1127_
timestamp 1701859473
transform 1 0 4910 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1129_
timestamp 1701859473
transform 1 0 5190 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1131_
timestamp 1701859473
transform -1 0 5750 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1133_
timestamp 1701859473
transform -1 0 5650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1135_
timestamp 1701859473
transform -1 0 5790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1137_
timestamp 1701859473
transform -1 0 5630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1140_
timestamp 1701859473
transform -1 0 5290 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1142_
timestamp 1701859473
transform 1 0 5010 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1144_
timestamp 1701859473
transform -1 0 5390 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1146_
timestamp 1701859473
transform 1 0 5350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1148_
timestamp 1701859473
transform -1 0 5810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1150_
timestamp 1701859473
transform 1 0 4970 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1152_
timestamp 1701859473
transform 1 0 5890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1154_
timestamp 1701859473
transform -1 0 5770 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1156_
timestamp 1701859473
transform 1 0 5130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1158_
timestamp 1701859473
transform -1 0 5750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1160_
timestamp 1701859473
transform -1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1163_
timestamp 1701859473
transform -1 0 5750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1165_
timestamp 1701859473
transform -1 0 4110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1167_
timestamp 1701859473
transform -1 0 4370 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1169_
timestamp 1701859473
transform 1 0 4490 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1171_
timestamp 1701859473
transform 1 0 5150 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1173_
timestamp 1701859473
transform 1 0 5310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1175_
timestamp 1701859473
transform 1 0 5570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1177_
timestamp 1701859473
transform 1 0 5290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1179_
timestamp 1701859473
transform -1 0 4810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1181_
timestamp 1701859473
transform -1 0 5030 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1183_
timestamp 1701859473
transform -1 0 4670 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1186_
timestamp 1701859473
transform -1 0 3870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1188_
timestamp 1701859473
transform -1 0 3330 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1190_
timestamp 1701859473
transform -1 0 3950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1192_
timestamp 1701859473
transform 1 0 4010 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1194_
timestamp 1701859473
transform -1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1196_
timestamp 1701859473
transform -1 0 5150 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1198_
timestamp 1701859473
transform -1 0 5290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1200_
timestamp 1701859473
transform -1 0 4990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1202_
timestamp 1701859473
transform 1 0 4710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1204_
timestamp 1701859473
transform -1 0 4870 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1206_
timestamp 1701859473
transform -1 0 5590 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1209_
timestamp 1701859473
transform 1 0 4110 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1211_
timestamp 1701859473
transform -1 0 4510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1213_
timestamp 1701859473
transform 1 0 4810 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1215_
timestamp 1701859473
transform 1 0 5090 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1217_
timestamp 1701859473
transform 1 0 4670 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1219_
timestamp 1701859473
transform -1 0 5270 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1221_
timestamp 1701859473
transform -1 0 3530 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1223_
timestamp 1701859473
transform 1 0 3130 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1225_
timestamp 1701859473
transform -1 0 3570 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1227_
timestamp 1701859473
transform -1 0 3470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1230_
timestamp 1701859473
transform -1 0 3590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1232_
timestamp 1701859473
transform -1 0 4210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1234_
timestamp 1701859473
transform -1 0 4590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1236_
timestamp 1701859473
transform 1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1238_
timestamp 1701859473
transform -1 0 4550 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1240_
timestamp 1701859473
transform 1 0 4990 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1242_
timestamp 1701859473
transform 1 0 4910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1244_
timestamp 1701859473
transform -1 0 4310 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1246_
timestamp 1701859473
transform 1 0 5630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1248_
timestamp 1701859473
transform -1 0 4850 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1250_
timestamp 1701859473
transform 1 0 5670 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1253_
timestamp 1701859473
transform 1 0 5350 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1255_
timestamp 1701859473
transform 1 0 5850 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1257_
timestamp 1701859473
transform 1 0 5530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1259_
timestamp 1701859473
transform 1 0 5830 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1261_
timestamp 1701859473
transform 1 0 5350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1263_
timestamp 1701859473
transform 1 0 5990 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1265_
timestamp 1701859473
transform 1 0 5470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1267_
timestamp 1701859473
transform -1 0 5730 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1269_
timestamp 1701859473
transform -1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1271_
timestamp 1701859473
transform 1 0 2530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1273_
timestamp 1701859473
transform 1 0 1570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1276_
timestamp 1701859473
transform -1 0 2190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1278_
timestamp 1701859473
transform 1 0 790 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1280_
timestamp 1701859473
transform 1 0 1110 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1282_
timestamp 1701859473
transform 1 0 1210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1284_
timestamp 1701859473
transform 1 0 5430 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1286_
timestamp 1701859473
transform -1 0 5470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1288_
timestamp 1701859473
transform -1 0 5150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1290_
timestamp 1701859473
transform 1 0 4830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1292_
timestamp 1701859473
transform -1 0 3850 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1294_
timestamp 1701859473
transform 1 0 4850 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1296_
timestamp 1701859473
transform 1 0 4650 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1299_
timestamp 1701859473
transform 1 0 5190 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1301_
timestamp 1701859473
transform -1 0 3990 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1303_
timestamp 1701859473
transform -1 0 3950 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1305_
timestamp 1701859473
transform 1 0 3690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1307_
timestamp 1701859473
transform 1 0 4450 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1309_
timestamp 1701859473
transform -1 0 3430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1311_
timestamp 1701859473
transform 1 0 2910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1313_
timestamp 1701859473
transform 1 0 2710 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1315_
timestamp 1701859473
transform -1 0 2430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1317_
timestamp 1701859473
transform 1 0 3170 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1319_
timestamp 1701859473
transform 1 0 2550 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1322_
timestamp 1701859473
transform 1 0 3330 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1324_
timestamp 1701859473
transform -1 0 3150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1326_
timestamp 1701859473
transform -1 0 2990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1328_
timestamp 1701859473
transform -1 0 4110 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1330_
timestamp 1701859473
transform -1 0 4650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1332_
timestamp 1701859473
transform 1 0 3810 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1334_
timestamp 1701859473
transform -1 0 3910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1336_
timestamp 1701859473
transform 1 0 3790 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1338_
timestamp 1701859473
transform 1 0 5510 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1340_
timestamp 1701859473
transform 1 0 3630 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1343_
timestamp 1701859473
transform 1 0 4230 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1345_
timestamp 1701859473
transform 1 0 4350 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1347_
timestamp 1701859473
transform 1 0 4510 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1349_
timestamp 1701859473
transform -1 0 4550 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1351_
timestamp 1701859473
transform 1 0 5890 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1353_
timestamp 1701859473
transform -1 0 3970 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1355_
timestamp 1701859473
transform 1 0 3510 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1357_
timestamp 1701859473
transform -1 0 2750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1359_
timestamp 1701859473
transform -1 0 2950 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1361_
timestamp 1701859473
transform -1 0 2790 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1363_
timestamp 1701859473
transform -1 0 1290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1366_
timestamp 1701859473
transform -1 0 3510 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1368_
timestamp 1701859473
transform -1 0 3390 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1370_
timestamp 1701859473
transform -1 0 3110 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1372_
timestamp 1701859473
transform -1 0 3570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1374_
timestamp 1701859473
transform -1 0 3390 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1376_
timestamp 1701859473
transform -1 0 3050 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1378_
timestamp 1701859473
transform -1 0 3190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1380_
timestamp 1701859473
transform 1 0 3270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1382_
timestamp 1701859473
transform -1 0 2990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1384_
timestamp 1701859473
transform 1 0 3310 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1386_
timestamp 1701859473
transform 1 0 2630 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1389_
timestamp 1701859473
transform 1 0 2090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1391_
timestamp 1701859473
transform 1 0 2230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1393_
timestamp 1701859473
transform 1 0 2270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1395_
timestamp 1701859473
transform -1 0 3110 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1397_
timestamp 1701859473
transform -1 0 2830 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1399_
timestamp 1701859473
transform -1 0 2650 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1401_
timestamp 1701859473
transform -1 0 2410 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1403_
timestamp 1701859473
transform -1 0 2350 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1405_
timestamp 1701859473
transform -1 0 3670 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1407_
timestamp 1701859473
transform -1 0 2950 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1409_
timestamp 1701859473
transform -1 0 2790 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1412_
timestamp 1701859473
transform -1 0 2650 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1414_
timestamp 1701859473
transform -1 0 3230 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1416_
timestamp 1701859473
transform -1 0 3350 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1418_
timestamp 1701859473
transform -1 0 3810 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1420_
timestamp 1701859473
transform 1 0 2030 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1422_
timestamp 1701859473
transform -1 0 2850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1424_
timestamp 1701859473
transform -1 0 2590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1426_
timestamp 1701859473
transform -1 0 2370 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1428_
timestamp 1701859473
transform 1 0 790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1430_
timestamp 1701859473
transform -1 0 3470 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1432_
timestamp 1701859473
transform -1 0 1050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1435_
timestamp 1701859473
transform -1 0 550 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1437_
timestamp 1701859473
transform 1 0 1890 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1439_
timestamp 1701859473
transform 1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1441_
timestamp 1701859473
transform -1 0 2190 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1443_
timestamp 1701859473
transform -1 0 1710 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1445_
timestamp 1701859473
transform 1 0 2090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1447_
timestamp 1701859473
transform 1 0 1690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1449_
timestamp 1701859473
transform -1 0 1550 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1451_
timestamp 1701859473
transform 1 0 1610 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1453_
timestamp 1701859473
transform 1 0 1350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1455_
timestamp 1701859473
transform 1 0 1710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1458_
timestamp 1701859473
transform 1 0 1430 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1460_
timestamp 1701859473
transform -1 0 1290 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1462_
timestamp 1701859473
transform -1 0 2530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1464_
timestamp 1701859473
transform 1 0 1530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1466_
timestamp 1701859473
transform 1 0 1130 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1468_
timestamp 1701859473
transform -1 0 1750 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1470_
timestamp 1701859473
transform -1 0 2210 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1472_
timestamp 1701859473
transform -1 0 2370 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1474_
timestamp 1701859473
transform -1 0 2170 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1476_
timestamp 1701859473
transform -1 0 2430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1479_
timestamp 1701859473
transform -1 0 2070 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1481_
timestamp 1701859473
transform 1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1483_
timestamp 1701859473
transform -1 0 1350 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1485_
timestamp 1701859473
transform -1 0 930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1487_
timestamp 1701859473
transform -1 0 350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1489_
timestamp 1701859473
transform -1 0 90 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1491_
timestamp 1701859473
transform 1 0 2210 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1493_
timestamp 1701859473
transform 1 0 1910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1495_
timestamp 1701859473
transform 1 0 1370 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1497_
timestamp 1701859473
transform 1 0 1550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1499_
timestamp 1701859473
transform -1 0 1510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1502_
timestamp 1701859473
transform -1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1504_
timestamp 1701859473
transform -1 0 470 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1506_
timestamp 1701859473
transform -1 0 990 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1508_
timestamp 1701859473
transform -1 0 770 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1510_
timestamp 1701859473
transform 1 0 1030 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1512_
timestamp 1701859473
transform 1 0 770 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1514_
timestamp 1701859473
transform 1 0 2110 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1516_
timestamp 1701859473
transform -1 0 1910 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1518_
timestamp 1701859473
transform -1 0 810 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1520_
timestamp 1701859473
transform -1 0 2010 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1522_
timestamp 1701859473
transform -1 0 2270 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1525_
timestamp 1701859473
transform 1 0 70 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1527_
timestamp 1701859473
transform -1 0 4550 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1529_
timestamp 1701859473
transform 1 0 4390 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1531_
timestamp 1701859473
transform -1 0 930 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1533_
timestamp 1701859473
transform 1 0 330 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1535_
timestamp 1701859473
transform -1 0 1410 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1537_
timestamp 1701859473
transform -1 0 390 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1539_
timestamp 1701859473
transform -1 0 1770 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1541_
timestamp 1701859473
transform -1 0 1110 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1543_
timestamp 1701859473
transform -1 0 1130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1545_
timestamp 1701859473
transform -1 0 1110 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1548_
timestamp 1701859473
transform -1 0 630 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1550_
timestamp 1701859473
transform 1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1552_
timestamp 1701859473
transform -1 0 4710 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1554_
timestamp 1701859473
transform -1 0 1330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1556_
timestamp 1701859473
transform 1 0 910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1558_
timestamp 1701859473
transform 1 0 910 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1560_
timestamp 1701859473
transform -1 0 1350 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1562_
timestamp 1701859473
transform 1 0 70 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1564_
timestamp 1701859473
transform -1 0 1190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1566_
timestamp 1701859473
transform -1 0 1430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1568_
timestamp 1701859473
transform -1 0 1270 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1571_
timestamp 1701859473
transform -1 0 770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1573_
timestamp 1701859473
transform -1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1575_
timestamp 1701859473
transform 1 0 5010 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1577_
timestamp 1701859473
transform -1 0 4730 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1579_
timestamp 1701859473
transform 1 0 70 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1581_
timestamp 1701859473
transform 1 0 170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1583_
timestamp 1701859473
transform -1 0 890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1585_
timestamp 1701859473
transform -1 0 690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1587_
timestamp 1701859473
transform -1 0 4910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1589_
timestamp 1701859473
transform -1 0 1530 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1592_
timestamp 1701859473
transform 1 0 170 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1594_
timestamp 1701859473
transform -1 0 2710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1596_
timestamp 1701859473
transform 1 0 3490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1598_
timestamp 1701859473
transform 1 0 2330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1600_
timestamp 1701859473
transform 1 0 3590 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1602_
timestamp 1701859473
transform 1 0 2870 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1604_
timestamp 1701859473
transform 1 0 2730 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1606_
timestamp 1701859473
transform 1 0 1910 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1608_
timestamp 1701859473
transform 1 0 1570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1637_
timestamp 1701859473
transform -1 0 4370 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1639_
timestamp 1701859473
transform 1 0 3970 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1642_
timestamp 1701859473
transform -1 0 3230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1644_
timestamp 1701859473
transform -1 0 4110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1646_
timestamp 1701859473
transform -1 0 4250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1648_
timestamp 1701859473
transform -1 0 4250 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1650_
timestamp 1701859473
transform -1 0 3970 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1652_
timestamp 1701859473
transform 1 0 3690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1654_
timestamp 1701859473
transform -1 0 4650 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1656_
timestamp 1701859473
transform 1 0 1490 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1658_
timestamp 1701859473
transform 1 0 3270 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1660_
timestamp 1701859473
transform 1 0 3570 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1662_
timestamp 1701859473
transform 1 0 3570 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1665_
timestamp 1701859473
transform -1 0 4010 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1667_
timestamp 1701859473
transform -1 0 3730 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1669_
timestamp 1701859473
transform -1 0 3550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1671_
timestamp 1701859473
transform -1 0 3110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1673_
timestamp 1701859473
transform -1 0 2930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1675_
timestamp 1701859473
transform -1 0 4430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1677_
timestamp 1701859473
transform 1 0 3830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1679_
timestamp 1701859473
transform 1 0 4630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1681_
timestamp 1701859473
transform 1 0 3930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1683_
timestamp 1701859473
transform 1 0 3990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1685_
timestamp 1701859473
transform -1 0 2870 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1688_
timestamp 1701859473
transform -1 0 2190 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1690_
timestamp 1701859473
transform 1 0 2710 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1692_
timestamp 1701859473
transform -1 0 3030 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1694_
timestamp 1701859473
transform 1 0 3190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1696_
timestamp 1701859473
transform 1 0 3450 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1698_
timestamp 1701859473
transform -1 0 3170 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1700_
timestamp 1701859473
transform 1 0 2290 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1702_
timestamp 1701859473
transform 1 0 2070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1704_
timestamp 1701859473
transform -1 0 1270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1706_
timestamp 1701859473
transform -1 0 2490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1708_
timestamp 1701859473
transform -1 0 1910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1711_
timestamp 1701859473
transform 1 0 2910 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1713_
timestamp 1701859473
transform -1 0 2770 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1715_
timestamp 1701859473
transform 1 0 2730 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1717_
timestamp 1701859473
transform -1 0 2630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1719_
timestamp 1701859473
transform 1 0 2090 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1721_
timestamp 1701859473
transform 1 0 1630 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1723_
timestamp 1701859473
transform 1 0 1770 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1725_
timestamp 1701859473
transform 1 0 2010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1727_
timestamp 1701859473
transform -1 0 1030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1729_
timestamp 1701859473
transform 1 0 1930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1731_
timestamp 1701859473
transform -1 0 2290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1734_
timestamp 1701859473
transform -1 0 1790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1736_
timestamp 1701859473
transform 1 0 1670 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1738_
timestamp 1701859473
transform -1 0 1170 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1740_
timestamp 1701859473
transform -1 0 1290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1742_
timestamp 1701859473
transform -1 0 2350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1744_
timestamp 1701859473
transform 1 0 2770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1746_
timestamp 1701859473
transform -1 0 2930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1748_
timestamp 1701859473
transform -1 0 1530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1750_
timestamp 1701859473
transform -1 0 870 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1752_
timestamp 1701859473
transform -1 0 450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1755_
timestamp 1701859473
transform -1 0 670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1757_
timestamp 1701859473
transform 1 0 1970 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1759_
timestamp 1701859473
transform -1 0 2310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1761_
timestamp 1701859473
transform 1 0 1690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1763_
timestamp 1701859473
transform -1 0 1370 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1765_
timestamp 1701859473
transform -1 0 770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1767_
timestamp 1701859473
transform 1 0 1170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1769_
timestamp 1701859473
transform -1 0 1550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1771_
timestamp 1701859473
transform -1 0 710 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1773_
timestamp 1701859473
transform 1 0 790 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1775_
timestamp 1701859473
transform 1 0 70 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1778_
timestamp 1701859473
transform 1 0 2770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1780_
timestamp 1701859473
transform -1 0 3550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1782_
timestamp 1701859473
transform 1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1784_
timestamp 1701859473
transform -1 0 1370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1786_
timestamp 1701859473
transform -1 0 1030 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1788_
timestamp 1701859473
transform 1 0 650 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1790_
timestamp 1701859473
transform -1 0 490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1792_
timestamp 1701859473
transform -1 0 1790 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1794_
timestamp 1701859473
transform 1 0 650 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1796_
timestamp 1701859473
transform 1 0 290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1798_
timestamp 1701859473
transform -1 0 710 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1801_
timestamp 1701859473
transform -1 0 250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1803_
timestamp 1701859473
transform 1 0 850 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1805_
timestamp 1701859473
transform 1 0 850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1807_
timestamp 1701859473
transform -1 0 90 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1809_
timestamp 1701859473
transform -1 0 1210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1811_
timestamp 1701859473
transform -1 0 210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1813_
timestamp 1701859473
transform -1 0 90 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1815_
timestamp 1701859473
transform -1 0 370 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1817_
timestamp 1701859473
transform -1 0 230 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1819_
timestamp 1701859473
transform -1 0 210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1821_
timestamp 1701859473
transform 1 0 570 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1824_
timestamp 1701859473
transform 1 0 70 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1826_
timestamp 1701859473
transform 1 0 1110 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert0
timestamp 1701859473
transform -1 0 2830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert2
timestamp 1701859473
transform 1 0 3490 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert4
timestamp 1701859473
transform -1 0 4590 0 1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert6
timestamp 1701859473
transform 1 0 4630 0 1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert14
timestamp 1701859473
transform 1 0 2730 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert16
timestamp 1701859473
transform -1 0 1890 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert18
timestamp 1701859473
transform 1 0 3350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert21
timestamp 1701859473
transform -1 0 90 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert23
timestamp 1701859473
transform 1 0 3550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert25
timestamp 1701859473
transform -1 0 3050 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert27
timestamp 1701859473
transform 1 0 2590 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert29
timestamp 1701859473
transform 1 0 2590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert31
timestamp 1701859473
transform 1 0 2950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert33
timestamp 1701859473
transform 1 0 3350 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert35
timestamp 1701859473
transform -1 0 4010 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert37
timestamp 1701859473
transform -1 0 3850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert39
timestamp 1701859473
transform -1 0 4550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert41
timestamp 1701859473
transform -1 0 2650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert8
timestamp 1701859473
transform 1 0 2210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 70 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert12
timestamp 1701859473
transform 1 0 70 0 -1 2350
box -12 -8 32 272
<< labels >>
flabel metal1 s 6243 2 6303 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 977 6297 983 6303 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 3977 6297 3983 6303 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 537 6297 543 6303 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal2 s 57 -23 63 -17 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 137 -23 143 -17 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 217 -23 223 -17 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 337 -23 343 -17 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 637 -23 643 -17 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal2 s 1137 -23 1143 -17 7 FreeSans 16 270 0 0 Done_o
port 18 nsew
rlabel metal2 4616 6296 4623 6303 0 ABCmd_i[2]
port 7 nsew
flabel metal2 s 4417 6297 4423 6303 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal2 s 4117 6297 4123 6303 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 1877 6297 1883 6303 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
rlabel metal3 -63 4648 -55 4656 0 LoadA_i
port 19 nsew
rlabel metal3 -63 4496 -55 4504 0 LoadB_i
port 20 nsew
flabel metal3 s -63 3976 -55 3984 7 FreeSans 16 0 0 0 reset
port 23 nsew
flabel metal3 s -63 3776 -55 3784 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -63 2736 -55 2744 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal3 s -63 2678 -55 2686 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal3 s -63 2476 -55 2484 7 FreeSans 16 0 0 0 clk
port 22 nsew
flabel metal3 s 6295 5416 6303 5424 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
rlabel metal2 4356 6295 4363 6302 0 ABCmd_i[0]
port 9 nsew
<< properties >>
string FIXED_BBOX -40 -40 6280 6300
<< end >>
