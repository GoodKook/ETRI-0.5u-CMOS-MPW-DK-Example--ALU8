VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_wrapper
  CLASS BLOCK ;
  FOREIGN ALU_wrapper ;
  ORIGIN 6.000 0.000 ;
  SIZE 960.000 BY 945.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 948.450 899.700 957.450 938.700 ;
        RECT 0.600 897.300 957.450 899.700 ;
        RECT 948.450 821.700 957.450 897.300 ;
        RECT 0.600 819.300 957.450 821.700 ;
        RECT 948.450 743.700 957.450 819.300 ;
        RECT 0.600 741.300 957.450 743.700 ;
        RECT 948.450 665.700 957.450 741.300 ;
        RECT 0.600 663.300 957.450 665.700 ;
        RECT 948.450 587.700 957.450 663.300 ;
        RECT 0.600 585.300 957.450 587.700 ;
        RECT 948.450 509.700 957.450 585.300 ;
        RECT 0.600 507.300 957.450 509.700 ;
        RECT 948.450 431.700 957.450 507.300 ;
        RECT 0.600 429.300 957.450 431.700 ;
        RECT 948.450 353.700 957.450 429.300 ;
        RECT 0.600 351.300 957.450 353.700 ;
        RECT 948.450 275.700 957.450 351.300 ;
        RECT 0.600 273.300 957.450 275.700 ;
        RECT 948.450 197.700 957.450 273.300 ;
        RECT 0.600 195.300 957.450 197.700 ;
        RECT 948.450 119.700 957.450 195.300 ;
        RECT 0.600 117.300 957.450 119.700 ;
        RECT 948.450 41.700 957.450 117.300 ;
        RECT 0.600 39.300 957.450 41.700 ;
        RECT 948.450 0.300 957.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 397.950 938.700 400.050 940.050 ;
        RECT 487.950 938.700 490.050 940.050 ;
        RECT 514.950 938.700 517.050 940.050 ;
        RECT 604.950 938.700 607.050 940.050 ;
        RECT 769.950 938.700 772.050 940.050 ;
        RECT -9.450 936.300 947.400 938.700 ;
        RECT -9.450 860.700 -0.450 936.300 ;
        RECT -9.450 858.300 947.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT 514.950 856.950 517.050 858.300 ;
        RECT 595.950 856.950 598.050 858.300 ;
        RECT 724.950 856.950 727.050 858.300 ;
        RECT 913.950 856.950 916.050 858.300 ;
        RECT -9.450 780.300 947.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 436.950 778.950 439.050 780.300 ;
        RECT 673.950 778.950 676.050 780.300 ;
        RECT 823.950 778.950 826.050 780.300 ;
        RECT 844.950 778.950 847.050 780.300 ;
        RECT -9.450 702.300 947.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 388.950 700.950 391.050 702.300 ;
        RECT 499.950 700.950 502.050 702.300 ;
        RECT 547.950 700.950 550.050 702.300 ;
        RECT 493.950 626.700 496.500 628.050 ;
        RECT -9.450 624.300 947.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 376.950 622.950 379.050 624.300 ;
        RECT 415.950 622.950 418.050 624.300 ;
        RECT 580.950 622.950 583.050 624.300 ;
        RECT 583.950 622.950 586.050 624.300 ;
        RECT 670.950 622.950 673.050 624.300 ;
        RECT 709.950 621.450 712.050 622.050 ;
        RECT 716.550 621.450 717.450 624.300 ;
        RECT 709.950 620.550 717.450 621.450 ;
        RECT 709.950 619.950 712.050 620.550 ;
        RECT -9.450 546.300 947.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT -9.450 468.300 947.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 370.950 466.950 373.050 468.300 ;
        RECT 434.550 466.050 435.450 468.300 ;
        RECT 493.950 466.950 496.050 468.300 ;
        RECT 430.950 464.550 435.450 466.050 ;
        RECT 430.950 463.950 435.000 464.550 ;
        RECT -9.450 390.300 947.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT -9.450 312.300 947.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT -9.450 234.300 947.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT -9.450 156.300 947.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT -9.450 78.300 947.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 947.400 2.700 ;
      LAYER metal2 ;
        RECT 397.950 937.950 400.050 940.050 ;
        RECT 487.950 937.950 490.050 940.050 ;
        RECT 514.950 937.950 517.050 940.050 ;
        RECT 604.950 937.950 607.050 940.050 ;
        RECT 769.950 937.950 772.050 940.050 ;
        RECT 398.400 915.450 399.450 937.950 ;
        RECT 401.400 915.450 402.600 916.650 ;
        RECT 398.400 914.400 402.600 915.450 ;
        RECT 488.400 915.450 489.450 937.950 ;
        RECT 491.400 915.450 492.600 916.650 ;
        RECT 488.400 914.400 492.600 915.450 ;
        RECT 512.400 915.450 513.600 916.650 ;
        RECT 515.400 915.450 516.450 937.950 ;
        RECT 512.400 914.400 516.450 915.450 ;
        RECT 602.400 915.450 603.600 916.650 ;
        RECT 605.400 915.450 606.450 937.950 ;
        RECT 602.400 914.400 606.450 915.450 ;
        RECT 770.400 915.450 771.450 937.950 ;
        RECT 773.400 915.450 774.600 916.650 ;
        RECT 770.400 914.400 774.600 915.450 ;
        RECT 689.400 875.400 690.600 877.650 ;
        RECT 689.400 859.050 690.450 875.400 ;
        RECT 502.950 856.950 505.050 859.050 ;
        RECT 511.950 856.950 517.050 859.050 ;
        RECT 595.950 856.950 598.050 859.050 ;
        RECT 688.950 856.950 691.050 859.050 ;
        RECT 724.950 856.950 730.050 859.050 ;
        RECT 913.950 856.950 916.050 859.050 ;
        RECT 503.400 816.450 504.450 856.950 ;
        RECT 596.400 838.050 597.450 856.950 ;
        RECT 595.950 835.950 598.050 838.050 ;
        RECT 635.400 837.900 636.600 838.650 ;
        RECT 836.400 837.900 837.600 838.650 ;
        RECT 914.400 838.050 915.450 856.950 ;
        RECT 634.950 835.800 637.050 837.900 ;
        RECT 835.950 835.800 838.050 837.900 ;
        RECT 913.950 835.950 916.050 838.050 ;
        RECT 500.400 815.400 504.450 816.450 ;
        RECT 500.400 804.600 501.450 815.400 ;
        RECT 500.400 802.350 501.600 804.600 ;
        RECT 821.400 804.450 822.600 804.600 ;
        RECT 818.400 803.400 822.600 804.450 ;
        RECT 818.400 793.050 819.450 803.400 ;
        RECT 821.400 802.350 822.600 803.400 ;
        RECT 842.400 804.450 843.600 804.600 ;
        RECT 842.400 803.400 846.450 804.450 ;
        RECT 842.400 802.350 843.600 803.400 ;
        RECT 817.950 790.950 820.050 793.050 ;
        RECT 823.950 790.950 826.050 793.050 ;
        RECT 824.400 781.050 825.450 790.950 ;
        RECT 845.400 781.050 846.450 803.400 ;
        RECT 436.950 778.950 439.050 781.050 ;
        RECT 673.950 778.950 676.050 781.050 ;
        RECT 823.950 778.950 826.050 781.050 ;
        RECT 844.950 778.950 847.050 781.050 ;
        RECT 437.400 763.050 438.450 778.950 ;
        RECT 436.800 760.950 438.900 763.050 ;
        RECT 464.400 759.900 465.600 760.650 ;
        RECT 463.950 757.800 466.050 759.900 ;
        RECT 581.400 758.400 582.600 760.650 ;
        RECT 499.950 709.950 502.050 712.050 ;
        RECT 511.950 709.950 514.050 712.050 ;
        RECT 500.400 703.050 501.450 709.950 ;
        RECT 388.950 700.950 391.050 703.050 ;
        RECT 499.950 700.950 502.050 703.050 ;
        RECT 377.400 680.400 378.600 682.650 ;
        RECT 377.400 673.050 378.450 680.400 ;
        RECT 389.400 673.050 390.450 700.950 ;
        RECT 440.400 681.000 441.600 682.650 ;
        RECT 512.400 682.050 513.450 709.950 ;
        RECT 581.400 706.050 582.450 758.400 ;
        RECT 674.400 726.600 675.450 778.950 ;
        RECT 674.400 724.350 675.600 726.600 ;
        RECT 547.950 700.950 550.050 706.050 ;
        RECT 580.950 703.950 583.050 706.050 ;
        RECT 439.950 676.950 442.050 681.000 ;
        RECT 511.950 679.950 514.050 682.050 ;
        RECT 674.400 680.400 675.600 682.650 ;
        RECT 695.400 680.400 696.600 682.650 ;
        RECT 376.950 670.950 379.050 673.050 ;
        RECT 388.950 670.950 391.050 673.050 ;
        RECT 674.400 658.050 675.450 680.400 ;
        RECT 695.400 658.050 696.450 680.400 ;
        RECT 664.950 655.950 667.050 658.050 ;
        RECT 673.950 655.950 676.050 658.050 ;
        RECT 694.950 655.950 697.050 658.050 ;
        RECT 709.950 655.950 712.050 658.050 ;
        RECT 412.950 647.100 415.050 649.200 ;
        RECT 584.400 648.450 585.600 648.600 ;
        RECT 581.400 647.400 585.600 648.450 ;
        RECT 413.400 646.350 414.600 647.100 ;
        RECT 415.800 640.950 417.900 643.050 ;
        RECT 416.400 625.050 417.450 640.950 ;
        RECT 493.950 625.950 496.050 628.050 ;
        RECT 376.950 622.950 379.050 625.050 ;
        RECT 415.950 622.950 418.050 625.050 ;
        RECT 377.400 598.050 378.450 622.950 ;
        RECT 494.400 603.450 495.450 625.950 ;
        RECT 581.400 625.050 582.450 647.400 ;
        RECT 584.400 646.350 585.600 647.400 ;
        RECT 665.400 625.050 666.450 655.950 ;
        RECT 580.950 622.950 583.050 625.050 ;
        RECT 583.950 622.950 586.050 625.050 ;
        RECT 664.950 622.950 667.050 625.050 ;
        RECT 670.950 622.950 673.050 628.050 ;
        RECT 497.400 603.450 498.600 604.650 ;
        RECT 566.400 603.900 567.600 604.650 ;
        RECT 584.400 604.050 585.450 622.950 ;
        RECT 710.400 622.050 711.450 655.950 ;
        RECT 709.950 619.950 712.050 622.050 ;
        RECT 494.400 602.400 498.600 603.450 ;
        RECT 376.950 595.950 379.050 598.050 ;
        RECT 388.950 595.950 391.050 598.050 ;
        RECT 389.400 570.600 390.450 595.950 ;
        RECT 494.400 589.050 495.450 602.400 ;
        RECT 565.950 601.800 568.050 603.900 ;
        RECT 583.950 601.950 586.050 604.050 ;
        RECT 475.950 586.950 478.050 589.050 ;
        RECT 493.950 586.950 496.050 589.050 ;
        RECT 476.400 570.600 477.450 586.950 ;
        RECT 389.400 568.350 390.600 570.600 ;
        RECT 476.400 568.350 477.600 570.600 ;
        RECT 389.400 524.400 390.600 526.650 ;
        RECT 431.400 524.400 432.600 526.650 ;
        RECT 500.400 524.400 501.600 526.650 ;
        RECT 389.400 499.050 390.450 524.400 ;
        RECT 361.950 496.950 364.050 499.050 ;
        RECT 388.950 496.950 391.050 499.050 ;
        RECT 362.400 484.050 363.450 496.950 ;
        RECT 361.950 481.950 364.050 484.050 ;
        RECT 370.950 481.800 373.050 483.900 ;
        RECT 371.400 469.050 372.450 481.800 ;
        RECT 370.950 466.950 373.050 469.050 ;
        RECT 431.400 466.050 432.450 524.400 ;
        RECT 500.400 495.450 501.450 524.400 ;
        RECT 500.400 494.400 504.450 495.450 ;
        RECT 503.400 469.050 504.450 494.400 ;
        RECT 493.950 466.950 499.050 469.050 ;
        RECT 502.950 466.950 505.050 469.050 ;
        RECT 430.950 463.950 433.050 466.050 ;
      LAYER metal3 ;
        RECT 502.950 858.600 505.050 859.050 ;
        RECT 511.950 858.600 514.050 859.050 ;
        RECT 502.950 857.400 514.050 858.600 ;
        RECT 502.950 856.950 505.050 857.400 ;
        RECT 511.950 856.950 514.050 857.400 ;
        RECT 688.950 858.600 691.050 859.050 ;
        RECT 727.950 858.600 730.050 859.050 ;
        RECT 688.950 857.400 730.050 858.600 ;
        RECT 688.950 856.950 691.050 857.400 ;
        RECT 727.950 856.950 730.050 857.400 ;
        RECT 595.950 837.600 598.050 838.050 ;
        RECT 634.950 837.600 637.050 837.900 ;
        RECT 595.950 836.400 637.050 837.600 ;
        RECT 595.950 835.950 598.050 836.400 ;
        RECT 634.950 835.800 637.050 836.400 ;
        RECT 835.950 837.600 838.050 837.900 ;
        RECT 913.950 837.600 916.050 838.050 ;
        RECT 835.950 836.400 916.050 837.600 ;
        RECT 835.950 835.800 838.050 836.400 ;
        RECT 913.950 835.950 916.050 836.400 ;
        RECT 817.950 792.600 820.050 793.050 ;
        RECT 823.950 792.600 826.050 793.050 ;
        RECT 817.950 791.400 826.050 792.600 ;
        RECT 817.950 790.950 820.050 791.400 ;
        RECT 823.950 790.950 826.050 791.400 ;
        RECT 436.800 762.000 438.900 763.050 ;
        RECT 436.800 760.950 439.050 762.000 ;
        RECT 436.950 759.600 439.050 760.950 ;
        RECT 463.950 759.600 466.050 759.900 ;
        RECT 436.950 759.000 466.050 759.600 ;
        RECT 437.250 758.400 466.050 759.000 ;
        RECT 463.950 757.800 466.050 758.400 ;
        RECT 499.950 711.600 502.050 712.050 ;
        RECT 511.950 711.600 514.050 712.050 ;
        RECT 499.950 710.400 514.050 711.600 ;
        RECT 499.950 709.950 502.050 710.400 ;
        RECT 511.950 709.950 514.050 710.400 ;
        RECT 547.950 705.600 550.050 706.050 ;
        RECT 580.950 705.600 583.050 706.050 ;
        RECT 547.950 704.400 583.050 705.600 ;
        RECT 547.950 703.950 550.050 704.400 ;
        RECT 580.950 703.950 583.050 704.400 ;
        RECT 511.950 681.600 514.050 682.050 ;
        RECT 503.400 680.400 514.050 681.600 ;
        RECT 439.950 678.600 442.050 679.050 ;
        RECT 503.400 678.600 504.600 680.400 ;
        RECT 511.950 679.950 514.050 680.400 ;
        RECT 439.950 677.400 504.600 678.600 ;
        RECT 439.950 676.950 442.050 677.400 ;
        RECT 376.950 672.600 379.050 673.050 ;
        RECT 388.950 672.600 391.050 673.050 ;
        RECT 376.950 671.400 391.050 672.600 ;
        RECT 376.950 670.950 379.050 671.400 ;
        RECT 388.950 670.950 391.050 671.400 ;
        RECT 664.950 657.600 667.050 658.050 ;
        RECT 673.950 657.600 676.050 658.050 ;
        RECT 664.950 656.400 676.050 657.600 ;
        RECT 664.950 655.950 667.050 656.400 ;
        RECT 673.950 655.950 676.050 656.400 ;
        RECT 694.950 657.600 697.050 658.050 ;
        RECT 709.950 657.600 712.050 658.050 ;
        RECT 694.950 656.400 712.050 657.600 ;
        RECT 694.950 655.950 697.050 656.400 ;
        RECT 709.950 655.950 712.050 656.400 ;
        RECT 412.950 648.600 415.050 649.200 ;
        RECT 412.950 647.400 417.450 648.600 ;
        RECT 412.950 647.100 415.050 647.400 ;
        RECT 416.250 643.050 417.450 647.400 ;
        RECT 415.800 640.950 417.900 643.050 ;
        RECT 664.950 624.600 667.050 625.050 ;
        RECT 670.950 624.600 673.050 628.050 ;
        RECT 664.950 624.000 673.050 624.600 ;
        RECT 664.950 623.400 672.600 624.000 ;
        RECT 664.950 622.950 667.050 623.400 ;
        RECT 565.950 603.600 568.050 603.900 ;
        RECT 583.950 603.600 586.050 604.050 ;
        RECT 565.950 602.400 586.050 603.600 ;
        RECT 565.950 601.800 568.050 602.400 ;
        RECT 583.950 601.950 586.050 602.400 ;
        RECT 376.950 597.600 379.050 598.050 ;
        RECT 388.950 597.600 391.050 598.050 ;
        RECT 376.950 596.400 391.050 597.600 ;
        RECT 376.950 595.950 379.050 596.400 ;
        RECT 388.950 595.950 391.050 596.400 ;
        RECT 475.950 588.600 478.050 589.050 ;
        RECT 493.950 588.600 496.050 589.050 ;
        RECT 475.950 587.400 496.050 588.600 ;
        RECT 475.950 586.950 478.050 587.400 ;
        RECT 493.950 586.950 496.050 587.400 ;
        RECT 361.950 498.600 364.050 499.050 ;
        RECT 388.950 498.600 391.050 499.050 ;
        RECT 361.950 497.400 391.050 498.600 ;
        RECT 361.950 496.950 364.050 497.400 ;
        RECT 388.950 496.950 391.050 497.400 ;
        RECT 361.950 483.600 364.050 484.050 ;
        RECT 370.950 483.600 373.050 483.900 ;
        RECT 361.950 482.400 373.050 483.600 ;
        RECT 361.950 481.950 364.050 482.400 ;
        RECT 370.950 481.800 373.050 482.400 ;
        RECT 496.950 468.600 499.050 469.050 ;
        RECT 502.950 468.600 505.050 469.050 ;
        RECT 496.950 467.400 505.050 468.600 ;
        RECT 496.950 466.950 499.050 467.400 ;
        RECT 502.950 466.950 505.050 467.400 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal1 ;
        RECT 346.950 831.450 349.050 832.050 ;
        RECT 355.950 831.450 358.050 831.900 ;
        RECT 346.950 830.550 358.050 831.450 ;
        RECT 346.950 829.950 349.050 830.550 ;
        RECT 355.950 829.800 358.050 830.550 ;
        RECT 394.950 825.450 397.050 829.050 ;
        RECT 400.950 825.450 403.050 826.050 ;
        RECT 394.950 825.000 403.050 825.450 ;
        RECT 395.550 824.550 403.050 825.000 ;
        RECT 400.950 823.950 403.050 824.550 ;
        RECT 886.950 765.450 889.050 766.050 ;
        RECT 901.950 765.450 904.050 766.050 ;
        RECT 886.950 764.550 904.050 765.450 ;
        RECT 886.950 763.950 889.050 764.550 ;
        RECT 901.950 763.950 904.050 764.550 ;
        RECT 358.950 759.450 363.000 760.050 ;
        RECT 358.950 757.950 363.450 759.450 ;
        RECT 362.550 757.050 363.450 757.950 ;
        RECT 362.550 755.550 367.050 757.050 ;
        RECT 363.000 754.950 367.050 755.550 ;
        RECT 685.950 714.450 688.050 715.050 ;
        RECT 691.950 714.450 694.050 715.050 ;
        RECT 685.950 713.550 694.050 714.450 ;
        RECT 685.950 712.950 688.050 713.550 ;
        RECT 691.950 712.950 694.050 713.550 ;
      LAYER metal2 ;
        RECT 293.400 918.450 294.450 945.450 ;
        RECT 295.950 918.450 298.050 919.200 ;
        RECT 293.400 917.400 298.050 918.450 ;
        RECT 295.950 917.100 298.050 917.400 ;
        RECT 310.950 917.100 313.050 919.200 ;
        RECT 296.400 916.350 297.600 917.100 ;
        RECT 311.400 895.050 312.450 917.100 ;
        RECT 301.950 892.950 304.050 895.050 ;
        RECT 310.950 892.950 313.050 895.050 ;
        RECT 328.950 892.950 331.050 895.050 ;
        RECT 302.400 885.600 303.450 892.950 ;
        RECT 302.400 883.350 303.600 885.600 ;
        RECT 329.400 841.050 330.450 892.950 ;
        RECT 328.950 838.950 331.050 841.050 ;
        RECT 347.400 834.900 348.600 835.650 ;
        RECT 346.800 834.000 348.900 834.900 ;
        RECT 346.800 832.800 349.050 834.000 ;
        RECT 346.950 829.950 349.050 832.800 ;
        RECT 355.950 829.800 358.050 831.900 ;
        RECT 356.400 826.050 357.450 829.800 ;
        RECT 355.950 823.950 358.050 826.050 ;
        RECT 388.950 823.950 391.050 826.050 ;
        RECT 394.950 823.950 397.050 829.050 ;
        RECT 400.950 823.950 403.050 826.050 ;
        RECT 389.400 778.050 390.450 823.950 ;
        RECT 401.400 807.600 402.450 823.950 ;
        RECT 401.400 805.350 402.600 807.600 ;
        RECT 358.950 775.950 361.050 778.050 ;
        RECT 388.950 775.950 391.050 778.050 ;
        RECT 359.400 760.050 360.450 775.950 ;
        RECT 811.950 769.950 814.050 772.050 ;
        RECT 886.950 769.950 889.050 772.050 ;
        RECT 812.400 766.050 813.450 769.950 ;
        RECT 887.400 766.050 888.450 769.950 ;
        RECT 811.950 763.950 814.050 766.050 ;
        RECT 886.950 763.950 889.050 766.050 ;
        RECT 787.950 761.100 790.050 763.200 ;
        RECT 788.400 760.350 789.600 761.100 ;
        RECT 793.950 760.800 796.050 762.900 ;
        RECT 901.950 762.000 904.050 766.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 368.400 757.050 369.600 757.650 ;
        RECT 364.950 755.400 369.600 757.050 ;
        RECT 364.950 754.950 369.000 755.400 ;
        RECT 365.400 735.450 366.450 754.950 ;
        RECT 794.400 751.050 795.450 760.800 ;
        RECT 902.400 760.350 903.600 762.000 ;
        RECT 739.950 748.950 742.050 751.050 ;
        RECT 793.950 748.950 796.050 751.050 ;
        RECT 362.400 734.400 366.450 735.450 ;
        RECT 362.400 730.050 363.450 734.400 ;
        RECT 379.950 733.950 382.050 736.050 ;
        RECT 427.950 733.950 430.050 736.050 ;
        RECT 361.950 727.950 364.050 730.050 ;
        RECT 368.400 723.900 369.600 724.650 ;
        RECT 367.950 721.800 370.050 723.900 ;
        RECT 368.400 712.050 369.450 721.800 ;
        RECT 380.400 712.050 381.450 733.950 ;
        RECT 367.950 709.950 370.050 712.050 ;
        RECT 379.950 709.950 382.050 712.050 ;
        RECT 428.400 703.050 429.450 733.950 ;
        RECT 587.400 722.400 588.600 724.650 ;
        RECT 587.400 715.050 588.450 722.400 ;
        RECT 740.400 715.050 741.450 748.950 ;
        RECT 586.950 712.950 589.050 715.050 ;
        RECT 682.950 712.950 688.050 715.050 ;
        RECT 691.950 712.950 697.050 715.050 ;
        RECT 739.950 712.950 742.050 715.050 ;
        RECT 757.950 712.950 760.050 715.050 ;
        RECT 427.950 700.950 430.050 703.050 ;
        RECT 436.950 700.950 439.050 703.050 ;
        RECT 437.400 691.050 438.450 700.950 ;
        RECT 587.400 697.050 588.450 712.950 ;
        RECT 526.950 694.950 529.050 697.050 ;
        RECT 586.950 694.950 589.050 697.050 ;
        RECT 527.400 691.050 528.450 694.950 ;
        RECT 436.950 688.950 439.050 691.050 ;
        RECT 526.950 688.950 529.050 691.050 ;
        RECT 758.400 625.050 759.450 712.950 ;
        RECT 757.950 622.950 760.050 625.050 ;
        RECT 808.950 619.950 811.050 622.050 ;
        RECT 886.950 619.950 889.050 622.050 ;
        RECT 809.400 573.450 810.450 619.950 ;
        RECT 887.400 606.600 888.450 619.950 ;
        RECT 887.400 604.350 888.600 606.600 ;
        RECT 806.400 572.400 810.450 573.450 ;
        RECT 806.400 565.050 807.450 572.400 ;
        RECT 875.400 567.000 876.600 568.650 ;
        RECT 805.950 562.950 808.050 565.050 ;
        RECT 874.950 562.950 877.050 567.000 ;
        RECT 806.400 547.050 807.450 562.950 ;
        RECT 538.950 544.950 541.050 547.050 ;
        RECT 805.950 544.950 808.050 547.050 ;
        RECT 539.400 538.050 540.450 544.950 ;
        RECT 806.400 538.050 807.450 544.950 ;
        RECT 481.950 535.950 484.050 538.050 ;
        RECT 538.950 535.950 541.050 538.050 ;
        RECT 799.950 535.950 802.050 538.050 ;
        RECT 805.950 535.950 808.050 538.050 ;
        RECT 482.400 532.050 483.450 535.950 ;
        RECT 469.950 529.950 472.050 532.050 ;
        RECT 481.950 529.950 484.050 532.050 ;
        RECT 470.400 511.050 471.450 529.950 ;
        RECT 800.400 528.600 801.450 535.950 ;
        RECT 800.400 526.350 801.600 528.600 ;
        RECT 424.950 508.950 427.050 511.050 ;
        RECT 469.950 508.950 472.050 511.050 ;
        RECT 425.400 478.050 426.450 508.950 ;
        RECT 331.950 475.950 334.050 478.050 ;
        RECT 352.950 475.950 355.050 478.050 ;
        RECT 424.950 475.950 427.050 478.050 ;
        RECT 329.400 450.450 330.600 450.600 ;
        RECT 332.400 450.450 333.450 475.950 ;
        RECT 329.400 449.400 333.450 450.450 ;
        RECT 329.400 448.350 330.600 449.400 ;
        RECT 353.400 421.050 354.450 475.950 ;
        RECT 352.950 418.950 355.050 421.050 ;
        RECT 370.950 418.950 373.050 421.050 ;
        RECT 185.400 411.000 186.600 412.650 ;
        RECT 344.400 411.000 345.600 412.650 ;
        RECT 365.400 411.000 366.600 412.650 ;
        RECT 184.950 406.950 187.050 411.000 ;
        RECT 268.950 408.450 273.000 409.050 ;
        RECT 268.950 406.950 273.450 408.450 ;
        RECT 301.950 406.950 304.050 409.050 ;
        RECT 343.950 406.950 346.050 411.000 ;
        RECT 364.950 406.950 367.050 411.000 ;
        RECT 371.400 409.050 372.450 418.950 ;
        RECT 370.950 406.950 373.050 409.050 ;
        RECT 272.400 397.050 273.450 406.950 ;
        RECT 302.400 397.050 303.450 406.950 ;
        RECT 271.950 394.950 274.050 397.050 ;
        RECT 301.950 394.950 304.050 397.050 ;
      LAYER metal3 ;
        RECT 295.950 918.750 298.050 919.200 ;
        RECT 310.950 918.750 313.050 919.200 ;
        RECT 295.950 917.550 313.050 918.750 ;
        RECT 295.950 917.100 298.050 917.550 ;
        RECT 310.950 917.100 313.050 917.550 ;
        RECT 301.950 894.600 304.050 895.050 ;
        RECT 310.950 894.600 313.050 895.050 ;
        RECT 328.950 894.600 331.050 895.050 ;
        RECT 301.950 893.400 331.050 894.600 ;
        RECT 301.950 892.950 304.050 893.400 ;
        RECT 310.950 892.950 313.050 893.400 ;
        RECT 328.950 892.950 331.050 893.400 ;
        RECT 328.950 837.600 331.050 841.050 ;
        RECT 328.950 837.000 333.600 837.600 ;
        RECT 329.400 836.400 333.600 837.000 ;
        RECT 332.400 834.600 333.600 836.400 ;
        RECT 346.800 834.600 348.900 834.900 ;
        RECT 332.400 833.400 348.900 834.600 ;
        RECT 346.800 832.800 348.900 833.400 ;
        RECT 355.950 825.600 358.050 826.050 ;
        RECT 388.950 825.600 391.050 826.050 ;
        RECT 394.950 825.600 397.050 826.050 ;
        RECT 355.950 824.400 397.050 825.600 ;
        RECT 355.950 823.950 358.050 824.400 ;
        RECT 388.950 823.950 391.050 824.400 ;
        RECT 394.950 823.950 397.050 824.400 ;
        RECT 358.950 777.600 361.050 778.050 ;
        RECT 388.950 777.600 391.050 778.050 ;
        RECT 358.950 776.400 391.050 777.600 ;
        RECT 358.950 775.950 361.050 776.400 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 811.950 771.600 814.050 772.050 ;
        RECT 886.950 771.600 889.050 772.050 ;
        RECT 811.950 770.400 889.050 771.600 ;
        RECT 811.950 769.950 814.050 770.400 ;
        RECT 886.950 769.950 889.050 770.400 ;
        RECT 810.000 765.600 814.050 766.050 ;
        RECT 809.400 763.950 814.050 765.600 ;
        RECT 787.950 762.750 790.050 763.200 ;
        RECT 793.950 762.750 796.050 762.900 ;
        RECT 787.950 762.600 796.050 762.750 ;
        RECT 809.400 762.600 810.600 763.950 ;
        RECT 787.950 761.550 810.600 762.600 ;
        RECT 787.950 761.100 790.050 761.550 ;
        RECT 793.950 761.400 810.600 761.550 ;
        RECT 793.950 760.800 796.050 761.400 ;
        RECT 739.950 750.600 742.050 751.050 ;
        RECT 793.950 750.600 796.050 751.050 ;
        RECT 739.950 749.400 796.050 750.600 ;
        RECT 739.950 748.950 742.050 749.400 ;
        RECT 793.950 748.950 796.050 749.400 ;
        RECT 379.950 735.600 382.050 736.050 ;
        RECT 427.950 735.600 430.050 736.050 ;
        RECT 379.950 734.400 430.050 735.600 ;
        RECT 379.950 733.950 382.050 734.400 ;
        RECT 427.950 733.950 430.050 734.400 ;
        RECT 361.950 726.600 364.050 730.050 ;
        RECT 361.950 726.000 369.600 726.600 ;
        RECT 362.400 725.400 369.600 726.000 ;
        RECT 368.400 723.900 369.600 725.400 ;
        RECT 367.950 721.800 370.050 723.900 ;
        RECT 586.950 714.600 589.050 715.050 ;
        RECT 682.950 714.600 685.050 715.050 ;
        RECT 586.950 713.400 685.050 714.600 ;
        RECT 586.950 712.950 589.050 713.400 ;
        RECT 682.950 712.950 685.050 713.400 ;
        RECT 694.950 714.600 697.050 715.050 ;
        RECT 739.950 714.600 742.050 715.050 ;
        RECT 757.950 714.600 760.050 715.050 ;
        RECT 694.950 713.400 760.050 714.600 ;
        RECT 694.950 712.950 697.050 713.400 ;
        RECT 739.950 712.950 742.050 713.400 ;
        RECT 757.950 712.950 760.050 713.400 ;
        RECT 367.950 711.600 370.050 712.050 ;
        RECT 379.950 711.600 382.050 712.050 ;
        RECT 367.950 710.400 382.050 711.600 ;
        RECT 367.950 709.950 370.050 710.400 ;
        RECT 379.950 709.950 382.050 710.400 ;
        RECT 427.950 702.600 430.050 703.050 ;
        RECT 436.950 702.600 439.050 703.050 ;
        RECT 427.950 701.400 439.050 702.600 ;
        RECT 427.950 700.950 430.050 701.400 ;
        RECT 436.950 700.950 439.050 701.400 ;
        RECT 526.950 696.600 529.050 697.050 ;
        RECT 586.950 696.600 589.050 697.050 ;
        RECT 526.950 695.400 589.050 696.600 ;
        RECT 526.950 694.950 529.050 695.400 ;
        RECT 586.950 694.950 589.050 695.400 ;
        RECT 436.950 690.600 439.050 691.050 ;
        RECT 526.950 690.600 529.050 691.050 ;
        RECT 436.950 689.400 529.050 690.600 ;
        RECT 436.950 688.950 439.050 689.400 ;
        RECT 526.950 688.950 529.050 689.400 ;
        RECT 757.950 624.600 760.050 625.050 ;
        RECT 757.950 623.400 780.600 624.600 ;
        RECT 757.950 622.950 760.050 623.400 ;
        RECT 779.400 621.600 780.600 623.400 ;
        RECT 808.950 621.600 811.050 622.050 ;
        RECT 886.950 621.600 889.050 622.050 ;
        RECT 779.400 620.400 889.050 621.600 ;
        RECT 808.950 619.950 811.050 620.400 ;
        RECT 886.950 619.950 889.050 620.400 ;
        RECT 805.950 564.600 808.050 565.050 ;
        RECT 874.950 564.600 877.050 565.050 ;
        RECT 805.950 563.400 877.050 564.600 ;
        RECT 805.950 562.950 808.050 563.400 ;
        RECT 874.950 562.950 877.050 563.400 ;
        RECT 538.950 546.600 541.050 547.050 ;
        RECT 805.950 546.600 808.050 547.050 ;
        RECT 538.950 545.400 808.050 546.600 ;
        RECT 538.950 544.950 541.050 545.400 ;
        RECT 805.950 544.950 808.050 545.400 ;
        RECT 481.950 537.600 484.050 538.050 ;
        RECT 538.950 537.600 541.050 538.050 ;
        RECT 481.950 536.400 541.050 537.600 ;
        RECT 481.950 535.950 484.050 536.400 ;
        RECT 538.950 535.950 541.050 536.400 ;
        RECT 799.950 537.600 802.050 538.050 ;
        RECT 805.950 537.600 808.050 538.050 ;
        RECT 799.950 536.400 808.050 537.600 ;
        RECT 799.950 535.950 802.050 536.400 ;
        RECT 805.950 535.950 808.050 536.400 ;
        RECT 469.950 531.600 472.050 532.050 ;
        RECT 481.950 531.600 484.050 532.050 ;
        RECT 469.950 530.400 484.050 531.600 ;
        RECT 469.950 529.950 472.050 530.400 ;
        RECT 481.950 529.950 484.050 530.400 ;
        RECT 424.950 510.600 427.050 511.050 ;
        RECT 469.950 510.600 472.050 511.050 ;
        RECT 424.950 509.400 472.050 510.600 ;
        RECT 424.950 508.950 427.050 509.400 ;
        RECT 469.950 508.950 472.050 509.400 ;
        RECT 331.950 477.600 334.050 478.050 ;
        RECT 352.950 477.600 355.050 478.050 ;
        RECT 424.950 477.600 427.050 478.050 ;
        RECT 331.950 476.400 427.050 477.600 ;
        RECT 331.950 475.950 334.050 476.400 ;
        RECT 352.950 475.950 355.050 476.400 ;
        RECT 424.950 475.950 427.050 476.400 ;
        RECT 352.950 420.600 355.050 421.050 ;
        RECT 370.950 420.600 373.050 421.050 ;
        RECT 352.950 419.400 373.050 420.600 ;
        RECT 352.950 418.950 355.050 419.400 ;
        RECT 370.950 418.950 373.050 419.400 ;
        RECT 184.950 408.600 187.050 409.050 ;
        RECT 268.950 408.600 271.050 409.050 ;
        RECT 184.950 407.400 271.050 408.600 ;
        RECT 184.950 406.950 187.050 407.400 ;
        RECT 268.950 406.950 271.050 407.400 ;
        RECT 301.950 408.600 304.050 409.050 ;
        RECT 343.950 408.600 346.050 409.050 ;
        RECT 364.950 408.600 367.050 409.050 ;
        RECT 370.950 408.600 373.050 409.050 ;
        RECT 301.950 407.400 373.050 408.600 ;
        RECT 301.950 406.950 304.050 407.400 ;
        RECT 343.950 406.950 346.050 407.400 ;
        RECT 364.950 406.950 367.050 407.400 ;
        RECT 370.950 406.950 373.050 407.400 ;
        RECT 271.950 396.600 274.050 397.050 ;
        RECT 301.950 396.600 304.050 397.050 ;
        RECT 271.950 395.400 304.050 396.600 ;
        RECT 271.950 394.950 274.050 395.400 ;
        RECT 301.950 394.950 304.050 395.400 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal2 ;
        RECT 254.400 940.050 255.450 945.450 ;
        RECT 253.950 937.950 256.050 940.050 ;
        RECT 268.950 937.950 271.050 940.050 ;
        RECT 242.400 878.400 243.600 880.650 ;
        RECT 263.400 878.400 264.600 880.650 ;
        RECT 242.400 865.050 243.450 878.400 ;
        RECT 263.400 865.050 264.450 878.400 ;
        RECT 269.400 865.050 270.450 937.950 ;
        RECT 241.950 862.950 244.050 865.050 ;
        RECT 262.950 862.950 265.050 865.050 ;
        RECT 268.950 862.950 271.050 865.050 ;
        RECT 331.950 862.950 334.050 865.050 ;
        RECT 332.400 856.050 333.450 862.950 ;
        RECT 331.950 853.950 334.050 856.050 ;
        RECT 442.950 853.950 445.050 856.050 ;
        RECT 332.400 808.200 333.450 853.950 ;
        RECT 325.950 806.100 328.050 808.200 ;
        RECT 331.950 806.100 334.050 808.200 ;
        RECT 440.400 807.450 441.600 807.600 ;
        RECT 443.400 807.450 444.450 853.950 ;
        RECT 440.400 806.400 444.450 807.450 ;
        RECT 317.400 801.900 318.600 802.650 ;
        RECT 326.400 802.050 327.450 806.100 ;
        RECT 332.400 805.350 333.600 806.100 ;
        RECT 440.400 805.350 441.600 806.400 ;
        RECT 316.950 799.800 319.050 801.900 ;
        RECT 325.950 799.950 328.050 802.050 ;
      LAYER metal3 ;
        RECT 253.950 939.600 256.050 940.050 ;
        RECT 268.950 939.600 271.050 940.050 ;
        RECT 253.950 938.400 271.050 939.600 ;
        RECT 253.950 937.950 256.050 938.400 ;
        RECT 268.950 937.950 271.050 938.400 ;
        RECT 241.950 864.600 244.050 865.050 ;
        RECT 262.950 864.600 265.050 865.050 ;
        RECT 268.950 864.600 271.050 865.050 ;
        RECT 331.950 864.600 334.050 865.050 ;
        RECT 241.950 863.400 334.050 864.600 ;
        RECT 241.950 862.950 244.050 863.400 ;
        RECT 262.950 862.950 265.050 863.400 ;
        RECT 268.950 862.950 271.050 863.400 ;
        RECT 331.950 862.950 334.050 863.400 ;
        RECT 331.950 855.600 334.050 856.050 ;
        RECT 442.950 855.600 445.050 856.050 ;
        RECT 331.950 854.400 445.050 855.600 ;
        RECT 331.950 853.950 334.050 854.400 ;
        RECT 442.950 853.950 445.050 854.400 ;
        RECT 325.950 807.750 328.050 808.200 ;
        RECT 331.950 807.750 334.050 808.200 ;
        RECT 325.950 806.550 334.050 807.750 ;
        RECT 325.950 806.100 328.050 806.550 ;
        RECT 331.950 806.100 334.050 806.550 ;
        RECT 316.950 801.600 319.050 801.900 ;
        RECT 325.950 801.600 328.050 802.050 ;
        RECT 316.950 800.400 328.050 801.600 ;
        RECT 316.950 799.800 319.050 800.400 ;
        RECT 325.950 799.950 328.050 800.400 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal1 ;
        RECT 19.950 609.450 22.050 610.050 ;
        RECT 25.950 609.450 28.050 609.900 ;
        RECT 19.950 608.550 28.050 609.450 ;
        RECT 19.950 607.950 22.050 608.550 ;
        RECT 25.950 607.800 28.050 608.550 ;
        RECT 318.000 495.450 322.050 496.050 ;
        RECT 317.550 493.950 322.050 495.450 ;
        RECT 317.550 490.050 318.450 493.950 ;
        RECT 313.950 488.550 318.450 490.050 ;
        RECT 313.950 487.950 318.000 488.550 ;
      LAYER metal2 ;
        RECT 70.950 709.950 73.050 712.050 ;
        RECT 112.950 709.950 115.050 712.050 ;
        RECT 181.950 709.950 184.050 712.050 ;
        RECT 232.950 709.950 235.050 712.050 ;
        RECT 71.400 691.050 72.450 709.950 ;
        RECT 113.400 694.050 114.450 709.950 ;
        RECT 182.400 694.050 183.450 709.950 ;
        RECT 112.950 691.950 115.050 694.050 ;
        RECT 157.950 691.950 160.050 694.050 ;
        RECT 181.950 691.950 184.050 694.050 ;
        RECT 31.950 688.950 34.050 691.050 ;
        RECT 43.950 688.950 46.050 691.050 ;
        RECT 70.950 688.950 73.050 691.050 ;
        RECT 32.400 684.600 33.450 688.950 ;
        RECT 32.400 682.350 33.600 684.600 ;
        RECT 44.400 663.450 45.450 688.950 ;
        RECT 158.400 685.050 159.450 691.950 ;
        RECT 182.400 687.450 183.450 691.950 ;
        RECT 182.400 686.400 186.450 687.450 ;
        RECT 157.950 682.950 160.050 685.050 ;
        RECT 185.400 684.600 186.450 686.400 ;
        RECT 233.400 684.600 234.450 709.950 ;
        RECT 185.400 682.350 186.600 684.600 ;
        RECT 233.400 682.350 234.600 684.600 ;
        RECT 157.950 676.950 160.050 679.050 ;
        RECT 44.400 662.400 48.450 663.450 ;
        RECT 47.400 628.050 48.450 662.400 ;
        RECT 56.400 644.400 57.600 646.650 ;
        RECT 56.400 628.050 57.450 644.400 ;
        RECT 19.950 625.950 22.050 628.050 ;
        RECT 46.950 625.950 49.050 628.050 ;
        RECT 55.950 625.950 58.050 628.050 ;
        RECT 20.400 610.050 21.450 625.950 ;
        RECT 158.400 625.050 159.450 676.950 ;
        RECT 157.950 622.950 160.050 625.050 ;
        RECT 187.950 622.950 190.050 625.050 ;
        RECT 19.950 606.000 22.050 610.050 ;
        RECT 25.950 607.800 28.050 609.900 ;
        RECT 158.400 609.450 159.450 622.950 ;
        RECT 155.400 608.400 159.450 609.450 ;
        RECT 20.400 604.350 21.600 606.000 ;
        RECT 26.400 580.050 27.450 607.800 ;
        RECT 155.400 606.600 156.450 608.400 ;
        RECT 155.400 604.350 156.600 606.600 ;
        RECT 1.950 577.950 4.050 580.050 ;
        RECT 25.950 577.950 28.050 580.050 ;
        RECT 188.400 579.450 189.450 622.950 ;
        RECT 287.400 600.450 288.600 601.650 ;
        RECT 284.400 599.400 288.600 600.450 ;
        RECT 284.400 592.050 285.450 599.400 ;
        RECT 283.950 589.950 286.050 592.050 ;
        RECT 316.950 589.950 319.050 592.050 ;
        RECT 188.400 579.000 192.450 579.450 ;
        RECT 188.400 578.400 193.050 579.000 ;
        RECT 2.400 535.050 3.450 577.950 ;
        RECT 190.950 574.950 193.050 578.400 ;
        RECT 284.400 577.050 285.450 589.950 ;
        RECT 283.950 574.950 286.050 577.050 ;
        RECT 317.400 570.450 318.450 589.950 ;
        RECT 317.400 569.400 321.450 570.450 ;
        RECT 1.950 532.950 4.050 535.050 ;
        RECT 2.400 502.050 3.450 532.950 ;
        RECT 1.950 499.950 4.050 502.050 ;
        RECT 19.950 499.950 22.050 502.050 ;
        RECT 2.400 489.900 3.450 499.950 ;
        RECT 20.400 495.600 21.450 499.950 ;
        RECT 320.400 496.050 321.450 569.400 ;
        RECT 20.400 493.350 21.600 495.600 ;
        RECT 319.950 493.950 322.050 496.050 ;
        RECT 56.400 489.900 57.600 490.650 ;
        RECT 1.950 487.800 4.050 489.900 ;
        RECT 55.950 487.800 58.050 489.900 ;
        RECT 313.950 487.950 316.050 490.050 ;
        RECT 56.400 460.050 57.450 487.800 ;
        RECT 314.400 460.050 315.450 487.950 ;
        RECT 55.950 457.950 58.050 460.050 ;
        RECT 76.950 457.800 79.050 459.900 ;
        RECT 274.950 457.950 277.050 460.050 ;
        RECT 313.950 457.950 316.050 460.050 ;
        RECT 77.400 450.600 78.450 457.800 ;
        RECT 275.400 450.600 276.450 457.950 ;
        RECT 77.400 448.350 78.600 450.600 ;
        RECT 275.400 448.350 276.600 450.600 ;
      LAYER metal3 ;
        RECT 70.950 711.600 73.050 712.050 ;
        RECT 112.950 711.600 115.050 712.050 ;
        RECT 70.950 710.400 115.050 711.600 ;
        RECT 70.950 709.950 73.050 710.400 ;
        RECT 112.950 709.950 115.050 710.400 ;
        RECT 181.950 711.600 184.050 712.050 ;
        RECT 232.950 711.600 235.050 712.050 ;
        RECT 181.950 710.400 235.050 711.600 ;
        RECT 181.950 709.950 184.050 710.400 ;
        RECT 232.950 709.950 235.050 710.400 ;
        RECT 112.950 693.600 115.050 694.050 ;
        RECT 157.950 693.600 160.050 694.050 ;
        RECT 181.950 693.600 184.050 694.050 ;
        RECT 112.950 692.400 184.050 693.600 ;
        RECT 112.950 691.950 115.050 692.400 ;
        RECT 157.950 691.950 160.050 692.400 ;
        RECT 181.950 691.950 184.050 692.400 ;
        RECT 31.950 690.600 34.050 691.050 ;
        RECT 43.950 690.600 46.050 691.050 ;
        RECT 70.950 690.600 73.050 691.050 ;
        RECT 31.950 689.400 73.050 690.600 ;
        RECT 31.950 688.950 34.050 689.400 ;
        RECT 43.950 688.950 46.050 689.400 ;
        RECT 70.950 688.950 73.050 689.400 ;
        RECT 157.950 682.950 160.050 685.050 ;
        RECT 158.400 679.050 159.600 682.950 ;
        RECT 157.950 676.950 160.050 679.050 ;
        RECT 19.950 627.600 22.050 628.050 ;
        RECT 46.950 627.600 49.050 628.050 ;
        RECT 55.950 627.600 58.050 628.050 ;
        RECT 19.950 626.400 58.050 627.600 ;
        RECT 19.950 625.950 22.050 626.400 ;
        RECT 46.950 625.950 49.050 626.400 ;
        RECT 55.950 625.950 58.050 626.400 ;
        RECT 157.950 624.600 160.050 625.050 ;
        RECT 187.950 624.600 190.050 625.050 ;
        RECT 157.950 623.400 190.050 624.600 ;
        RECT 157.950 622.950 160.050 623.400 ;
        RECT 187.950 622.950 190.050 623.400 ;
        RECT 283.950 591.600 286.050 592.050 ;
        RECT 316.950 591.600 319.050 592.050 ;
        RECT 283.950 590.400 319.050 591.600 ;
        RECT 283.950 589.950 286.050 590.400 ;
        RECT 316.950 589.950 319.050 590.400 ;
        RECT 1.950 579.600 4.050 580.050 ;
        RECT 25.950 579.600 28.050 580.050 ;
        RECT 1.950 578.400 28.050 579.600 ;
        RECT 1.950 577.950 4.050 578.400 ;
        RECT 25.950 577.950 28.050 578.400 ;
        RECT 190.950 576.600 193.050 577.050 ;
        RECT 283.950 576.600 286.050 577.050 ;
        RECT 190.950 575.400 286.050 576.600 ;
        RECT 190.950 574.950 193.050 575.400 ;
        RECT 283.950 574.950 286.050 575.400 ;
        RECT 1.950 534.600 4.050 535.050 ;
        RECT -3.600 533.400 4.050 534.600 ;
        RECT 1.950 532.950 4.050 533.400 ;
        RECT 1.950 501.600 4.050 502.050 ;
        RECT 19.950 501.600 22.050 502.050 ;
        RECT 1.950 500.400 22.050 501.600 ;
        RECT 1.950 499.950 4.050 500.400 ;
        RECT 19.950 499.950 22.050 500.400 ;
        RECT 1.950 489.450 4.050 489.900 ;
        RECT 55.950 489.450 58.050 489.900 ;
        RECT 1.950 488.250 58.050 489.450 ;
        RECT 1.950 487.800 4.050 488.250 ;
        RECT 55.950 487.800 58.050 488.250 ;
        RECT 55.950 459.600 58.050 460.050 ;
        RECT 76.950 459.600 79.050 459.900 ;
        RECT 55.950 458.400 79.050 459.600 ;
        RECT 55.950 457.950 58.050 458.400 ;
        RECT 76.950 457.800 79.050 458.400 ;
        RECT 274.950 459.600 277.050 460.050 ;
        RECT 313.950 459.600 316.050 460.050 ;
        RECT 274.950 458.400 316.050 459.600 ;
        RECT 274.950 457.950 277.050 458.400 ;
        RECT 313.950 457.950 316.050 458.400 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal2 ;
        RECT 7.950 605.100 10.050 607.200 ;
        RECT 13.950 605.100 16.050 607.200 ;
        RECT 8.400 574.200 9.450 605.100 ;
        RECT 14.400 604.350 15.600 605.100 ;
        RECT 7.950 572.100 10.050 574.200 ;
        RECT 16.950 572.100 19.050 574.200 ;
        RECT 8.400 529.050 9.450 572.100 ;
        RECT 17.400 571.350 18.600 572.100 ;
        RECT 7.950 526.950 10.050 529.050 ;
        RECT 13.950 527.100 16.050 529.200 ;
        RECT 14.400 526.350 15.600 527.100 ;
      LAYER metal3 ;
        RECT 7.950 606.750 10.050 607.200 ;
        RECT 13.950 606.750 16.050 607.200 ;
        RECT 7.950 605.550 16.050 606.750 ;
        RECT 7.950 605.100 10.050 605.550 ;
        RECT 13.950 605.100 16.050 605.550 ;
        RECT 7.950 573.750 10.050 574.200 ;
        RECT 16.950 573.750 19.050 574.200 ;
        RECT 7.950 572.550 19.050 573.750 ;
        RECT 7.950 572.100 10.050 572.550 ;
        RECT 16.950 572.100 19.050 572.550 ;
        RECT 7.950 528.600 10.050 529.050 ;
        RECT 13.950 528.600 16.050 529.200 ;
        RECT -3.600 527.400 16.050 528.600 ;
        RECT 7.950 526.950 10.050 527.400 ;
        RECT 13.950 527.100 16.050 527.400 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal1 ;
        RECT 79.950 687.450 82.050 688.050 ;
        RECT 91.950 687.450 94.050 688.050 ;
        RECT 79.950 686.550 94.050 687.450 ;
        RECT 79.950 685.950 82.050 686.550 ;
        RECT 91.950 685.950 94.050 686.550 ;
      LAYER metal2 ;
        RECT 91.950 694.950 94.050 697.050 ;
        RECT 130.950 694.950 133.050 697.050 ;
        RECT 10.950 691.950 13.050 694.050 ;
        RECT 79.950 691.950 82.050 694.050 ;
        RECT 11.400 685.200 12.450 691.950 ;
        RECT 80.400 688.050 81.450 691.950 ;
        RECT 92.400 688.050 93.450 694.950 ;
        RECT 79.950 685.950 82.050 688.050 ;
        RECT 91.950 685.950 94.050 688.050 ;
        RECT 10.950 683.100 13.050 685.200 ;
        RECT 11.400 682.350 12.600 683.100 ;
        RECT 131.400 673.050 132.450 694.950 ;
        RECT 161.400 677.400 162.600 679.650 ;
        RECT 161.400 673.050 162.450 677.400 ;
        RECT 130.950 670.950 133.050 673.050 ;
        RECT 160.950 670.950 163.050 673.050 ;
      LAYER metal3 ;
        RECT 91.950 696.600 94.050 697.050 ;
        RECT 130.950 696.600 133.050 697.050 ;
        RECT 91.950 695.400 133.050 696.600 ;
        RECT 91.950 694.950 94.050 695.400 ;
        RECT 130.950 694.950 133.050 695.400 ;
        RECT 10.950 693.600 13.050 694.050 ;
        RECT 79.950 693.600 82.050 694.050 ;
        RECT 10.950 692.400 82.050 693.600 ;
        RECT 10.950 691.950 13.050 692.400 ;
        RECT 79.950 691.950 82.050 692.400 ;
        RECT 10.950 684.600 13.050 685.200 ;
        RECT -3.600 683.400 13.050 684.600 ;
        RECT 10.950 683.100 13.050 683.400 ;
        RECT 130.950 672.600 133.050 673.050 ;
        RECT 160.950 672.600 163.050 673.050 ;
        RECT 130.950 671.400 163.050 672.600 ;
        RECT 130.950 670.950 133.050 671.400 ;
        RECT 160.950 670.950 163.050 671.400 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal2 ;
        RECT 44.400 729.450 45.600 729.600 ;
        RECT 155.400 729.450 156.600 729.600 ;
        RECT 44.400 728.400 48.450 729.450 ;
        RECT 44.400 727.350 45.600 728.400 ;
        RECT 47.400 700.050 48.450 728.400 ;
        RECT 155.400 728.400 159.450 729.450 ;
        RECT 155.400 727.350 156.600 728.400 ;
        RECT 158.400 700.050 159.450 728.400 ;
        RECT 1.950 697.950 4.050 700.050 ;
        RECT 46.950 697.950 49.050 700.050 ;
        RECT 151.950 697.950 154.050 700.050 ;
        RECT 157.950 697.950 160.050 700.050 ;
        RECT 2.400 652.050 3.450 697.950 ;
        RECT 1.950 649.950 4.050 652.050 ;
        RECT 13.950 650.100 16.050 652.200 ;
        RECT 152.400 651.600 153.450 697.950 ;
        RECT 14.400 649.350 15.600 650.100 ;
        RECT 152.400 649.350 153.600 651.600 ;
      LAYER metal3 ;
        RECT 1.950 699.600 4.050 700.050 ;
        RECT 46.950 699.600 49.050 700.050 ;
        RECT 151.950 699.600 154.050 700.050 ;
        RECT 157.950 699.600 160.050 700.050 ;
        RECT 1.950 698.400 160.050 699.600 ;
        RECT 1.950 697.950 4.050 698.400 ;
        RECT 46.950 697.950 49.050 698.400 ;
        RECT 151.950 697.950 154.050 698.400 ;
        RECT 157.950 697.950 160.050 698.400 ;
        RECT 1.950 651.600 4.050 652.050 ;
        RECT 13.950 651.600 16.050 652.200 ;
        RECT -3.600 650.400 16.050 651.600 ;
        RECT 1.950 649.950 4.050 650.400 ;
        RECT 13.950 650.100 16.050 650.400 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal2 ;
        RECT 166.950 449.100 169.050 451.200 ;
        RECT 167.400 448.350 168.600 449.100 ;
        RECT 175.950 448.950 178.050 451.050 ;
        RECT 176.400 444.900 177.450 448.950 ;
        RECT 185.400 444.900 186.600 445.650 ;
        RECT 175.950 442.800 178.050 444.900 ;
        RECT 184.950 442.800 187.050 444.900 ;
        RECT 1.950 436.950 4.050 439.050 ;
        RECT 25.950 436.950 28.050 439.050 ;
        RECT 2.400 418.050 3.450 436.950 ;
        RECT 1.950 415.950 4.050 418.050 ;
        RECT 26.400 417.600 27.450 436.950 ;
        RECT 176.400 436.050 177.450 442.800 ;
        RECT 103.950 433.950 106.050 436.050 ;
        RECT 175.950 433.950 178.050 436.050 ;
        RECT 26.400 415.350 27.600 417.600 ;
        RECT 92.400 411.900 93.600 412.650 ;
        RECT 104.400 411.900 105.450 433.950 ;
        RECT 91.950 409.800 94.050 411.900 ;
        RECT 103.950 409.800 106.050 411.900 ;
      LAYER metal3 ;
        RECT 166.950 450.600 169.050 451.200 ;
        RECT 175.950 450.600 178.050 451.050 ;
        RECT 166.950 449.400 178.050 450.600 ;
        RECT 166.950 449.100 169.050 449.400 ;
        RECT 175.950 448.950 178.050 449.400 ;
        RECT 175.950 444.450 178.050 444.900 ;
        RECT 184.950 444.450 187.050 444.900 ;
        RECT 175.950 443.250 187.050 444.450 ;
        RECT 175.950 442.800 178.050 443.250 ;
        RECT 184.950 442.800 187.050 443.250 ;
        RECT 1.950 438.600 4.050 439.050 ;
        RECT 25.950 438.600 28.050 439.050 ;
        RECT 1.950 437.400 105.600 438.600 ;
        RECT 1.950 436.950 4.050 437.400 ;
        RECT 25.950 436.950 28.050 437.400 ;
        RECT 104.400 436.050 105.600 437.400 ;
        RECT 103.950 435.600 106.050 436.050 ;
        RECT 175.950 435.600 178.050 436.050 ;
        RECT 103.950 434.400 178.050 435.600 ;
        RECT 103.950 433.950 106.050 434.400 ;
        RECT 175.950 433.950 178.050 434.400 ;
        RECT 1.950 417.600 4.050 418.050 ;
        RECT -3.600 416.400 4.050 417.600 ;
        RECT 1.950 415.950 4.050 416.400 ;
        RECT 91.950 411.450 94.050 411.900 ;
        RECT 103.950 411.450 106.050 411.900 ;
        RECT 91.950 410.250 106.050 411.450 ;
        RECT 91.950 409.800 94.050 410.250 ;
        RECT 103.950 409.800 106.050 410.250 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal1 ;
        RECT 124.950 564.450 127.050 565.050 ;
        RECT 133.950 564.450 136.050 565.050 ;
        RECT 124.950 563.550 136.050 564.450 ;
        RECT 124.950 562.950 127.050 563.550 ;
        RECT 133.950 562.950 136.050 563.550 ;
        RECT 217.950 561.450 220.050 562.050 ;
        RECT 217.950 561.000 225.450 561.450 ;
        RECT 217.950 560.550 226.050 561.000 ;
        RECT 217.950 559.950 220.050 560.550 ;
        RECT 223.950 559.050 226.050 560.550 ;
        RECT 223.800 558.000 226.050 559.050 ;
        RECT 223.800 556.950 225.900 558.000 ;
        RECT 229.950 456.450 232.050 457.050 ;
        RECT 244.950 456.450 247.050 457.050 ;
        RECT 229.950 455.550 247.050 456.450 ;
        RECT 229.950 454.950 232.050 455.550 ;
        RECT 244.950 454.950 247.050 455.550 ;
      LAYER metal2 ;
        RECT 124.950 572.100 127.050 574.200 ;
        RECT 139.800 572.100 141.900 574.200 ;
        RECT 298.950 572.100 301.050 574.200 ;
        RECT 304.950 572.100 307.050 574.200 ;
        RECT 74.400 567.000 75.600 568.650 ;
        RECT 73.950 562.950 76.050 567.000 ;
        RECT 125.400 565.050 126.450 572.100 ;
        RECT 140.400 571.350 141.600 572.100 ;
        RECT 109.950 562.950 112.050 565.050 ;
        RECT 124.950 562.950 127.050 565.050 ;
        RECT 110.400 505.050 111.450 562.950 ;
        RECT 133.950 562.050 136.050 565.050 ;
        RECT 299.400 562.050 300.450 572.100 ;
        RECT 305.400 571.350 306.600 572.100 ;
        RECT 133.950 561.000 139.050 562.050 ;
        RECT 134.400 560.400 139.050 561.000 ;
        RECT 135.000 559.950 139.050 560.400 ;
        RECT 214.950 559.950 220.050 562.050 ;
        RECT 223.950 559.050 226.050 562.050 ;
        RECT 298.950 559.950 301.050 562.050 ;
        RECT 223.800 558.000 226.050 559.050 ;
        RECT 223.800 556.950 225.900 558.000 ;
        RECT 109.950 502.950 112.050 505.050 ;
        RECT 118.950 502.950 121.050 505.050 ;
        RECT 119.400 487.050 120.450 502.950 ;
        RECT 152.400 489.000 153.600 490.650 ;
        RECT 118.950 484.950 121.050 487.050 ;
        RECT 151.950 484.950 154.050 489.000 ;
        RECT 119.400 481.050 120.450 484.950 ;
        RECT 73.950 478.950 76.050 481.050 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 74.400 457.050 75.450 478.950 ;
        RECT 1.950 454.950 4.050 457.050 ;
        RECT 73.950 454.950 76.050 457.050 ;
        RECT 2.400 445.050 3.450 454.950 ;
        RECT 152.400 454.050 153.450 484.950 ;
        RECT 226.950 454.950 232.050 457.050 ;
        RECT 244.950 454.950 247.050 457.050 ;
        RECT 151.950 451.950 154.050 454.050 ;
        RECT 1.950 442.950 4.050 445.050 ;
        RECT 11.400 444.900 12.600 445.650 ;
        RECT 10.950 442.800 13.050 444.900 ;
        RECT 11.400 411.450 12.450 442.800 ;
        RECT 245.400 420.450 246.450 454.950 ;
        RECT 242.400 419.400 246.450 420.450 ;
        RECT 242.400 417.600 243.450 419.400 ;
        RECT 242.400 415.350 243.600 417.600 ;
        RECT 14.400 411.450 15.600 412.650 ;
        RECT 11.400 410.400 15.600 411.450 ;
      LAYER metal3 ;
        RECT 124.950 573.750 127.050 574.200 ;
        RECT 139.800 573.750 141.900 574.200 ;
        RECT 124.950 572.550 141.900 573.750 ;
        RECT 124.950 572.100 127.050 572.550 ;
        RECT 139.800 572.100 141.900 572.550 ;
        RECT 298.950 573.750 301.050 574.200 ;
        RECT 304.950 573.750 307.050 574.200 ;
        RECT 298.950 572.550 307.050 573.750 ;
        RECT 298.950 572.100 301.050 572.550 ;
        RECT 304.950 572.100 307.050 572.550 ;
        RECT 73.950 564.600 76.050 565.050 ;
        RECT 109.950 564.600 112.050 565.050 ;
        RECT 124.950 564.600 127.050 565.050 ;
        RECT 73.950 563.400 127.050 564.600 ;
        RECT 73.950 562.950 76.050 563.400 ;
        RECT 109.950 562.950 112.050 563.400 ;
        RECT 124.950 562.950 127.050 563.400 ;
        RECT 136.950 561.600 139.050 562.050 ;
        RECT 214.950 561.600 217.050 562.050 ;
        RECT 136.950 560.400 217.050 561.600 ;
        RECT 136.950 559.950 139.050 560.400 ;
        RECT 214.950 559.950 217.050 560.400 ;
        RECT 223.950 561.600 226.050 562.050 ;
        RECT 298.950 561.600 301.050 562.050 ;
        RECT 223.950 560.400 301.050 561.600 ;
        RECT 223.950 559.950 226.050 560.400 ;
        RECT 298.950 559.950 301.050 560.400 ;
        RECT 109.950 504.600 112.050 505.050 ;
        RECT 118.950 504.600 121.050 505.050 ;
        RECT 109.950 503.400 121.050 504.600 ;
        RECT 109.950 502.950 112.050 503.400 ;
        RECT 118.950 502.950 121.050 503.400 ;
        RECT 118.950 486.600 121.050 487.050 ;
        RECT 151.950 486.600 154.050 487.050 ;
        RECT 118.950 485.400 154.050 486.600 ;
        RECT 118.950 484.950 121.050 485.400 ;
        RECT 151.950 484.950 154.050 485.400 ;
        RECT 73.950 480.600 76.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 73.950 479.400 121.050 480.600 ;
        RECT 73.950 478.950 76.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 1.950 456.600 4.050 457.050 ;
        RECT 73.950 456.600 76.050 457.050 ;
        RECT 226.950 456.600 229.050 457.050 ;
        RECT 1.950 455.400 76.050 456.600 ;
        RECT 1.950 454.950 4.050 455.400 ;
        RECT 73.950 454.950 76.050 455.400 ;
        RECT 221.400 455.400 229.050 456.600 ;
        RECT 151.950 453.600 154.050 454.050 ;
        RECT 221.400 453.600 222.600 455.400 ;
        RECT 226.950 454.950 229.050 455.400 ;
        RECT 151.950 452.400 222.600 453.600 ;
        RECT 151.950 451.950 154.050 452.400 ;
        RECT 1.950 444.600 4.050 445.050 ;
        RECT 10.950 444.600 13.050 444.900 ;
        RECT -3.600 443.400 13.050 444.600 ;
        RECT 1.950 442.950 4.050 443.400 ;
        RECT 10.950 442.800 13.050 443.400 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal2 ;
        RECT 761.400 940.050 762.450 945.450 ;
        RECT 754.950 937.950 757.050 940.050 ;
        RECT 760.950 937.950 763.050 940.050 ;
        RECT 755.400 928.050 756.450 937.950 ;
        RECT 754.950 925.950 757.050 928.050 ;
        RECT 757.950 919.950 760.050 922.050 ;
        RECT 758.400 916.050 759.450 919.950 ;
        RECT 757.950 913.950 760.050 916.050 ;
        RECT 769.950 910.950 772.050 913.050 ;
        RECT 770.400 900.450 771.450 910.950 ;
        RECT 767.400 899.400 771.450 900.450 ;
        RECT 767.400 862.050 768.450 899.400 ;
        RECT 757.950 859.950 760.050 862.050 ;
        RECT 766.950 859.950 769.050 862.050 ;
        RECT 758.400 832.050 759.450 859.950 ;
        RECT 751.950 829.950 754.050 832.050 ;
        RECT 757.950 829.950 760.050 832.050 ;
        RECT 752.400 799.050 753.450 829.950 ;
        RECT 751.950 796.950 754.050 799.050 ;
        RECT 757.950 796.950 760.050 799.050 ;
        RECT 758.400 762.600 759.450 796.950 ;
        RECT 758.400 760.350 759.600 762.600 ;
      LAYER metal3 ;
        RECT 754.950 939.600 757.050 940.050 ;
        RECT 760.950 939.600 763.050 940.050 ;
        RECT 754.950 938.400 763.050 939.600 ;
        RECT 754.950 937.950 757.050 938.400 ;
        RECT 760.950 937.950 763.050 938.400 ;
        RECT 753.000 927.600 757.050 928.050 ;
        RECT 752.400 925.950 757.050 927.600 ;
        RECT 752.400 921.600 753.600 925.950 ;
        RECT 757.950 921.600 760.050 922.050 ;
        RECT 752.400 920.400 760.050 921.600 ;
        RECT 757.950 919.950 760.050 920.400 ;
        RECT 757.950 912.600 760.050 916.050 ;
        RECT 769.950 912.600 772.050 913.050 ;
        RECT 757.950 912.000 772.050 912.600 ;
        RECT 758.400 911.400 772.050 912.000 ;
        RECT 769.950 910.950 772.050 911.400 ;
        RECT 757.950 861.600 760.050 862.050 ;
        RECT 766.950 861.600 769.050 862.050 ;
        RECT 757.950 860.400 769.050 861.600 ;
        RECT 757.950 859.950 760.050 860.400 ;
        RECT 766.950 859.950 769.050 860.400 ;
        RECT 751.950 831.600 754.050 832.050 ;
        RECT 757.950 831.600 760.050 832.050 ;
        RECT 751.950 830.400 760.050 831.600 ;
        RECT 751.950 829.950 754.050 830.400 ;
        RECT 757.950 829.950 760.050 830.400 ;
        RECT 751.950 798.600 754.050 799.050 ;
        RECT 757.950 798.600 760.050 799.050 ;
        RECT 751.950 797.400 760.050 798.600 ;
        RECT 751.950 796.950 754.050 797.400 ;
        RECT 757.950 796.950 760.050 797.400 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal2 ;
        RECT 686.400 944.400 690.450 945.450 ;
        RECT 686.400 918.600 687.450 944.400 ;
        RECT 686.400 916.350 687.600 918.600 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal2 ;
        RECT 731.400 944.400 735.450 945.450 ;
        RECT 734.400 915.450 735.450 944.400 ;
        RECT 731.400 914.400 735.450 915.450 ;
        RECT 731.400 889.050 732.450 914.400 ;
        RECT 730.950 886.950 733.050 889.050 ;
        RECT 733.950 874.950 736.050 877.050 ;
        RECT 734.400 853.050 735.450 874.950 ;
        RECT 727.950 850.950 730.050 853.050 ;
        RECT 733.950 850.950 736.050 853.050 ;
        RECT 728.400 840.600 729.450 850.950 ;
        RECT 728.400 838.350 729.600 840.600 ;
      LAYER metal3 ;
        RECT 730.950 886.950 733.050 889.050 ;
        RECT 731.400 877.050 732.600 886.950 ;
        RECT 731.400 875.400 736.050 877.050 ;
        RECT 732.000 874.950 736.050 875.400 ;
        RECT 727.950 852.600 730.050 853.050 ;
        RECT 733.950 852.600 736.050 853.050 ;
        RECT 727.950 851.400 736.050 852.600 ;
        RECT 727.950 850.950 730.050 851.400 ;
        RECT 733.950 850.950 736.050 851.400 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal2 ;
        RECT 428.400 944.400 432.450 945.450 ;
        RECT 431.400 918.600 432.450 944.400 ;
        RECT 431.400 916.350 432.600 918.600 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal2 ;
        RECT 935.400 801.900 936.600 802.650 ;
        RECT 934.950 799.800 937.050 801.900 ;
      LAYER metal3 ;
        RECT 934.950 801.600 937.050 801.900 ;
        RECT 934.950 800.400 954.600 801.600 ;
        RECT 934.950 799.800 937.050 800.400 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal2 ;
        RECT 587.400 944.400 591.450 945.450 ;
        RECT 590.400 918.600 591.450 944.400 ;
        RECT 590.400 916.350 591.600 918.600 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal2 ;
        RECT 317.400 944.400 321.450 945.450 ;
        RECT 317.400 918.600 318.450 944.400 ;
        RECT 317.400 916.350 318.600 918.600 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal2 ;
        RECT 710.400 944.400 714.450 945.450 ;
        RECT 713.400 918.600 714.450 944.400 ;
        RECT 713.400 916.350 714.600 918.600 ;
    END
  END ACC_o[0]
  PIN Done_LED
    PORT
      LAYER metal2 ;
        RECT 935.400 879.900 936.600 880.650 ;
        RECT 934.950 877.800 937.050 879.900 ;
      LAYER metal3 ;
        RECT 934.950 879.600 937.050 879.900 ;
        RECT 934.950 878.400 954.600 879.600 ;
        RECT 934.950 877.800 937.050 878.400 ;
    END
  END Done_LED
  PIN Done_o
    PORT
      LAYER metal2 ;
        RECT 928.950 839.100 931.050 841.200 ;
        RECT 929.400 838.350 930.600 839.100 ;
      LAYER metal3 ;
        RECT 928.950 840.600 931.050 841.200 ;
        RECT 928.950 839.400 954.600 840.600 ;
        RECT 928.950 839.100 931.050 839.400 ;
    END
  END Done_o
  PIN LoadA_i
    PORT
      LAYER metal2 ;
        RECT 875.400 944.400 879.450 945.450 ;
        RECT 875.400 919.050 876.450 944.400 ;
        RECT 874.950 916.950 877.050 919.050 ;
        RECT 842.400 912.900 843.600 913.650 ;
        RECT 857.400 912.900 858.600 913.650 ;
        RECT 878.400 912.900 879.600 913.650 ;
        RECT 841.950 910.800 844.050 912.900 ;
        RECT 856.950 910.800 859.050 912.900 ;
        RECT 877.950 910.800 880.050 912.900 ;
      LAYER metal3 ;
        RECT 874.950 916.950 877.050 919.050 ;
        RECT 841.950 912.600 844.050 912.900 ;
        RECT 856.950 912.600 859.050 912.900 ;
        RECT 875.400 912.600 876.600 916.950 ;
        RECT 877.950 912.600 880.050 912.900 ;
        RECT 841.950 911.400 880.050 912.600 ;
        RECT 841.950 910.800 844.050 911.400 ;
        RECT 856.950 910.800 859.050 911.400 ;
        RECT 877.950 910.800 880.050 911.400 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal2 ;
        RECT 854.400 931.050 855.450 945.450 ;
        RECT 853.950 930.450 856.050 931.050 ;
        RECT 851.400 929.400 856.050 930.450 ;
        RECT 851.400 907.050 852.450 929.400 ;
        RECT 853.950 928.950 856.050 929.400 ;
        RECT 859.950 928.950 862.050 931.050 ;
        RECT 904.950 928.950 907.050 931.050 ;
        RECT 860.400 918.600 861.450 928.950 ;
        RECT 905.400 919.200 906.450 928.950 ;
        RECT 860.400 916.350 861.600 918.600 ;
        RECT 904.950 917.100 907.050 919.200 ;
        RECT 905.400 916.350 906.600 917.100 ;
        RECT 910.950 916.950 913.050 919.050 ;
        RECT 799.950 904.950 802.050 907.050 ;
        RECT 850.950 904.950 853.050 907.050 ;
        RECT 800.400 885.600 801.450 904.950 ;
        RECT 911.400 885.600 912.450 916.950 ;
        RECT 800.400 883.350 801.600 885.600 ;
        RECT 911.400 883.350 912.600 885.600 ;
      LAYER metal3 ;
        RECT 853.950 930.600 856.050 931.050 ;
        RECT 859.950 930.600 862.050 931.050 ;
        RECT 904.950 930.600 907.050 931.050 ;
        RECT 853.950 929.400 907.050 930.600 ;
        RECT 853.950 928.950 856.050 929.400 ;
        RECT 859.950 928.950 862.050 929.400 ;
        RECT 904.950 928.950 907.050 929.400 ;
        RECT 904.950 918.600 907.050 919.200 ;
        RECT 910.950 918.600 913.050 919.050 ;
        RECT 904.950 917.400 913.050 918.600 ;
        RECT 904.950 917.100 907.050 917.400 ;
        RECT 910.950 916.950 913.050 917.400 ;
        RECT 799.950 906.600 802.050 907.050 ;
        RECT 850.950 906.600 853.050 907.050 ;
        RECT 799.950 905.400 853.050 906.600 ;
        RECT 799.950 904.950 802.050 905.400 ;
        RECT 850.950 904.950 853.050 905.400 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal2 ;
        RECT 926.400 912.900 927.600 913.650 ;
        RECT 941.400 912.900 942.600 913.650 ;
        RECT 925.950 910.800 928.050 912.900 ;
        RECT 940.950 910.800 943.050 912.900 ;
      LAYER metal3 ;
        RECT 925.950 912.600 928.050 912.900 ;
        RECT 940.950 912.600 943.050 912.900 ;
        RECT 953.400 912.600 954.600 918.600 ;
        RECT 925.950 911.400 954.600 912.600 ;
        RECT 925.950 910.800 928.050 911.400 ;
        RECT 940.950 910.800 943.050 911.400 ;
    END
  END LoadCmd_i
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 500.400 940.050 501.450 945.450 ;
        RECT 499.950 937.950 502.050 940.050 ;
        RECT 550.950 937.950 553.050 940.050 ;
        RECT 551.400 910.050 552.450 937.950 ;
        RECT 508.950 907.950 511.050 910.050 ;
        RECT 550.950 907.950 553.050 910.050 ;
        RECT 509.400 841.200 510.450 907.950 ;
        RECT 508.950 839.100 511.050 841.200 ;
        RECT 514.950 839.100 517.050 841.200 ;
        RECT 509.400 838.350 510.600 839.100 ;
        RECT 515.400 829.050 516.450 839.100 ;
        RECT 514.950 826.950 517.050 829.050 ;
        RECT 598.950 826.950 601.050 829.050 ;
        RECT 599.400 775.050 600.450 826.950 ;
        RECT 725.400 800.400 726.600 802.650 ;
        RECT 725.400 775.050 726.450 800.400 ;
        RECT 598.950 772.950 601.050 775.050 ;
        RECT 685.950 772.950 688.050 775.050 ;
        RECT 724.950 772.950 727.050 775.050 ;
        RECT 599.400 763.050 600.450 772.950 ;
        RECT 598.950 760.950 601.050 763.050 ;
        RECT 686.400 762.600 687.450 772.950 ;
        RECT 686.400 760.350 687.600 762.600 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 584.400 691.050 585.450 757.950 ;
        RECT 532.950 688.950 535.050 691.050 ;
        RECT 571.950 688.950 574.050 691.050 ;
        RECT 583.950 688.950 586.050 691.050 ;
        RECT 533.400 684.600 534.450 688.950 ;
        RECT 572.400 684.600 573.450 688.950 ;
        RECT 533.400 682.350 534.600 684.600 ;
        RECT 572.400 682.350 573.600 684.600 ;
      LAYER metal3 ;
        RECT 499.950 939.600 502.050 940.050 ;
        RECT 550.950 939.600 553.050 940.050 ;
        RECT 499.950 938.400 553.050 939.600 ;
        RECT 499.950 937.950 502.050 938.400 ;
        RECT 550.950 937.950 553.050 938.400 ;
        RECT 508.950 909.600 511.050 910.050 ;
        RECT 550.950 909.600 553.050 910.050 ;
        RECT 508.950 908.400 553.050 909.600 ;
        RECT 508.950 907.950 511.050 908.400 ;
        RECT 550.950 907.950 553.050 908.400 ;
        RECT 508.950 840.750 511.050 841.200 ;
        RECT 514.950 840.750 517.050 841.200 ;
        RECT 508.950 839.550 517.050 840.750 ;
        RECT 508.950 839.100 511.050 839.550 ;
        RECT 514.950 839.100 517.050 839.550 ;
        RECT 514.950 828.600 517.050 829.050 ;
        RECT 598.950 828.600 601.050 829.050 ;
        RECT 514.950 827.400 601.050 828.600 ;
        RECT 514.950 826.950 517.050 827.400 ;
        RECT 598.950 826.950 601.050 827.400 ;
        RECT 598.950 774.600 601.050 775.050 ;
        RECT 685.950 774.600 688.050 775.050 ;
        RECT 724.950 774.600 727.050 775.050 ;
        RECT 598.950 773.400 727.050 774.600 ;
        RECT 598.950 772.950 601.050 773.400 ;
        RECT 685.950 772.950 688.050 773.400 ;
        RECT 724.950 772.950 727.050 773.400 ;
        RECT 598.950 762.600 601.050 763.050 ;
        RECT 584.400 762.000 601.050 762.600 ;
        RECT 583.950 761.400 601.050 762.000 ;
        RECT 583.950 757.950 586.050 761.400 ;
        RECT 598.950 760.950 601.050 761.400 ;
        RECT 532.950 690.600 535.050 691.050 ;
        RECT 571.950 690.600 574.050 691.050 ;
        RECT 583.950 690.600 586.050 691.050 ;
        RECT 532.950 689.400 586.050 690.600 ;
        RECT 532.950 688.950 535.050 689.400 ;
        RECT 571.950 688.950 574.050 689.400 ;
        RECT 583.950 688.950 586.050 689.400 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 434.400 944.400 438.450 945.450 ;
        RECT 434.400 916.050 435.450 944.400 ;
        RECT 433.950 913.950 436.050 916.050 ;
        RECT 439.950 913.950 442.050 916.050 ;
        RECT 440.400 885.600 441.450 913.950 ;
        RECT 440.400 883.350 441.600 885.600 ;
      LAYER metal3 ;
        RECT 433.950 915.600 436.050 916.050 ;
        RECT 439.950 915.600 442.050 916.050 ;
        RECT 433.950 914.400 442.050 915.600 ;
        RECT 433.950 913.950 436.050 914.400 ;
        RECT 439.950 913.950 442.050 914.400 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 14.100 929.400 15.900 936.000 ;
        RECT 17.100 929.400 18.900 935.400 ;
        RECT 14.100 916.050 15.900 917.850 ;
        RECT 17.100 916.050 18.300 929.400 ;
        RECT 32.100 924.300 33.900 935.400 ;
        RECT 35.100 925.500 36.900 936.000 ;
        RECT 32.100 923.400 36.600 924.300 ;
        RECT 39.600 923.400 41.400 935.400 ;
        RECT 44.100 925.500 45.900 936.000 ;
        RECT 47.100 924.600 48.900 935.400 ;
        RECT 62.100 929.400 63.900 936.000 ;
        RECT 65.100 929.400 66.900 935.400 ;
        RECT 68.100 930.000 69.900 936.000 ;
        RECT 65.400 929.100 66.900 929.400 ;
        RECT 71.100 929.400 72.900 935.400 ;
        RECT 83.100 929.400 84.900 936.000 ;
        RECT 86.100 929.400 87.900 935.400 ;
        RECT 89.100 930.000 90.900 936.000 ;
        RECT 71.100 929.100 72.000 929.400 ;
        RECT 65.400 928.200 72.000 929.100 ;
        RECT 86.400 929.100 87.900 929.400 ;
        RECT 92.100 929.400 93.900 935.400 ;
        RECT 107.100 929.400 108.900 936.000 ;
        RECT 110.100 929.400 111.900 935.400 ;
        RECT 113.100 929.400 114.900 936.000 ;
        RECT 128.100 929.400 129.900 936.000 ;
        RECT 131.100 929.400 132.900 935.400 ;
        RECT 143.100 929.400 144.900 936.000 ;
        RECT 146.100 929.400 147.900 935.400 ;
        RECT 149.100 930.000 150.900 936.000 ;
        RECT 92.100 929.100 93.000 929.400 ;
        RECT 86.400 928.200 93.000 929.100 ;
        RECT 34.500 921.300 36.600 923.400 ;
        RECT 40.200 922.050 41.400 923.400 ;
        RECT 44.100 923.400 48.900 924.600 ;
        RECT 44.100 922.500 46.200 923.400 ;
        RECT 40.200 921.000 41.700 922.050 ;
        RECT 37.800 919.500 39.900 919.800 ;
        RECT 36.000 917.700 39.900 919.500 ;
        RECT 40.800 919.050 41.700 921.000 ;
        RECT 40.800 916.950 42.900 919.050 ;
        RECT 40.800 916.800 42.300 916.950 ;
        RECT 37.200 916.050 39.000 916.500 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 32.100 914.700 39.000 916.050 ;
        RECT 39.900 915.900 42.300 916.800 ;
        RECT 46.800 916.050 48.600 917.850 ;
        RECT 65.100 916.050 66.900 917.850 ;
        RECT 71.100 916.050 72.000 928.200 ;
        RECT 76.950 921.450 79.050 922.050 ;
        RECT 88.950 921.450 91.050 922.050 ;
        RECT 76.950 920.550 91.050 921.450 ;
        RECT 76.950 919.950 79.050 920.550 ;
        RECT 88.950 919.950 91.050 920.550 ;
        RECT 86.100 916.050 87.900 917.850 ;
        RECT 92.100 916.050 93.000 928.200 ;
        RECT 110.100 916.050 111.300 929.400 ;
        RECT 128.100 916.050 129.900 917.850 ;
        RECT 131.100 916.050 132.300 929.400 ;
        RECT 146.400 929.100 147.900 929.400 ;
        RECT 152.100 929.400 153.900 935.400 ;
        RECT 164.100 929.400 165.900 936.000 ;
        RECT 167.100 929.400 168.900 935.400 ;
        RECT 170.100 929.400 171.900 936.000 ;
        RECT 185.700 929.400 187.500 936.000 ;
        RECT 152.100 929.100 153.000 929.400 ;
        RECT 146.400 928.200 153.000 929.100 ;
        RECT 133.950 918.450 138.000 919.050 ;
        RECT 133.950 916.950 138.450 918.450 ;
        RECT 32.100 913.950 34.200 914.700 ;
        RECT 17.100 903.600 18.300 913.950 ;
        RECT 32.400 912.150 34.200 913.950 ;
        RECT 37.200 911.400 39.000 913.200 ;
        RECT 36.900 909.300 39.000 911.400 ;
        RECT 32.700 908.400 39.000 909.300 ;
        RECT 39.900 910.200 41.100 915.900 ;
        RECT 42.300 913.200 44.100 915.000 ;
        RECT 46.800 913.950 48.900 916.050 ;
        RECT 61.950 913.950 64.050 916.050 ;
        RECT 64.950 913.950 67.050 916.050 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 82.950 913.950 85.050 916.050 ;
        RECT 85.950 913.950 88.050 916.050 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 106.950 913.950 109.050 916.050 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 127.950 913.950 130.050 916.050 ;
        RECT 130.950 913.950 133.050 916.050 ;
        RECT 42.000 911.100 44.100 913.200 ;
        RECT 62.100 912.150 63.900 913.950 ;
        RECT 68.100 912.150 69.900 913.950 ;
        RECT 71.100 910.200 72.000 913.950 ;
        RECT 83.100 912.150 84.900 913.950 ;
        RECT 89.100 912.150 90.900 913.950 ;
        RECT 92.100 910.200 93.000 913.950 ;
        RECT 107.250 912.150 109.050 913.950 ;
        RECT 32.700 906.600 33.900 908.400 ;
        RECT 39.900 908.100 42.900 910.200 ;
        RECT 39.900 906.600 41.100 908.100 ;
        RECT 44.100 907.500 46.200 908.700 ;
        RECT 44.100 906.600 48.900 907.500 ;
        RECT 14.100 900.000 15.900 903.600 ;
        RECT 17.100 900.600 18.900 903.600 ;
        RECT 32.100 900.600 33.900 906.600 ;
        RECT 35.100 900.000 36.900 905.700 ;
        RECT 39.600 900.600 41.400 906.600 ;
        RECT 44.100 900.000 45.900 905.700 ;
        RECT 47.100 900.600 48.900 906.600 ;
        RECT 62.100 900.000 63.900 909.600 ;
        RECT 68.700 909.000 72.000 910.200 ;
        RECT 68.700 900.600 70.500 909.000 ;
        RECT 83.100 900.000 84.900 909.600 ;
        RECT 89.700 909.000 93.000 910.200 ;
        RECT 89.700 900.600 91.500 909.000 ;
        RECT 110.100 908.700 111.300 913.950 ;
        RECT 113.100 912.150 114.900 913.950 ;
        RECT 110.100 907.800 114.300 908.700 ;
        RECT 107.400 900.000 109.200 906.600 ;
        RECT 112.500 900.600 114.300 907.800 ;
        RECT 131.100 903.600 132.300 913.950 ;
        RECT 137.550 912.450 138.450 916.950 ;
        RECT 146.100 916.050 147.900 917.850 ;
        RECT 152.100 916.050 153.000 928.200 ;
        RECT 167.700 916.050 168.900 929.400 ;
        RECT 186.000 926.100 187.800 927.900 ;
        RECT 188.700 924.900 190.500 935.400 ;
        RECT 188.100 923.400 190.500 924.900 ;
        RECT 193.800 923.400 195.600 936.000 ;
        RECT 209.100 929.400 210.900 936.000 ;
        RECT 212.100 929.400 213.900 935.400 ;
        RECT 215.100 929.400 216.900 936.000 ;
        RECT 227.100 929.400 228.900 936.000 ;
        RECT 230.100 929.400 231.900 935.400 ;
        RECT 233.100 930.000 234.900 936.000 ;
        RECT 188.100 916.050 189.300 923.400 ;
        RECT 199.950 918.450 202.050 919.050 ;
        RECT 205.950 918.450 208.050 919.050 ;
        RECT 194.100 916.050 195.900 917.850 ;
        RECT 199.950 917.550 208.050 918.450 ;
        RECT 199.950 916.950 202.050 917.550 ;
        RECT 205.950 916.950 208.050 917.550 ;
        RECT 212.100 916.050 213.300 929.400 ;
        RECT 230.400 929.100 231.900 929.400 ;
        RECT 236.100 929.400 237.900 935.400 ;
        RECT 251.100 929.400 252.900 936.000 ;
        RECT 254.100 929.400 255.900 935.400 ;
        RECT 257.100 930.000 258.900 936.000 ;
        RECT 236.100 929.100 237.000 929.400 ;
        RECT 230.400 928.200 237.000 929.100 ;
        RECT 254.400 929.100 255.900 929.400 ;
        RECT 260.100 929.400 261.900 935.400 ;
        RECT 275.100 929.400 276.900 936.000 ;
        RECT 278.100 929.400 279.900 935.400 ;
        RECT 281.100 929.400 282.900 936.000 ;
        RECT 260.100 929.100 261.000 929.400 ;
        RECT 254.400 928.200 261.000 929.100 ;
        RECT 230.100 916.050 231.900 917.850 ;
        RECT 236.100 916.050 237.000 928.200 ;
        RECT 254.100 916.050 255.900 917.850 ;
        RECT 260.100 916.050 261.000 928.200 ;
        RECT 278.700 916.050 279.900 929.400 ;
        RECT 296.100 923.400 297.900 935.400 ;
        RECT 300.600 923.400 302.400 936.000 ;
        RECT 303.600 924.900 305.400 935.400 ;
        RECT 303.600 923.400 306.000 924.900 ;
        RECT 296.100 921.900 297.300 923.400 ;
        RECT 296.100 920.700 303.900 921.900 ;
        RECT 302.100 920.100 303.900 920.700 ;
        RECT 300.000 916.050 301.800 917.850 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 148.950 913.950 151.050 916.050 ;
        RECT 151.950 913.950 154.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 166.950 913.950 169.050 916.050 ;
        RECT 169.950 913.950 172.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 190.950 913.950 193.050 916.050 ;
        RECT 193.950 913.950 196.050 916.050 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 211.950 913.950 214.050 916.050 ;
        RECT 214.950 913.950 217.050 916.050 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 235.950 913.950 238.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 256.950 913.950 259.050 916.050 ;
        RECT 259.950 913.950 262.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 280.950 913.950 283.050 916.050 ;
        RECT 296.100 913.950 298.200 916.050 ;
        RECT 299.400 913.950 301.500 916.050 ;
        RECT 137.550 912.000 141.450 912.450 ;
        RECT 143.100 912.150 144.900 913.950 ;
        RECT 149.100 912.150 150.900 913.950 ;
        RECT 137.550 911.550 142.050 912.000 ;
        RECT 139.950 907.950 142.050 911.550 ;
        RECT 152.100 910.200 153.000 913.950 ;
        RECT 164.100 912.150 165.900 913.950 ;
        RECT 133.950 906.900 138.000 907.050 ;
        RECT 133.950 904.950 139.050 906.900 ;
        RECT 136.950 904.800 139.050 904.950 ;
        RECT 128.100 900.000 129.900 903.600 ;
        RECT 131.100 900.600 132.900 903.600 ;
        RECT 143.100 900.000 144.900 909.600 ;
        RECT 149.700 909.000 153.000 910.200 ;
        RECT 149.700 900.600 151.500 909.000 ;
        RECT 167.700 908.700 168.900 913.950 ;
        RECT 169.950 912.150 171.750 913.950 ;
        RECT 185.100 912.150 186.900 913.950 ;
        RECT 188.100 909.600 189.300 913.950 ;
        RECT 191.100 912.150 192.900 913.950 ;
        RECT 209.250 912.150 211.050 913.950 ;
        RECT 164.700 907.800 168.900 908.700 ;
        RECT 185.700 908.700 189.300 909.600 ;
        RECT 212.100 908.700 213.300 913.950 ;
        RECT 215.100 912.150 216.900 913.950 ;
        RECT 227.100 912.150 228.900 913.950 ;
        RECT 233.100 912.150 234.900 913.950 ;
        RECT 236.100 910.200 237.000 913.950 ;
        RECT 238.950 912.450 241.050 913.050 ;
        RECT 244.950 912.450 247.050 913.050 ;
        RECT 238.950 911.550 247.050 912.450 ;
        RECT 251.100 912.150 252.900 913.950 ;
        RECT 257.100 912.150 258.900 913.950 ;
        RECT 238.950 910.950 241.050 911.550 ;
        RECT 244.950 910.950 247.050 911.550 ;
        RECT 260.100 910.200 261.000 913.950 ;
        RECT 275.100 912.150 276.900 913.950 ;
        RECT 164.700 900.600 166.500 907.800 ;
        RECT 185.700 906.600 186.900 908.700 ;
        RECT 212.100 907.800 216.300 908.700 ;
        RECT 169.800 900.000 171.600 906.600 ;
        RECT 185.100 900.600 186.900 906.600 ;
        RECT 188.100 905.700 195.900 907.050 ;
        RECT 188.100 900.600 189.900 905.700 ;
        RECT 191.100 900.000 192.900 904.800 ;
        RECT 194.100 900.600 195.900 905.700 ;
        RECT 209.400 900.000 211.200 906.600 ;
        RECT 214.500 900.600 216.300 907.800 ;
        RECT 227.100 900.000 228.900 909.600 ;
        RECT 233.700 909.000 237.000 910.200 ;
        RECT 233.700 900.600 235.500 909.000 ;
        RECT 251.100 900.000 252.900 909.600 ;
        RECT 257.700 909.000 261.000 910.200 ;
        RECT 257.700 900.600 259.500 909.000 ;
        RECT 278.700 908.700 279.900 913.950 ;
        RECT 280.950 912.150 282.750 913.950 ;
        RECT 296.400 912.150 298.200 913.950 ;
        RECT 302.700 909.600 303.600 920.100 ;
        RECT 304.800 916.050 306.000 923.400 ;
        RECT 317.100 923.400 318.900 935.400 ;
        RECT 320.100 925.200 321.900 936.000 ;
        RECT 323.100 929.400 324.900 935.400 ;
        RECT 338.100 929.400 339.900 936.000 ;
        RECT 341.100 929.400 342.900 935.400 ;
        RECT 344.700 929.400 346.500 936.000 ;
        RECT 347.700 929.400 349.500 935.400 ;
        RECT 351.000 929.400 352.800 936.000 ;
        RECT 354.000 929.400 355.800 935.400 ;
        RECT 357.000 929.400 358.800 936.000 ;
        RECT 360.000 929.400 361.800 935.400 ;
        RECT 363.000 929.400 364.800 936.000 ;
        RECT 366.000 932.400 367.800 935.400 ;
        RECT 369.000 932.400 370.800 935.400 ;
        RECT 372.000 932.400 373.800 935.400 ;
        RECT 365.700 930.300 367.800 932.400 ;
        RECT 368.700 930.300 370.800 932.400 ;
        RECT 371.700 930.300 373.800 932.400 ;
        RECT 375.000 929.400 376.800 935.400 ;
        RECT 378.000 929.400 379.800 936.000 ;
        RECT 317.100 916.050 318.300 923.400 ;
        RECT 323.700 922.500 324.900 929.400 ;
        RECT 319.200 921.600 324.900 922.500 ;
        RECT 319.200 920.700 321.000 921.600 ;
        RECT 304.800 913.950 306.900 916.050 ;
        RECT 302.700 908.700 304.800 909.600 ;
        RECT 275.700 907.800 279.900 908.700 ;
        RECT 299.400 907.800 304.800 908.700 ;
        RECT 275.700 900.600 277.500 907.800 ;
        RECT 280.800 900.000 282.600 906.600 ;
        RECT 299.400 903.600 300.300 907.800 ;
        RECT 306.000 906.600 306.900 913.950 ;
        RECT 296.100 900.600 297.900 903.600 ;
        RECT 299.100 900.600 300.900 903.600 ;
        RECT 296.100 900.000 297.300 900.600 ;
        RECT 302.100 900.000 303.900 906.000 ;
        RECT 305.100 900.600 306.900 906.600 ;
        RECT 317.100 913.950 319.200 916.050 ;
        RECT 317.100 906.600 318.300 913.950 ;
        RECT 320.100 909.300 321.000 920.700 ;
        RECT 322.800 916.050 324.600 917.850 ;
        RECT 338.100 916.050 339.900 917.850 ;
        RECT 341.100 916.050 342.300 929.400 ;
        RECT 348.000 919.050 349.500 929.400 ;
        RECT 354.000 928.500 355.200 929.400 ;
        RECT 347.100 916.950 349.500 919.050 ;
        RECT 322.500 913.950 324.600 916.050 ;
        RECT 337.950 913.950 340.050 916.050 ;
        RECT 340.950 913.950 343.050 916.050 ;
        RECT 319.200 908.400 321.000 909.300 ;
        RECT 319.200 907.500 324.900 908.400 ;
        RECT 317.100 900.600 318.900 906.600 ;
        RECT 320.100 900.000 321.900 906.600 ;
        RECT 323.700 903.600 324.900 907.500 ;
        RECT 341.100 903.600 342.300 913.950 ;
        RECT 348.000 903.600 349.500 916.950 ;
        RECT 323.100 900.600 324.900 903.600 ;
        RECT 338.100 900.000 339.900 903.600 ;
        RECT 341.100 900.600 342.900 903.600 ;
        RECT 344.700 900.000 346.500 903.600 ;
        RECT 347.700 900.600 349.500 903.600 ;
        RECT 351.300 927.600 355.200 928.500 ;
        RECT 351.300 924.300 352.200 927.600 ;
        RECT 356.100 926.400 357.900 927.000 ;
        RECT 360.600 926.400 361.800 929.400 ;
        RECT 368.700 928.500 370.800 929.400 ;
        RECT 362.700 927.300 370.800 928.500 ;
        RECT 362.700 926.700 364.500 927.300 ;
        RECT 356.100 925.200 361.800 926.400 ;
        RECT 374.100 925.500 376.800 929.400 ;
        RECT 381.000 927.900 382.800 935.400 ;
        RECT 384.900 929.400 386.700 936.000 ;
        RECT 387.900 929.400 389.700 935.400 ;
        RECT 390.900 932.400 392.700 935.400 ;
        RECT 393.900 932.400 395.700 935.400 ;
        RECT 390.600 930.300 392.700 932.400 ;
        RECT 393.600 930.300 395.700 932.400 ;
        RECT 397.500 929.400 399.300 936.000 ;
        RECT 379.500 925.800 382.800 927.900 ;
        RECT 388.200 927.300 390.300 929.400 ;
        RECT 400.500 926.400 402.300 935.400 ;
        RECT 403.500 929.400 405.300 936.000 ;
        RECT 406.500 930.300 408.300 935.400 ;
        RECT 406.500 929.400 408.600 930.300 ;
        RECT 409.500 929.400 411.300 936.000 ;
        RECT 425.100 929.400 426.900 935.400 ;
        RECT 407.700 928.500 408.600 929.400 ;
        RECT 407.700 927.600 411.300 928.500 ;
        RECT 405.000 926.400 406.800 926.700 ;
        RECT 365.700 924.300 367.800 925.500 ;
        RECT 351.300 923.400 367.800 924.300 ;
        RECT 371.100 924.600 373.200 925.500 ;
        RECT 387.600 925.200 406.800 926.400 ;
        RECT 387.600 924.600 388.800 925.200 ;
        RECT 405.000 924.900 406.800 925.200 ;
        RECT 371.100 923.400 388.800 924.600 ;
        RECT 391.500 923.700 393.600 924.300 ;
        RECT 401.700 923.700 403.500 924.300 ;
        RECT 351.300 906.600 352.200 923.400 ;
        RECT 391.500 922.500 403.500 923.700 ;
        RECT 353.100 921.300 388.800 922.500 ;
        RECT 391.500 922.200 393.600 922.500 ;
        RECT 353.100 920.700 354.900 921.300 ;
        RECT 387.600 920.700 388.800 921.300 ;
        RECT 356.100 916.950 358.200 919.050 ;
        RECT 356.700 914.100 358.200 916.950 ;
        RECT 360.300 916.800 365.400 918.600 ;
        RECT 364.500 915.300 365.400 916.800 ;
        RECT 368.100 918.300 369.900 920.100 ;
        RECT 374.100 919.800 376.200 920.100 ;
        RECT 387.600 919.800 401.100 920.700 ;
        RECT 368.100 917.100 369.000 918.300 ;
        RECT 374.100 918.000 378.000 919.800 ;
        RECT 379.500 918.300 381.600 919.200 ;
        RECT 399.300 919.050 401.100 919.800 ;
        RECT 379.500 917.100 390.600 918.300 ;
        RECT 399.300 917.250 403.200 919.050 ;
        RECT 368.100 916.200 381.600 917.100 ;
        RECT 388.800 916.500 390.600 917.100 ;
        RECT 401.100 916.950 403.200 917.250 ;
        RECT 407.100 916.950 409.200 919.050 ;
        RECT 407.100 915.300 408.900 916.950 ;
        RECT 364.500 914.100 408.900 915.300 ;
        RECT 356.700 912.600 363.300 914.100 ;
        RECT 353.100 909.900 360.900 911.700 ;
        RECT 361.800 911.100 378.900 912.600 ;
        RECT 376.800 910.500 378.900 911.100 ;
        RECT 383.100 912.000 385.200 913.050 ;
        RECT 383.100 911.100 388.200 912.000 ;
        RECT 391.800 911.400 393.600 913.200 ;
        RECT 410.100 911.400 411.300 927.600 ;
        RECT 425.100 922.500 426.300 929.400 ;
        RECT 428.100 925.200 429.900 936.000 ;
        RECT 431.100 923.400 432.900 935.400 ;
        RECT 434.700 929.400 436.500 936.000 ;
        RECT 437.700 929.400 439.500 935.400 ;
        RECT 441.000 929.400 442.800 936.000 ;
        RECT 444.000 929.400 445.800 935.400 ;
        RECT 447.000 929.400 448.800 936.000 ;
        RECT 450.000 929.400 451.800 935.400 ;
        RECT 453.000 929.400 454.800 936.000 ;
        RECT 456.000 932.400 457.800 935.400 ;
        RECT 459.000 932.400 460.800 935.400 ;
        RECT 462.000 932.400 463.800 935.400 ;
        RECT 455.700 930.300 457.800 932.400 ;
        RECT 458.700 930.300 460.800 932.400 ;
        RECT 461.700 930.300 463.800 932.400 ;
        RECT 465.000 929.400 466.800 935.400 ;
        RECT 468.000 929.400 469.800 936.000 ;
        RECT 425.100 921.600 430.800 922.500 ;
        RECT 429.000 920.700 430.800 921.600 ;
        RECT 425.400 916.050 427.200 917.850 ;
        RECT 425.400 913.950 427.500 916.050 ;
        RECT 383.100 910.950 385.200 911.100 ;
        RECT 359.400 906.600 360.900 909.900 ;
        RECT 377.100 908.700 378.900 910.500 ;
        RECT 386.400 910.200 388.200 911.100 ;
        RECT 392.700 908.400 393.600 911.400 ;
        RECT 394.500 910.200 411.300 911.400 ;
        RECT 394.500 909.300 396.600 910.200 ;
        RECT 405.300 908.700 407.100 909.300 ;
        RECT 365.100 906.600 371.700 908.400 ;
        RECT 386.400 907.200 393.600 908.400 ;
        RECT 398.700 907.500 407.100 908.700 ;
        RECT 386.400 906.600 387.300 907.200 ;
        RECT 389.400 906.600 391.200 907.200 ;
        RECT 398.700 906.600 400.200 907.500 ;
        RECT 410.100 906.600 411.300 910.200 ;
        RECT 429.000 909.300 429.900 920.700 ;
        RECT 431.700 916.050 432.900 923.400 ;
        RECT 438.000 919.050 439.500 929.400 ;
        RECT 444.000 928.500 445.200 929.400 ;
        RECT 437.100 916.950 439.500 919.050 ;
        RECT 430.800 913.950 432.900 916.050 ;
        RECT 429.000 908.400 430.800 909.300 ;
        RECT 351.300 900.600 353.100 906.600 ;
        RECT 356.700 900.000 358.500 906.600 ;
        RECT 359.400 905.400 363.600 906.600 ;
        RECT 361.800 900.600 363.600 905.400 ;
        RECT 365.700 903.600 367.800 905.700 ;
        RECT 368.700 903.600 370.800 905.700 ;
        RECT 371.700 903.600 373.800 905.700 ;
        RECT 374.700 903.600 376.800 905.700 ;
        RECT 380.100 904.500 382.800 906.600 ;
        RECT 384.600 905.400 387.300 906.600 ;
        RECT 384.600 904.500 386.400 905.400 ;
        RECT 366.000 900.600 367.800 903.600 ;
        RECT 369.000 900.600 370.800 903.600 ;
        RECT 372.000 900.600 373.800 903.600 ;
        RECT 375.000 900.600 376.800 903.600 ;
        RECT 378.000 900.000 379.800 903.600 ;
        RECT 381.000 900.600 382.800 904.500 ;
        RECT 388.200 903.600 390.300 905.700 ;
        RECT 391.200 903.600 393.300 905.700 ;
        RECT 394.200 903.600 396.300 905.700 ;
        RECT 385.500 900.000 387.300 903.600 ;
        RECT 388.500 900.600 390.300 903.600 ;
        RECT 391.500 900.600 393.300 903.600 ;
        RECT 394.500 900.600 396.300 903.600 ;
        RECT 398.700 900.600 400.500 906.600 ;
        RECT 404.100 900.000 405.900 906.600 ;
        RECT 409.500 900.600 411.300 906.600 ;
        RECT 425.100 907.500 430.800 908.400 ;
        RECT 425.100 903.600 426.300 907.500 ;
        RECT 431.700 906.600 432.900 913.950 ;
        RECT 425.100 900.600 426.900 903.600 ;
        RECT 428.100 900.000 429.900 906.600 ;
        RECT 431.100 900.600 432.900 906.600 ;
        RECT 438.000 903.600 439.500 916.950 ;
        RECT 434.700 900.000 436.500 903.600 ;
        RECT 437.700 900.600 439.500 903.600 ;
        RECT 441.300 927.600 445.200 928.500 ;
        RECT 441.300 924.300 442.200 927.600 ;
        RECT 446.100 926.400 447.900 927.000 ;
        RECT 450.600 926.400 451.800 929.400 ;
        RECT 458.700 928.500 460.800 929.400 ;
        RECT 452.700 927.300 460.800 928.500 ;
        RECT 452.700 926.700 454.500 927.300 ;
        RECT 446.100 925.200 451.800 926.400 ;
        RECT 464.100 925.500 466.800 929.400 ;
        RECT 471.000 927.900 472.800 935.400 ;
        RECT 474.900 929.400 476.700 936.000 ;
        RECT 477.900 929.400 479.700 935.400 ;
        RECT 480.900 932.400 482.700 935.400 ;
        RECT 483.900 932.400 485.700 935.400 ;
        RECT 480.600 930.300 482.700 932.400 ;
        RECT 483.600 930.300 485.700 932.400 ;
        RECT 487.500 929.400 489.300 936.000 ;
        RECT 469.500 925.800 472.800 927.900 ;
        RECT 478.200 927.300 480.300 929.400 ;
        RECT 490.500 926.400 492.300 935.400 ;
        RECT 493.500 929.400 495.300 936.000 ;
        RECT 496.500 930.300 498.300 935.400 ;
        RECT 496.500 929.400 498.600 930.300 ;
        RECT 499.500 929.400 501.300 936.000 ;
        RECT 503.700 929.400 505.500 936.000 ;
        RECT 506.700 930.300 508.500 935.400 ;
        RECT 506.400 929.400 508.500 930.300 ;
        RECT 509.700 929.400 511.500 936.000 ;
        RECT 497.700 928.500 498.600 929.400 ;
        RECT 506.400 928.500 507.300 929.400 ;
        RECT 497.700 927.600 501.300 928.500 ;
        RECT 495.000 926.400 496.800 926.700 ;
        RECT 455.700 924.300 457.800 925.500 ;
        RECT 441.300 923.400 457.800 924.300 ;
        RECT 461.100 924.600 463.200 925.500 ;
        RECT 477.600 925.200 496.800 926.400 ;
        RECT 477.600 924.600 478.800 925.200 ;
        RECT 495.000 924.900 496.800 925.200 ;
        RECT 461.100 923.400 478.800 924.600 ;
        RECT 481.500 923.700 483.600 924.300 ;
        RECT 491.700 923.700 493.500 924.300 ;
        RECT 441.300 906.600 442.200 923.400 ;
        RECT 481.500 922.500 493.500 923.700 ;
        RECT 443.100 921.300 478.800 922.500 ;
        RECT 481.500 922.200 483.600 922.500 ;
        RECT 443.100 920.700 444.900 921.300 ;
        RECT 477.600 920.700 478.800 921.300 ;
        RECT 446.100 916.950 448.200 919.050 ;
        RECT 446.700 914.100 448.200 916.950 ;
        RECT 450.300 916.800 455.400 918.600 ;
        RECT 454.500 915.300 455.400 916.800 ;
        RECT 458.100 918.300 459.900 920.100 ;
        RECT 464.100 919.800 466.200 920.100 ;
        RECT 477.600 919.800 491.100 920.700 ;
        RECT 458.100 917.100 459.000 918.300 ;
        RECT 464.100 918.000 468.000 919.800 ;
        RECT 469.500 918.300 471.600 919.200 ;
        RECT 489.300 919.050 491.100 919.800 ;
        RECT 469.500 917.100 480.600 918.300 ;
        RECT 489.300 917.250 493.200 919.050 ;
        RECT 458.100 916.200 471.600 917.100 ;
        RECT 478.800 916.500 480.600 917.100 ;
        RECT 491.100 916.950 493.200 917.250 ;
        RECT 497.100 916.950 499.200 919.050 ;
        RECT 497.100 915.300 498.900 916.950 ;
        RECT 454.500 914.100 498.900 915.300 ;
        RECT 446.700 912.600 453.300 914.100 ;
        RECT 443.100 909.900 450.900 911.700 ;
        RECT 451.800 911.100 468.900 912.600 ;
        RECT 466.800 910.500 468.900 911.100 ;
        RECT 473.100 912.000 475.200 913.050 ;
        RECT 473.100 911.100 478.200 912.000 ;
        RECT 481.800 911.400 483.600 913.200 ;
        RECT 500.100 911.400 501.300 927.600 ;
        RECT 473.100 910.950 475.200 911.100 ;
        RECT 449.400 906.600 450.900 909.900 ;
        RECT 467.100 908.700 468.900 910.500 ;
        RECT 476.400 910.200 478.200 911.100 ;
        RECT 482.700 908.400 483.600 911.400 ;
        RECT 484.500 910.200 501.300 911.400 ;
        RECT 484.500 909.300 486.600 910.200 ;
        RECT 495.300 908.700 497.100 909.300 ;
        RECT 455.100 906.600 461.700 908.400 ;
        RECT 476.400 907.200 483.600 908.400 ;
        RECT 488.700 907.500 497.100 908.700 ;
        RECT 476.400 906.600 477.300 907.200 ;
        RECT 479.400 906.600 481.200 907.200 ;
        RECT 488.700 906.600 490.200 907.500 ;
        RECT 500.100 906.600 501.300 910.200 ;
        RECT 441.300 900.600 443.100 906.600 ;
        RECT 446.700 900.000 448.500 906.600 ;
        RECT 449.400 905.400 453.600 906.600 ;
        RECT 451.800 900.600 453.600 905.400 ;
        RECT 455.700 903.600 457.800 905.700 ;
        RECT 458.700 903.600 460.800 905.700 ;
        RECT 461.700 903.600 463.800 905.700 ;
        RECT 464.700 903.600 466.800 905.700 ;
        RECT 470.100 904.500 472.800 906.600 ;
        RECT 474.600 905.400 477.300 906.600 ;
        RECT 474.600 904.500 476.400 905.400 ;
        RECT 456.000 900.600 457.800 903.600 ;
        RECT 459.000 900.600 460.800 903.600 ;
        RECT 462.000 900.600 463.800 903.600 ;
        RECT 465.000 900.600 466.800 903.600 ;
        RECT 468.000 900.000 469.800 903.600 ;
        RECT 471.000 900.600 472.800 904.500 ;
        RECT 478.200 903.600 480.300 905.700 ;
        RECT 481.200 903.600 483.300 905.700 ;
        RECT 484.200 903.600 486.300 905.700 ;
        RECT 475.500 900.000 477.300 903.600 ;
        RECT 478.500 900.600 480.300 903.600 ;
        RECT 481.500 900.600 483.300 903.600 ;
        RECT 484.500 900.600 486.300 903.600 ;
        RECT 488.700 900.600 490.500 906.600 ;
        RECT 494.100 900.000 495.900 906.600 ;
        RECT 499.500 900.600 501.300 906.600 ;
        RECT 503.700 927.600 507.300 928.500 ;
        RECT 503.700 911.400 504.900 927.600 ;
        RECT 508.200 926.400 510.000 926.700 ;
        RECT 512.700 926.400 514.500 935.400 ;
        RECT 515.700 929.400 517.500 936.000 ;
        RECT 519.300 932.400 521.100 935.400 ;
        RECT 522.300 932.400 524.100 935.400 ;
        RECT 519.300 930.300 521.400 932.400 ;
        RECT 522.300 930.300 524.400 932.400 ;
        RECT 525.300 929.400 527.100 935.400 ;
        RECT 528.300 929.400 530.100 936.000 ;
        RECT 524.700 927.300 526.800 929.400 ;
        RECT 532.200 927.900 534.000 935.400 ;
        RECT 535.200 929.400 537.000 936.000 ;
        RECT 538.200 929.400 540.000 935.400 ;
        RECT 541.200 932.400 543.000 935.400 ;
        RECT 544.200 932.400 546.000 935.400 ;
        RECT 547.200 932.400 549.000 935.400 ;
        RECT 541.200 930.300 543.300 932.400 ;
        RECT 544.200 930.300 546.300 932.400 ;
        RECT 547.200 930.300 549.300 932.400 ;
        RECT 550.200 929.400 552.000 936.000 ;
        RECT 553.200 929.400 555.000 935.400 ;
        RECT 556.200 929.400 558.000 936.000 ;
        RECT 559.200 929.400 561.000 935.400 ;
        RECT 562.200 929.400 564.000 936.000 ;
        RECT 565.500 929.400 567.300 935.400 ;
        RECT 568.500 929.400 570.300 936.000 ;
        RECT 584.100 929.400 585.900 935.400 ;
        RECT 508.200 925.200 527.400 926.400 ;
        RECT 532.200 925.800 535.500 927.900 ;
        RECT 538.200 925.500 540.900 929.400 ;
        RECT 544.200 928.500 546.300 929.400 ;
        RECT 544.200 927.300 552.300 928.500 ;
        RECT 550.500 926.700 552.300 927.300 ;
        RECT 553.200 926.400 554.400 929.400 ;
        RECT 559.800 928.500 561.000 929.400 ;
        RECT 559.800 927.600 563.700 928.500 ;
        RECT 557.100 926.400 558.900 927.000 ;
        RECT 508.200 924.900 510.000 925.200 ;
        RECT 526.200 924.600 527.400 925.200 ;
        RECT 541.800 924.600 543.900 925.500 ;
        RECT 511.500 923.700 513.300 924.300 ;
        RECT 521.400 923.700 523.500 924.300 ;
        RECT 511.500 922.500 523.500 923.700 ;
        RECT 526.200 923.400 543.900 924.600 ;
        RECT 547.200 924.300 549.300 925.500 ;
        RECT 553.200 925.200 558.900 926.400 ;
        RECT 562.800 924.300 563.700 927.600 ;
        RECT 547.200 923.400 563.700 924.300 ;
        RECT 521.400 922.200 523.500 922.500 ;
        RECT 526.200 921.300 561.900 922.500 ;
        RECT 526.200 920.700 527.400 921.300 ;
        RECT 560.100 920.700 561.900 921.300 ;
        RECT 513.900 919.800 527.400 920.700 ;
        RECT 538.800 919.800 540.900 920.100 ;
        RECT 513.900 919.050 515.700 919.800 ;
        RECT 505.800 916.950 507.900 919.050 ;
        RECT 511.800 917.250 515.700 919.050 ;
        RECT 533.400 918.300 535.500 919.200 ;
        RECT 511.800 916.950 513.900 917.250 ;
        RECT 524.400 917.100 535.500 918.300 ;
        RECT 537.000 918.000 540.900 919.800 ;
        RECT 545.100 918.300 546.900 920.100 ;
        RECT 546.000 917.100 546.900 918.300 ;
        RECT 506.100 915.300 507.900 916.950 ;
        RECT 524.400 916.500 526.200 917.100 ;
        RECT 533.400 916.200 546.900 917.100 ;
        RECT 549.600 916.800 554.700 918.600 ;
        RECT 556.800 916.950 558.900 919.050 ;
        RECT 549.600 915.300 550.500 916.800 ;
        RECT 506.100 914.100 550.500 915.300 ;
        RECT 556.800 914.100 558.300 916.950 ;
        RECT 521.400 911.400 523.200 913.200 ;
        RECT 529.800 912.000 531.900 913.050 ;
        RECT 551.700 912.600 558.300 914.100 ;
        RECT 503.700 910.200 520.500 911.400 ;
        RECT 503.700 906.600 504.900 910.200 ;
        RECT 518.400 909.300 520.500 910.200 ;
        RECT 507.900 908.700 509.700 909.300 ;
        RECT 507.900 907.500 516.300 908.700 ;
        RECT 514.800 906.600 516.300 907.500 ;
        RECT 521.400 908.400 522.300 911.400 ;
        RECT 526.800 911.100 531.900 912.000 ;
        RECT 526.800 910.200 528.600 911.100 ;
        RECT 529.800 910.950 531.900 911.100 ;
        RECT 536.100 911.100 553.200 912.600 ;
        RECT 536.100 910.500 538.200 911.100 ;
        RECT 536.100 908.700 537.900 910.500 ;
        RECT 554.100 909.900 561.900 911.700 ;
        RECT 521.400 907.200 528.600 908.400 ;
        RECT 523.800 906.600 525.600 907.200 ;
        RECT 527.700 906.600 528.600 907.200 ;
        RECT 543.300 906.600 549.900 908.400 ;
        RECT 554.100 906.600 555.600 909.900 ;
        RECT 562.800 906.600 563.700 923.400 ;
        RECT 503.700 900.600 505.500 906.600 ;
        RECT 509.100 900.000 510.900 906.600 ;
        RECT 514.500 900.600 516.300 906.600 ;
        RECT 518.700 903.600 520.800 905.700 ;
        RECT 521.700 903.600 523.800 905.700 ;
        RECT 524.700 903.600 526.800 905.700 ;
        RECT 527.700 905.400 530.400 906.600 ;
        RECT 528.600 904.500 530.400 905.400 ;
        RECT 532.200 904.500 534.900 906.600 ;
        RECT 518.700 900.600 520.500 903.600 ;
        RECT 521.700 900.600 523.500 903.600 ;
        RECT 524.700 900.600 526.500 903.600 ;
        RECT 527.700 900.000 529.500 903.600 ;
        RECT 532.200 900.600 534.000 904.500 ;
        RECT 538.200 903.600 540.300 905.700 ;
        RECT 541.200 903.600 543.300 905.700 ;
        RECT 544.200 903.600 546.300 905.700 ;
        RECT 547.200 903.600 549.300 905.700 ;
        RECT 551.400 905.400 555.600 906.600 ;
        RECT 535.200 900.000 537.000 903.600 ;
        RECT 538.200 900.600 540.000 903.600 ;
        RECT 541.200 900.600 543.000 903.600 ;
        RECT 544.200 900.600 546.000 903.600 ;
        RECT 547.200 900.600 549.000 903.600 ;
        RECT 551.400 900.600 553.200 905.400 ;
        RECT 556.500 900.000 558.300 906.600 ;
        RECT 561.900 900.600 563.700 906.600 ;
        RECT 565.500 919.050 567.000 929.400 ;
        RECT 584.100 922.500 585.300 929.400 ;
        RECT 587.100 925.200 588.900 936.000 ;
        RECT 590.100 923.400 591.900 935.400 ;
        RECT 593.700 929.400 595.500 936.000 ;
        RECT 596.700 930.300 598.500 935.400 ;
        RECT 596.400 929.400 598.500 930.300 ;
        RECT 599.700 929.400 601.500 936.000 ;
        RECT 596.400 928.500 597.300 929.400 ;
        RECT 584.100 921.600 589.800 922.500 ;
        RECT 588.000 920.700 589.800 921.600 ;
        RECT 565.500 916.950 567.900 919.050 ;
        RECT 565.500 903.600 567.000 916.950 ;
        RECT 584.400 916.050 586.200 917.850 ;
        RECT 584.400 913.950 586.500 916.050 ;
        RECT 588.000 909.300 588.900 920.700 ;
        RECT 590.700 916.050 591.900 923.400 ;
        RECT 589.800 913.950 591.900 916.050 ;
        RECT 588.000 908.400 589.800 909.300 ;
        RECT 584.100 907.500 589.800 908.400 ;
        RECT 584.100 903.600 585.300 907.500 ;
        RECT 590.700 906.600 591.900 913.950 ;
        RECT 565.500 900.600 567.300 903.600 ;
        RECT 568.500 900.000 570.300 903.600 ;
        RECT 584.100 900.600 585.900 903.600 ;
        RECT 587.100 900.000 588.900 906.600 ;
        RECT 590.100 900.600 591.900 906.600 ;
        RECT 593.700 927.600 597.300 928.500 ;
        RECT 593.700 911.400 594.900 927.600 ;
        RECT 598.200 926.400 600.000 926.700 ;
        RECT 602.700 926.400 604.500 935.400 ;
        RECT 605.700 929.400 607.500 936.000 ;
        RECT 609.300 932.400 611.100 935.400 ;
        RECT 612.300 932.400 614.100 935.400 ;
        RECT 609.300 930.300 611.400 932.400 ;
        RECT 612.300 930.300 614.400 932.400 ;
        RECT 615.300 929.400 617.100 935.400 ;
        RECT 618.300 929.400 620.100 936.000 ;
        RECT 614.700 927.300 616.800 929.400 ;
        RECT 622.200 927.900 624.000 935.400 ;
        RECT 625.200 929.400 627.000 936.000 ;
        RECT 628.200 929.400 630.000 935.400 ;
        RECT 631.200 932.400 633.000 935.400 ;
        RECT 634.200 932.400 636.000 935.400 ;
        RECT 637.200 932.400 639.000 935.400 ;
        RECT 631.200 930.300 633.300 932.400 ;
        RECT 634.200 930.300 636.300 932.400 ;
        RECT 637.200 930.300 639.300 932.400 ;
        RECT 640.200 929.400 642.000 936.000 ;
        RECT 643.200 929.400 645.000 935.400 ;
        RECT 646.200 929.400 648.000 936.000 ;
        RECT 649.200 929.400 651.000 935.400 ;
        RECT 652.200 929.400 654.000 936.000 ;
        RECT 655.500 929.400 657.300 935.400 ;
        RECT 658.500 929.400 660.300 936.000 ;
        RECT 671.100 929.400 672.900 936.000 ;
        RECT 674.100 929.400 675.900 935.400 ;
        RECT 598.200 925.200 617.400 926.400 ;
        RECT 622.200 925.800 625.500 927.900 ;
        RECT 628.200 925.500 630.900 929.400 ;
        RECT 634.200 928.500 636.300 929.400 ;
        RECT 634.200 927.300 642.300 928.500 ;
        RECT 640.500 926.700 642.300 927.300 ;
        RECT 643.200 926.400 644.400 929.400 ;
        RECT 649.800 928.500 651.000 929.400 ;
        RECT 649.800 927.600 653.700 928.500 ;
        RECT 647.100 926.400 648.900 927.000 ;
        RECT 598.200 924.900 600.000 925.200 ;
        RECT 616.200 924.600 617.400 925.200 ;
        RECT 631.800 924.600 633.900 925.500 ;
        RECT 601.500 923.700 603.300 924.300 ;
        RECT 611.400 923.700 613.500 924.300 ;
        RECT 601.500 922.500 613.500 923.700 ;
        RECT 616.200 923.400 633.900 924.600 ;
        RECT 637.200 924.300 639.300 925.500 ;
        RECT 643.200 925.200 648.900 926.400 ;
        RECT 652.800 924.300 653.700 927.600 ;
        RECT 637.200 923.400 653.700 924.300 ;
        RECT 611.400 922.200 613.500 922.500 ;
        RECT 616.200 921.300 651.900 922.500 ;
        RECT 616.200 920.700 617.400 921.300 ;
        RECT 650.100 920.700 651.900 921.300 ;
        RECT 603.900 919.800 617.400 920.700 ;
        RECT 628.800 919.800 630.900 920.100 ;
        RECT 603.900 919.050 605.700 919.800 ;
        RECT 595.800 916.950 597.900 919.050 ;
        RECT 601.800 917.250 605.700 919.050 ;
        RECT 623.400 918.300 625.500 919.200 ;
        RECT 601.800 916.950 603.900 917.250 ;
        RECT 614.400 917.100 625.500 918.300 ;
        RECT 627.000 918.000 630.900 919.800 ;
        RECT 635.100 918.300 636.900 920.100 ;
        RECT 636.000 917.100 636.900 918.300 ;
        RECT 596.100 915.300 597.900 916.950 ;
        RECT 614.400 916.500 616.200 917.100 ;
        RECT 623.400 916.200 636.900 917.100 ;
        RECT 639.600 916.800 644.700 918.600 ;
        RECT 646.800 916.950 648.900 919.050 ;
        RECT 639.600 915.300 640.500 916.800 ;
        RECT 596.100 914.100 640.500 915.300 ;
        RECT 646.800 914.100 648.300 916.950 ;
        RECT 611.400 911.400 613.200 913.200 ;
        RECT 619.800 912.000 621.900 913.050 ;
        RECT 641.700 912.600 648.300 914.100 ;
        RECT 593.700 910.200 610.500 911.400 ;
        RECT 593.700 906.600 594.900 910.200 ;
        RECT 608.400 909.300 610.500 910.200 ;
        RECT 597.900 908.700 599.700 909.300 ;
        RECT 597.900 907.500 606.300 908.700 ;
        RECT 604.800 906.600 606.300 907.500 ;
        RECT 611.400 908.400 612.300 911.400 ;
        RECT 616.800 911.100 621.900 912.000 ;
        RECT 616.800 910.200 618.600 911.100 ;
        RECT 619.800 910.950 621.900 911.100 ;
        RECT 626.100 911.100 643.200 912.600 ;
        RECT 626.100 910.500 628.200 911.100 ;
        RECT 626.100 908.700 627.900 910.500 ;
        RECT 644.100 909.900 651.900 911.700 ;
        RECT 611.400 907.200 618.600 908.400 ;
        RECT 613.800 906.600 615.600 907.200 ;
        RECT 617.700 906.600 618.600 907.200 ;
        RECT 633.300 906.600 639.900 908.400 ;
        RECT 644.100 906.600 645.600 909.900 ;
        RECT 652.800 906.600 653.700 923.400 ;
        RECT 593.700 900.600 595.500 906.600 ;
        RECT 599.100 900.000 600.900 906.600 ;
        RECT 604.500 900.600 606.300 906.600 ;
        RECT 608.700 903.600 610.800 905.700 ;
        RECT 611.700 903.600 613.800 905.700 ;
        RECT 614.700 903.600 616.800 905.700 ;
        RECT 617.700 905.400 620.400 906.600 ;
        RECT 618.600 904.500 620.400 905.400 ;
        RECT 622.200 904.500 624.900 906.600 ;
        RECT 608.700 900.600 610.500 903.600 ;
        RECT 611.700 900.600 613.500 903.600 ;
        RECT 614.700 900.600 616.500 903.600 ;
        RECT 617.700 900.000 619.500 903.600 ;
        RECT 622.200 900.600 624.000 904.500 ;
        RECT 628.200 903.600 630.300 905.700 ;
        RECT 631.200 903.600 633.300 905.700 ;
        RECT 634.200 903.600 636.300 905.700 ;
        RECT 637.200 903.600 639.300 905.700 ;
        RECT 641.400 905.400 645.600 906.600 ;
        RECT 625.200 900.000 627.000 903.600 ;
        RECT 628.200 900.600 630.000 903.600 ;
        RECT 631.200 900.600 633.000 903.600 ;
        RECT 634.200 900.600 636.000 903.600 ;
        RECT 637.200 900.600 639.000 903.600 ;
        RECT 641.400 900.600 643.200 905.400 ;
        RECT 646.500 900.000 648.300 906.600 ;
        RECT 651.900 900.600 653.700 906.600 ;
        RECT 655.500 919.050 657.000 929.400 ;
        RECT 655.500 916.950 657.900 919.050 ;
        RECT 655.500 903.600 657.000 916.950 ;
        RECT 671.100 916.050 672.900 917.850 ;
        RECT 674.100 916.050 675.300 929.400 ;
        RECT 686.100 923.400 687.900 935.400 ;
        RECT 689.100 925.200 690.900 936.000 ;
        RECT 692.100 929.400 693.900 935.400 ;
        RECT 686.100 916.050 687.300 923.400 ;
        RECT 692.700 922.500 693.900 929.400 ;
        RECT 688.200 921.600 693.900 922.500 ;
        RECT 707.100 929.400 708.900 935.400 ;
        RECT 707.100 922.500 708.300 929.400 ;
        RECT 710.100 925.200 711.900 936.000 ;
        RECT 713.100 923.400 714.900 935.400 ;
        RECT 716.700 929.400 718.500 936.000 ;
        RECT 719.700 929.400 721.500 935.400 ;
        RECT 723.000 929.400 724.800 936.000 ;
        RECT 726.000 929.400 727.800 935.400 ;
        RECT 729.000 929.400 730.800 936.000 ;
        RECT 732.000 929.400 733.800 935.400 ;
        RECT 735.000 929.400 736.800 936.000 ;
        RECT 738.000 932.400 739.800 935.400 ;
        RECT 741.000 932.400 742.800 935.400 ;
        RECT 744.000 932.400 745.800 935.400 ;
        RECT 737.700 930.300 739.800 932.400 ;
        RECT 740.700 930.300 742.800 932.400 ;
        RECT 743.700 930.300 745.800 932.400 ;
        RECT 747.000 929.400 748.800 935.400 ;
        RECT 750.000 929.400 751.800 936.000 ;
        RECT 707.100 921.600 712.800 922.500 ;
        RECT 688.200 920.700 690.000 921.600 ;
        RECT 670.950 913.950 673.050 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 686.100 913.950 688.200 916.050 ;
        RECT 674.100 903.600 675.300 913.950 ;
        RECT 686.100 906.600 687.300 913.950 ;
        RECT 689.100 909.300 690.000 920.700 ;
        RECT 711.000 920.700 712.800 921.600 ;
        RECT 691.800 916.050 693.600 917.850 ;
        RECT 691.500 913.950 693.600 916.050 ;
        RECT 707.400 916.050 709.200 917.850 ;
        RECT 707.400 913.950 709.500 916.050 ;
        RECT 688.200 908.400 690.000 909.300 ;
        RECT 711.000 909.300 711.900 920.700 ;
        RECT 713.700 916.050 714.900 923.400 ;
        RECT 720.000 919.050 721.500 929.400 ;
        RECT 726.000 928.500 727.200 929.400 ;
        RECT 719.100 916.950 721.500 919.050 ;
        RECT 712.800 913.950 714.900 916.050 ;
        RECT 711.000 908.400 712.800 909.300 ;
        RECT 688.200 907.500 693.900 908.400 ;
        RECT 655.500 900.600 657.300 903.600 ;
        RECT 658.500 900.000 660.300 903.600 ;
        RECT 671.100 900.000 672.900 903.600 ;
        RECT 674.100 900.600 675.900 903.600 ;
        RECT 686.100 900.600 687.900 906.600 ;
        RECT 689.100 900.000 690.900 906.600 ;
        RECT 692.700 903.600 693.900 907.500 ;
        RECT 692.100 900.600 693.900 903.600 ;
        RECT 707.100 907.500 712.800 908.400 ;
        RECT 707.100 903.600 708.300 907.500 ;
        RECT 713.700 906.600 714.900 913.950 ;
        RECT 707.100 900.600 708.900 903.600 ;
        RECT 710.100 900.000 711.900 906.600 ;
        RECT 713.100 900.600 714.900 906.600 ;
        RECT 720.000 903.600 721.500 916.950 ;
        RECT 716.700 900.000 718.500 903.600 ;
        RECT 719.700 900.600 721.500 903.600 ;
        RECT 723.300 927.600 727.200 928.500 ;
        RECT 723.300 924.300 724.200 927.600 ;
        RECT 728.100 926.400 729.900 927.000 ;
        RECT 732.600 926.400 733.800 929.400 ;
        RECT 740.700 928.500 742.800 929.400 ;
        RECT 734.700 927.300 742.800 928.500 ;
        RECT 734.700 926.700 736.500 927.300 ;
        RECT 728.100 925.200 733.800 926.400 ;
        RECT 746.100 925.500 748.800 929.400 ;
        RECT 753.000 927.900 754.800 935.400 ;
        RECT 756.900 929.400 758.700 936.000 ;
        RECT 759.900 929.400 761.700 935.400 ;
        RECT 762.900 932.400 764.700 935.400 ;
        RECT 765.900 932.400 767.700 935.400 ;
        RECT 762.600 930.300 764.700 932.400 ;
        RECT 765.600 930.300 767.700 932.400 ;
        RECT 769.500 929.400 771.300 936.000 ;
        RECT 751.500 925.800 754.800 927.900 ;
        RECT 760.200 927.300 762.300 929.400 ;
        RECT 772.500 926.400 774.300 935.400 ;
        RECT 775.500 929.400 777.300 936.000 ;
        RECT 778.500 930.300 780.300 935.400 ;
        RECT 778.500 929.400 780.600 930.300 ;
        RECT 781.500 929.400 783.300 936.000 ;
        RECT 779.700 928.500 780.600 929.400 ;
        RECT 779.700 927.600 783.300 928.500 ;
        RECT 777.000 926.400 778.800 926.700 ;
        RECT 737.700 924.300 739.800 925.500 ;
        RECT 723.300 923.400 739.800 924.300 ;
        RECT 743.100 924.600 745.200 925.500 ;
        RECT 759.600 925.200 778.800 926.400 ;
        RECT 759.600 924.600 760.800 925.200 ;
        RECT 777.000 924.900 778.800 925.200 ;
        RECT 743.100 923.400 760.800 924.600 ;
        RECT 763.500 923.700 765.600 924.300 ;
        RECT 773.700 923.700 775.500 924.300 ;
        RECT 723.300 906.600 724.200 923.400 ;
        RECT 763.500 922.500 775.500 923.700 ;
        RECT 725.100 921.300 760.800 922.500 ;
        RECT 763.500 922.200 765.600 922.500 ;
        RECT 725.100 920.700 726.900 921.300 ;
        RECT 759.600 920.700 760.800 921.300 ;
        RECT 728.100 916.950 730.200 919.050 ;
        RECT 728.700 914.100 730.200 916.950 ;
        RECT 732.300 916.800 737.400 918.600 ;
        RECT 736.500 915.300 737.400 916.800 ;
        RECT 740.100 918.300 741.900 920.100 ;
        RECT 746.100 919.800 748.200 920.100 ;
        RECT 759.600 919.800 773.100 920.700 ;
        RECT 740.100 917.100 741.000 918.300 ;
        RECT 746.100 918.000 750.000 919.800 ;
        RECT 751.500 918.300 753.600 919.200 ;
        RECT 771.300 919.050 773.100 919.800 ;
        RECT 751.500 917.100 762.600 918.300 ;
        RECT 771.300 917.250 775.200 919.050 ;
        RECT 740.100 916.200 753.600 917.100 ;
        RECT 760.800 916.500 762.600 917.100 ;
        RECT 773.100 916.950 775.200 917.250 ;
        RECT 779.100 916.950 781.200 919.050 ;
        RECT 779.100 915.300 780.900 916.950 ;
        RECT 736.500 914.100 780.900 915.300 ;
        RECT 728.700 912.600 735.300 914.100 ;
        RECT 725.100 909.900 732.900 911.700 ;
        RECT 733.800 911.100 750.900 912.600 ;
        RECT 748.800 910.500 750.900 911.100 ;
        RECT 755.100 912.000 757.200 913.050 ;
        RECT 755.100 911.100 760.200 912.000 ;
        RECT 763.800 911.400 765.600 913.200 ;
        RECT 782.100 911.400 783.300 927.600 ;
        RECT 795.600 924.900 797.400 935.400 ;
        RECT 795.000 923.400 797.400 924.900 ;
        RECT 798.600 923.400 800.400 936.000 ;
        RECT 803.100 923.400 804.900 935.400 ;
        RECT 815.700 929.400 817.500 936.000 ;
        RECT 816.000 926.100 817.800 927.900 ;
        RECT 818.700 924.900 820.500 935.400 ;
        RECT 795.000 916.050 796.200 923.400 ;
        RECT 803.700 921.900 804.900 923.400 ;
        RECT 797.100 920.700 804.900 921.900 ;
        RECT 818.100 923.400 820.500 924.900 ;
        RECT 823.800 923.400 825.600 936.000 ;
        RECT 839.100 929.400 840.900 935.400 ;
        RECT 842.100 929.400 843.900 936.000 ;
        RECT 797.100 920.100 798.900 920.700 ;
        RECT 755.100 910.950 757.200 911.100 ;
        RECT 731.400 906.600 732.900 909.900 ;
        RECT 749.100 908.700 750.900 910.500 ;
        RECT 758.400 910.200 760.200 911.100 ;
        RECT 764.700 908.400 765.600 911.400 ;
        RECT 766.500 910.200 783.300 911.400 ;
        RECT 766.500 909.300 768.600 910.200 ;
        RECT 777.300 908.700 779.100 909.300 ;
        RECT 737.100 906.600 743.700 908.400 ;
        RECT 758.400 907.200 765.600 908.400 ;
        RECT 770.700 907.500 779.100 908.700 ;
        RECT 758.400 906.600 759.300 907.200 ;
        RECT 761.400 906.600 763.200 907.200 ;
        RECT 770.700 906.600 772.200 907.500 ;
        RECT 782.100 906.600 783.300 910.200 ;
        RECT 723.300 900.600 725.100 906.600 ;
        RECT 728.700 900.000 730.500 906.600 ;
        RECT 731.400 905.400 735.600 906.600 ;
        RECT 733.800 900.600 735.600 905.400 ;
        RECT 737.700 903.600 739.800 905.700 ;
        RECT 740.700 903.600 742.800 905.700 ;
        RECT 743.700 903.600 745.800 905.700 ;
        RECT 746.700 903.600 748.800 905.700 ;
        RECT 752.100 904.500 754.800 906.600 ;
        RECT 756.600 905.400 759.300 906.600 ;
        RECT 756.600 904.500 758.400 905.400 ;
        RECT 738.000 900.600 739.800 903.600 ;
        RECT 741.000 900.600 742.800 903.600 ;
        RECT 744.000 900.600 745.800 903.600 ;
        RECT 747.000 900.600 748.800 903.600 ;
        RECT 750.000 900.000 751.800 903.600 ;
        RECT 753.000 900.600 754.800 904.500 ;
        RECT 760.200 903.600 762.300 905.700 ;
        RECT 763.200 903.600 765.300 905.700 ;
        RECT 766.200 903.600 768.300 905.700 ;
        RECT 757.500 900.000 759.300 903.600 ;
        RECT 760.500 900.600 762.300 903.600 ;
        RECT 763.500 900.600 765.300 903.600 ;
        RECT 766.500 900.600 768.300 903.600 ;
        RECT 770.700 900.600 772.500 906.600 ;
        RECT 776.100 900.000 777.900 906.600 ;
        RECT 781.500 900.600 783.300 906.600 ;
        RECT 794.100 913.950 796.200 916.050 ;
        RECT 794.100 906.600 795.000 913.950 ;
        RECT 797.400 909.600 798.300 920.100 ;
        RECT 805.950 918.450 808.050 919.050 ;
        RECT 811.950 918.450 814.050 919.050 ;
        RECT 799.200 916.050 801.000 917.850 ;
        RECT 805.950 917.550 814.050 918.450 ;
        RECT 805.950 916.950 808.050 917.550 ;
        RECT 811.950 916.950 814.050 917.550 ;
        RECT 818.100 916.050 819.300 923.400 ;
        RECT 824.100 916.050 825.900 917.850 ;
        RECT 839.700 916.050 840.900 929.400 ;
        RECT 857.400 923.400 859.200 936.000 ;
        RECT 862.500 924.900 864.300 935.400 ;
        RECT 865.500 929.400 867.300 936.000 ;
        RECT 865.200 926.100 867.000 927.900 ;
        RECT 862.500 923.400 864.900 924.900 ;
        RECT 878.100 923.400 879.900 936.000 ;
        RECT 883.200 924.600 885.000 935.400 ;
        RECT 881.400 923.400 885.000 924.600 ;
        RECT 896.400 923.400 898.200 936.000 ;
        RECT 901.500 924.900 903.300 935.400 ;
        RECT 904.500 929.400 906.300 936.000 ;
        RECT 904.200 926.100 906.000 927.900 ;
        RECT 901.500 923.400 903.900 924.900 ;
        RECT 921.000 924.600 922.800 935.400 ;
        RECT 921.000 923.400 924.600 924.600 ;
        RECT 926.100 923.400 927.900 936.000 ;
        RECT 938.100 929.400 939.900 935.400 ;
        RECT 941.100 929.400 942.900 936.000 ;
        RECT 842.100 916.050 843.900 917.850 ;
        RECT 857.100 916.050 858.900 917.850 ;
        RECT 863.700 916.050 864.900 923.400 ;
        RECT 871.950 921.450 874.050 922.050 ;
        RECT 877.950 921.450 880.050 922.050 ;
        RECT 871.950 920.550 880.050 921.450 ;
        RECT 871.950 919.950 874.050 920.550 ;
        RECT 877.950 919.950 880.050 920.550 ;
        RECT 878.250 916.050 880.050 917.850 ;
        RECT 881.400 916.050 882.300 923.400 ;
        RECT 884.100 916.050 885.900 917.850 ;
        RECT 896.100 916.050 897.900 917.850 ;
        RECT 902.700 916.050 903.900 923.400 ;
        RECT 920.100 916.050 921.900 917.850 ;
        RECT 923.700 916.050 924.600 923.400 ;
        RECT 925.950 916.050 927.750 917.850 ;
        RECT 938.700 916.050 939.900 929.400 ;
        RECT 941.100 916.050 942.900 917.850 ;
        RECT 799.500 913.950 801.600 916.050 ;
        RECT 802.800 913.950 804.900 916.050 ;
        RECT 814.950 913.950 817.050 916.050 ;
        RECT 817.950 913.950 820.050 916.050 ;
        RECT 820.950 913.950 823.050 916.050 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 838.950 913.950 841.050 916.050 ;
        RECT 841.950 913.950 844.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 859.950 913.950 862.050 916.050 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 865.950 913.950 868.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 880.950 913.950 883.050 916.050 ;
        RECT 883.950 913.950 886.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 901.950 913.950 904.050 916.050 ;
        RECT 904.950 913.950 907.050 916.050 ;
        RECT 919.950 913.950 922.050 916.050 ;
        RECT 922.950 913.950 925.050 916.050 ;
        RECT 925.950 913.950 928.050 916.050 ;
        RECT 937.950 913.950 940.050 916.050 ;
        RECT 940.950 913.950 943.050 916.050 ;
        RECT 802.800 912.150 804.600 913.950 ;
        RECT 815.100 912.150 816.900 913.950 ;
        RECT 818.100 909.600 819.300 913.950 ;
        RECT 821.100 912.150 822.900 913.950 ;
        RECT 796.200 908.700 798.300 909.600 ;
        RECT 815.700 908.700 819.300 909.600 ;
        RECT 796.200 907.800 801.600 908.700 ;
        RECT 794.100 900.600 795.900 906.600 ;
        RECT 797.100 900.000 798.900 906.000 ;
        RECT 800.700 903.600 801.600 907.800 ;
        RECT 815.700 906.600 816.900 908.700 ;
        RECT 800.100 900.600 801.900 903.600 ;
        RECT 803.100 900.600 804.900 903.600 ;
        RECT 815.100 900.600 816.900 906.600 ;
        RECT 818.100 905.700 825.900 907.050 ;
        RECT 818.100 900.600 819.900 905.700 ;
        RECT 803.700 900.000 804.900 900.600 ;
        RECT 821.100 900.000 822.900 904.800 ;
        RECT 824.100 900.600 825.900 905.700 ;
        RECT 839.700 903.600 840.900 913.950 ;
        RECT 860.100 912.150 861.900 913.950 ;
        RECT 863.700 909.600 864.900 913.950 ;
        RECT 866.100 912.150 867.900 913.950 ;
        RECT 863.700 908.700 867.300 909.600 ;
        RECT 857.100 905.700 864.900 907.050 ;
        RECT 839.100 900.600 840.900 903.600 ;
        RECT 842.100 900.000 843.900 903.600 ;
        RECT 857.100 900.600 858.900 905.700 ;
        RECT 860.100 900.000 861.900 904.800 ;
        RECT 863.100 900.600 864.900 905.700 ;
        RECT 866.100 906.600 867.300 908.700 ;
        RECT 866.100 900.600 867.900 906.600 ;
        RECT 881.400 903.600 882.300 913.950 ;
        RECT 899.100 912.150 900.900 913.950 ;
        RECT 902.700 909.600 903.900 913.950 ;
        RECT 905.100 912.150 906.900 913.950 ;
        RECT 902.700 908.700 906.300 909.600 ;
        RECT 896.100 905.700 903.900 907.050 ;
        RECT 878.100 900.000 879.900 903.600 ;
        RECT 881.100 900.600 882.900 903.600 ;
        RECT 884.100 900.000 885.900 903.600 ;
        RECT 896.100 900.600 897.900 905.700 ;
        RECT 899.100 900.000 900.900 904.800 ;
        RECT 902.100 900.600 903.900 905.700 ;
        RECT 905.100 906.600 906.300 908.700 ;
        RECT 905.100 900.600 906.900 906.600 ;
        RECT 923.700 903.600 924.600 913.950 ;
        RECT 938.700 903.600 939.900 913.950 ;
        RECT 920.100 900.000 921.900 903.600 ;
        RECT 923.100 900.600 924.900 903.600 ;
        RECT 926.100 900.000 927.900 903.600 ;
        RECT 938.100 900.600 939.900 903.600 ;
        RECT 941.100 900.000 942.900 903.600 ;
        RECT 14.100 893.400 15.900 897.000 ;
        RECT 17.100 893.400 18.900 896.400 ;
        RECT 20.100 893.400 21.900 897.000 ;
        RECT 32.700 893.400 34.500 897.000 ;
        RECT 17.400 883.050 18.300 893.400 ;
        RECT 35.700 891.600 37.500 896.400 ;
        RECT 32.400 890.400 37.500 891.600 ;
        RECT 40.200 890.400 42.000 897.000 ;
        RECT 56.100 893.400 57.900 897.000 ;
        RECT 59.100 893.400 60.900 896.400 ;
        RECT 32.400 883.050 33.300 890.400 ;
        RECT 34.950 883.050 36.750 884.850 ;
        RECT 41.100 883.050 42.900 884.850 ;
        RECT 59.100 883.050 60.300 893.400 ;
        RECT 74.700 889.200 76.500 896.400 ;
        RECT 79.800 890.400 81.600 897.000 ;
        RECT 92.100 890.400 93.900 896.400 ;
        RECT 74.700 888.300 78.900 889.200 ;
        RECT 74.100 883.050 75.900 884.850 ;
        RECT 77.700 883.050 78.900 888.300 ;
        RECT 92.700 888.300 93.900 890.400 ;
        RECT 95.100 891.300 96.900 896.400 ;
        RECT 98.100 892.200 99.900 897.000 ;
        RECT 101.100 891.300 102.900 896.400 ;
        RECT 95.100 889.950 102.900 891.300 ;
        RECT 113.700 889.200 115.500 896.400 ;
        RECT 118.800 890.400 120.600 897.000 ;
        RECT 113.700 888.300 117.900 889.200 ;
        RECT 92.700 887.400 96.300 888.300 ;
        RECT 79.950 883.050 81.750 884.850 ;
        RECT 92.100 883.050 93.900 884.850 ;
        RECT 95.100 883.050 96.300 887.400 ;
        RECT 98.100 883.050 99.900 884.850 ;
        RECT 113.100 883.050 114.900 884.850 ;
        RECT 116.700 883.050 117.900 888.300 ;
        RECT 131.100 887.400 132.900 897.000 ;
        RECT 137.700 888.000 139.500 896.400 ;
        RECT 155.400 890.400 157.200 897.000 ;
        RECT 160.500 889.200 162.300 896.400 ;
        RECT 158.100 888.300 162.300 889.200 ;
        RECT 173.700 889.200 175.500 896.400 ;
        RECT 178.800 890.400 180.600 897.000 ;
        RECT 194.700 889.200 196.500 896.400 ;
        RECT 199.800 890.400 201.600 897.000 ;
        RECT 173.700 888.300 177.900 889.200 ;
        RECT 194.700 888.300 198.900 889.200 ;
        RECT 137.700 886.800 141.000 888.000 ;
        RECT 126.000 885.450 130.050 886.050 ;
        RECT 118.950 883.050 120.750 884.850 ;
        RECT 125.550 883.950 130.050 885.450 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 19.950 880.950 22.050 883.050 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 73.950 880.950 76.050 883.050 ;
        RECT 76.950 880.950 79.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 91.950 880.950 94.050 883.050 ;
        RECT 94.950 880.950 97.050 883.050 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 100.950 880.950 103.050 883.050 ;
        RECT 112.950 880.950 115.050 883.050 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 118.950 880.950 121.050 883.050 ;
        RECT 14.250 879.150 16.050 880.950 ;
        RECT 17.400 873.600 18.300 880.950 ;
        RECT 20.100 879.150 21.900 880.950 ;
        RECT 19.950 876.450 22.050 877.050 ;
        RECT 25.950 876.450 28.050 877.050 ;
        RECT 19.950 875.550 28.050 876.450 ;
        RECT 19.950 874.950 22.050 875.550 ;
        RECT 25.950 874.950 28.050 875.550 ;
        RECT 32.400 873.600 33.300 880.950 ;
        RECT 37.950 879.150 39.750 880.950 ;
        RECT 56.100 879.150 57.900 880.950 ;
        RECT 14.100 861.000 15.900 873.600 ;
        RECT 17.400 872.400 21.000 873.600 ;
        RECT 19.200 861.600 21.000 872.400 ;
        RECT 32.100 861.600 33.900 873.600 ;
        RECT 35.100 872.700 42.900 873.600 ;
        RECT 35.100 861.600 36.900 872.700 ;
        RECT 38.100 861.000 39.900 871.800 ;
        RECT 41.100 861.600 42.900 872.700 ;
        RECT 59.100 867.600 60.300 880.950 ;
        RECT 77.700 867.600 78.900 880.950 ;
        RECT 95.100 873.600 96.300 880.950 ;
        RECT 101.100 879.150 102.900 880.950 ;
        RECT 95.100 872.100 97.500 873.600 ;
        RECT 93.000 869.100 94.800 870.900 ;
        RECT 56.100 861.000 57.900 867.600 ;
        RECT 59.100 861.600 60.900 867.600 ;
        RECT 74.100 861.000 75.900 867.600 ;
        RECT 77.100 861.600 78.900 867.600 ;
        RECT 80.100 861.000 81.900 867.600 ;
        RECT 92.700 861.000 94.500 867.600 ;
        RECT 95.700 861.600 97.500 872.100 ;
        RECT 100.800 861.000 102.600 873.600 ;
        RECT 116.700 867.600 117.900 880.950 ;
        RECT 125.550 880.050 126.450 883.950 ;
        RECT 131.100 883.050 132.900 884.850 ;
        RECT 137.100 883.050 138.900 884.850 ;
        RECT 140.100 883.050 141.000 886.800 ;
        RECT 155.250 883.050 157.050 884.850 ;
        RECT 158.100 883.050 159.300 888.300 ;
        RECT 161.100 883.050 162.900 884.850 ;
        RECT 173.100 883.050 174.900 884.850 ;
        RECT 176.700 883.050 177.900 888.300 ;
        RECT 178.950 883.050 180.750 884.850 ;
        RECT 194.100 883.050 195.900 884.850 ;
        RECT 197.700 883.050 198.900 888.300 ;
        RECT 212.100 887.400 213.900 897.000 ;
        RECT 218.700 888.000 220.500 896.400 ;
        RECT 236.700 889.200 238.500 896.400 ;
        RECT 241.800 890.400 243.600 897.000 ;
        RECT 236.700 888.300 240.900 889.200 ;
        RECT 218.700 886.800 222.000 888.000 ;
        RECT 199.950 883.050 201.750 884.850 ;
        RECT 212.100 883.050 213.900 884.850 ;
        RECT 218.100 883.050 219.900 884.850 ;
        RECT 221.100 883.050 222.000 886.800 ;
        RECT 236.100 883.050 237.900 884.850 ;
        RECT 239.700 883.050 240.900 888.300 ;
        RECT 256.500 888.000 258.300 896.400 ;
        RECT 255.000 886.800 258.300 888.000 ;
        RECT 263.100 887.400 264.900 897.000 ;
        RECT 278.100 893.400 279.900 897.000 ;
        RECT 281.100 893.400 282.900 896.400 ;
        RECT 284.100 893.400 285.900 897.000 ;
        RECT 296.100 893.400 297.900 897.000 ;
        RECT 299.100 893.400 300.900 896.400 ;
        RECT 302.100 893.400 303.900 897.000 ;
        RECT 317.100 893.400 318.900 897.000 ;
        RECT 320.100 893.400 321.900 896.400 ;
        RECT 323.100 893.400 324.900 897.000 ;
        RECT 241.950 883.050 243.750 884.850 ;
        RECT 255.000 883.050 255.900 886.800 ;
        RECT 257.100 883.050 258.900 884.850 ;
        RECT 263.100 883.050 264.900 884.850 ;
        RECT 281.400 883.050 282.300 893.400 ;
        RECT 283.950 888.450 286.050 889.050 ;
        RECT 289.950 888.450 292.050 889.050 ;
        RECT 283.950 887.550 292.050 888.450 ;
        RECT 283.950 886.950 286.050 887.550 ;
        RECT 289.950 886.950 292.050 887.550 ;
        RECT 299.700 883.050 300.600 893.400 ;
        RECT 320.400 883.050 321.300 893.400 ;
        RECT 335.100 887.400 336.900 897.000 ;
        RECT 341.700 888.000 343.500 896.400 ;
        RECT 361.500 890.400 363.300 897.000 ;
        RECT 366.000 890.400 367.800 896.400 ;
        RECT 370.500 890.400 372.300 897.000 ;
        RECT 386.100 893.400 387.900 896.400 ;
        RECT 389.100 893.400 390.900 897.000 ;
        RECT 341.700 886.800 345.000 888.000 ;
        RECT 335.100 883.050 336.900 884.850 ;
        RECT 341.100 883.050 342.900 884.850 ;
        RECT 344.100 883.050 345.000 886.800 ;
        RECT 359.100 883.050 360.900 884.850 ;
        RECT 365.700 883.050 366.900 890.400 ;
        RECT 370.950 883.050 372.750 884.850 ;
        RECT 386.700 883.050 387.900 893.400 ;
        RECT 404.700 890.400 406.500 897.000 ;
        RECT 409.200 890.400 411.000 896.400 ;
        RECT 413.700 890.400 415.500 897.000 ;
        RECT 431.100 890.400 432.900 897.000 ;
        RECT 434.100 890.400 435.900 896.400 ;
        RECT 437.100 890.400 438.900 897.000 ;
        RECT 440.100 890.400 441.900 896.400 ;
        RECT 443.100 890.400 444.900 897.000 ;
        RECT 458.100 890.400 459.900 896.400 ;
        RECT 461.100 890.400 462.900 897.000 ;
        RECT 464.100 893.400 465.900 896.400 ;
        RECT 404.250 883.050 406.050 884.850 ;
        RECT 410.100 883.050 411.300 890.400 ;
        RECT 434.700 889.500 435.900 890.400 ;
        RECT 440.700 889.500 441.900 890.400 ;
        RECT 434.700 888.300 441.900 889.500 ;
        RECT 416.100 883.050 417.900 884.850 ;
        RECT 434.700 883.050 435.900 888.300 ;
        RECT 458.100 883.050 459.300 890.400 ;
        RECT 464.700 889.500 465.900 893.400 ;
        RECT 476.100 891.300 477.900 896.400 ;
        RECT 479.100 892.200 480.900 897.000 ;
        RECT 482.100 891.300 483.900 896.400 ;
        RECT 476.100 889.950 483.900 891.300 ;
        RECT 485.100 890.400 486.900 896.400 ;
        RECT 497.100 893.400 498.900 896.400 ;
        RECT 460.200 888.600 465.900 889.500 ;
        RECT 460.200 887.700 462.000 888.600 ;
        RECT 485.100 888.300 486.300 890.400 ;
        RECT 497.100 889.500 498.300 893.400 ;
        RECT 500.100 890.400 501.900 897.000 ;
        RECT 503.100 890.400 504.900 896.400 ;
        RECT 515.100 890.400 516.900 896.400 ;
        RECT 497.100 888.600 502.800 889.500 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 154.950 880.950 157.050 883.050 ;
        RECT 157.950 880.950 160.050 883.050 ;
        RECT 160.950 880.950 163.050 883.050 ;
        RECT 172.950 880.950 175.050 883.050 ;
        RECT 175.950 880.950 178.050 883.050 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 211.950 880.950 214.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 217.950 880.950 220.050 883.050 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 277.950 880.950 280.050 883.050 ;
        RECT 280.950 880.950 283.050 883.050 ;
        RECT 283.950 880.950 286.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 301.950 880.950 304.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 361.950 880.950 364.050 883.050 ;
        RECT 364.950 880.950 367.050 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 403.950 880.950 406.050 883.050 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 433.800 880.950 435.900 883.050 ;
        RECT 439.800 880.950 441.900 883.050 ;
        RECT 121.950 878.550 126.450 880.050 ;
        RECT 134.100 879.150 135.900 880.950 ;
        RECT 121.950 877.950 126.000 878.550 ;
        RECT 140.100 868.800 141.000 880.950 ;
        RECT 134.400 867.900 141.000 868.800 ;
        RECT 134.400 867.600 135.900 867.900 ;
        RECT 113.100 861.000 114.900 867.600 ;
        RECT 116.100 861.600 117.900 867.600 ;
        RECT 119.100 861.000 120.900 867.600 ;
        RECT 131.100 861.000 132.900 867.600 ;
        RECT 134.100 861.600 135.900 867.600 ;
        RECT 140.100 867.600 141.000 867.900 ;
        RECT 158.100 867.600 159.300 880.950 ;
        RECT 176.700 867.600 177.900 880.950 ;
        RECT 197.700 867.600 198.900 880.950 ;
        RECT 215.100 879.150 216.900 880.950 ;
        RECT 199.950 873.450 202.050 874.050 ;
        RECT 211.950 873.450 214.050 874.050 ;
        RECT 199.950 872.550 214.050 873.450 ;
        RECT 199.950 871.950 202.050 872.550 ;
        RECT 211.950 871.950 214.050 872.550 ;
        RECT 221.100 868.800 222.000 880.950 ;
        RECT 215.400 867.900 222.000 868.800 ;
        RECT 215.400 867.600 216.900 867.900 ;
        RECT 137.100 861.000 138.900 867.000 ;
        RECT 140.100 861.600 141.900 867.600 ;
        RECT 155.100 861.000 156.900 867.600 ;
        RECT 158.100 861.600 159.900 867.600 ;
        RECT 161.100 861.000 162.900 867.600 ;
        RECT 173.100 861.000 174.900 867.600 ;
        RECT 176.100 861.600 177.900 867.600 ;
        RECT 179.100 861.000 180.900 867.600 ;
        RECT 194.100 861.000 195.900 867.600 ;
        RECT 197.100 861.600 198.900 867.600 ;
        RECT 200.100 861.000 201.900 867.600 ;
        RECT 212.100 861.000 213.900 867.600 ;
        RECT 215.100 861.600 216.900 867.600 ;
        RECT 221.100 867.600 222.000 867.900 ;
        RECT 239.700 867.600 240.900 880.950 ;
        RECT 255.000 868.800 255.900 880.950 ;
        RECT 260.100 879.150 261.900 880.950 ;
        RECT 278.250 879.150 280.050 880.950 ;
        RECT 281.400 873.600 282.300 880.950 ;
        RECT 284.100 879.150 285.900 880.950 ;
        RECT 296.100 879.150 297.900 880.950 ;
        RECT 299.700 873.600 300.600 880.950 ;
        RECT 301.950 879.150 303.750 880.950 ;
        RECT 317.250 879.150 319.050 880.950 ;
        RECT 320.400 873.600 321.300 880.950 ;
        RECT 323.100 879.150 324.900 880.950 ;
        RECT 338.100 879.150 339.900 880.950 ;
        RECT 255.000 867.900 261.600 868.800 ;
        RECT 255.000 867.600 255.900 867.900 ;
        RECT 218.100 861.000 219.900 867.000 ;
        RECT 221.100 861.600 222.900 867.600 ;
        RECT 236.100 861.000 237.900 867.600 ;
        RECT 239.100 861.600 240.900 867.600 ;
        RECT 242.100 861.000 243.900 867.600 ;
        RECT 254.100 861.600 255.900 867.600 ;
        RECT 260.100 867.600 261.600 867.900 ;
        RECT 257.100 861.000 258.900 867.000 ;
        RECT 260.100 861.600 261.900 867.600 ;
        RECT 263.100 861.000 264.900 867.600 ;
        RECT 278.100 861.000 279.900 873.600 ;
        RECT 281.400 872.400 285.000 873.600 ;
        RECT 283.200 861.600 285.000 872.400 ;
        RECT 297.000 872.400 300.600 873.600 ;
        RECT 297.000 861.600 298.800 872.400 ;
        RECT 302.100 861.000 303.900 873.600 ;
        RECT 317.100 861.000 318.900 873.600 ;
        RECT 320.400 872.400 324.000 873.600 ;
        RECT 322.200 861.600 324.000 872.400 ;
        RECT 344.100 868.800 345.000 880.950 ;
        RECT 362.100 879.150 363.900 880.950 ;
        RECT 366.000 875.400 366.900 880.950 ;
        RECT 367.950 879.150 369.750 880.950 ;
        RECT 362.100 874.500 366.900 875.400 ;
        RECT 338.400 867.900 345.000 868.800 ;
        RECT 338.400 867.600 339.900 867.900 ;
        RECT 335.100 861.000 336.900 867.600 ;
        RECT 338.100 861.600 339.900 867.600 ;
        RECT 344.100 867.600 345.000 867.900 ;
        RECT 341.100 861.000 342.900 867.000 ;
        RECT 344.100 861.600 345.900 867.600 ;
        RECT 359.100 862.500 360.900 873.600 ;
        RECT 362.100 863.400 363.900 874.500 ;
        RECT 365.100 872.400 372.900 873.300 ;
        RECT 365.100 862.500 366.900 872.400 ;
        RECT 359.100 861.600 366.900 862.500 ;
        RECT 368.100 861.000 369.900 871.500 ;
        RECT 371.100 861.600 372.900 872.400 ;
        RECT 386.700 867.600 387.900 880.950 ;
        RECT 389.100 879.150 390.900 880.950 ;
        RECT 407.250 879.150 409.050 880.950 ;
        RECT 410.100 875.400 411.000 880.950 ;
        RECT 413.100 879.150 414.900 880.950 ;
        RECT 434.700 875.400 435.900 880.950 ;
        RECT 440.100 879.150 441.900 880.950 ;
        RECT 458.100 880.950 460.200 883.050 ;
        RECT 410.100 874.500 414.900 875.400 ;
        RECT 404.100 872.400 411.900 873.300 ;
        RECT 386.100 861.600 387.900 867.600 ;
        RECT 389.100 861.000 390.900 867.600 ;
        RECT 404.100 861.600 405.900 872.400 ;
        RECT 407.100 861.000 408.900 871.500 ;
        RECT 410.100 862.500 411.900 872.400 ;
        RECT 413.100 863.400 414.900 874.500 ;
        RECT 434.700 874.500 441.900 875.400 ;
        RECT 434.700 873.600 435.900 874.500 ;
        RECT 416.100 862.500 417.900 873.600 ;
        RECT 410.100 861.600 417.900 862.500 ;
        RECT 431.100 861.000 432.900 873.600 ;
        RECT 434.100 861.600 435.900 873.600 ;
        RECT 437.100 861.000 438.900 873.600 ;
        RECT 440.100 861.600 441.900 874.500 ;
        RECT 458.100 873.600 459.300 880.950 ;
        RECT 461.100 876.300 462.000 887.700 ;
        RECT 482.700 887.400 486.300 888.300 ;
        RECT 501.000 887.700 502.800 888.600 ;
        RECT 479.100 883.050 480.900 884.850 ;
        RECT 482.700 883.050 483.900 887.400 ;
        RECT 485.100 883.050 486.900 884.850 ;
        RECT 463.500 880.950 465.600 883.050 ;
        RECT 475.950 880.950 478.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 481.950 880.950 484.050 883.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 497.400 880.950 499.500 883.050 ;
        RECT 463.800 879.150 465.600 880.950 ;
        RECT 476.100 879.150 477.900 880.950 ;
        RECT 460.200 875.400 462.000 876.300 ;
        RECT 460.200 874.500 465.900 875.400 ;
        RECT 443.100 861.000 444.900 873.600 ;
        RECT 458.100 861.600 459.900 873.600 ;
        RECT 461.100 861.000 462.900 871.800 ;
        RECT 464.700 867.600 465.900 874.500 ;
        RECT 482.700 873.600 483.900 880.950 ;
        RECT 497.400 879.150 499.200 880.950 ;
        RECT 501.000 876.300 501.900 887.700 ;
        RECT 503.700 883.050 504.900 890.400 ;
        RECT 515.700 888.300 516.900 890.400 ;
        RECT 518.100 891.300 519.900 896.400 ;
        RECT 521.100 892.200 522.900 897.000 ;
        RECT 524.100 891.300 525.900 896.400 ;
        RECT 536.100 893.400 537.900 897.000 ;
        RECT 539.100 893.400 540.900 896.400 ;
        RECT 542.100 893.400 543.900 897.000 ;
        RECT 554.100 893.400 555.900 896.400 ;
        RECT 557.100 893.400 558.900 897.000 ;
        RECT 518.100 889.950 525.900 891.300 ;
        RECT 515.700 887.400 519.300 888.300 ;
        RECT 515.100 883.050 516.900 884.850 ;
        RECT 518.100 883.050 519.300 887.400 ;
        RECT 521.100 883.050 522.900 884.850 ;
        RECT 539.400 883.050 540.300 893.400 ;
        RECT 554.700 883.050 555.900 893.400 ;
        RECT 572.100 890.400 573.900 896.400 ;
        RECT 572.700 888.300 573.900 890.400 ;
        RECT 575.100 891.300 576.900 896.400 ;
        RECT 578.100 892.200 579.900 897.000 ;
        RECT 581.100 891.300 582.900 896.400 ;
        RECT 596.100 893.400 597.900 896.400 ;
        RECT 599.100 893.400 600.900 897.000 ;
        RECT 575.100 889.950 582.900 891.300 ;
        RECT 572.700 887.400 576.300 888.300 ;
        RECT 572.100 883.050 573.900 884.850 ;
        RECT 575.100 883.050 576.300 887.400 ;
        RECT 578.100 883.050 579.900 884.850 ;
        RECT 596.700 883.050 597.900 893.400 ;
        RECT 614.100 890.400 615.900 896.400 ;
        RECT 614.700 888.300 615.900 890.400 ;
        RECT 617.100 891.300 618.900 896.400 ;
        RECT 620.100 892.200 621.900 897.000 ;
        RECT 623.100 891.300 624.900 896.400 ;
        RECT 626.700 893.400 628.500 897.000 ;
        RECT 629.700 893.400 631.500 896.400 ;
        RECT 617.100 889.950 624.900 891.300 ;
        RECT 614.700 887.400 618.300 888.300 ;
        RECT 614.100 883.050 615.900 884.850 ;
        RECT 617.100 883.050 618.300 887.400 ;
        RECT 620.100 883.050 621.900 884.850 ;
        RECT 502.800 880.950 504.900 883.050 ;
        RECT 514.950 880.950 517.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 571.950 880.950 574.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 501.000 875.400 502.800 876.300 ;
        RECT 464.100 861.600 465.900 867.600 ;
        RECT 476.400 861.000 478.200 873.600 ;
        RECT 481.500 872.100 483.900 873.600 ;
        RECT 497.100 874.500 502.800 875.400 ;
        RECT 481.500 861.600 483.300 872.100 ;
        RECT 484.200 869.100 486.000 870.900 ;
        RECT 497.100 867.600 498.300 874.500 ;
        RECT 503.700 873.600 504.900 880.950 ;
        RECT 484.500 861.000 486.300 867.600 ;
        RECT 497.100 861.600 498.900 867.600 ;
        RECT 500.100 861.000 501.900 871.800 ;
        RECT 503.100 861.600 504.900 873.600 ;
        RECT 518.100 873.600 519.300 880.950 ;
        RECT 524.100 879.150 525.900 880.950 ;
        RECT 536.250 879.150 538.050 880.950 ;
        RECT 539.400 873.600 540.300 880.950 ;
        RECT 542.100 879.150 543.900 880.950 ;
        RECT 518.100 872.100 520.500 873.600 ;
        RECT 516.000 869.100 517.800 870.900 ;
        RECT 515.700 861.000 517.500 867.600 ;
        RECT 518.700 861.600 520.500 872.100 ;
        RECT 523.800 861.000 525.600 873.600 ;
        RECT 536.100 861.000 537.900 873.600 ;
        RECT 539.400 872.400 543.000 873.600 ;
        RECT 541.200 861.600 543.000 872.400 ;
        RECT 554.700 867.600 555.900 880.950 ;
        RECT 557.100 879.150 558.900 880.950 ;
        RECT 575.100 873.600 576.300 880.950 ;
        RECT 581.100 879.150 582.900 880.950 ;
        RECT 575.100 872.100 577.500 873.600 ;
        RECT 573.000 869.100 574.800 870.900 ;
        RECT 554.100 861.600 555.900 867.600 ;
        RECT 557.100 861.000 558.900 867.600 ;
        RECT 572.700 861.000 574.500 867.600 ;
        RECT 575.700 861.600 577.500 872.100 ;
        RECT 580.800 861.000 582.600 873.600 ;
        RECT 596.700 867.600 597.900 880.950 ;
        RECT 599.100 879.150 600.900 880.950 ;
        RECT 617.100 873.600 618.300 880.950 ;
        RECT 623.100 879.150 624.900 880.950 ;
        RECT 630.000 880.050 631.500 893.400 ;
        RECT 629.100 877.950 631.500 880.050 ;
        RECT 617.100 872.100 619.500 873.600 ;
        RECT 615.000 869.100 616.800 870.900 ;
        RECT 596.100 861.600 597.900 867.600 ;
        RECT 599.100 861.000 600.900 867.600 ;
        RECT 614.700 861.000 616.500 867.600 ;
        RECT 617.700 861.600 619.500 872.100 ;
        RECT 622.800 861.000 624.600 873.600 ;
        RECT 630.000 867.600 631.500 877.950 ;
        RECT 633.300 890.400 635.100 896.400 ;
        RECT 638.700 890.400 640.500 897.000 ;
        RECT 643.800 891.600 645.600 896.400 ;
        RECT 648.000 893.400 649.800 896.400 ;
        RECT 651.000 893.400 652.800 896.400 ;
        RECT 654.000 893.400 655.800 896.400 ;
        RECT 657.000 893.400 658.800 896.400 ;
        RECT 660.000 893.400 661.800 897.000 ;
        RECT 641.400 890.400 645.600 891.600 ;
        RECT 647.700 891.300 649.800 893.400 ;
        RECT 650.700 891.300 652.800 893.400 ;
        RECT 653.700 891.300 655.800 893.400 ;
        RECT 656.700 891.300 658.800 893.400 ;
        RECT 663.000 892.500 664.800 896.400 ;
        RECT 667.500 893.400 669.300 897.000 ;
        RECT 670.500 893.400 672.300 896.400 ;
        RECT 673.500 893.400 675.300 896.400 ;
        RECT 676.500 893.400 678.300 896.400 ;
        RECT 662.100 890.400 664.800 892.500 ;
        RECT 666.600 891.600 668.400 892.500 ;
        RECT 666.600 890.400 669.300 891.600 ;
        RECT 670.200 891.300 672.300 893.400 ;
        RECT 673.200 891.300 675.300 893.400 ;
        RECT 676.200 891.300 678.300 893.400 ;
        RECT 680.700 890.400 682.500 896.400 ;
        RECT 686.100 890.400 687.900 897.000 ;
        RECT 691.500 890.400 693.300 896.400 ;
        RECT 707.400 890.400 709.200 897.000 ;
        RECT 633.300 873.600 634.200 890.400 ;
        RECT 641.400 887.100 642.900 890.400 ;
        RECT 647.100 888.600 653.700 890.400 ;
        RECT 668.400 889.800 669.300 890.400 ;
        RECT 671.400 889.800 673.200 890.400 ;
        RECT 668.400 888.600 675.600 889.800 ;
        RECT 635.100 885.300 642.900 887.100 ;
        RECT 659.100 886.500 660.900 888.300 ;
        RECT 658.800 885.900 660.900 886.500 ;
        RECT 643.800 884.400 660.900 885.900 ;
        RECT 665.100 885.900 667.200 886.050 ;
        RECT 668.400 885.900 670.200 886.800 ;
        RECT 665.100 885.000 670.200 885.900 ;
        RECT 674.700 885.600 675.600 888.600 ;
        RECT 680.700 889.500 682.200 890.400 ;
        RECT 680.700 888.300 689.100 889.500 ;
        RECT 687.300 887.700 689.100 888.300 ;
        RECT 676.500 886.800 678.600 887.700 ;
        RECT 692.100 886.800 693.300 890.400 ;
        RECT 712.500 889.200 714.300 896.400 ;
        RECT 725.700 890.400 727.500 897.000 ;
        RECT 730.200 890.400 732.000 896.400 ;
        RECT 734.700 890.400 736.500 897.000 ;
        RECT 752.100 890.400 753.900 896.400 ;
        RECT 676.500 885.600 693.300 886.800 ;
        RECT 638.700 882.900 645.300 884.400 ;
        RECT 665.100 883.950 667.200 885.000 ;
        RECT 673.800 883.800 675.600 885.600 ;
        RECT 638.700 880.050 640.200 882.900 ;
        RECT 646.500 881.700 690.900 882.900 ;
        RECT 646.500 880.200 647.400 881.700 ;
        RECT 638.100 877.950 640.200 880.050 ;
        RECT 642.300 878.400 647.400 880.200 ;
        RECT 650.100 879.900 663.600 880.800 ;
        RECT 670.800 879.900 672.600 880.500 ;
        RECT 689.100 880.050 690.900 881.700 ;
        RECT 650.100 878.700 651.000 879.900 ;
        RECT 650.100 876.900 651.900 878.700 ;
        RECT 656.100 877.200 660.000 879.000 ;
        RECT 661.500 878.700 672.600 879.900 ;
        RECT 683.100 879.750 685.200 880.050 ;
        RECT 661.500 877.800 663.600 878.700 ;
        RECT 681.300 877.950 685.200 879.750 ;
        RECT 689.100 877.950 691.200 880.050 ;
        RECT 681.300 877.200 683.100 877.950 ;
        RECT 656.100 876.900 658.200 877.200 ;
        RECT 669.600 876.300 683.100 877.200 ;
        RECT 635.100 875.700 636.900 876.300 ;
        RECT 669.600 875.700 670.800 876.300 ;
        RECT 635.100 874.500 670.800 875.700 ;
        RECT 673.500 874.500 675.600 874.800 ;
        RECT 633.300 872.700 649.800 873.600 ;
        RECT 633.300 869.400 634.200 872.700 ;
        RECT 638.100 870.600 643.800 871.800 ;
        RECT 647.700 871.500 649.800 872.700 ;
        RECT 653.100 872.400 670.800 873.600 ;
        RECT 673.500 873.300 685.500 874.500 ;
        RECT 673.500 872.700 675.600 873.300 ;
        RECT 683.700 872.700 685.500 873.300 ;
        RECT 653.100 871.500 655.200 872.400 ;
        RECT 669.600 871.800 670.800 872.400 ;
        RECT 687.000 871.800 688.800 872.100 ;
        RECT 638.100 870.000 639.900 870.600 ;
        RECT 633.300 868.500 637.200 869.400 ;
        RECT 636.000 867.600 637.200 868.500 ;
        RECT 642.600 867.600 643.800 870.600 ;
        RECT 644.700 869.700 646.500 870.300 ;
        RECT 644.700 868.500 652.800 869.700 ;
        RECT 650.700 867.600 652.800 868.500 ;
        RECT 656.100 867.600 658.800 871.500 ;
        RECT 661.500 869.100 664.800 871.200 ;
        RECT 669.600 870.600 688.800 871.800 ;
        RECT 626.700 861.000 628.500 867.600 ;
        RECT 629.700 861.600 631.500 867.600 ;
        RECT 633.000 861.000 634.800 867.600 ;
        RECT 636.000 861.600 637.800 867.600 ;
        RECT 639.000 861.000 640.800 867.600 ;
        RECT 642.000 861.600 643.800 867.600 ;
        RECT 645.000 861.000 646.800 867.600 ;
        RECT 647.700 864.600 649.800 866.700 ;
        RECT 650.700 864.600 652.800 866.700 ;
        RECT 653.700 864.600 655.800 866.700 ;
        RECT 648.000 861.600 649.800 864.600 ;
        RECT 651.000 861.600 652.800 864.600 ;
        RECT 654.000 861.600 655.800 864.600 ;
        RECT 657.000 861.600 658.800 867.600 ;
        RECT 660.000 861.000 661.800 867.600 ;
        RECT 663.000 861.600 664.800 869.100 ;
        RECT 670.200 867.600 672.300 869.700 ;
        RECT 666.900 861.000 668.700 867.600 ;
        RECT 669.900 861.600 671.700 867.600 ;
        RECT 672.600 864.600 674.700 866.700 ;
        RECT 675.600 864.600 677.700 866.700 ;
        RECT 672.900 861.600 674.700 864.600 ;
        RECT 675.900 861.600 677.700 864.600 ;
        RECT 679.500 861.000 681.300 867.600 ;
        RECT 682.500 861.600 684.300 870.600 ;
        RECT 687.000 870.300 688.800 870.600 ;
        RECT 692.100 869.400 693.300 885.600 ;
        RECT 710.100 888.300 714.300 889.200 ;
        RECT 707.250 883.050 709.050 884.850 ;
        RECT 710.100 883.050 711.300 888.300 ;
        RECT 713.100 883.050 714.900 884.850 ;
        RECT 725.250 883.050 727.050 884.850 ;
        RECT 731.100 883.050 732.300 890.400 ;
        RECT 752.700 888.300 753.900 890.400 ;
        RECT 755.100 891.300 756.900 896.400 ;
        RECT 758.100 892.200 759.900 897.000 ;
        RECT 761.100 891.300 762.900 896.400 ;
        RECT 755.100 889.950 762.900 891.300 ;
        RECT 752.700 887.400 756.300 888.300 ;
        RECT 773.100 887.400 774.900 897.000 ;
        RECT 779.700 888.000 781.500 896.400 ;
        RECT 797.100 893.400 798.900 896.400 ;
        RECT 800.100 893.400 801.900 897.000 ;
        RECT 815.100 895.500 822.900 896.400 ;
        RECT 737.100 883.050 738.900 884.850 ;
        RECT 752.100 883.050 753.900 884.850 ;
        RECT 755.100 883.050 756.300 887.400 ;
        RECT 779.700 886.800 783.000 888.000 ;
        RECT 758.100 883.050 759.900 884.850 ;
        RECT 773.100 883.050 774.900 884.850 ;
        RECT 779.100 883.050 780.900 884.850 ;
        RECT 782.100 883.050 783.000 886.800 ;
        RECT 784.950 885.450 789.000 886.050 ;
        RECT 784.950 883.950 789.450 885.450 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 736.950 880.950 739.050 883.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 689.700 868.500 693.300 869.400 ;
        RECT 689.700 867.600 690.600 868.500 ;
        RECT 710.100 867.600 711.300 880.950 ;
        RECT 728.250 879.150 730.050 880.950 ;
        RECT 731.100 875.400 732.000 880.950 ;
        RECT 734.100 879.150 735.900 880.950 ;
        RECT 731.100 874.500 735.900 875.400 ;
        RECT 725.100 872.400 732.900 873.300 ;
        RECT 685.500 861.000 687.300 867.600 ;
        RECT 688.500 866.700 690.600 867.600 ;
        RECT 688.500 861.600 690.300 866.700 ;
        RECT 691.500 861.000 693.300 867.600 ;
        RECT 707.100 861.000 708.900 867.600 ;
        RECT 710.100 861.600 711.900 867.600 ;
        RECT 713.100 861.000 714.900 867.600 ;
        RECT 725.100 861.600 726.900 872.400 ;
        RECT 728.100 861.000 729.900 871.500 ;
        RECT 731.100 862.500 732.900 872.400 ;
        RECT 734.100 863.400 735.900 874.500 ;
        RECT 755.100 873.600 756.300 880.950 ;
        RECT 761.100 879.150 762.900 880.950 ;
        RECT 776.100 879.150 777.900 880.950 ;
        RECT 737.100 862.500 738.900 873.600 ;
        RECT 755.100 872.100 757.500 873.600 ;
        RECT 753.000 869.100 754.800 870.900 ;
        RECT 731.100 861.600 738.900 862.500 ;
        RECT 752.700 861.000 754.500 867.600 ;
        RECT 755.700 861.600 757.500 872.100 ;
        RECT 760.800 861.000 762.600 873.600 ;
        RECT 782.100 868.800 783.000 880.950 ;
        RECT 788.550 880.050 789.450 883.950 ;
        RECT 797.700 883.050 798.900 893.400 ;
        RECT 815.100 890.400 816.900 895.500 ;
        RECT 818.100 890.400 819.900 894.600 ;
        RECT 821.100 891.000 822.900 895.500 ;
        RECT 824.100 891.900 825.900 897.000 ;
        RECT 827.100 891.000 828.900 896.400 ;
        RECT 842.100 893.400 843.900 897.000 ;
        RECT 845.100 893.400 846.900 896.400 ;
        RECT 818.700 888.900 819.600 890.400 ;
        RECT 821.100 890.100 828.900 891.000 ;
        RECT 818.700 887.700 823.050 888.900 ;
        RECT 818.250 883.050 820.050 884.850 ;
        RECT 822.000 883.050 823.050 887.700 ;
        RECT 829.950 888.450 832.050 889.050 ;
        RECT 841.950 888.450 844.050 889.200 ;
        RECT 829.950 887.550 844.050 888.450 ;
        RECT 829.950 886.950 832.050 887.550 ;
        RECT 841.950 887.100 844.050 887.550 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 799.950 880.950 802.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 817.950 880.950 820.050 883.050 ;
        RECT 820.950 880.950 823.050 883.050 ;
        RECT 823.950 883.050 825.750 884.850 ;
        RECT 845.100 883.050 846.300 893.400 ;
        RECT 861.600 892.200 863.400 896.400 ;
        RECT 860.700 890.400 863.400 892.200 ;
        RECT 864.600 890.400 866.400 897.000 ;
        RECT 860.700 883.050 861.600 890.400 ;
        RECT 862.500 888.600 864.300 889.500 ;
        RECT 869.100 888.600 870.900 896.400 ;
        RECT 886.500 890.400 888.300 897.000 ;
        RECT 891.000 890.400 892.800 896.400 ;
        RECT 895.500 890.400 897.300 897.000 ;
        RECT 911.100 893.400 912.900 897.000 ;
        RECT 914.100 893.400 915.900 896.400 ;
        RECT 917.100 893.400 918.900 897.000 ;
        RECT 929.100 893.400 930.900 896.400 ;
        RECT 862.500 887.700 870.900 888.600 ;
        RECT 823.950 880.950 826.050 883.050 ;
        RECT 826.950 880.950 829.050 883.050 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 844.950 880.950 847.050 883.050 ;
        RECT 860.100 880.950 862.200 883.050 ;
        RECT 863.400 880.950 865.500 883.050 ;
        RECT 784.950 878.550 789.450 880.050 ;
        RECT 784.950 877.950 789.000 878.550 ;
        RECT 776.400 867.900 783.000 868.800 ;
        RECT 776.400 867.600 777.900 867.900 ;
        RECT 773.100 861.000 774.900 867.600 ;
        RECT 776.100 861.600 777.900 867.600 ;
        RECT 782.100 867.600 783.000 867.900 ;
        RECT 797.700 867.600 798.900 880.950 ;
        RECT 800.100 879.150 801.900 880.950 ;
        RECT 815.250 879.150 817.050 880.950 ;
        RECT 822.000 873.600 823.050 880.950 ;
        RECT 827.100 879.150 828.900 880.950 ;
        RECT 842.100 879.150 843.900 880.950 ;
        RECT 779.100 861.000 780.900 867.000 ;
        RECT 782.100 861.600 783.900 867.600 ;
        RECT 797.100 861.600 798.900 867.600 ;
        RECT 800.100 861.000 801.900 867.600 ;
        RECT 816.600 861.000 818.400 873.600 ;
        RECT 821.100 861.600 824.400 873.600 ;
        RECT 827.100 861.000 828.900 873.600 ;
        RECT 845.100 867.600 846.300 880.950 ;
        RECT 860.700 873.600 861.600 880.950 ;
        RECT 864.000 879.150 865.800 880.950 ;
        RECT 842.100 861.000 843.900 867.600 ;
        RECT 845.100 861.600 846.900 867.600 ;
        RECT 860.100 861.600 861.900 873.600 ;
        RECT 863.100 861.000 864.900 873.000 ;
        RECT 867.000 867.600 867.900 887.700 ;
        RECT 868.950 883.050 870.750 884.850 ;
        RECT 884.100 883.050 885.900 884.850 ;
        RECT 890.700 883.050 891.900 890.400 ;
        RECT 895.950 883.050 897.750 884.850 ;
        RECT 914.400 883.050 915.300 893.400 ;
        RECT 929.100 889.500 930.300 893.400 ;
        RECT 932.100 890.400 933.900 897.000 ;
        RECT 935.100 890.400 936.900 896.400 ;
        RECT 929.100 888.600 934.800 889.500 ;
        RECT 933.000 887.700 934.800 888.600 ;
        RECT 868.800 880.950 870.900 883.050 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 886.950 880.950 889.050 883.050 ;
        RECT 889.950 880.950 892.050 883.050 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 910.950 880.950 913.050 883.050 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 929.400 880.950 931.500 883.050 ;
        RECT 887.100 879.150 888.900 880.950 ;
        RECT 891.000 875.400 891.900 880.950 ;
        RECT 892.950 879.150 894.750 880.950 ;
        RECT 911.250 879.150 913.050 880.950 ;
        RECT 887.100 874.500 891.900 875.400 ;
        RECT 866.100 861.600 867.900 867.600 ;
        RECT 869.100 861.000 870.900 867.600 ;
        RECT 884.100 862.500 885.900 873.600 ;
        RECT 887.100 863.400 888.900 874.500 ;
        RECT 914.400 873.600 915.300 880.950 ;
        RECT 917.100 879.150 918.900 880.950 ;
        RECT 929.400 879.150 931.200 880.950 ;
        RECT 933.000 876.300 933.900 887.700 ;
        RECT 935.700 883.050 936.900 890.400 ;
        RECT 934.800 880.950 936.900 883.050 ;
        RECT 933.000 875.400 934.800 876.300 ;
        RECT 929.100 874.500 934.800 875.400 ;
        RECT 890.100 872.400 897.900 873.300 ;
        RECT 890.100 862.500 891.900 872.400 ;
        RECT 884.100 861.600 891.900 862.500 ;
        RECT 893.100 861.000 894.900 871.500 ;
        RECT 896.100 861.600 897.900 872.400 ;
        RECT 911.100 861.000 912.900 873.600 ;
        RECT 914.400 872.400 918.000 873.600 ;
        RECT 916.200 861.600 918.000 872.400 ;
        RECT 929.100 867.600 930.300 874.500 ;
        RECT 935.700 873.600 936.900 880.950 ;
        RECT 929.100 861.600 930.900 867.600 ;
        RECT 932.100 861.000 933.900 871.800 ;
        RECT 935.100 861.600 936.900 873.600 ;
        RECT 14.400 845.400 16.200 858.000 ;
        RECT 19.500 846.900 21.300 857.400 ;
        RECT 22.500 851.400 24.300 858.000 ;
        RECT 35.700 851.400 37.500 858.000 ;
        RECT 22.200 848.100 24.000 849.900 ;
        RECT 36.000 848.100 37.800 849.900 ;
        RECT 38.700 846.900 40.500 857.400 ;
        RECT 19.500 845.400 21.900 846.900 ;
        RECT 14.100 838.050 15.900 839.850 ;
        RECT 20.700 838.050 21.900 845.400 ;
        RECT 38.100 845.400 40.500 846.900 ;
        RECT 43.800 845.400 45.600 858.000 ;
        RECT 59.700 851.400 61.500 858.000 ;
        RECT 60.000 848.100 61.800 849.900 ;
        RECT 62.700 846.900 64.500 857.400 ;
        RECT 62.100 845.400 64.500 846.900 ;
        RECT 67.800 845.400 69.600 858.000 ;
        RECT 83.700 851.400 85.500 858.000 ;
        RECT 84.000 848.100 85.800 849.900 ;
        RECT 86.700 846.900 88.500 857.400 ;
        RECT 86.100 845.400 88.500 846.900 ;
        RECT 91.800 845.400 93.600 858.000 ;
        RECT 104.100 851.400 105.900 858.000 ;
        RECT 107.100 851.400 108.900 857.400 ;
        RECT 110.100 851.400 111.900 858.000 ;
        RECT 122.700 851.400 124.500 858.000 ;
        RECT 25.950 838.950 34.050 841.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 22.950 835.950 25.050 838.050 ;
        RECT 17.100 834.150 18.900 835.950 ;
        RECT 20.700 831.600 21.900 835.950 ;
        RECT 23.100 834.150 24.900 835.950 ;
        RECT 29.550 835.050 30.450 838.950 ;
        RECT 38.100 838.050 39.300 845.400 ;
        RECT 52.950 843.450 55.050 844.050 ;
        RECT 58.950 843.450 61.050 844.050 ;
        RECT 52.950 842.550 61.050 843.450 ;
        RECT 52.950 841.950 55.050 842.550 ;
        RECT 58.950 841.950 61.050 842.550 ;
        RECT 44.100 838.050 45.900 839.850 ;
        RECT 62.100 838.050 63.300 845.400 ;
        RECT 68.100 838.050 69.900 839.850 ;
        RECT 86.100 838.050 87.300 845.400 ;
        RECT 92.100 838.050 93.900 839.850 ;
        RECT 107.100 838.050 108.300 851.400 ;
        RECT 123.000 848.100 124.800 849.900 ;
        RECT 125.700 846.900 127.500 857.400 ;
        RECT 125.100 845.400 127.500 846.900 ;
        RECT 130.800 845.400 132.600 858.000 ;
        RECT 146.100 851.400 147.900 858.000 ;
        RECT 149.100 851.400 150.900 857.400 ;
        RECT 117.000 840.450 121.050 841.050 ;
        RECT 116.550 838.950 121.050 840.450 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 43.950 835.950 46.050 838.050 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 88.950 835.950 91.050 838.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 29.550 833.550 34.050 835.050 ;
        RECT 35.100 834.150 36.900 835.950 ;
        RECT 30.000 832.950 34.050 833.550 ;
        RECT 20.700 830.700 24.300 831.600 ;
        RECT 14.100 827.700 21.900 829.050 ;
        RECT 14.100 822.600 15.900 827.700 ;
        RECT 17.100 822.000 18.900 826.800 ;
        RECT 20.100 822.600 21.900 827.700 ;
        RECT 23.100 828.600 24.300 830.700 ;
        RECT 28.950 829.050 31.050 832.050 ;
        RECT 38.100 831.600 39.300 835.950 ;
        RECT 41.100 834.150 42.900 835.950 ;
        RECT 59.100 834.150 60.900 835.950 ;
        RECT 62.100 831.600 63.300 835.950 ;
        RECT 65.100 834.150 66.900 835.950 ;
        RECT 83.100 834.150 84.900 835.950 ;
        RECT 86.100 831.600 87.300 835.950 ;
        RECT 89.100 834.150 90.900 835.950 ;
        RECT 104.250 834.150 106.050 835.950 ;
        RECT 35.700 830.700 39.300 831.600 ;
        RECT 59.700 830.700 63.300 831.600 ;
        RECT 83.700 830.700 87.300 831.600 ;
        RECT 107.100 830.700 108.300 835.950 ;
        RECT 110.100 834.150 111.900 835.950 ;
        RECT 116.550 835.050 117.450 838.950 ;
        RECT 125.100 838.050 126.300 845.400 ;
        RECT 131.100 838.050 132.900 839.850 ;
        RECT 146.100 838.050 147.900 839.850 ;
        RECT 149.100 838.050 150.300 851.400 ;
        RECT 161.100 846.600 162.900 857.400 ;
        RECT 164.100 847.500 165.900 858.000 ;
        RECT 161.100 845.400 165.900 846.600 ;
        RECT 163.800 844.500 165.900 845.400 ;
        RECT 168.600 845.400 170.400 857.400 ;
        RECT 173.100 847.500 174.900 858.000 ;
        RECT 176.100 846.300 177.900 857.400 ;
        RECT 188.100 851.400 189.900 858.000 ;
        RECT 191.100 851.400 192.900 857.400 ;
        RECT 173.400 845.400 177.900 846.300 ;
        RECT 168.600 844.050 169.800 845.400 ;
        RECT 168.300 843.000 169.800 844.050 ;
        RECT 173.400 843.300 175.500 845.400 ;
        RECT 168.300 841.050 169.200 843.000 ;
        RECT 161.400 838.050 163.200 839.850 ;
        RECT 167.100 838.950 169.200 841.050 ;
        RECT 170.100 841.500 172.200 841.800 ;
        RECT 170.100 839.700 174.000 841.500 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 130.950 835.950 133.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 148.950 835.950 151.050 838.050 ;
        RECT 161.100 835.950 163.200 838.050 ;
        RECT 167.700 838.800 169.200 838.950 ;
        RECT 167.700 837.900 170.100 838.800 ;
        RECT 112.950 833.550 117.450 835.050 ;
        RECT 122.100 834.150 123.900 835.950 ;
        RECT 112.950 832.950 117.000 833.550 ;
        RECT 125.100 831.600 126.300 835.950 ;
        RECT 128.100 834.150 129.900 835.950 ;
        RECT 122.700 830.700 126.300 831.600 ;
        RECT 28.950 828.900 33.000 829.050 ;
        RECT 23.100 822.600 24.900 828.600 ;
        RECT 28.950 828.000 34.050 828.900 ;
        RECT 35.700 828.600 36.900 830.700 ;
        RECT 29.550 827.550 34.050 828.000 ;
        RECT 30.000 826.950 34.050 827.550 ;
        RECT 31.950 826.800 34.050 826.950 ;
        RECT 35.100 822.600 36.900 828.600 ;
        RECT 38.100 827.700 45.900 829.050 ;
        RECT 59.700 828.600 60.900 830.700 ;
        RECT 38.100 822.600 39.900 827.700 ;
        RECT 41.100 822.000 42.900 826.800 ;
        RECT 44.100 822.600 45.900 827.700 ;
        RECT 59.100 822.600 60.900 828.600 ;
        RECT 62.100 827.700 69.900 829.050 ;
        RECT 83.700 828.600 84.900 830.700 ;
        RECT 107.100 829.800 111.300 830.700 ;
        RECT 62.100 822.600 63.900 827.700 ;
        RECT 65.100 822.000 66.900 826.800 ;
        RECT 68.100 822.600 69.900 827.700 ;
        RECT 83.100 822.600 84.900 828.600 ;
        RECT 86.100 827.700 93.900 829.050 ;
        RECT 86.100 822.600 87.900 827.700 ;
        RECT 89.100 822.000 90.900 826.800 ;
        RECT 92.100 822.600 93.900 827.700 ;
        RECT 104.400 822.000 106.200 828.600 ;
        RECT 109.500 822.600 111.300 829.800 ;
        RECT 122.700 828.600 123.900 830.700 ;
        RECT 122.100 822.600 123.900 828.600 ;
        RECT 125.100 827.700 132.900 829.050 ;
        RECT 125.100 822.600 126.900 827.700 ;
        RECT 128.100 822.000 129.900 826.800 ;
        RECT 131.100 822.600 132.900 827.700 ;
        RECT 149.100 825.600 150.300 835.950 ;
        RECT 165.900 835.200 167.700 837.000 ;
        RECT 165.900 833.100 168.000 835.200 ;
        RECT 168.900 832.200 170.100 837.900 ;
        RECT 171.000 838.050 172.800 838.500 ;
        RECT 188.100 838.050 189.900 839.850 ;
        RECT 191.100 838.050 192.300 851.400 ;
        RECT 206.100 845.400 207.900 857.400 ;
        RECT 209.100 846.300 210.900 857.400 ;
        RECT 212.100 847.200 213.900 858.000 ;
        RECT 215.100 846.300 216.900 857.400 ;
        RECT 230.100 851.400 231.900 858.000 ;
        RECT 233.100 851.400 234.900 857.400 ;
        RECT 209.100 845.400 216.900 846.300 ;
        RECT 206.400 838.050 207.300 845.400 ;
        RECT 211.950 838.050 213.750 839.850 ;
        RECT 230.100 838.050 231.900 839.850 ;
        RECT 233.100 838.050 234.300 851.400 ;
        RECT 248.100 846.600 249.900 857.400 ;
        RECT 251.100 847.500 252.900 858.000 ;
        RECT 248.100 845.400 252.900 846.600 ;
        RECT 250.800 844.500 252.900 845.400 ;
        RECT 255.600 845.400 257.400 857.400 ;
        RECT 260.100 847.500 261.900 858.000 ;
        RECT 263.100 846.300 264.900 857.400 ;
        RECT 260.400 845.400 264.900 846.300 ;
        RECT 279.000 846.600 280.800 857.400 ;
        RECT 279.000 845.400 282.600 846.600 ;
        RECT 284.100 845.400 285.900 858.000 ;
        RECT 296.100 851.400 297.900 858.000 ;
        RECT 299.100 851.400 300.900 857.400 ;
        RECT 255.600 844.050 256.800 845.400 ;
        RECT 255.300 843.000 256.800 844.050 ;
        RECT 260.400 843.300 262.500 845.400 ;
        RECT 255.300 841.050 256.200 843.000 ;
        RECT 248.400 838.050 250.200 839.850 ;
        RECT 254.100 838.950 256.200 841.050 ;
        RECT 257.100 841.500 259.200 841.800 ;
        RECT 257.100 839.700 261.000 841.500 ;
        RECT 171.000 836.700 177.900 838.050 ;
        RECT 175.800 835.950 177.900 836.700 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 248.100 835.950 250.200 838.050 ;
        RECT 254.700 838.800 256.200 838.950 ;
        RECT 254.700 837.900 257.100 838.800 ;
        RECT 163.800 829.500 165.900 830.700 ;
        RECT 167.100 830.100 170.100 832.200 ;
        RECT 171.000 833.400 172.800 835.200 ;
        RECT 175.800 834.150 177.600 835.950 ;
        RECT 171.000 831.300 173.100 833.400 ;
        RECT 171.000 830.400 177.300 831.300 ;
        RECT 161.100 828.600 165.900 829.500 ;
        RECT 168.900 828.600 170.100 830.100 ;
        RECT 176.100 828.600 177.300 830.400 ;
        RECT 146.100 822.000 147.900 825.600 ;
        RECT 149.100 822.600 150.900 825.600 ;
        RECT 161.100 822.600 162.900 828.600 ;
        RECT 164.100 822.000 165.900 827.700 ;
        RECT 168.600 822.600 170.400 828.600 ;
        RECT 173.100 822.000 174.900 827.700 ;
        RECT 176.100 822.600 177.900 828.600 ;
        RECT 191.100 825.600 192.300 835.950 ;
        RECT 206.400 828.600 207.300 835.950 ;
        RECT 208.950 834.150 210.750 835.950 ;
        RECT 215.100 834.150 216.900 835.950 ;
        RECT 206.400 827.400 211.500 828.600 ;
        RECT 188.100 822.000 189.900 825.600 ;
        RECT 191.100 822.600 192.900 825.600 ;
        RECT 206.700 822.000 208.500 825.600 ;
        RECT 209.700 822.600 211.500 827.400 ;
        RECT 214.200 822.000 216.000 828.600 ;
        RECT 233.100 825.600 234.300 835.950 ;
        RECT 252.900 835.200 254.700 837.000 ;
        RECT 252.900 833.100 255.000 835.200 ;
        RECT 255.900 832.200 257.100 837.900 ;
        RECT 258.000 838.050 259.800 838.500 ;
        RECT 278.100 838.050 279.900 839.850 ;
        RECT 281.700 838.050 282.600 845.400 ;
        RECT 283.950 838.050 285.750 839.850 ;
        RECT 258.000 836.700 264.900 838.050 ;
        RECT 262.800 835.950 264.900 836.700 ;
        RECT 277.950 835.950 280.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 296.100 835.950 298.200 838.050 ;
        RECT 250.800 829.500 252.900 830.700 ;
        RECT 254.100 830.100 257.100 832.200 ;
        RECT 258.000 833.400 259.800 835.200 ;
        RECT 262.800 834.150 264.600 835.950 ;
        RECT 258.000 831.300 260.100 833.400 ;
        RECT 258.000 830.400 264.300 831.300 ;
        RECT 248.100 828.600 252.900 829.500 ;
        RECT 255.900 828.600 257.100 830.100 ;
        RECT 263.100 828.600 264.300 830.400 ;
        RECT 230.100 822.000 231.900 825.600 ;
        RECT 233.100 822.600 234.900 825.600 ;
        RECT 248.100 822.600 249.900 828.600 ;
        RECT 251.100 822.000 252.900 827.700 ;
        RECT 255.600 822.600 257.400 828.600 ;
        RECT 260.100 822.000 261.900 827.700 ;
        RECT 263.100 822.600 264.900 828.600 ;
        RECT 268.950 828.450 271.050 829.050 ;
        RECT 277.950 828.450 280.050 829.050 ;
        RECT 268.950 827.550 280.050 828.450 ;
        RECT 268.950 826.950 271.050 827.550 ;
        RECT 277.950 826.950 280.050 827.550 ;
        RECT 281.700 825.600 282.600 835.950 ;
        RECT 296.250 834.150 298.050 835.950 ;
        RECT 299.100 831.300 300.000 851.400 ;
        RECT 302.100 846.000 303.900 858.000 ;
        RECT 305.100 845.400 306.900 857.400 ;
        RECT 320.100 851.400 321.900 858.000 ;
        RECT 323.100 851.400 324.900 857.400 ;
        RECT 326.100 851.400 327.900 858.000 ;
        RECT 301.200 838.050 303.000 839.850 ;
        RECT 305.400 838.050 306.300 845.400 ;
        RECT 323.100 838.050 324.300 851.400 ;
        RECT 342.000 846.600 343.800 857.400 ;
        RECT 342.000 845.400 345.600 846.600 ;
        RECT 347.100 845.400 348.900 858.000 ;
        RECT 362.100 846.300 363.900 857.400 ;
        RECT 365.100 847.200 366.900 858.000 ;
        RECT 368.100 846.300 369.900 857.400 ;
        RECT 362.100 845.400 369.900 846.300 ;
        RECT 371.100 845.400 372.900 857.400 ;
        RECT 383.100 845.400 384.900 858.000 ;
        RECT 388.200 846.600 390.000 857.400 ;
        RECT 386.400 845.400 390.000 846.600 ;
        RECT 404.100 845.400 405.900 858.000 ;
        RECT 409.200 846.600 411.000 857.400 ;
        RECT 407.400 845.400 411.000 846.600 ;
        RECT 425.100 846.600 426.900 857.400 ;
        RECT 428.100 847.500 429.900 858.000 ;
        RECT 431.100 856.500 438.900 857.400 ;
        RECT 431.100 846.600 432.900 856.500 ;
        RECT 425.100 845.700 432.900 846.600 ;
        RECT 341.100 838.050 342.900 839.850 ;
        RECT 344.700 838.050 345.600 845.400 ;
        RECT 346.950 838.050 348.750 839.850 ;
        RECT 365.250 838.050 367.050 839.850 ;
        RECT 371.700 838.050 372.600 845.400 ;
        RECT 383.250 838.050 385.050 839.850 ;
        RECT 386.400 838.050 387.300 845.400 ;
        RECT 389.100 838.050 390.900 839.850 ;
        RECT 404.250 838.050 406.050 839.850 ;
        RECT 407.400 838.050 408.300 845.400 ;
        RECT 434.100 844.500 435.900 855.600 ;
        RECT 437.100 845.400 438.900 856.500 ;
        RECT 452.100 851.400 453.900 858.000 ;
        RECT 455.100 851.400 456.900 857.400 ;
        RECT 470.100 851.400 471.900 857.400 ;
        RECT 473.100 851.400 474.900 858.000 ;
        RECT 431.100 843.600 435.900 844.500 ;
        RECT 420.000 840.450 424.050 841.050 ;
        RECT 410.100 838.050 411.900 839.850 ;
        RECT 419.550 838.950 424.050 840.450 ;
        RECT 301.500 835.950 303.600 838.050 ;
        RECT 304.800 835.950 306.900 838.050 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 296.100 830.400 304.500 831.300 ;
        RECT 278.100 822.000 279.900 825.600 ;
        RECT 281.100 822.600 282.900 825.600 ;
        RECT 284.100 822.000 285.900 825.600 ;
        RECT 296.100 822.600 297.900 830.400 ;
        RECT 302.700 829.500 304.500 830.400 ;
        RECT 305.400 828.600 306.300 835.950 ;
        RECT 320.250 834.150 322.050 835.950 ;
        RECT 323.100 830.700 324.300 835.950 ;
        RECT 326.100 834.150 327.900 835.950 ;
        RECT 323.100 829.800 327.300 830.700 ;
        RECT 300.600 822.000 302.400 828.600 ;
        RECT 303.600 826.800 306.300 828.600 ;
        RECT 303.600 822.600 305.400 826.800 ;
        RECT 320.400 822.000 322.200 828.600 ;
        RECT 325.500 822.600 327.300 829.800 ;
        RECT 344.700 825.600 345.600 835.950 ;
        RECT 362.100 834.150 363.900 835.950 ;
        RECT 368.250 834.150 370.050 835.950 ;
        RECT 371.700 828.600 372.600 835.950 ;
        RECT 341.100 822.000 342.900 825.600 ;
        RECT 344.100 822.600 345.900 825.600 ;
        RECT 347.100 822.000 348.900 825.600 ;
        RECT 363.000 822.000 364.800 828.600 ;
        RECT 367.500 827.400 372.600 828.600 ;
        RECT 367.500 822.600 369.300 827.400 ;
        RECT 386.400 825.600 387.300 835.950 ;
        RECT 388.950 831.450 391.050 832.050 ;
        RECT 397.950 831.450 400.050 832.050 ;
        RECT 388.950 830.550 400.050 831.450 ;
        RECT 388.950 829.950 391.050 830.550 ;
        RECT 397.950 829.950 400.050 830.550 ;
        RECT 407.400 825.600 408.300 835.950 ;
        RECT 419.550 834.450 420.450 838.950 ;
        RECT 428.250 838.050 430.050 839.850 ;
        RECT 431.100 838.050 432.000 843.600 ;
        RECT 439.950 840.450 442.050 841.050 ;
        RECT 445.950 840.450 448.050 841.050 ;
        RECT 434.100 838.050 435.900 839.850 ;
        RECT 439.950 839.550 448.050 840.450 ;
        RECT 439.950 838.950 442.050 839.550 ;
        RECT 445.950 838.950 448.050 839.550 ;
        RECT 452.100 838.050 453.900 839.850 ;
        RECT 455.100 838.050 456.300 851.400 ;
        RECT 470.700 838.050 471.900 851.400 ;
        RECT 488.100 845.400 489.900 858.000 ;
        RECT 491.100 844.500 492.900 857.400 ;
        RECT 494.100 845.400 495.900 858.000 ;
        RECT 497.100 844.500 498.900 857.400 ;
        RECT 500.100 845.400 501.900 858.000 ;
        RECT 503.100 844.500 504.900 857.400 ;
        RECT 506.100 845.400 507.900 858.000 ;
        RECT 509.100 844.500 510.900 857.400 ;
        RECT 512.100 845.400 513.900 858.000 ;
        RECT 527.100 851.400 528.900 858.000 ;
        RECT 530.100 851.400 531.900 857.400 ;
        RECT 542.100 851.400 543.900 857.400 ;
        RECT 490.050 843.300 492.900 844.500 ;
        RECT 495.000 843.300 498.900 844.500 ;
        RECT 501.000 843.300 504.900 844.500 ;
        RECT 507.000 843.300 510.900 844.500 ;
        RECT 473.100 838.050 474.900 839.850 ;
        RECT 490.050 838.050 491.100 843.300 ;
        RECT 424.950 835.950 427.050 838.050 ;
        RECT 427.950 835.950 430.050 838.050 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 451.950 835.950 454.050 838.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 469.950 835.950 472.050 838.050 ;
        RECT 472.950 835.950 475.050 838.050 ;
        RECT 490.050 835.950 493.200 838.050 ;
        RECT 413.550 833.550 420.450 834.450 ;
        RECT 425.250 834.150 427.050 835.950 ;
        RECT 413.550 832.050 414.450 833.550 ;
        RECT 411.000 831.750 414.450 832.050 ;
        RECT 409.950 830.550 414.450 831.750 ;
        RECT 415.950 831.450 418.050 832.050 ;
        RECT 427.950 831.450 430.050 831.750 ;
        RECT 415.950 830.550 430.050 831.450 ;
        RECT 409.950 829.950 414.000 830.550 ;
        RECT 415.950 829.950 418.050 830.550 ;
        RECT 409.950 829.650 412.050 829.950 ;
        RECT 427.950 829.650 430.050 830.550 ;
        RECT 431.100 828.600 432.300 835.950 ;
        RECT 437.100 834.150 438.900 835.950 ;
        RECT 370.500 822.000 372.300 825.600 ;
        RECT 383.100 822.000 384.900 825.600 ;
        RECT 386.100 822.600 387.900 825.600 ;
        RECT 389.100 822.000 390.900 825.600 ;
        RECT 404.100 822.000 405.900 825.600 ;
        RECT 407.100 822.600 408.900 825.600 ;
        RECT 410.100 822.000 411.900 825.600 ;
        RECT 425.700 822.000 427.500 828.600 ;
        RECT 430.200 822.600 432.000 828.600 ;
        RECT 434.700 822.000 436.500 828.600 ;
        RECT 455.100 825.600 456.300 835.950 ;
        RECT 470.700 825.600 471.900 835.950 ;
        RECT 490.050 830.700 491.100 835.950 ;
        RECT 492.000 832.800 493.800 833.400 ;
        RECT 495.000 832.800 496.200 843.300 ;
        RECT 492.000 831.600 496.200 832.800 ;
        RECT 498.000 832.800 499.800 833.400 ;
        RECT 501.000 832.800 502.200 843.300 ;
        RECT 498.000 831.600 502.200 832.800 ;
        RECT 504.000 832.800 505.800 833.400 ;
        RECT 507.000 832.800 508.200 843.300 ;
        RECT 527.100 838.050 528.900 839.850 ;
        RECT 530.100 838.050 531.300 851.400 ;
        RECT 542.100 844.500 543.300 851.400 ;
        RECT 545.100 847.200 546.900 858.000 ;
        RECT 548.100 845.400 549.900 857.400 ;
        RECT 563.100 851.400 564.900 858.000 ;
        RECT 566.100 851.400 567.900 857.400 ;
        RECT 569.100 851.400 570.900 858.000 ;
        RECT 542.100 843.600 547.800 844.500 ;
        RECT 546.000 842.700 547.800 843.600 ;
        RECT 542.400 838.050 544.200 839.850 ;
        RECT 509.100 835.950 511.200 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 542.400 835.950 544.500 838.050 ;
        RECT 509.400 834.150 511.200 835.950 ;
        RECT 504.000 831.600 508.200 832.800 ;
        RECT 495.000 830.700 496.200 831.600 ;
        RECT 501.000 830.700 502.200 831.600 ;
        RECT 507.000 830.700 508.200 831.600 ;
        RECT 490.050 829.500 492.900 830.700 ;
        RECT 495.000 829.500 498.900 830.700 ;
        RECT 501.000 829.500 504.900 830.700 ;
        RECT 507.000 829.500 510.900 830.700 ;
        RECT 452.100 822.000 453.900 825.600 ;
        RECT 455.100 822.600 456.900 825.600 ;
        RECT 470.100 822.600 471.900 825.600 ;
        RECT 473.100 822.000 474.900 825.600 ;
        RECT 488.100 822.000 489.900 828.600 ;
        RECT 491.100 822.600 492.900 829.500 ;
        RECT 494.100 822.000 495.900 828.600 ;
        RECT 497.100 822.600 498.900 829.500 ;
        RECT 500.100 822.000 501.900 828.600 ;
        RECT 503.100 822.600 504.900 829.500 ;
        RECT 506.100 822.000 507.900 828.600 ;
        RECT 509.100 822.600 510.900 829.500 ;
        RECT 512.100 822.000 513.900 828.600 ;
        RECT 530.100 825.600 531.300 835.950 ;
        RECT 546.000 831.300 546.900 842.700 ;
        RECT 548.700 838.050 549.900 845.400 ;
        RECT 553.950 843.450 556.050 844.050 ;
        RECT 562.950 843.450 565.050 844.050 ;
        RECT 553.950 842.550 565.050 843.450 ;
        RECT 553.950 841.950 556.050 842.550 ;
        RECT 562.950 841.950 565.050 842.550 ;
        RECT 566.100 838.050 567.300 851.400 ;
        RECT 582.000 846.600 583.800 857.400 ;
        RECT 582.000 845.400 585.600 846.600 ;
        RECT 587.100 845.400 588.900 858.000 ;
        RECT 602.100 851.400 603.900 857.400 ;
        RECT 605.100 851.400 606.900 858.000 ;
        RECT 571.950 840.450 576.000 841.050 ;
        RECT 571.950 838.950 576.450 840.450 ;
        RECT 547.800 835.950 549.900 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 546.000 830.400 547.800 831.300 ;
        RECT 542.100 829.500 547.800 830.400 ;
        RECT 542.100 825.600 543.300 829.500 ;
        RECT 548.700 828.600 549.900 835.950 ;
        RECT 563.250 834.150 565.050 835.950 ;
        RECT 566.100 830.700 567.300 835.950 ;
        RECT 569.100 834.150 570.900 835.950 ;
        RECT 575.550 835.050 576.450 838.950 ;
        RECT 581.100 838.050 582.900 839.850 ;
        RECT 584.700 838.050 585.600 845.400 ;
        RECT 586.950 838.050 588.750 839.850 ;
        RECT 602.700 838.050 603.900 851.400 ;
        RECT 618.000 846.600 619.800 857.400 ;
        RECT 618.000 845.400 621.600 846.600 ;
        RECT 623.100 845.400 624.900 858.000 ;
        RECT 626.700 851.400 628.500 858.000 ;
        RECT 629.700 852.300 631.500 857.400 ;
        RECT 629.400 851.400 631.500 852.300 ;
        RECT 632.700 851.400 634.500 858.000 ;
        RECT 629.400 850.500 630.300 851.400 ;
        RECT 626.700 849.600 630.300 850.500 ;
        RECT 612.000 840.450 616.050 841.050 ;
        RECT 605.100 838.050 606.900 839.850 ;
        RECT 611.550 838.950 616.050 840.450 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 571.950 833.550 576.450 835.050 ;
        RECT 571.950 832.950 576.000 833.550 ;
        RECT 566.100 829.800 570.300 830.700 ;
        RECT 527.100 822.000 528.900 825.600 ;
        RECT 530.100 822.600 531.900 825.600 ;
        RECT 542.100 822.600 543.900 825.600 ;
        RECT 545.100 822.000 546.900 828.600 ;
        RECT 548.100 822.600 549.900 828.600 ;
        RECT 563.400 822.000 565.200 828.600 ;
        RECT 568.500 822.600 570.300 829.800 ;
        RECT 584.700 825.600 585.600 835.950 ;
        RECT 602.700 825.600 603.900 835.950 ;
        RECT 611.550 835.050 612.450 838.950 ;
        RECT 617.100 838.050 618.900 839.850 ;
        RECT 620.700 838.050 621.600 845.400 ;
        RECT 622.950 838.050 624.750 839.850 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 611.550 833.550 616.050 835.050 ;
        RECT 612.000 832.950 616.050 833.550 ;
        RECT 620.700 825.600 621.600 835.950 ;
        RECT 626.700 833.400 627.900 849.600 ;
        RECT 631.200 848.400 633.000 848.700 ;
        RECT 635.700 848.400 637.500 857.400 ;
        RECT 638.700 851.400 640.500 858.000 ;
        RECT 642.300 854.400 644.100 857.400 ;
        RECT 645.300 854.400 647.100 857.400 ;
        RECT 642.300 852.300 644.400 854.400 ;
        RECT 645.300 852.300 647.400 854.400 ;
        RECT 648.300 851.400 650.100 857.400 ;
        RECT 651.300 851.400 653.100 858.000 ;
        RECT 647.700 849.300 649.800 851.400 ;
        RECT 655.200 849.900 657.000 857.400 ;
        RECT 658.200 851.400 660.000 858.000 ;
        RECT 661.200 851.400 663.000 857.400 ;
        RECT 664.200 854.400 666.000 857.400 ;
        RECT 667.200 854.400 669.000 857.400 ;
        RECT 670.200 854.400 672.000 857.400 ;
        RECT 664.200 852.300 666.300 854.400 ;
        RECT 667.200 852.300 669.300 854.400 ;
        RECT 670.200 852.300 672.300 854.400 ;
        RECT 673.200 851.400 675.000 858.000 ;
        RECT 676.200 851.400 678.000 857.400 ;
        RECT 679.200 851.400 681.000 858.000 ;
        RECT 682.200 851.400 684.000 857.400 ;
        RECT 685.200 851.400 687.000 858.000 ;
        RECT 688.500 851.400 690.300 857.400 ;
        RECT 691.500 851.400 693.300 858.000 ;
        RECT 707.100 851.400 708.900 858.000 ;
        RECT 710.100 851.400 711.900 857.400 ;
        RECT 713.100 851.400 714.900 858.000 ;
        RECT 631.200 847.200 650.400 848.400 ;
        RECT 655.200 847.800 658.500 849.900 ;
        RECT 661.200 847.500 663.900 851.400 ;
        RECT 667.200 850.500 669.300 851.400 ;
        RECT 667.200 849.300 675.300 850.500 ;
        RECT 673.500 848.700 675.300 849.300 ;
        RECT 676.200 848.400 677.400 851.400 ;
        RECT 682.800 850.500 684.000 851.400 ;
        RECT 682.800 849.600 686.700 850.500 ;
        RECT 680.100 848.400 681.900 849.000 ;
        RECT 631.200 846.900 633.000 847.200 ;
        RECT 649.200 846.600 650.400 847.200 ;
        RECT 664.800 846.600 666.900 847.500 ;
        RECT 634.500 845.700 636.300 846.300 ;
        RECT 644.400 845.700 646.500 846.300 ;
        RECT 634.500 844.500 646.500 845.700 ;
        RECT 649.200 845.400 666.900 846.600 ;
        RECT 670.200 846.300 672.300 847.500 ;
        RECT 676.200 847.200 681.900 848.400 ;
        RECT 685.800 846.300 686.700 849.600 ;
        RECT 670.200 845.400 686.700 846.300 ;
        RECT 644.400 844.200 646.500 844.500 ;
        RECT 649.200 843.300 684.900 844.500 ;
        RECT 649.200 842.700 650.400 843.300 ;
        RECT 683.100 842.700 684.900 843.300 ;
        RECT 636.900 841.800 650.400 842.700 ;
        RECT 661.800 841.800 663.900 842.100 ;
        RECT 636.900 841.050 638.700 841.800 ;
        RECT 628.800 838.950 630.900 841.050 ;
        RECT 634.800 839.250 638.700 841.050 ;
        RECT 656.400 840.300 658.500 841.200 ;
        RECT 634.800 838.950 636.900 839.250 ;
        RECT 647.400 839.100 658.500 840.300 ;
        RECT 660.000 840.000 663.900 841.800 ;
        RECT 668.100 840.300 669.900 842.100 ;
        RECT 669.000 839.100 669.900 840.300 ;
        RECT 629.100 837.300 630.900 838.950 ;
        RECT 647.400 838.500 649.200 839.100 ;
        RECT 656.400 838.200 669.900 839.100 ;
        RECT 672.600 838.800 677.700 840.600 ;
        RECT 679.800 838.950 681.900 841.050 ;
        RECT 672.600 837.300 673.500 838.800 ;
        RECT 629.100 836.100 673.500 837.300 ;
        RECT 679.800 836.100 681.300 838.950 ;
        RECT 644.400 833.400 646.200 835.200 ;
        RECT 652.800 834.000 654.900 835.050 ;
        RECT 674.700 834.600 681.300 836.100 ;
        RECT 626.700 832.200 643.500 833.400 ;
        RECT 626.700 828.600 627.900 832.200 ;
        RECT 641.400 831.300 643.500 832.200 ;
        RECT 630.900 830.700 632.700 831.300 ;
        RECT 630.900 829.500 639.300 830.700 ;
        RECT 637.800 828.600 639.300 829.500 ;
        RECT 644.400 830.400 645.300 833.400 ;
        RECT 649.800 833.100 654.900 834.000 ;
        RECT 649.800 832.200 651.600 833.100 ;
        RECT 652.800 832.950 654.900 833.100 ;
        RECT 659.100 833.100 676.200 834.600 ;
        RECT 659.100 832.500 661.200 833.100 ;
        RECT 659.100 830.700 660.900 832.500 ;
        RECT 677.100 831.900 684.900 833.700 ;
        RECT 644.400 829.200 651.600 830.400 ;
        RECT 646.800 828.600 648.600 829.200 ;
        RECT 650.700 828.600 651.600 829.200 ;
        RECT 666.300 828.600 672.900 830.400 ;
        RECT 677.100 828.600 678.600 831.900 ;
        RECT 685.800 828.600 686.700 845.400 ;
        RECT 581.100 822.000 582.900 825.600 ;
        RECT 584.100 822.600 585.900 825.600 ;
        RECT 587.100 822.000 588.900 825.600 ;
        RECT 602.100 822.600 603.900 825.600 ;
        RECT 605.100 822.000 606.900 825.600 ;
        RECT 617.100 822.000 618.900 825.600 ;
        RECT 620.100 822.600 621.900 825.600 ;
        RECT 623.100 822.000 624.900 825.600 ;
        RECT 626.700 822.600 628.500 828.600 ;
        RECT 632.100 822.000 633.900 828.600 ;
        RECT 637.500 822.600 639.300 828.600 ;
        RECT 641.700 825.600 643.800 827.700 ;
        RECT 644.700 825.600 646.800 827.700 ;
        RECT 647.700 825.600 649.800 827.700 ;
        RECT 650.700 827.400 653.400 828.600 ;
        RECT 651.600 826.500 653.400 827.400 ;
        RECT 655.200 826.500 657.900 828.600 ;
        RECT 641.700 822.600 643.500 825.600 ;
        RECT 644.700 822.600 646.500 825.600 ;
        RECT 647.700 822.600 649.500 825.600 ;
        RECT 650.700 822.000 652.500 825.600 ;
        RECT 655.200 822.600 657.000 826.500 ;
        RECT 661.200 825.600 663.300 827.700 ;
        RECT 664.200 825.600 666.300 827.700 ;
        RECT 667.200 825.600 669.300 827.700 ;
        RECT 670.200 825.600 672.300 827.700 ;
        RECT 674.400 827.400 678.600 828.600 ;
        RECT 658.200 822.000 660.000 825.600 ;
        RECT 661.200 822.600 663.000 825.600 ;
        RECT 664.200 822.600 666.000 825.600 ;
        RECT 667.200 822.600 669.000 825.600 ;
        RECT 670.200 822.600 672.000 825.600 ;
        RECT 674.400 822.600 676.200 827.400 ;
        RECT 679.500 822.000 681.300 828.600 ;
        RECT 684.900 822.600 686.700 828.600 ;
        RECT 688.500 841.050 690.000 851.400 ;
        RECT 694.950 843.450 697.050 844.050 ;
        RECT 700.950 843.450 703.050 844.050 ;
        RECT 706.950 843.450 709.050 844.050 ;
        RECT 694.950 842.550 709.050 843.450 ;
        RECT 694.950 841.950 697.050 842.550 ;
        RECT 700.950 841.950 703.050 842.550 ;
        RECT 706.950 841.950 709.050 842.550 ;
        RECT 688.500 838.950 690.900 841.050 ;
        RECT 688.500 825.600 690.000 838.950 ;
        RECT 710.700 838.050 711.900 851.400 ;
        RECT 728.100 845.400 729.900 857.400 ;
        RECT 731.100 847.200 732.900 858.000 ;
        RECT 734.100 851.400 735.900 857.400 ;
        RECT 749.100 851.400 750.900 858.000 ;
        RECT 752.100 851.400 753.900 857.400 ;
        RECT 728.100 838.050 729.300 845.400 ;
        RECT 734.700 844.500 735.900 851.400 ;
        RECT 730.200 843.600 735.900 844.500 ;
        RECT 730.200 842.700 732.000 843.600 ;
        RECT 706.950 835.950 709.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 728.100 835.950 730.200 838.050 ;
        RECT 707.100 834.150 708.900 835.950 ;
        RECT 710.700 830.700 711.900 835.950 ;
        RECT 712.950 834.150 714.750 835.950 ;
        RECT 707.700 829.800 711.900 830.700 ;
        RECT 688.500 822.600 690.300 825.600 ;
        RECT 691.500 822.000 693.300 825.600 ;
        RECT 707.700 822.600 709.500 829.800 ;
        RECT 728.100 828.600 729.300 835.950 ;
        RECT 731.100 831.300 732.000 842.700 ;
        RECT 733.800 838.050 735.600 839.850 ;
        RECT 749.100 838.050 750.900 839.850 ;
        RECT 752.100 838.050 753.300 851.400 ;
        RECT 767.100 846.300 768.900 857.400 ;
        RECT 770.100 847.200 771.900 858.000 ;
        RECT 773.100 846.300 774.900 857.400 ;
        RECT 767.100 845.400 774.900 846.300 ;
        RECT 776.100 845.400 777.900 857.400 ;
        RECT 779.700 851.400 781.500 858.000 ;
        RECT 782.700 851.400 784.500 857.400 ;
        RECT 786.000 851.400 787.800 858.000 ;
        RECT 789.000 851.400 790.800 857.400 ;
        RECT 792.000 851.400 793.800 858.000 ;
        RECT 795.000 851.400 796.800 857.400 ;
        RECT 798.000 851.400 799.800 858.000 ;
        RECT 801.000 854.400 802.800 857.400 ;
        RECT 804.000 854.400 805.800 857.400 ;
        RECT 807.000 854.400 808.800 857.400 ;
        RECT 800.700 852.300 802.800 854.400 ;
        RECT 803.700 852.300 805.800 854.400 ;
        RECT 806.700 852.300 808.800 854.400 ;
        RECT 810.000 851.400 811.800 857.400 ;
        RECT 813.000 851.400 814.800 858.000 ;
        RECT 770.250 838.050 772.050 839.850 ;
        RECT 776.700 838.050 777.600 845.400 ;
        RECT 783.000 841.050 784.500 851.400 ;
        RECT 789.000 850.500 790.200 851.400 ;
        RECT 782.100 838.950 784.500 841.050 ;
        RECT 733.500 835.950 735.600 838.050 ;
        RECT 748.950 835.950 751.050 838.050 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 772.950 835.950 775.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 730.200 830.400 732.000 831.300 ;
        RECT 730.200 829.500 735.900 830.400 ;
        RECT 712.800 822.000 714.600 828.600 ;
        RECT 728.100 822.600 729.900 828.600 ;
        RECT 731.100 822.000 732.900 828.600 ;
        RECT 734.700 825.600 735.900 829.500 ;
        RECT 752.100 825.600 753.300 835.950 ;
        RECT 767.100 834.150 768.900 835.950 ;
        RECT 773.250 834.150 775.050 835.950 ;
        RECT 776.700 828.600 777.600 835.950 ;
        RECT 734.100 822.600 735.900 825.600 ;
        RECT 749.100 822.000 750.900 825.600 ;
        RECT 752.100 822.600 753.900 825.600 ;
        RECT 768.000 822.000 769.800 828.600 ;
        RECT 772.500 827.400 777.600 828.600 ;
        RECT 772.500 822.600 774.300 827.400 ;
        RECT 783.000 825.600 784.500 838.950 ;
        RECT 775.500 822.000 777.300 825.600 ;
        RECT 779.700 822.000 781.500 825.600 ;
        RECT 782.700 822.600 784.500 825.600 ;
        RECT 786.300 849.600 790.200 850.500 ;
        RECT 786.300 846.300 787.200 849.600 ;
        RECT 791.100 848.400 792.900 849.000 ;
        RECT 795.600 848.400 796.800 851.400 ;
        RECT 803.700 850.500 805.800 851.400 ;
        RECT 797.700 849.300 805.800 850.500 ;
        RECT 797.700 848.700 799.500 849.300 ;
        RECT 791.100 847.200 796.800 848.400 ;
        RECT 809.100 847.500 811.800 851.400 ;
        RECT 816.000 849.900 817.800 857.400 ;
        RECT 819.900 851.400 821.700 858.000 ;
        RECT 822.900 851.400 824.700 857.400 ;
        RECT 825.900 854.400 827.700 857.400 ;
        RECT 828.900 854.400 830.700 857.400 ;
        RECT 825.600 852.300 827.700 854.400 ;
        RECT 828.600 852.300 830.700 854.400 ;
        RECT 832.500 851.400 834.300 858.000 ;
        RECT 814.500 847.800 817.800 849.900 ;
        RECT 823.200 849.300 825.300 851.400 ;
        RECT 835.500 848.400 837.300 857.400 ;
        RECT 838.500 851.400 840.300 858.000 ;
        RECT 841.500 852.300 843.300 857.400 ;
        RECT 841.500 851.400 843.600 852.300 ;
        RECT 844.500 851.400 846.300 858.000 ;
        RECT 857.700 851.400 859.500 858.000 ;
        RECT 842.700 850.500 843.600 851.400 ;
        RECT 842.700 849.600 846.300 850.500 ;
        RECT 840.000 848.400 841.800 848.700 ;
        RECT 800.700 846.300 802.800 847.500 ;
        RECT 786.300 845.400 802.800 846.300 ;
        RECT 806.100 846.600 808.200 847.500 ;
        RECT 822.600 847.200 841.800 848.400 ;
        RECT 822.600 846.600 823.800 847.200 ;
        RECT 840.000 846.900 841.800 847.200 ;
        RECT 806.100 845.400 823.800 846.600 ;
        RECT 826.500 845.700 828.600 846.300 ;
        RECT 836.700 845.700 838.500 846.300 ;
        RECT 786.300 828.600 787.200 845.400 ;
        RECT 826.500 844.500 838.500 845.700 ;
        RECT 788.100 843.300 823.800 844.500 ;
        RECT 826.500 844.200 828.600 844.500 ;
        RECT 788.100 842.700 789.900 843.300 ;
        RECT 822.600 842.700 823.800 843.300 ;
        RECT 791.100 838.950 793.200 841.050 ;
        RECT 791.700 836.100 793.200 838.950 ;
        RECT 795.300 838.800 800.400 840.600 ;
        RECT 799.500 837.300 800.400 838.800 ;
        RECT 803.100 840.300 804.900 842.100 ;
        RECT 809.100 841.800 811.200 842.100 ;
        RECT 822.600 841.800 836.100 842.700 ;
        RECT 803.100 839.100 804.000 840.300 ;
        RECT 809.100 840.000 813.000 841.800 ;
        RECT 814.500 840.300 816.600 841.200 ;
        RECT 834.300 841.050 836.100 841.800 ;
        RECT 814.500 839.100 825.600 840.300 ;
        RECT 834.300 839.250 838.200 841.050 ;
        RECT 803.100 838.200 816.600 839.100 ;
        RECT 823.800 838.500 825.600 839.100 ;
        RECT 836.100 838.950 838.200 839.250 ;
        RECT 842.100 838.950 844.200 841.050 ;
        RECT 842.100 837.300 843.900 838.950 ;
        RECT 799.500 836.100 843.900 837.300 ;
        RECT 791.700 834.600 798.300 836.100 ;
        RECT 788.100 831.900 795.900 833.700 ;
        RECT 796.800 833.100 813.900 834.600 ;
        RECT 811.800 832.500 813.900 833.100 ;
        RECT 818.100 834.000 820.200 835.050 ;
        RECT 818.100 833.100 823.200 834.000 ;
        RECT 826.800 833.400 828.600 835.200 ;
        RECT 845.100 833.400 846.300 849.600 ;
        RECT 858.000 848.100 859.800 849.900 ;
        RECT 860.700 846.900 862.500 857.400 ;
        RECT 860.100 845.400 862.500 846.900 ;
        RECT 865.800 845.400 867.600 858.000 ;
        RECT 881.400 845.400 883.200 858.000 ;
        RECT 886.500 846.900 888.300 857.400 ;
        RECT 889.500 851.400 891.300 858.000 ;
        RECT 905.100 851.400 906.900 857.400 ;
        RECT 908.100 851.400 909.900 858.000 ;
        RECT 923.100 851.400 924.900 857.400 ;
        RECT 889.200 848.100 891.000 849.900 ;
        RECT 886.500 845.400 888.900 846.900 ;
        RECT 860.100 838.050 861.300 845.400 ;
        RECT 866.100 838.050 867.900 839.850 ;
        RECT 881.100 838.050 882.900 839.850 ;
        RECT 887.700 838.050 888.900 845.400 ;
        RECT 905.700 838.050 906.900 851.400 ;
        RECT 923.100 844.500 924.300 851.400 ;
        RECT 926.100 847.200 927.900 858.000 ;
        RECT 929.100 845.400 930.900 857.400 ;
        RECT 923.100 843.600 928.800 844.500 ;
        RECT 927.000 842.700 928.800 843.600 ;
        RECT 908.100 838.050 909.900 839.850 ;
        RECT 923.400 838.050 925.200 839.850 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 907.950 835.950 910.050 838.050 ;
        RECT 923.400 835.950 925.500 838.050 ;
        RECT 857.100 834.150 858.900 835.950 ;
        RECT 818.100 832.950 820.200 833.100 ;
        RECT 794.400 828.600 795.900 831.900 ;
        RECT 812.100 830.700 813.900 832.500 ;
        RECT 821.400 832.200 823.200 833.100 ;
        RECT 827.700 830.400 828.600 833.400 ;
        RECT 829.500 832.200 846.300 833.400 ;
        RECT 829.500 831.300 831.600 832.200 ;
        RECT 840.300 830.700 842.100 831.300 ;
        RECT 800.100 828.600 806.700 830.400 ;
        RECT 821.400 829.200 828.600 830.400 ;
        RECT 833.700 829.500 842.100 830.700 ;
        RECT 821.400 828.600 822.300 829.200 ;
        RECT 824.400 828.600 826.200 829.200 ;
        RECT 833.700 828.600 835.200 829.500 ;
        RECT 845.100 828.600 846.300 832.200 ;
        RECT 860.100 831.600 861.300 835.950 ;
        RECT 863.100 834.150 864.900 835.950 ;
        RECT 884.100 834.150 885.900 835.950 ;
        RECT 857.700 830.700 861.300 831.600 ;
        RECT 887.700 831.600 888.900 835.950 ;
        RECT 890.100 834.150 891.900 835.950 ;
        RECT 887.700 830.700 891.300 831.600 ;
        RECT 857.700 828.600 858.900 830.700 ;
        RECT 786.300 822.600 788.100 828.600 ;
        RECT 791.700 822.000 793.500 828.600 ;
        RECT 794.400 827.400 798.600 828.600 ;
        RECT 796.800 822.600 798.600 827.400 ;
        RECT 800.700 825.600 802.800 827.700 ;
        RECT 803.700 825.600 805.800 827.700 ;
        RECT 806.700 825.600 808.800 827.700 ;
        RECT 809.700 825.600 811.800 827.700 ;
        RECT 815.100 826.500 817.800 828.600 ;
        RECT 819.600 827.400 822.300 828.600 ;
        RECT 819.600 826.500 821.400 827.400 ;
        RECT 801.000 822.600 802.800 825.600 ;
        RECT 804.000 822.600 805.800 825.600 ;
        RECT 807.000 822.600 808.800 825.600 ;
        RECT 810.000 822.600 811.800 825.600 ;
        RECT 813.000 822.000 814.800 825.600 ;
        RECT 816.000 822.600 817.800 826.500 ;
        RECT 823.200 825.600 825.300 827.700 ;
        RECT 826.200 825.600 828.300 827.700 ;
        RECT 829.200 825.600 831.300 827.700 ;
        RECT 820.500 822.000 822.300 825.600 ;
        RECT 823.500 822.600 825.300 825.600 ;
        RECT 826.500 822.600 828.300 825.600 ;
        RECT 829.500 822.600 831.300 825.600 ;
        RECT 833.700 822.600 835.500 828.600 ;
        RECT 839.100 822.000 840.900 828.600 ;
        RECT 844.500 822.600 846.300 828.600 ;
        RECT 857.100 822.600 858.900 828.600 ;
        RECT 860.100 827.700 867.900 829.050 ;
        RECT 860.100 822.600 861.900 827.700 ;
        RECT 863.100 822.000 864.900 826.800 ;
        RECT 866.100 822.600 867.900 827.700 ;
        RECT 881.100 827.700 888.900 829.050 ;
        RECT 881.100 822.600 882.900 827.700 ;
        RECT 884.100 822.000 885.900 826.800 ;
        RECT 887.100 822.600 888.900 827.700 ;
        RECT 890.100 828.600 891.300 830.700 ;
        RECT 890.100 822.600 891.900 828.600 ;
        RECT 905.700 825.600 906.900 835.950 ;
        RECT 927.000 831.300 927.900 842.700 ;
        RECT 929.700 838.050 930.900 845.400 ;
        RECT 928.800 835.950 930.900 838.050 ;
        RECT 927.000 830.400 928.800 831.300 ;
        RECT 923.100 829.500 928.800 830.400 ;
        RECT 923.100 825.600 924.300 829.500 ;
        RECT 929.700 828.600 930.900 835.950 ;
        RECT 905.100 822.600 906.900 825.600 ;
        RECT 908.100 822.000 909.900 825.600 ;
        RECT 923.100 822.600 924.900 825.600 ;
        RECT 926.100 822.000 927.900 828.600 ;
        RECT 929.100 822.600 930.900 828.600 ;
        RECT 14.100 812.400 15.900 818.400 ;
        RECT 14.700 810.300 15.900 812.400 ;
        RECT 17.100 813.300 18.900 818.400 ;
        RECT 20.100 814.200 21.900 819.000 ;
        RECT 23.100 813.300 24.900 818.400 ;
        RECT 17.100 811.950 24.900 813.300 ;
        RECT 39.000 812.400 40.800 819.000 ;
        RECT 43.500 813.600 45.300 818.400 ;
        RECT 46.500 815.400 48.300 819.000 ;
        RECT 43.500 812.400 48.600 813.600 ;
        RECT 62.100 812.400 63.900 818.400 ;
        RECT 65.100 813.300 66.900 819.000 ;
        RECT 69.600 812.400 71.400 818.400 ;
        RECT 74.100 813.300 75.900 819.000 ;
        RECT 77.100 812.400 78.900 818.400 ;
        RECT 14.700 809.400 18.300 810.300 ;
        RECT 14.100 805.050 15.900 806.850 ;
        RECT 17.100 805.050 18.300 809.400 ;
        RECT 20.100 805.050 21.900 806.850 ;
        RECT 38.100 805.050 39.900 806.850 ;
        RECT 44.250 805.050 46.050 806.850 ;
        RECT 47.700 805.050 48.600 812.400 ;
        RECT 62.700 810.600 63.900 812.400 ;
        RECT 69.900 810.900 71.100 812.400 ;
        RECT 74.100 811.500 78.900 812.400 ;
        RECT 89.100 813.300 90.900 818.400 ;
        RECT 92.100 814.200 93.900 819.000 ;
        RECT 95.100 813.300 96.900 818.400 ;
        RECT 89.100 811.950 96.900 813.300 ;
        RECT 98.100 812.400 99.900 818.400 ;
        RECT 113.100 813.300 114.900 818.400 ;
        RECT 116.100 814.200 117.900 819.000 ;
        RECT 134.100 818.400 135.300 819.000 ;
        RECT 119.100 813.300 120.900 818.400 ;
        RECT 62.700 809.700 69.000 810.600 ;
        RECT 66.900 807.600 69.000 809.700 ;
        RECT 62.400 805.050 64.200 806.850 ;
        RECT 67.200 805.800 69.000 807.600 ;
        RECT 69.900 808.800 72.900 810.900 ;
        RECT 74.100 810.300 76.200 811.500 ;
        RECT 98.100 810.300 99.300 812.400 ;
        RECT 113.100 811.950 120.900 813.300 ;
        RECT 122.100 812.400 123.900 818.400 ;
        RECT 134.100 815.400 135.900 818.400 ;
        RECT 137.100 815.400 138.900 818.400 ;
        RECT 122.100 810.300 123.300 812.400 ;
        RECT 137.400 811.200 138.300 815.400 ;
        RECT 140.100 813.000 141.900 819.000 ;
        RECT 143.100 812.400 144.900 818.400 ;
        RECT 158.700 812.400 160.500 819.000 ;
        RECT 163.200 812.400 165.000 818.400 ;
        RECT 167.700 812.400 169.500 819.000 ;
        RECT 185.100 813.300 186.900 818.400 ;
        RECT 188.100 814.200 189.900 819.000 ;
        RECT 191.100 813.300 192.900 818.400 ;
        RECT 137.400 810.300 142.800 811.200 ;
        RECT 95.700 809.400 99.300 810.300 ;
        RECT 119.700 809.400 123.300 810.300 ;
        RECT 140.700 809.400 142.800 810.300 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 62.100 804.300 64.200 805.050 ;
        RECT 62.100 802.950 69.000 804.300 ;
        RECT 17.100 795.600 18.300 802.950 ;
        RECT 23.100 801.150 24.900 802.950 ;
        RECT 41.250 801.150 43.050 802.950 ;
        RECT 19.950 798.450 22.050 799.050 ;
        RECT 25.950 798.450 28.050 799.050 ;
        RECT 31.950 798.450 34.050 799.050 ;
        RECT 43.950 798.450 46.050 799.050 ;
        RECT 19.950 797.550 46.050 798.450 ;
        RECT 19.950 796.950 22.050 797.550 ;
        RECT 25.950 796.950 28.050 797.550 ;
        RECT 31.950 796.950 34.050 797.550 ;
        RECT 43.950 796.950 46.050 797.550 ;
        RECT 47.700 795.600 48.600 802.950 ;
        RECT 67.200 802.500 69.000 802.950 ;
        RECT 69.900 803.100 71.100 808.800 ;
        RECT 72.000 805.800 74.100 807.900 ;
        RECT 72.300 804.000 74.100 805.800 ;
        RECT 92.100 805.050 93.900 806.850 ;
        RECT 95.700 805.050 96.900 809.400 ;
        RECT 98.100 805.050 99.900 806.850 ;
        RECT 116.100 805.050 117.900 806.850 ;
        RECT 119.700 805.050 120.900 809.400 ;
        RECT 122.100 805.050 123.900 806.850 ;
        RECT 134.400 805.050 136.200 806.850 ;
        RECT 69.900 802.200 72.300 803.100 ;
        RECT 70.800 802.050 72.300 802.200 ;
        RECT 76.800 802.950 78.900 805.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 134.100 802.950 136.200 805.050 ;
        RECT 137.400 802.950 139.500 805.050 ;
        RECT 66.000 799.500 69.900 801.300 ;
        RECT 67.800 799.200 69.900 799.500 ;
        RECT 70.800 799.950 72.900 802.050 ;
        RECT 76.800 801.150 78.600 802.950 ;
        RECT 89.100 801.150 90.900 802.950 ;
        RECT 70.800 798.000 71.700 799.950 ;
        RECT 64.500 795.600 66.600 797.700 ;
        RECT 70.200 796.950 71.700 798.000 ;
        RECT 70.200 795.600 71.400 796.950 ;
        RECT 17.100 794.100 19.500 795.600 ;
        RECT 15.000 791.100 16.800 792.900 ;
        RECT 14.700 783.000 16.500 789.600 ;
        RECT 17.700 783.600 19.500 794.100 ;
        RECT 22.800 783.000 24.600 795.600 ;
        RECT 38.100 794.700 45.900 795.600 ;
        RECT 38.100 783.600 39.900 794.700 ;
        RECT 41.100 783.000 42.900 793.800 ;
        RECT 44.100 783.600 45.900 794.700 ;
        RECT 47.100 783.600 48.900 795.600 ;
        RECT 62.100 794.700 66.600 795.600 ;
        RECT 62.100 783.600 63.900 794.700 ;
        RECT 65.100 783.000 66.900 793.500 ;
        RECT 69.600 783.600 71.400 795.600 ;
        RECT 74.100 795.600 76.200 796.500 ;
        RECT 95.700 795.600 96.900 802.950 ;
        RECT 113.100 801.150 114.900 802.950 ;
        RECT 109.950 798.450 112.050 799.050 ;
        RECT 115.950 798.450 118.050 799.050 ;
        RECT 109.950 797.550 118.050 798.450 ;
        RECT 109.950 796.950 112.050 797.550 ;
        RECT 115.950 796.950 118.050 797.550 ;
        RECT 119.700 795.600 120.900 802.950 ;
        RECT 138.000 801.150 139.800 802.950 ;
        RECT 140.700 798.900 141.600 809.400 ;
        RECT 144.000 805.050 144.900 812.400 ;
        RECT 158.250 805.050 160.050 806.850 ;
        RECT 164.100 805.050 165.300 812.400 ;
        RECT 185.100 811.950 192.900 813.300 ;
        RECT 194.100 812.400 195.900 818.400 ;
        RECT 206.100 813.300 207.900 818.400 ;
        RECT 209.100 814.200 210.900 819.000 ;
        RECT 212.100 813.300 213.900 818.400 ;
        RECT 194.100 810.300 195.300 812.400 ;
        RECT 206.100 811.950 213.900 813.300 ;
        RECT 215.100 812.400 216.900 818.400 ;
        RECT 230.100 813.300 231.900 818.400 ;
        RECT 233.100 814.200 234.900 819.000 ;
        RECT 236.100 813.300 237.900 818.400 ;
        RECT 215.100 810.300 216.300 812.400 ;
        RECT 230.100 811.950 237.900 813.300 ;
        RECT 239.100 812.400 240.900 818.400 ;
        RECT 251.100 815.400 252.900 819.000 ;
        RECT 254.100 815.400 255.900 818.400 ;
        RECT 239.100 810.300 240.300 812.400 ;
        RECT 191.700 809.400 195.300 810.300 ;
        RECT 212.700 809.400 216.300 810.300 ;
        RECT 236.700 809.400 240.300 810.300 ;
        RECT 170.100 805.050 171.900 806.850 ;
        RECT 188.100 805.050 189.900 806.850 ;
        RECT 191.700 805.050 192.900 809.400 ;
        RECT 194.100 805.050 195.900 806.850 ;
        RECT 209.100 805.050 210.900 806.850 ;
        RECT 212.700 805.050 213.900 809.400 ;
        RECT 215.100 805.050 216.900 806.850 ;
        RECT 233.100 805.050 234.900 806.850 ;
        RECT 236.700 805.050 237.900 809.400 ;
        RECT 239.100 805.050 240.900 806.850 ;
        RECT 254.100 805.050 255.300 815.400 ;
        RECT 269.100 812.400 270.900 818.400 ;
        RECT 269.700 810.300 270.900 812.400 ;
        RECT 272.100 813.300 273.900 818.400 ;
        RECT 275.100 814.200 276.900 819.000 ;
        RECT 278.100 813.300 279.900 818.400 ;
        RECT 272.100 811.950 279.900 813.300 ;
        RECT 293.400 812.400 295.200 819.000 ;
        RECT 298.500 811.200 300.300 818.400 ;
        RECT 296.100 810.300 300.300 811.200 ;
        RECT 311.700 811.200 313.500 818.400 ;
        RECT 316.800 812.400 318.600 819.000 ;
        RECT 332.100 815.400 333.900 819.000 ;
        RECT 335.100 815.400 336.900 818.400 ;
        RECT 311.700 810.300 315.900 811.200 ;
        RECT 269.700 809.400 273.300 810.300 ;
        RECT 269.100 805.050 270.900 806.850 ;
        RECT 272.100 805.050 273.300 809.400 ;
        RECT 275.100 805.050 276.900 806.850 ;
        RECT 293.250 805.050 295.050 806.850 ;
        RECT 296.100 805.050 297.300 810.300 ;
        RECT 299.100 805.050 300.900 806.850 ;
        RECT 311.100 805.050 312.900 806.850 ;
        RECT 314.700 805.050 315.900 810.300 ;
        RECT 316.950 805.050 318.750 806.850 ;
        RECT 335.100 805.050 336.300 815.400 ;
        RECT 347.100 812.400 348.900 818.400 ;
        RECT 347.700 810.300 348.900 812.400 ;
        RECT 350.100 813.300 351.900 818.400 ;
        RECT 353.100 814.200 354.900 819.000 ;
        RECT 356.100 813.300 357.900 818.400 ;
        RECT 350.100 811.950 357.900 813.300 ;
        RECT 372.000 812.400 373.800 819.000 ;
        RECT 376.500 813.600 378.300 818.400 ;
        RECT 379.500 815.400 381.300 819.000 ;
        RECT 395.100 815.400 396.900 819.000 ;
        RECT 398.100 815.400 399.900 818.400 ;
        RECT 401.100 815.400 402.900 819.000 ;
        RECT 376.500 812.400 381.600 813.600 ;
        RECT 347.700 809.400 351.300 810.300 ;
        RECT 347.100 805.050 348.900 806.850 ;
        RECT 350.100 805.050 351.300 809.400 ;
        RECT 353.100 805.050 354.900 806.850 ;
        RECT 371.100 805.050 372.900 806.850 ;
        RECT 377.250 805.050 379.050 806.850 ;
        RECT 380.700 805.050 381.600 812.400 ;
        RECT 398.700 805.050 399.600 815.400 ;
        RECT 414.000 812.400 415.800 819.000 ;
        RECT 418.500 813.600 420.300 818.400 ;
        RECT 421.500 815.400 423.300 819.000 ;
        RECT 437.100 815.400 438.900 818.400 ;
        RECT 440.100 815.400 441.900 819.000 ;
        RECT 443.700 815.400 445.500 819.000 ;
        RECT 446.700 815.400 448.500 818.400 ;
        RECT 418.500 812.400 423.600 813.600 ;
        RECT 413.100 805.050 414.900 806.850 ;
        RECT 419.250 805.050 421.050 806.850 ;
        RECT 422.700 805.050 423.600 812.400 ;
        RECT 437.700 805.050 438.900 815.400 ;
        RECT 142.800 802.950 144.900 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 166.950 802.950 169.050 805.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 184.950 802.950 187.050 805.050 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 205.950 802.950 208.050 805.050 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 292.950 802.950 295.050 805.050 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 298.950 802.950 301.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 313.950 802.950 316.050 805.050 ;
        RECT 316.950 802.950 319.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 140.100 798.300 141.900 798.900 ;
        RECT 74.100 794.400 78.900 795.600 ;
        RECT 74.100 783.000 75.900 793.500 ;
        RECT 77.100 783.600 78.900 794.400 ;
        RECT 89.400 783.000 91.200 795.600 ;
        RECT 94.500 794.100 96.900 795.600 ;
        RECT 94.500 783.600 96.300 794.100 ;
        RECT 97.200 791.100 99.000 792.900 ;
        RECT 97.500 783.000 99.300 789.600 ;
        RECT 113.400 783.000 115.200 795.600 ;
        RECT 118.500 794.100 120.900 795.600 ;
        RECT 134.100 797.100 141.900 798.300 ;
        RECT 134.100 795.600 135.300 797.100 ;
        RECT 142.800 795.600 144.000 802.950 ;
        RECT 161.250 801.150 163.050 802.950 ;
        RECT 164.100 797.400 165.000 802.950 ;
        RECT 167.100 801.150 168.900 802.950 ;
        RECT 185.100 801.150 186.900 802.950 ;
        RECT 164.100 796.500 168.900 797.400 ;
        RECT 118.500 783.600 120.300 794.100 ;
        RECT 121.200 791.100 123.000 792.900 ;
        RECT 121.500 783.000 123.300 789.600 ;
        RECT 134.100 783.600 135.900 795.600 ;
        RECT 138.600 783.000 140.400 795.600 ;
        RECT 141.600 794.100 144.000 795.600 ;
        RECT 158.100 794.400 165.900 795.300 ;
        RECT 141.600 783.600 143.400 794.100 ;
        RECT 158.100 783.600 159.900 794.400 ;
        RECT 161.100 783.000 162.900 793.500 ;
        RECT 164.100 784.500 165.900 794.400 ;
        RECT 167.100 785.400 168.900 796.500 ;
        RECT 191.700 795.600 192.900 802.950 ;
        RECT 206.100 801.150 207.900 802.950 ;
        RECT 212.700 795.600 213.900 802.950 ;
        RECT 230.100 801.150 231.900 802.950 ;
        RECT 236.700 795.600 237.900 802.950 ;
        RECT 251.100 801.150 252.900 802.950 ;
        RECT 170.100 784.500 171.900 795.600 ;
        RECT 164.100 783.600 171.900 784.500 ;
        RECT 185.400 783.000 187.200 795.600 ;
        RECT 190.500 794.100 192.900 795.600 ;
        RECT 190.500 783.600 192.300 794.100 ;
        RECT 193.200 791.100 195.000 792.900 ;
        RECT 193.500 783.000 195.300 789.600 ;
        RECT 206.400 783.000 208.200 795.600 ;
        RECT 211.500 794.100 213.900 795.600 ;
        RECT 211.500 783.600 213.300 794.100 ;
        RECT 214.200 791.100 216.000 792.900 ;
        RECT 214.500 783.000 216.300 789.600 ;
        RECT 230.400 783.000 232.200 795.600 ;
        RECT 235.500 794.100 237.900 795.600 ;
        RECT 235.500 783.600 237.300 794.100 ;
        RECT 238.200 791.100 240.000 792.900 ;
        RECT 254.100 789.600 255.300 802.950 ;
        RECT 272.100 795.600 273.300 802.950 ;
        RECT 278.100 801.150 279.900 802.950 ;
        RECT 272.100 794.100 274.500 795.600 ;
        RECT 270.000 791.100 271.800 792.900 ;
        RECT 238.500 783.000 240.300 789.600 ;
        RECT 251.100 783.000 252.900 789.600 ;
        RECT 254.100 783.600 255.900 789.600 ;
        RECT 269.700 783.000 271.500 789.600 ;
        RECT 272.700 783.600 274.500 794.100 ;
        RECT 277.800 783.000 279.600 795.600 ;
        RECT 296.100 789.600 297.300 802.950 ;
        RECT 314.700 789.600 315.900 802.950 ;
        RECT 332.100 801.150 333.900 802.950 ;
        RECT 335.100 789.600 336.300 802.950 ;
        RECT 350.100 795.600 351.300 802.950 ;
        RECT 356.100 801.150 357.900 802.950 ;
        RECT 374.250 801.150 376.050 802.950 ;
        RECT 380.700 795.600 381.600 802.950 ;
        RECT 395.100 801.150 396.900 802.950 ;
        RECT 398.700 795.600 399.600 802.950 ;
        RECT 400.950 801.150 402.750 802.950 ;
        RECT 416.250 801.150 418.050 802.950 ;
        RECT 422.700 795.600 423.600 802.950 ;
        RECT 350.100 794.100 352.500 795.600 ;
        RECT 348.000 791.100 349.800 792.900 ;
        RECT 293.100 783.000 294.900 789.600 ;
        RECT 296.100 783.600 297.900 789.600 ;
        RECT 299.100 783.000 300.900 789.600 ;
        RECT 311.100 783.000 312.900 789.600 ;
        RECT 314.100 783.600 315.900 789.600 ;
        RECT 317.100 783.000 318.900 789.600 ;
        RECT 332.100 783.000 333.900 789.600 ;
        RECT 335.100 783.600 336.900 789.600 ;
        RECT 347.700 783.000 349.500 789.600 ;
        RECT 350.700 783.600 352.500 794.100 ;
        RECT 355.800 783.000 357.600 795.600 ;
        RECT 371.100 794.700 378.900 795.600 ;
        RECT 371.100 783.600 372.900 794.700 ;
        RECT 374.100 783.000 375.900 793.800 ;
        RECT 377.100 783.600 378.900 794.700 ;
        RECT 380.100 783.600 381.900 795.600 ;
        RECT 396.000 794.400 399.600 795.600 ;
        RECT 396.000 783.600 397.800 794.400 ;
        RECT 401.100 783.000 402.900 795.600 ;
        RECT 413.100 794.700 420.900 795.600 ;
        RECT 413.100 783.600 414.900 794.700 ;
        RECT 416.100 783.000 417.900 793.800 ;
        RECT 419.100 783.600 420.900 794.700 ;
        RECT 422.100 783.600 423.900 795.600 ;
        RECT 437.700 789.600 438.900 802.950 ;
        RECT 440.100 801.150 441.900 802.950 ;
        RECT 447.000 802.050 448.500 815.400 ;
        RECT 446.100 799.950 448.500 802.050 ;
        RECT 447.000 789.600 448.500 799.950 ;
        RECT 450.300 812.400 452.100 818.400 ;
        RECT 455.700 812.400 457.500 819.000 ;
        RECT 460.800 813.600 462.600 818.400 ;
        RECT 465.000 815.400 466.800 818.400 ;
        RECT 468.000 815.400 469.800 818.400 ;
        RECT 471.000 815.400 472.800 818.400 ;
        RECT 474.000 815.400 475.800 818.400 ;
        RECT 477.000 815.400 478.800 819.000 ;
        RECT 458.400 812.400 462.600 813.600 ;
        RECT 464.700 813.300 466.800 815.400 ;
        RECT 467.700 813.300 469.800 815.400 ;
        RECT 470.700 813.300 472.800 815.400 ;
        RECT 473.700 813.300 475.800 815.400 ;
        RECT 480.000 814.500 481.800 818.400 ;
        RECT 484.500 815.400 486.300 819.000 ;
        RECT 487.500 815.400 489.300 818.400 ;
        RECT 490.500 815.400 492.300 818.400 ;
        RECT 493.500 815.400 495.300 818.400 ;
        RECT 479.100 812.400 481.800 814.500 ;
        RECT 483.600 813.600 485.400 814.500 ;
        RECT 483.600 812.400 486.300 813.600 ;
        RECT 487.200 813.300 489.300 815.400 ;
        RECT 490.200 813.300 492.300 815.400 ;
        RECT 493.200 813.300 495.300 815.400 ;
        RECT 497.700 812.400 499.500 818.400 ;
        RECT 503.100 812.400 504.900 819.000 ;
        RECT 508.500 812.400 510.300 818.400 ;
        RECT 450.300 795.600 451.200 812.400 ;
        RECT 458.400 809.100 459.900 812.400 ;
        RECT 464.100 810.600 470.700 812.400 ;
        RECT 485.400 811.800 486.300 812.400 ;
        RECT 488.400 811.800 490.200 812.400 ;
        RECT 485.400 810.600 492.600 811.800 ;
        RECT 452.100 807.300 459.900 809.100 ;
        RECT 476.100 808.500 477.900 810.300 ;
        RECT 475.800 807.900 477.900 808.500 ;
        RECT 460.800 806.400 477.900 807.900 ;
        RECT 482.100 807.900 484.200 808.050 ;
        RECT 485.400 807.900 487.200 808.800 ;
        RECT 482.100 807.000 487.200 807.900 ;
        RECT 491.700 807.600 492.600 810.600 ;
        RECT 497.700 811.500 499.200 812.400 ;
        RECT 497.700 810.300 506.100 811.500 ;
        RECT 504.300 809.700 506.100 810.300 ;
        RECT 493.500 808.800 495.600 809.700 ;
        RECT 509.100 808.800 510.300 812.400 ;
        RECT 524.100 813.300 525.900 818.400 ;
        RECT 527.100 814.200 528.900 819.000 ;
        RECT 530.100 813.300 531.900 818.400 ;
        RECT 524.100 811.950 531.900 813.300 ;
        RECT 533.100 812.400 534.900 818.400 ;
        RECT 545.400 812.400 547.200 819.000 ;
        RECT 533.100 810.300 534.300 812.400 ;
        RECT 550.500 811.200 552.300 818.400 ;
        RECT 493.500 807.600 510.300 808.800 ;
        RECT 530.700 809.400 534.300 810.300 ;
        RECT 548.100 810.300 552.300 811.200 ;
        RECT 563.700 811.200 565.500 818.400 ;
        RECT 568.800 812.400 570.600 819.000 ;
        RECT 584.100 815.400 585.900 818.400 ;
        RECT 584.100 811.500 585.300 815.400 ;
        RECT 587.100 812.400 588.900 819.000 ;
        RECT 590.100 812.400 591.900 818.400 ;
        RECT 563.700 810.300 567.900 811.200 ;
        RECT 584.100 810.600 589.800 811.500 ;
        RECT 455.700 804.900 462.300 806.400 ;
        RECT 482.100 805.950 484.200 807.000 ;
        RECT 490.800 805.800 492.600 807.600 ;
        RECT 455.700 802.050 457.200 804.900 ;
        RECT 463.500 803.700 507.900 804.900 ;
        RECT 463.500 802.200 464.400 803.700 ;
        RECT 455.100 799.950 457.200 802.050 ;
        RECT 459.300 800.400 464.400 802.200 ;
        RECT 467.100 801.900 480.600 802.800 ;
        RECT 487.800 801.900 489.600 802.500 ;
        RECT 506.100 802.050 507.900 803.700 ;
        RECT 467.100 800.700 468.000 801.900 ;
        RECT 467.100 798.900 468.900 800.700 ;
        RECT 473.100 799.200 477.000 801.000 ;
        RECT 478.500 800.700 489.600 801.900 ;
        RECT 500.100 801.750 502.200 802.050 ;
        RECT 478.500 799.800 480.600 800.700 ;
        RECT 498.300 799.950 502.200 801.750 ;
        RECT 506.100 799.950 508.200 802.050 ;
        RECT 498.300 799.200 500.100 799.950 ;
        RECT 473.100 798.900 475.200 799.200 ;
        RECT 486.600 798.300 500.100 799.200 ;
        RECT 452.100 797.700 453.900 798.300 ;
        RECT 486.600 797.700 487.800 798.300 ;
        RECT 452.100 796.500 487.800 797.700 ;
        RECT 490.500 796.500 492.600 796.800 ;
        RECT 450.300 794.700 466.800 795.600 ;
        RECT 450.300 791.400 451.200 794.700 ;
        RECT 455.100 792.600 460.800 793.800 ;
        RECT 464.700 793.500 466.800 794.700 ;
        RECT 470.100 794.400 487.800 795.600 ;
        RECT 490.500 795.300 502.500 796.500 ;
        RECT 490.500 794.700 492.600 795.300 ;
        RECT 500.700 794.700 502.500 795.300 ;
        RECT 470.100 793.500 472.200 794.400 ;
        RECT 486.600 793.800 487.800 794.400 ;
        RECT 504.000 793.800 505.800 794.100 ;
        RECT 455.100 792.000 456.900 792.600 ;
        RECT 450.300 790.500 454.200 791.400 ;
        RECT 453.000 789.600 454.200 790.500 ;
        RECT 459.600 789.600 460.800 792.600 ;
        RECT 461.700 791.700 463.500 792.300 ;
        RECT 461.700 790.500 469.800 791.700 ;
        RECT 467.700 789.600 469.800 790.500 ;
        RECT 473.100 789.600 475.800 793.500 ;
        RECT 478.500 791.100 481.800 793.200 ;
        RECT 486.600 792.600 505.800 793.800 ;
        RECT 437.100 783.600 438.900 789.600 ;
        RECT 440.100 783.000 441.900 789.600 ;
        RECT 443.700 783.000 445.500 789.600 ;
        RECT 446.700 783.600 448.500 789.600 ;
        RECT 450.000 783.000 451.800 789.600 ;
        RECT 453.000 783.600 454.800 789.600 ;
        RECT 456.000 783.000 457.800 789.600 ;
        RECT 459.000 783.600 460.800 789.600 ;
        RECT 462.000 783.000 463.800 789.600 ;
        RECT 464.700 786.600 466.800 788.700 ;
        RECT 467.700 786.600 469.800 788.700 ;
        RECT 470.700 786.600 472.800 788.700 ;
        RECT 465.000 783.600 466.800 786.600 ;
        RECT 468.000 783.600 469.800 786.600 ;
        RECT 471.000 783.600 472.800 786.600 ;
        RECT 474.000 783.600 475.800 789.600 ;
        RECT 477.000 783.000 478.800 789.600 ;
        RECT 480.000 783.600 481.800 791.100 ;
        RECT 487.200 789.600 489.300 791.700 ;
        RECT 483.900 783.000 485.700 789.600 ;
        RECT 486.900 783.600 488.700 789.600 ;
        RECT 489.600 786.600 491.700 788.700 ;
        RECT 492.600 786.600 494.700 788.700 ;
        RECT 489.900 783.600 491.700 786.600 ;
        RECT 492.900 783.600 494.700 786.600 ;
        RECT 496.500 783.000 498.300 789.600 ;
        RECT 499.500 783.600 501.300 792.600 ;
        RECT 504.000 792.300 505.800 792.600 ;
        RECT 509.100 791.400 510.300 807.600 ;
        RECT 519.000 807.450 523.050 808.050 ;
        RECT 518.550 805.950 523.050 807.450 ;
        RECT 518.550 802.050 519.450 805.950 ;
        RECT 527.100 805.050 528.900 806.850 ;
        RECT 530.700 805.050 531.900 809.400 ;
        RECT 535.950 807.450 540.000 808.050 ;
        RECT 533.100 805.050 534.900 806.850 ;
        RECT 535.950 805.950 540.450 807.450 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 529.950 802.950 532.050 805.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 518.550 800.550 523.050 802.050 ;
        RECT 524.100 801.150 525.900 802.950 ;
        RECT 519.000 799.950 523.050 800.550 ;
        RECT 511.950 798.450 514.050 799.050 ;
        RECT 526.950 798.450 529.050 798.750 ;
        RECT 511.950 797.550 529.050 798.450 ;
        RECT 511.950 796.950 514.050 797.550 ;
        RECT 526.950 796.650 529.050 797.550 ;
        RECT 530.700 795.600 531.900 802.950 ;
        RECT 539.550 798.900 540.450 805.950 ;
        RECT 545.250 805.050 547.050 806.850 ;
        RECT 548.100 805.050 549.300 810.300 ;
        RECT 551.100 805.050 552.900 806.850 ;
        RECT 563.100 805.050 564.900 806.850 ;
        RECT 566.700 805.050 567.900 810.300 ;
        RECT 588.000 809.700 589.800 810.600 ;
        RECT 571.950 807.450 576.000 808.050 ;
        RECT 568.950 805.050 570.750 806.850 ;
        RECT 571.950 805.950 576.450 807.450 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 568.950 802.950 571.050 805.050 ;
        RECT 538.950 796.800 541.050 798.900 ;
        RECT 506.700 790.500 510.300 791.400 ;
        RECT 506.700 789.600 507.600 790.500 ;
        RECT 502.500 783.000 504.300 789.600 ;
        RECT 505.500 788.700 507.600 789.600 ;
        RECT 505.500 783.600 507.300 788.700 ;
        RECT 508.500 783.000 510.300 789.600 ;
        RECT 524.400 783.000 526.200 795.600 ;
        RECT 529.500 794.100 531.900 795.600 ;
        RECT 529.500 783.600 531.300 794.100 ;
        RECT 532.200 791.100 534.000 792.900 ;
        RECT 548.100 789.600 549.300 802.950 ;
        RECT 566.700 789.600 567.900 802.950 ;
        RECT 575.550 799.050 576.450 805.950 ;
        RECT 584.400 802.950 586.500 805.050 ;
        RECT 584.400 801.150 586.200 802.950 ;
        RECT 575.550 798.900 579.000 799.050 ;
        RECT 575.550 797.550 580.050 798.900 ;
        RECT 576.000 796.950 580.050 797.550 ;
        RECT 588.000 798.300 588.900 809.700 ;
        RECT 590.700 805.050 591.900 812.400 ;
        RECT 589.800 802.950 591.900 805.050 ;
        RECT 588.000 797.400 589.800 798.300 ;
        RECT 577.950 796.800 580.050 796.950 ;
        RECT 584.100 796.500 589.800 797.400 ;
        RECT 584.100 789.600 585.300 796.500 ;
        RECT 590.700 795.600 591.900 802.950 ;
        RECT 532.500 783.000 534.300 789.600 ;
        RECT 545.100 783.000 546.900 789.600 ;
        RECT 548.100 783.600 549.900 789.600 ;
        RECT 551.100 783.000 552.900 789.600 ;
        RECT 563.100 783.000 564.900 789.600 ;
        RECT 566.100 783.600 567.900 789.600 ;
        RECT 569.100 783.000 570.900 789.600 ;
        RECT 584.100 783.600 585.900 789.600 ;
        RECT 587.100 783.000 588.900 793.800 ;
        RECT 590.100 783.600 591.900 795.600 ;
        RECT 602.100 812.400 603.900 818.400 ;
        RECT 605.100 812.400 606.900 819.000 ;
        RECT 608.100 815.400 609.900 818.400 ;
        RECT 623.700 815.400 625.500 819.000 ;
        RECT 602.100 805.050 603.300 812.400 ;
        RECT 608.700 811.500 609.900 815.400 ;
        RECT 626.700 813.600 628.500 818.400 ;
        RECT 604.200 810.600 609.900 811.500 ;
        RECT 623.400 812.400 628.500 813.600 ;
        RECT 631.200 812.400 633.000 819.000 ;
        RECT 647.400 812.400 649.200 819.000 ;
        RECT 604.200 809.700 606.000 810.600 ;
        RECT 602.100 802.950 604.200 805.050 ;
        RECT 602.100 795.600 603.300 802.950 ;
        RECT 605.100 798.300 606.000 809.700 ;
        RECT 623.400 805.050 624.300 812.400 ;
        RECT 652.500 811.200 654.300 818.400 ;
        RECT 667.500 812.400 669.300 819.000 ;
        RECT 672.000 812.400 673.800 818.400 ;
        RECT 676.500 812.400 678.300 819.000 ;
        RECT 689.100 815.400 690.900 818.400 ;
        RECT 692.100 815.400 693.900 819.000 ;
        RECT 650.100 810.300 654.300 811.200 ;
        RECT 625.950 805.050 627.750 806.850 ;
        RECT 632.100 805.050 633.900 806.850 ;
        RECT 647.250 805.050 649.050 806.850 ;
        RECT 650.100 805.050 651.300 810.300 ;
        RECT 655.950 807.450 658.050 811.050 ;
        RECT 661.950 807.450 664.050 808.050 ;
        RECT 655.950 807.000 664.050 807.450 ;
        RECT 653.100 805.050 654.900 806.850 ;
        RECT 656.550 806.550 664.050 807.000 ;
        RECT 661.950 805.950 664.050 806.550 ;
        RECT 665.100 805.050 666.900 806.850 ;
        RECT 671.700 805.050 672.900 812.400 ;
        RECT 676.950 805.050 678.750 806.850 ;
        RECT 689.700 805.050 690.900 815.400 ;
        RECT 704.100 812.400 705.900 819.000 ;
        RECT 707.100 812.400 708.900 818.400 ;
        RECT 710.100 812.400 711.900 819.000 ;
        RECT 722.100 812.400 723.900 819.000 ;
        RECT 704.400 805.050 706.200 806.850 ;
        RECT 707.400 805.050 708.450 812.400 ;
        RECT 725.100 811.500 726.900 818.400 ;
        RECT 728.100 812.400 729.900 819.000 ;
        RECT 731.100 811.500 732.900 818.400 ;
        RECT 734.100 812.400 735.900 819.000 ;
        RECT 737.100 811.500 738.900 818.400 ;
        RECT 740.100 812.400 741.900 819.000 ;
        RECT 743.100 811.500 744.900 818.400 ;
        RECT 746.100 812.400 747.900 819.000 ;
        RECT 758.100 815.400 759.900 819.000 ;
        RECT 761.100 815.400 762.900 818.400 ;
        RECT 764.700 815.400 766.500 819.000 ;
        RECT 767.700 815.400 769.500 818.400 ;
        RECT 725.100 810.300 729.000 811.500 ;
        RECT 731.100 810.300 735.000 811.500 ;
        RECT 737.100 810.300 741.000 811.500 ;
        RECT 743.100 810.300 745.950 811.500 ;
        RECT 727.800 809.400 729.000 810.300 ;
        RECT 733.800 809.400 735.000 810.300 ;
        RECT 739.800 809.400 741.000 810.300 ;
        RECT 727.800 808.200 732.000 809.400 ;
        RECT 724.800 805.050 726.600 806.850 ;
        RECT 607.500 802.950 609.600 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 704.400 802.950 706.500 805.050 ;
        RECT 707.400 802.950 711.600 805.050 ;
        RECT 724.800 802.950 726.900 805.050 ;
        RECT 607.800 801.150 609.600 802.950 ;
        RECT 604.200 797.400 606.000 798.300 ;
        RECT 604.200 796.500 609.900 797.400 ;
        RECT 602.100 783.600 603.900 795.600 ;
        RECT 605.100 783.000 606.900 793.800 ;
        RECT 608.700 789.600 609.900 796.500 ;
        RECT 623.400 795.600 624.300 802.950 ;
        RECT 628.950 801.150 630.750 802.950 ;
        RECT 608.100 783.600 609.900 789.600 ;
        RECT 623.100 783.600 624.900 795.600 ;
        RECT 626.100 794.700 633.900 795.600 ;
        RECT 626.100 783.600 627.900 794.700 ;
        RECT 629.100 783.000 630.900 793.800 ;
        RECT 632.100 783.600 633.900 794.700 ;
        RECT 650.100 789.600 651.300 802.950 ;
        RECT 668.100 801.150 669.900 802.950 ;
        RECT 672.000 797.400 672.900 802.950 ;
        RECT 673.950 801.150 675.750 802.950 ;
        RECT 668.100 796.500 672.900 797.400 ;
        RECT 647.100 783.000 648.900 789.600 ;
        RECT 650.100 783.600 651.900 789.600 ;
        RECT 653.100 783.000 654.900 789.600 ;
        RECT 665.100 784.500 666.900 795.600 ;
        RECT 668.100 785.400 669.900 796.500 ;
        RECT 671.100 794.400 678.900 795.300 ;
        RECT 671.100 784.500 672.900 794.400 ;
        RECT 665.100 783.600 672.900 784.500 ;
        RECT 674.100 783.000 675.900 793.500 ;
        RECT 677.100 783.600 678.900 794.400 ;
        RECT 689.700 789.600 690.900 802.950 ;
        RECT 692.100 801.150 693.900 802.950 ;
        RECT 707.400 795.600 708.450 802.950 ;
        RECT 727.800 797.700 729.000 808.200 ;
        RECT 730.200 807.600 732.000 808.200 ;
        RECT 733.800 808.200 738.000 809.400 ;
        RECT 733.800 797.700 735.000 808.200 ;
        RECT 736.200 807.600 738.000 808.200 ;
        RECT 739.800 808.200 744.000 809.400 ;
        RECT 739.800 797.700 741.000 808.200 ;
        RECT 742.200 807.600 744.000 808.200 ;
        RECT 744.900 805.050 745.950 810.300 ;
        RECT 761.100 805.050 762.300 815.400 ;
        RECT 742.800 802.950 745.950 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 744.900 797.700 745.950 802.950 ;
        RECT 758.100 801.150 759.900 802.950 ;
        RECT 725.100 796.500 729.000 797.700 ;
        RECT 731.100 796.500 735.000 797.700 ;
        RECT 737.100 796.500 741.000 797.700 ;
        RECT 743.100 796.500 745.950 797.700 ;
        RECT 689.100 783.600 690.900 789.600 ;
        RECT 692.100 783.000 693.900 789.600 ;
        RECT 704.100 783.000 705.900 795.600 ;
        RECT 707.100 783.600 708.900 795.600 ;
        RECT 710.100 783.000 711.900 795.600 ;
        RECT 722.100 783.000 723.900 795.600 ;
        RECT 725.100 783.600 726.900 796.500 ;
        RECT 728.100 783.000 729.900 795.600 ;
        RECT 731.100 783.600 732.900 796.500 ;
        RECT 734.100 783.000 735.900 795.600 ;
        RECT 737.100 783.600 738.900 796.500 ;
        RECT 740.100 783.000 741.900 795.600 ;
        RECT 743.100 783.600 744.900 796.500 ;
        RECT 746.100 783.000 747.900 795.600 ;
        RECT 761.100 789.600 762.300 802.950 ;
        RECT 768.000 802.050 769.500 815.400 ;
        RECT 767.100 799.950 769.500 802.050 ;
        RECT 768.000 789.600 769.500 799.950 ;
        RECT 771.300 812.400 773.100 818.400 ;
        RECT 776.700 812.400 778.500 819.000 ;
        RECT 781.800 813.600 783.600 818.400 ;
        RECT 786.000 815.400 787.800 818.400 ;
        RECT 789.000 815.400 790.800 818.400 ;
        RECT 792.000 815.400 793.800 818.400 ;
        RECT 795.000 815.400 796.800 818.400 ;
        RECT 798.000 815.400 799.800 819.000 ;
        RECT 779.400 812.400 783.600 813.600 ;
        RECT 785.700 813.300 787.800 815.400 ;
        RECT 788.700 813.300 790.800 815.400 ;
        RECT 791.700 813.300 793.800 815.400 ;
        RECT 794.700 813.300 796.800 815.400 ;
        RECT 801.000 814.500 802.800 818.400 ;
        RECT 805.500 815.400 807.300 819.000 ;
        RECT 808.500 815.400 810.300 818.400 ;
        RECT 811.500 815.400 813.300 818.400 ;
        RECT 814.500 815.400 816.300 818.400 ;
        RECT 800.100 812.400 802.800 814.500 ;
        RECT 804.600 813.600 806.400 814.500 ;
        RECT 804.600 812.400 807.300 813.600 ;
        RECT 808.200 813.300 810.300 815.400 ;
        RECT 811.200 813.300 813.300 815.400 ;
        RECT 814.200 813.300 816.300 815.400 ;
        RECT 818.700 812.400 820.500 818.400 ;
        RECT 824.100 812.400 825.900 819.000 ;
        RECT 829.500 812.400 831.300 818.400 ;
        RECT 771.300 795.600 772.200 812.400 ;
        RECT 779.400 809.100 780.900 812.400 ;
        RECT 785.100 810.600 791.700 812.400 ;
        RECT 806.400 811.800 807.300 812.400 ;
        RECT 809.400 811.800 811.200 812.400 ;
        RECT 806.400 810.600 813.600 811.800 ;
        RECT 773.100 807.300 780.900 809.100 ;
        RECT 797.100 808.500 798.900 810.300 ;
        RECT 796.800 807.900 798.900 808.500 ;
        RECT 781.800 806.400 798.900 807.900 ;
        RECT 803.100 807.900 805.200 808.050 ;
        RECT 806.400 807.900 808.200 808.800 ;
        RECT 803.100 807.000 808.200 807.900 ;
        RECT 812.700 807.600 813.600 810.600 ;
        RECT 818.700 811.500 820.200 812.400 ;
        RECT 818.700 810.300 827.100 811.500 ;
        RECT 825.300 809.700 827.100 810.300 ;
        RECT 814.500 808.800 816.600 809.700 ;
        RECT 830.100 808.800 831.300 812.400 ;
        RECT 814.500 807.600 831.300 808.800 ;
        RECT 776.700 804.900 783.300 806.400 ;
        RECT 803.100 805.950 805.200 807.000 ;
        RECT 811.800 805.800 813.600 807.600 ;
        RECT 776.700 802.050 778.200 804.900 ;
        RECT 784.500 803.700 828.900 804.900 ;
        RECT 784.500 802.200 785.400 803.700 ;
        RECT 776.100 799.950 778.200 802.050 ;
        RECT 780.300 800.400 785.400 802.200 ;
        RECT 788.100 801.900 801.600 802.800 ;
        RECT 808.800 801.900 810.600 802.500 ;
        RECT 827.100 802.050 828.900 803.700 ;
        RECT 788.100 800.700 789.000 801.900 ;
        RECT 788.100 798.900 789.900 800.700 ;
        RECT 794.100 799.200 798.000 801.000 ;
        RECT 799.500 800.700 810.600 801.900 ;
        RECT 821.100 801.750 823.200 802.050 ;
        RECT 799.500 799.800 801.600 800.700 ;
        RECT 819.300 799.950 823.200 801.750 ;
        RECT 827.100 799.950 829.200 802.050 ;
        RECT 819.300 799.200 821.100 799.950 ;
        RECT 794.100 798.900 796.200 799.200 ;
        RECT 807.600 798.300 821.100 799.200 ;
        RECT 773.100 797.700 774.900 798.300 ;
        RECT 807.600 797.700 808.800 798.300 ;
        RECT 773.100 796.500 808.800 797.700 ;
        RECT 811.500 796.500 813.600 796.800 ;
        RECT 771.300 794.700 787.800 795.600 ;
        RECT 771.300 791.400 772.200 794.700 ;
        RECT 776.100 792.600 781.800 793.800 ;
        RECT 785.700 793.500 787.800 794.700 ;
        RECT 791.100 794.400 808.800 795.600 ;
        RECT 811.500 795.300 823.500 796.500 ;
        RECT 811.500 794.700 813.600 795.300 ;
        RECT 821.700 794.700 823.500 795.300 ;
        RECT 791.100 793.500 793.200 794.400 ;
        RECT 807.600 793.800 808.800 794.400 ;
        RECT 825.000 793.800 826.800 794.100 ;
        RECT 776.100 792.000 777.900 792.600 ;
        RECT 771.300 790.500 775.200 791.400 ;
        RECT 774.000 789.600 775.200 790.500 ;
        RECT 780.600 789.600 781.800 792.600 ;
        RECT 782.700 791.700 784.500 792.300 ;
        RECT 782.700 790.500 790.800 791.700 ;
        RECT 788.700 789.600 790.800 790.500 ;
        RECT 794.100 789.600 796.800 793.500 ;
        RECT 799.500 791.100 802.800 793.200 ;
        RECT 807.600 792.600 826.800 793.800 ;
        RECT 758.100 783.000 759.900 789.600 ;
        RECT 761.100 783.600 762.900 789.600 ;
        RECT 764.700 783.000 766.500 789.600 ;
        RECT 767.700 783.600 769.500 789.600 ;
        RECT 771.000 783.000 772.800 789.600 ;
        RECT 774.000 783.600 775.800 789.600 ;
        RECT 777.000 783.000 778.800 789.600 ;
        RECT 780.000 783.600 781.800 789.600 ;
        RECT 783.000 783.000 784.800 789.600 ;
        RECT 785.700 786.600 787.800 788.700 ;
        RECT 788.700 786.600 790.800 788.700 ;
        RECT 791.700 786.600 793.800 788.700 ;
        RECT 786.000 783.600 787.800 786.600 ;
        RECT 789.000 783.600 790.800 786.600 ;
        RECT 792.000 783.600 793.800 786.600 ;
        RECT 795.000 783.600 796.800 789.600 ;
        RECT 798.000 783.000 799.800 789.600 ;
        RECT 801.000 783.600 802.800 791.100 ;
        RECT 808.200 789.600 810.300 791.700 ;
        RECT 804.900 783.000 806.700 789.600 ;
        RECT 807.900 783.600 809.700 789.600 ;
        RECT 810.600 786.600 812.700 788.700 ;
        RECT 813.600 786.600 815.700 788.700 ;
        RECT 810.900 783.600 812.700 786.600 ;
        RECT 813.900 783.600 815.700 786.600 ;
        RECT 817.500 783.000 819.300 789.600 ;
        RECT 820.500 783.600 822.300 792.600 ;
        RECT 825.000 792.300 826.800 792.600 ;
        RECT 830.100 791.400 831.300 807.600 ;
        RECT 827.700 790.500 831.300 791.400 ;
        RECT 833.700 812.400 835.500 818.400 ;
        RECT 839.100 812.400 840.900 819.000 ;
        RECT 844.500 812.400 846.300 818.400 ;
        RECT 848.700 815.400 850.500 818.400 ;
        RECT 851.700 815.400 853.500 818.400 ;
        RECT 854.700 815.400 856.500 818.400 ;
        RECT 857.700 815.400 859.500 819.000 ;
        RECT 848.700 813.300 850.800 815.400 ;
        RECT 851.700 813.300 853.800 815.400 ;
        RECT 854.700 813.300 856.800 815.400 ;
        RECT 862.200 814.500 864.000 818.400 ;
        RECT 865.200 815.400 867.000 819.000 ;
        RECT 868.200 815.400 870.000 818.400 ;
        RECT 871.200 815.400 873.000 818.400 ;
        RECT 874.200 815.400 876.000 818.400 ;
        RECT 877.200 815.400 879.000 818.400 ;
        RECT 858.600 813.600 860.400 814.500 ;
        RECT 857.700 812.400 860.400 813.600 ;
        RECT 862.200 812.400 864.900 814.500 ;
        RECT 868.200 813.300 870.300 815.400 ;
        RECT 871.200 813.300 873.300 815.400 ;
        RECT 874.200 813.300 876.300 815.400 ;
        RECT 877.200 813.300 879.300 815.400 ;
        RECT 881.400 813.600 883.200 818.400 ;
        RECT 881.400 812.400 885.600 813.600 ;
        RECT 886.500 812.400 888.300 819.000 ;
        RECT 891.900 812.400 893.700 818.400 ;
        RECT 833.700 808.800 834.900 812.400 ;
        RECT 844.800 811.500 846.300 812.400 ;
        RECT 853.800 811.800 855.600 812.400 ;
        RECT 857.700 811.800 858.600 812.400 ;
        RECT 837.900 810.300 846.300 811.500 ;
        RECT 851.400 810.600 858.600 811.800 ;
        RECT 873.300 810.600 879.900 812.400 ;
        RECT 837.900 809.700 839.700 810.300 ;
        RECT 848.400 808.800 850.500 809.700 ;
        RECT 833.700 807.600 850.500 808.800 ;
        RECT 851.400 807.600 852.300 810.600 ;
        RECT 856.800 807.900 858.600 808.800 ;
        RECT 866.100 808.500 867.900 810.300 ;
        RECT 884.100 809.100 885.600 812.400 ;
        RECT 859.800 807.900 861.900 808.050 ;
        RECT 833.700 791.400 834.900 807.600 ;
        RECT 851.400 805.800 853.200 807.600 ;
        RECT 856.800 807.000 861.900 807.900 ;
        RECT 859.800 805.950 861.900 807.000 ;
        RECT 866.100 807.900 868.200 808.500 ;
        RECT 866.100 806.400 883.200 807.900 ;
        RECT 884.100 807.300 891.900 809.100 ;
        RECT 881.700 804.900 888.300 806.400 ;
        RECT 836.100 803.700 880.500 804.900 ;
        RECT 836.100 802.050 837.900 803.700 ;
        RECT 835.800 799.950 837.900 802.050 ;
        RECT 841.800 801.750 843.900 802.050 ;
        RECT 854.400 801.900 856.200 802.500 ;
        RECT 863.400 801.900 876.900 802.800 ;
        RECT 841.800 799.950 845.700 801.750 ;
        RECT 854.400 800.700 865.500 801.900 ;
        RECT 843.900 799.200 845.700 799.950 ;
        RECT 863.400 799.800 865.500 800.700 ;
        RECT 867.000 799.200 870.900 801.000 ;
        RECT 876.000 800.700 876.900 801.900 ;
        RECT 843.900 798.300 857.400 799.200 ;
        RECT 868.800 798.900 870.900 799.200 ;
        RECT 875.100 798.900 876.900 800.700 ;
        RECT 879.600 802.200 880.500 803.700 ;
        RECT 879.600 800.400 884.700 802.200 ;
        RECT 886.800 802.050 888.300 804.900 ;
        RECT 886.800 799.950 888.900 802.050 ;
        RECT 856.200 797.700 857.400 798.300 ;
        RECT 890.100 797.700 891.900 798.300 ;
        RECT 851.400 796.500 853.500 796.800 ;
        RECT 856.200 796.500 891.900 797.700 ;
        RECT 841.500 795.300 853.500 796.500 ;
        RECT 892.800 795.600 893.700 812.400 ;
        RECT 841.500 794.700 843.300 795.300 ;
        RECT 851.400 794.700 853.500 795.300 ;
        RECT 856.200 794.400 873.900 795.600 ;
        RECT 838.200 793.800 840.000 794.100 ;
        RECT 856.200 793.800 857.400 794.400 ;
        RECT 838.200 792.600 857.400 793.800 ;
        RECT 871.800 793.500 873.900 794.400 ;
        RECT 877.200 794.700 893.700 795.600 ;
        RECT 877.200 793.500 879.300 794.700 ;
        RECT 838.200 792.300 840.000 792.600 ;
        RECT 833.700 790.500 837.300 791.400 ;
        RECT 827.700 789.600 828.600 790.500 ;
        RECT 836.400 789.600 837.300 790.500 ;
        RECT 823.500 783.000 825.300 789.600 ;
        RECT 826.500 788.700 828.600 789.600 ;
        RECT 826.500 783.600 828.300 788.700 ;
        RECT 829.500 783.000 831.300 789.600 ;
        RECT 833.700 783.000 835.500 789.600 ;
        RECT 836.400 788.700 838.500 789.600 ;
        RECT 836.700 783.600 838.500 788.700 ;
        RECT 839.700 783.000 841.500 789.600 ;
        RECT 842.700 783.600 844.500 792.600 ;
        RECT 854.700 789.600 856.800 791.700 ;
        RECT 862.200 791.100 865.500 793.200 ;
        RECT 845.700 783.000 847.500 789.600 ;
        RECT 849.300 786.600 851.400 788.700 ;
        RECT 852.300 786.600 854.400 788.700 ;
        RECT 849.300 783.600 851.100 786.600 ;
        RECT 852.300 783.600 854.100 786.600 ;
        RECT 855.300 783.600 857.100 789.600 ;
        RECT 858.300 783.000 860.100 789.600 ;
        RECT 862.200 783.600 864.000 791.100 ;
        RECT 868.200 789.600 870.900 793.500 ;
        RECT 883.200 792.600 888.900 793.800 ;
        RECT 880.500 791.700 882.300 792.300 ;
        RECT 874.200 790.500 882.300 791.700 ;
        RECT 874.200 789.600 876.300 790.500 ;
        RECT 883.200 789.600 884.400 792.600 ;
        RECT 887.100 792.000 888.900 792.600 ;
        RECT 892.800 791.400 893.700 794.700 ;
        RECT 889.800 790.500 893.700 791.400 ;
        RECT 895.500 815.400 897.300 818.400 ;
        RECT 898.500 815.400 900.300 819.000 ;
        RECT 914.100 815.400 915.900 819.000 ;
        RECT 917.100 815.400 918.900 818.400 ;
        RECT 929.100 815.400 930.900 818.400 ;
        RECT 895.500 802.050 897.000 815.400 ;
        RECT 917.100 805.050 918.300 815.400 ;
        RECT 929.100 811.500 930.300 815.400 ;
        RECT 932.100 812.400 933.900 819.000 ;
        RECT 935.100 812.400 936.900 818.400 ;
        RECT 929.100 810.600 934.800 811.500 ;
        RECT 933.000 809.700 934.800 810.600 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 929.400 802.950 931.500 805.050 ;
        RECT 895.500 799.950 897.900 802.050 ;
        RECT 914.100 801.150 915.900 802.950 ;
        RECT 889.800 789.600 891.000 790.500 ;
        RECT 895.500 789.600 897.000 799.950 ;
        RECT 917.100 789.600 918.300 802.950 ;
        RECT 929.400 801.150 931.200 802.950 ;
        RECT 933.000 798.300 933.900 809.700 ;
        RECT 935.700 805.050 936.900 812.400 ;
        RECT 934.800 802.950 936.900 805.050 ;
        RECT 933.000 797.400 934.800 798.300 ;
        RECT 929.100 796.500 934.800 797.400 ;
        RECT 929.100 789.600 930.300 796.500 ;
        RECT 935.700 795.600 936.900 802.950 ;
        RECT 865.200 783.000 867.000 789.600 ;
        RECT 868.200 783.600 870.000 789.600 ;
        RECT 871.200 786.600 873.300 788.700 ;
        RECT 874.200 786.600 876.300 788.700 ;
        RECT 877.200 786.600 879.300 788.700 ;
        RECT 871.200 783.600 873.000 786.600 ;
        RECT 874.200 783.600 876.000 786.600 ;
        RECT 877.200 783.600 879.000 786.600 ;
        RECT 880.200 783.000 882.000 789.600 ;
        RECT 883.200 783.600 885.000 789.600 ;
        RECT 886.200 783.000 888.000 789.600 ;
        RECT 889.200 783.600 891.000 789.600 ;
        RECT 892.200 783.000 894.000 789.600 ;
        RECT 895.500 783.600 897.300 789.600 ;
        RECT 898.500 783.000 900.300 789.600 ;
        RECT 914.100 783.000 915.900 789.600 ;
        RECT 917.100 783.600 918.900 789.600 ;
        RECT 929.100 783.600 930.900 789.600 ;
        RECT 932.100 783.000 933.900 793.800 ;
        RECT 935.100 783.600 936.900 795.600 ;
        RECT 11.100 767.400 12.900 779.400 ;
        RECT 14.100 768.300 15.900 779.400 ;
        RECT 17.100 769.200 18.900 780.000 ;
        RECT 20.100 768.300 21.900 779.400 ;
        RECT 35.100 773.400 36.900 779.400 ;
        RECT 38.100 773.400 39.900 780.000 ;
        RECT 14.100 767.400 21.900 768.300 ;
        RECT 11.400 760.050 12.300 767.400 ;
        RECT 16.950 760.050 18.750 761.850 ;
        RECT 35.700 760.050 36.900 773.400 ;
        RECT 53.400 767.400 55.200 780.000 ;
        RECT 58.500 768.900 60.300 779.400 ;
        RECT 61.500 773.400 63.300 780.000 ;
        RECT 61.200 770.100 63.000 771.900 ;
        RECT 58.500 767.400 60.900 768.900 ;
        RECT 74.100 767.400 75.900 779.400 ;
        RECT 77.100 768.300 78.900 779.400 ;
        RECT 80.100 769.200 81.900 780.000 ;
        RECT 83.100 768.300 84.900 779.400 ;
        RECT 77.100 767.400 84.900 768.300 ;
        RECT 98.100 768.300 99.900 779.400 ;
        RECT 101.100 769.200 102.900 780.000 ;
        RECT 104.100 768.300 105.900 779.400 ;
        RECT 98.100 767.400 105.900 768.300 ;
        RECT 107.100 767.400 108.900 779.400 ;
        RECT 119.700 773.400 121.500 780.000 ;
        RECT 120.000 770.100 121.800 771.900 ;
        RECT 122.700 768.900 124.500 779.400 ;
        RECT 122.100 767.400 124.500 768.900 ;
        RECT 127.800 767.400 129.600 780.000 ;
        RECT 140.400 767.400 142.200 780.000 ;
        RECT 145.500 768.900 147.300 779.400 ;
        RECT 148.500 773.400 150.300 780.000 ;
        RECT 148.200 770.100 150.000 771.900 ;
        RECT 145.500 767.400 147.900 768.900 ;
        RECT 164.100 767.400 165.900 779.400 ;
        RECT 167.100 768.300 168.900 779.400 ;
        RECT 170.100 769.200 171.900 780.000 ;
        RECT 173.100 768.300 174.900 779.400 ;
        RECT 167.100 767.400 174.900 768.300 ;
        RECT 188.400 767.400 190.200 780.000 ;
        RECT 193.500 768.900 195.300 779.400 ;
        RECT 196.500 773.400 198.300 780.000 ;
        RECT 196.200 770.100 198.000 771.900 ;
        RECT 193.500 767.400 195.900 768.900 ;
        RECT 212.400 767.400 214.200 780.000 ;
        RECT 217.500 768.900 219.300 779.400 ;
        RECT 220.500 773.400 222.300 780.000 ;
        RECT 236.700 773.400 238.500 780.000 ;
        RECT 220.200 770.100 222.000 771.900 ;
        RECT 237.000 770.100 238.800 771.900 ;
        RECT 239.700 768.900 241.500 779.400 ;
        RECT 217.500 767.400 219.900 768.900 ;
        RECT 38.100 760.050 39.900 761.850 ;
        RECT 53.100 760.050 54.900 761.850 ;
        RECT 59.700 760.050 60.900 767.400 ;
        RECT 74.400 760.050 75.300 767.400 ;
        RECT 93.000 762.450 97.050 763.050 ;
        RECT 79.950 760.050 81.750 761.850 ;
        RECT 92.550 760.950 97.050 762.450 ;
        RECT 10.950 757.950 13.050 760.050 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 11.400 750.600 12.300 757.950 ;
        RECT 13.950 756.150 15.750 757.950 ;
        RECT 20.100 756.150 21.900 757.950 ;
        RECT 13.950 753.450 16.050 754.050 ;
        RECT 25.950 753.450 28.050 754.050 ;
        RECT 13.950 752.550 28.050 753.450 ;
        RECT 13.950 751.950 16.050 752.550 ;
        RECT 25.950 751.950 28.050 752.550 ;
        RECT 11.400 749.400 16.500 750.600 ;
        RECT 11.700 744.000 13.500 747.600 ;
        RECT 14.700 744.600 16.500 749.400 ;
        RECT 19.200 744.000 21.000 750.600 ;
        RECT 35.700 747.600 36.900 757.950 ;
        RECT 56.100 756.150 57.900 757.950 ;
        RECT 59.700 753.600 60.900 757.950 ;
        RECT 62.100 756.150 63.900 757.950 ;
        RECT 59.700 752.700 63.300 753.600 ;
        RECT 53.100 749.700 60.900 751.050 ;
        RECT 35.100 744.600 36.900 747.600 ;
        RECT 38.100 744.000 39.900 747.600 ;
        RECT 53.100 744.600 54.900 749.700 ;
        RECT 56.100 744.000 57.900 748.800 ;
        RECT 59.100 744.600 60.900 749.700 ;
        RECT 62.100 750.600 63.300 752.700 ;
        RECT 74.400 750.600 75.300 757.950 ;
        RECT 76.950 756.150 78.750 757.950 ;
        RECT 83.100 756.150 84.900 757.950 ;
        RECT 92.550 753.450 93.450 760.950 ;
        RECT 101.250 760.050 103.050 761.850 ;
        RECT 107.700 760.050 108.600 767.400 ;
        RECT 114.000 762.450 118.050 763.050 ;
        RECT 113.550 760.950 118.050 762.450 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 98.100 756.150 99.900 757.950 ;
        RECT 104.250 756.150 106.050 757.950 ;
        RECT 97.950 753.450 100.050 754.050 ;
        RECT 92.550 752.550 100.050 753.450 ;
        RECT 97.950 751.950 100.050 752.550 ;
        RECT 107.700 750.600 108.600 757.950 ;
        RECT 113.550 757.050 114.450 760.950 ;
        RECT 122.100 760.050 123.300 767.400 ;
        RECT 135.000 762.450 139.050 763.050 ;
        RECT 128.100 760.050 129.900 761.850 ;
        RECT 134.550 760.950 139.050 762.450 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 127.950 757.950 130.050 760.050 ;
        RECT 113.550 755.550 118.050 757.050 ;
        RECT 119.100 756.150 120.900 757.950 ;
        RECT 114.000 754.950 118.050 755.550 ;
        RECT 122.100 753.600 123.300 757.950 ;
        RECT 125.100 756.150 126.900 757.950 ;
        RECT 134.550 757.050 135.450 760.950 ;
        RECT 140.100 760.050 141.900 761.850 ;
        RECT 146.700 760.050 147.900 767.400 ;
        RECT 164.400 760.050 165.300 767.400 ;
        RECT 169.950 760.050 171.750 761.850 ;
        RECT 188.100 760.050 189.900 761.850 ;
        RECT 194.700 760.050 195.900 767.400 ;
        RECT 212.100 760.050 213.900 761.850 ;
        RECT 218.700 760.050 219.900 767.400 ;
        RECT 239.100 767.400 241.500 768.900 ;
        RECT 244.800 767.400 246.600 780.000 ;
        RECT 260.100 768.300 261.900 779.400 ;
        RECT 263.100 769.500 264.900 780.000 ;
        RECT 267.600 768.300 269.400 779.400 ;
        RECT 271.800 769.500 273.900 780.000 ;
        RECT 275.100 768.600 276.900 779.400 ;
        RECT 239.100 760.050 240.300 767.400 ;
        RECT 260.100 767.100 264.900 768.300 ;
        RECT 267.600 767.400 270.900 768.300 ;
        RECT 262.800 766.200 264.900 767.100 ;
        RECT 262.800 765.300 268.200 766.200 ;
        RECT 266.400 763.500 268.200 765.300 ;
        RECT 269.700 763.050 270.900 767.400 ;
        RECT 271.800 767.400 276.900 768.600 ;
        RECT 287.100 767.400 288.900 779.400 ;
        RECT 290.100 768.300 291.900 779.400 ;
        RECT 293.100 769.200 294.900 780.000 ;
        RECT 296.100 768.300 297.900 779.400 ;
        RECT 290.100 767.400 297.900 768.300 ;
        RECT 311.100 767.400 312.900 779.400 ;
        RECT 314.100 768.300 315.900 779.400 ;
        RECT 317.100 769.200 318.900 780.000 ;
        RECT 320.100 768.300 321.900 779.400 ;
        RECT 335.100 773.400 336.900 780.000 ;
        RECT 338.100 773.400 339.900 779.400 ;
        RECT 350.100 773.400 351.900 779.400 ;
        RECT 314.100 767.400 321.900 768.300 ;
        RECT 271.800 766.500 273.900 767.400 ;
        RECT 269.100 762.300 271.200 763.050 ;
        RECT 245.100 760.050 246.900 761.850 ;
        RECT 264.900 760.200 266.700 762.000 ;
        RECT 268.200 760.950 271.200 762.300 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 172.950 757.950 175.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 220.950 757.950 223.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 130.950 755.550 135.450 757.050 ;
        RECT 143.100 756.150 144.900 757.950 ;
        RECT 130.950 754.950 135.000 755.550 ;
        RECT 119.700 752.700 123.300 753.600 ;
        RECT 146.700 753.600 147.900 757.950 ;
        RECT 149.100 756.150 150.900 757.950 ;
        RECT 146.700 752.700 150.300 753.600 ;
        RECT 119.700 750.600 120.900 752.700 ;
        RECT 62.100 744.600 63.900 750.600 ;
        RECT 74.400 749.400 79.500 750.600 ;
        RECT 74.700 744.000 76.500 747.600 ;
        RECT 77.700 744.600 79.500 749.400 ;
        RECT 82.200 744.000 84.000 750.600 ;
        RECT 99.000 744.000 100.800 750.600 ;
        RECT 103.500 749.400 108.600 750.600 ;
        RECT 103.500 744.600 105.300 749.400 ;
        RECT 106.500 744.000 108.300 747.600 ;
        RECT 119.100 744.600 120.900 750.600 ;
        RECT 122.100 749.700 129.900 751.050 ;
        RECT 122.100 744.600 123.900 749.700 ;
        RECT 125.100 744.000 126.900 748.800 ;
        RECT 128.100 744.600 129.900 749.700 ;
        RECT 140.100 749.700 147.900 751.050 ;
        RECT 140.100 744.600 141.900 749.700 ;
        RECT 143.100 744.000 144.900 748.800 ;
        RECT 146.100 744.600 147.900 749.700 ;
        RECT 149.100 750.600 150.300 752.700 ;
        RECT 164.400 750.600 165.300 757.950 ;
        RECT 166.950 756.150 168.750 757.950 ;
        RECT 173.100 756.150 174.900 757.950 ;
        RECT 191.100 756.150 192.900 757.950 ;
        RECT 194.700 753.600 195.900 757.950 ;
        RECT 197.100 756.150 198.900 757.950 ;
        RECT 215.100 756.150 216.900 757.950 ;
        RECT 218.700 753.600 219.900 757.950 ;
        RECT 221.100 756.150 222.900 757.950 ;
        RECT 236.100 756.150 237.900 757.950 ;
        RECT 239.100 753.600 240.300 757.950 ;
        RECT 242.100 756.150 243.900 757.950 ;
        RECT 260.100 757.800 262.200 760.050 ;
        RECT 264.900 758.100 267.000 760.200 ;
        RECT 260.400 757.200 262.200 757.800 ;
        RECT 260.400 756.000 267.000 757.200 ;
        RECT 264.900 755.100 267.000 756.000 ;
        RECT 194.700 752.700 198.300 753.600 ;
        RECT 218.700 752.700 222.300 753.600 ;
        RECT 149.100 744.600 150.900 750.600 ;
        RECT 164.400 749.400 169.500 750.600 ;
        RECT 164.700 744.000 166.500 747.600 ;
        RECT 167.700 744.600 169.500 749.400 ;
        RECT 172.200 744.000 174.000 750.600 ;
        RECT 188.100 749.700 195.900 751.050 ;
        RECT 188.100 744.600 189.900 749.700 ;
        RECT 191.100 744.000 192.900 748.800 ;
        RECT 194.100 744.600 195.900 749.700 ;
        RECT 197.100 750.600 198.300 752.700 ;
        RECT 197.100 744.600 198.900 750.600 ;
        RECT 212.100 749.700 219.900 751.050 ;
        RECT 212.100 744.600 213.900 749.700 ;
        RECT 215.100 744.000 216.900 748.800 ;
        RECT 218.100 744.600 219.900 749.700 ;
        RECT 221.100 750.600 222.300 752.700 ;
        RECT 236.700 752.700 240.300 753.600 ;
        RECT 262.500 753.000 264.600 753.600 ;
        RECT 265.500 753.300 267.300 755.100 ;
        RECT 268.200 754.200 269.100 760.950 ;
        RECT 274.800 760.050 276.600 761.850 ;
        RECT 287.400 760.050 288.300 767.400 ;
        RECT 298.950 762.450 303.000 763.050 ;
        RECT 292.950 760.050 294.750 761.850 ;
        RECT 298.950 760.950 303.450 762.450 ;
        RECT 270.000 758.100 271.800 759.900 ;
        RECT 270.000 756.000 272.100 758.100 ;
        RECT 274.800 757.950 276.900 760.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 236.700 750.600 237.900 752.700 ;
        RECT 260.100 751.500 264.600 753.000 ;
        RECT 268.200 752.100 271.200 754.200 ;
        RECT 221.100 744.600 222.900 750.600 ;
        RECT 236.100 744.600 237.900 750.600 ;
        RECT 239.100 749.700 246.900 751.050 ;
        RECT 239.100 744.600 240.900 749.700 ;
        RECT 242.100 744.000 243.900 748.800 ;
        RECT 245.100 744.600 246.900 749.700 ;
        RECT 260.100 750.600 261.600 751.500 ;
        RECT 260.100 744.600 261.900 750.600 ;
        RECT 268.200 750.000 269.100 752.100 ;
        RECT 272.400 751.500 274.500 753.900 ;
        RECT 272.400 750.600 276.900 751.500 ;
        RECT 263.100 744.000 264.900 749.700 ;
        RECT 267.300 744.600 269.100 750.000 ;
        RECT 271.800 744.000 273.600 749.700 ;
        RECT 275.100 744.600 276.900 750.600 ;
        RECT 287.400 750.600 288.300 757.950 ;
        RECT 289.950 756.150 291.750 757.950 ;
        RECT 296.100 756.150 297.900 757.950 ;
        RECT 302.550 756.450 303.450 760.950 ;
        RECT 311.400 760.050 312.300 767.400 ;
        RECT 313.950 765.450 316.050 766.050 ;
        RECT 334.950 765.450 337.050 766.050 ;
        RECT 313.950 764.550 337.050 765.450 ;
        RECT 313.950 763.950 316.050 764.550 ;
        RECT 334.950 763.950 337.050 764.550 ;
        RECT 316.950 760.050 318.750 761.850 ;
        RECT 335.100 760.050 336.900 761.850 ;
        RECT 338.100 760.050 339.300 773.400 ;
        RECT 350.100 766.500 351.300 773.400 ;
        RECT 353.100 769.200 354.900 780.000 ;
        RECT 356.100 767.400 357.900 779.400 ;
        RECT 368.100 767.400 369.900 780.000 ;
        RECT 373.200 768.600 375.000 779.400 ;
        RECT 371.400 767.400 375.000 768.600 ;
        RECT 387.000 768.600 388.800 779.400 ;
        RECT 387.000 767.400 390.600 768.600 ;
        RECT 392.100 767.400 393.900 780.000 ;
        RECT 404.100 773.400 405.900 780.000 ;
        RECT 407.100 773.400 408.900 779.400 ;
        RECT 410.100 773.400 411.900 780.000 ;
        RECT 425.700 773.400 427.500 780.000 ;
        RECT 350.100 765.600 355.800 766.500 ;
        RECT 354.000 764.700 355.800 765.600 ;
        RECT 350.400 760.050 352.200 761.850 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 313.950 757.950 316.050 760.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 350.400 757.950 352.500 760.050 ;
        RECT 307.950 756.450 310.050 757.050 ;
        RECT 302.550 755.550 310.050 756.450 ;
        RECT 307.950 754.950 310.050 755.550 ;
        RECT 311.400 750.600 312.300 757.950 ;
        RECT 313.950 756.150 315.750 757.950 ;
        RECT 320.100 756.150 321.900 757.950 ;
        RECT 287.400 749.400 292.500 750.600 ;
        RECT 287.700 744.000 289.500 747.600 ;
        RECT 290.700 744.600 292.500 749.400 ;
        RECT 295.200 744.000 297.000 750.600 ;
        RECT 311.400 749.400 316.500 750.600 ;
        RECT 311.700 744.000 313.500 747.600 ;
        RECT 314.700 744.600 316.500 749.400 ;
        RECT 319.200 744.000 321.000 750.600 ;
        RECT 338.100 747.600 339.300 757.950 ;
        RECT 354.000 753.300 354.900 764.700 ;
        RECT 356.700 760.050 357.900 767.400 ;
        RECT 368.250 760.050 370.050 761.850 ;
        RECT 371.400 760.050 372.300 767.400 ;
        RECT 384.000 765.450 388.050 766.050 ;
        RECT 383.550 763.950 388.050 765.450 ;
        RECT 383.550 762.450 384.450 763.950 ;
        RECT 374.100 760.050 375.900 761.850 ;
        RECT 380.550 761.550 384.450 762.450 ;
        RECT 355.800 757.950 357.900 760.050 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 354.000 752.400 355.800 753.300 ;
        RECT 350.100 751.500 355.800 752.400 ;
        RECT 350.100 747.600 351.300 751.500 ;
        RECT 356.700 750.600 357.900 757.950 ;
        RECT 335.100 744.000 336.900 747.600 ;
        RECT 338.100 744.600 339.900 747.600 ;
        RECT 350.100 744.600 351.900 747.600 ;
        RECT 353.100 744.000 354.900 750.600 ;
        RECT 356.100 744.600 357.900 750.600 ;
        RECT 371.400 747.600 372.300 757.950 ;
        RECT 380.550 757.050 381.450 761.550 ;
        RECT 386.100 760.050 387.900 761.850 ;
        RECT 389.700 760.050 390.600 767.400 ;
        RECT 397.950 763.950 400.050 766.050 ;
        RECT 391.950 760.050 393.750 761.850 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 380.550 755.550 385.050 757.050 ;
        RECT 381.000 754.950 385.050 755.550 ;
        RECT 389.700 747.600 390.600 757.950 ;
        RECT 398.550 757.050 399.450 763.950 ;
        RECT 407.700 760.050 408.900 773.400 ;
        RECT 426.000 770.100 427.800 771.900 ;
        RECT 428.700 768.900 430.500 779.400 ;
        RECT 428.100 767.400 430.500 768.900 ;
        RECT 433.800 767.400 435.600 780.000 ;
        RECT 446.100 773.400 447.900 780.000 ;
        RECT 449.100 773.400 450.900 779.400 ;
        RECT 452.100 773.400 453.900 780.000 ;
        RECT 455.700 773.400 457.500 780.000 ;
        RECT 458.700 774.300 460.500 779.400 ;
        RECT 458.400 773.400 460.500 774.300 ;
        RECT 461.700 773.400 463.500 780.000 ;
        RECT 409.950 765.450 412.050 766.050 ;
        RECT 418.950 765.450 421.050 766.050 ;
        RECT 409.950 764.550 421.050 765.450 ;
        RECT 409.950 763.950 412.050 764.550 ;
        RECT 418.950 763.950 421.050 764.550 ;
        RECT 428.100 760.050 429.300 767.400 ;
        RECT 441.000 762.450 445.050 763.050 ;
        RECT 434.100 760.050 435.900 761.850 ;
        RECT 440.550 760.950 445.050 762.450 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 427.950 757.950 430.050 760.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 394.950 755.550 399.450 757.050 ;
        RECT 404.100 756.150 405.900 757.950 ;
        RECT 394.950 754.950 399.000 755.550 ;
        RECT 407.700 752.700 408.900 757.950 ;
        RECT 409.950 756.150 411.750 757.950 ;
        RECT 425.100 756.150 426.900 757.950 ;
        RECT 428.100 753.600 429.300 757.950 ;
        RECT 431.100 756.150 432.900 757.950 ;
        RECT 440.550 757.050 441.450 760.950 ;
        RECT 449.700 760.050 450.900 773.400 ;
        RECT 458.400 772.500 459.300 773.400 ;
        RECT 455.700 771.600 459.300 772.500 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 436.950 755.550 441.450 757.050 ;
        RECT 446.100 756.150 447.900 757.950 ;
        RECT 436.950 754.950 441.000 755.550 ;
        RECT 404.700 751.800 408.900 752.700 ;
        RECT 425.700 752.700 429.300 753.600 ;
        RECT 449.700 752.700 450.900 757.950 ;
        RECT 451.950 756.150 453.750 757.950 ;
        RECT 368.100 744.000 369.900 747.600 ;
        RECT 371.100 744.600 372.900 747.600 ;
        RECT 374.100 744.000 375.900 747.600 ;
        RECT 386.100 744.000 387.900 747.600 ;
        RECT 389.100 744.600 390.900 747.600 ;
        RECT 392.100 744.000 393.900 747.600 ;
        RECT 404.700 744.600 406.500 751.800 ;
        RECT 425.700 750.600 426.900 752.700 ;
        RECT 446.700 751.800 450.900 752.700 ;
        RECT 455.700 755.400 456.900 771.600 ;
        RECT 460.200 770.400 462.000 770.700 ;
        RECT 464.700 770.400 466.500 779.400 ;
        RECT 467.700 773.400 469.500 780.000 ;
        RECT 471.300 776.400 473.100 779.400 ;
        RECT 474.300 776.400 476.100 779.400 ;
        RECT 471.300 774.300 473.400 776.400 ;
        RECT 474.300 774.300 476.400 776.400 ;
        RECT 477.300 773.400 479.100 779.400 ;
        RECT 480.300 773.400 482.100 780.000 ;
        RECT 476.700 771.300 478.800 773.400 ;
        RECT 484.200 771.900 486.000 779.400 ;
        RECT 487.200 773.400 489.000 780.000 ;
        RECT 490.200 773.400 492.000 779.400 ;
        RECT 493.200 776.400 495.000 779.400 ;
        RECT 496.200 776.400 498.000 779.400 ;
        RECT 499.200 776.400 501.000 779.400 ;
        RECT 493.200 774.300 495.300 776.400 ;
        RECT 496.200 774.300 498.300 776.400 ;
        RECT 499.200 774.300 501.300 776.400 ;
        RECT 502.200 773.400 504.000 780.000 ;
        RECT 505.200 773.400 507.000 779.400 ;
        RECT 508.200 773.400 510.000 780.000 ;
        RECT 511.200 773.400 513.000 779.400 ;
        RECT 514.200 773.400 516.000 780.000 ;
        RECT 517.500 773.400 519.300 779.400 ;
        RECT 520.500 773.400 522.300 780.000 ;
        RECT 524.700 773.400 526.500 780.000 ;
        RECT 527.700 773.400 529.500 779.400 ;
        RECT 531.000 773.400 532.800 780.000 ;
        RECT 534.000 773.400 535.800 779.400 ;
        RECT 537.000 773.400 538.800 780.000 ;
        RECT 540.000 773.400 541.800 779.400 ;
        RECT 543.000 773.400 544.800 780.000 ;
        RECT 546.000 776.400 547.800 779.400 ;
        RECT 549.000 776.400 550.800 779.400 ;
        RECT 552.000 776.400 553.800 779.400 ;
        RECT 545.700 774.300 547.800 776.400 ;
        RECT 548.700 774.300 550.800 776.400 ;
        RECT 551.700 774.300 553.800 776.400 ;
        RECT 555.000 773.400 556.800 779.400 ;
        RECT 558.000 773.400 559.800 780.000 ;
        RECT 460.200 769.200 479.400 770.400 ;
        RECT 484.200 769.800 487.500 771.900 ;
        RECT 490.200 769.500 492.900 773.400 ;
        RECT 496.200 772.500 498.300 773.400 ;
        RECT 496.200 771.300 504.300 772.500 ;
        RECT 502.500 770.700 504.300 771.300 ;
        RECT 505.200 770.400 506.400 773.400 ;
        RECT 511.800 772.500 513.000 773.400 ;
        RECT 511.800 771.600 515.700 772.500 ;
        RECT 509.100 770.400 510.900 771.000 ;
        RECT 460.200 768.900 462.000 769.200 ;
        RECT 478.200 768.600 479.400 769.200 ;
        RECT 493.800 768.600 495.900 769.500 ;
        RECT 463.500 767.700 465.300 768.300 ;
        RECT 473.400 767.700 475.500 768.300 ;
        RECT 463.500 766.500 475.500 767.700 ;
        RECT 478.200 767.400 495.900 768.600 ;
        RECT 499.200 768.300 501.300 769.500 ;
        RECT 505.200 769.200 510.900 770.400 ;
        RECT 514.800 768.300 515.700 771.600 ;
        RECT 499.200 767.400 515.700 768.300 ;
        RECT 473.400 766.200 475.500 766.500 ;
        RECT 478.200 765.300 513.900 766.500 ;
        RECT 478.200 764.700 479.400 765.300 ;
        RECT 512.100 764.700 513.900 765.300 ;
        RECT 465.900 763.800 479.400 764.700 ;
        RECT 490.800 763.800 492.900 764.100 ;
        RECT 465.900 763.050 467.700 763.800 ;
        RECT 457.800 760.950 459.900 763.050 ;
        RECT 463.800 761.250 467.700 763.050 ;
        RECT 485.400 762.300 487.500 763.200 ;
        RECT 463.800 760.950 465.900 761.250 ;
        RECT 476.400 761.100 487.500 762.300 ;
        RECT 489.000 762.000 492.900 763.800 ;
        RECT 497.100 762.300 498.900 764.100 ;
        RECT 498.000 761.100 498.900 762.300 ;
        RECT 458.100 759.300 459.900 760.950 ;
        RECT 476.400 760.500 478.200 761.100 ;
        RECT 485.400 760.200 498.900 761.100 ;
        RECT 501.600 760.800 506.700 762.600 ;
        RECT 508.800 760.950 510.900 763.050 ;
        RECT 501.600 759.300 502.500 760.800 ;
        RECT 458.100 758.100 502.500 759.300 ;
        RECT 508.800 758.100 510.300 760.950 ;
        RECT 473.400 755.400 475.200 757.200 ;
        RECT 481.800 756.000 483.900 757.050 ;
        RECT 503.700 756.600 510.300 758.100 ;
        RECT 455.700 754.200 472.500 755.400 ;
        RECT 409.800 744.000 411.600 750.600 ;
        RECT 425.100 744.600 426.900 750.600 ;
        RECT 428.100 749.700 435.900 751.050 ;
        RECT 428.100 744.600 429.900 749.700 ;
        RECT 431.100 744.000 432.900 748.800 ;
        RECT 434.100 744.600 435.900 749.700 ;
        RECT 446.700 744.600 448.500 751.800 ;
        RECT 455.700 750.600 456.900 754.200 ;
        RECT 470.400 753.300 472.500 754.200 ;
        RECT 459.900 752.700 461.700 753.300 ;
        RECT 459.900 751.500 468.300 752.700 ;
        RECT 466.800 750.600 468.300 751.500 ;
        RECT 473.400 752.400 474.300 755.400 ;
        RECT 478.800 755.100 483.900 756.000 ;
        RECT 478.800 754.200 480.600 755.100 ;
        RECT 481.800 754.950 483.900 755.100 ;
        RECT 488.100 755.100 505.200 756.600 ;
        RECT 488.100 754.500 490.200 755.100 ;
        RECT 488.100 752.700 489.900 754.500 ;
        RECT 506.100 753.900 513.900 755.700 ;
        RECT 473.400 751.200 480.600 752.400 ;
        RECT 475.800 750.600 477.600 751.200 ;
        RECT 479.700 750.600 480.600 751.200 ;
        RECT 495.300 750.600 501.900 752.400 ;
        RECT 506.100 750.600 507.600 753.900 ;
        RECT 514.800 750.600 515.700 767.400 ;
        RECT 451.800 744.000 453.600 750.600 ;
        RECT 455.700 744.600 457.500 750.600 ;
        RECT 461.100 744.000 462.900 750.600 ;
        RECT 466.500 744.600 468.300 750.600 ;
        RECT 470.700 747.600 472.800 749.700 ;
        RECT 473.700 747.600 475.800 749.700 ;
        RECT 476.700 747.600 478.800 749.700 ;
        RECT 479.700 749.400 482.400 750.600 ;
        RECT 480.600 748.500 482.400 749.400 ;
        RECT 484.200 748.500 486.900 750.600 ;
        RECT 470.700 744.600 472.500 747.600 ;
        RECT 473.700 744.600 475.500 747.600 ;
        RECT 476.700 744.600 478.500 747.600 ;
        RECT 479.700 744.000 481.500 747.600 ;
        RECT 484.200 744.600 486.000 748.500 ;
        RECT 490.200 747.600 492.300 749.700 ;
        RECT 493.200 747.600 495.300 749.700 ;
        RECT 496.200 747.600 498.300 749.700 ;
        RECT 499.200 747.600 501.300 749.700 ;
        RECT 503.400 749.400 507.600 750.600 ;
        RECT 487.200 744.000 489.000 747.600 ;
        RECT 490.200 744.600 492.000 747.600 ;
        RECT 493.200 744.600 495.000 747.600 ;
        RECT 496.200 744.600 498.000 747.600 ;
        RECT 499.200 744.600 501.000 747.600 ;
        RECT 503.400 744.600 505.200 749.400 ;
        RECT 508.500 744.000 510.300 750.600 ;
        RECT 513.900 744.600 515.700 750.600 ;
        RECT 517.500 763.050 519.000 773.400 ;
        RECT 528.000 763.050 529.500 773.400 ;
        RECT 534.000 772.500 535.200 773.400 ;
        RECT 517.500 760.950 519.900 763.050 ;
        RECT 527.100 760.950 529.500 763.050 ;
        RECT 517.500 747.600 519.000 760.950 ;
        RECT 528.000 747.600 529.500 760.950 ;
        RECT 517.500 744.600 519.300 747.600 ;
        RECT 520.500 744.000 522.300 747.600 ;
        RECT 524.700 744.000 526.500 747.600 ;
        RECT 527.700 744.600 529.500 747.600 ;
        RECT 531.300 771.600 535.200 772.500 ;
        RECT 531.300 768.300 532.200 771.600 ;
        RECT 536.100 770.400 537.900 771.000 ;
        RECT 540.600 770.400 541.800 773.400 ;
        RECT 548.700 772.500 550.800 773.400 ;
        RECT 542.700 771.300 550.800 772.500 ;
        RECT 542.700 770.700 544.500 771.300 ;
        RECT 536.100 769.200 541.800 770.400 ;
        RECT 554.100 769.500 556.800 773.400 ;
        RECT 561.000 771.900 562.800 779.400 ;
        RECT 564.900 773.400 566.700 780.000 ;
        RECT 567.900 773.400 569.700 779.400 ;
        RECT 570.900 776.400 572.700 779.400 ;
        RECT 573.900 776.400 575.700 779.400 ;
        RECT 570.600 774.300 572.700 776.400 ;
        RECT 573.600 774.300 575.700 776.400 ;
        RECT 577.500 773.400 579.300 780.000 ;
        RECT 559.500 769.800 562.800 771.900 ;
        RECT 568.200 771.300 570.300 773.400 ;
        RECT 580.500 770.400 582.300 779.400 ;
        RECT 583.500 773.400 585.300 780.000 ;
        RECT 586.500 774.300 588.300 779.400 ;
        RECT 586.500 773.400 588.600 774.300 ;
        RECT 589.500 773.400 591.300 780.000 ;
        RECT 602.100 773.400 603.900 780.000 ;
        RECT 605.100 773.400 606.900 779.400 ;
        RECT 587.700 772.500 588.600 773.400 ;
        RECT 587.700 771.600 591.300 772.500 ;
        RECT 585.000 770.400 586.800 770.700 ;
        RECT 545.700 768.300 547.800 769.500 ;
        RECT 531.300 767.400 547.800 768.300 ;
        RECT 551.100 768.600 553.200 769.500 ;
        RECT 567.600 769.200 586.800 770.400 ;
        RECT 567.600 768.600 568.800 769.200 ;
        RECT 585.000 768.900 586.800 769.200 ;
        RECT 551.100 767.400 568.800 768.600 ;
        RECT 571.500 767.700 573.600 768.300 ;
        RECT 581.700 767.700 583.500 768.300 ;
        RECT 531.300 750.600 532.200 767.400 ;
        RECT 571.500 766.500 583.500 767.700 ;
        RECT 533.100 765.300 568.800 766.500 ;
        RECT 571.500 766.200 573.600 766.500 ;
        RECT 533.100 764.700 534.900 765.300 ;
        RECT 567.600 764.700 568.800 765.300 ;
        RECT 536.100 760.950 538.200 763.050 ;
        RECT 536.700 758.100 538.200 760.950 ;
        RECT 540.300 760.800 545.400 762.600 ;
        RECT 544.500 759.300 545.400 760.800 ;
        RECT 548.100 762.300 549.900 764.100 ;
        RECT 554.100 763.800 556.200 764.100 ;
        RECT 567.600 763.800 581.100 764.700 ;
        RECT 548.100 761.100 549.000 762.300 ;
        RECT 554.100 762.000 558.000 763.800 ;
        RECT 559.500 762.300 561.600 763.200 ;
        RECT 579.300 763.050 581.100 763.800 ;
        RECT 559.500 761.100 570.600 762.300 ;
        RECT 579.300 761.250 583.200 763.050 ;
        RECT 548.100 760.200 561.600 761.100 ;
        RECT 568.800 760.500 570.600 761.100 ;
        RECT 581.100 760.950 583.200 761.250 ;
        RECT 587.100 760.950 589.200 763.050 ;
        RECT 587.100 759.300 588.900 760.950 ;
        RECT 544.500 758.100 588.900 759.300 ;
        RECT 536.700 756.600 543.300 758.100 ;
        RECT 533.100 753.900 540.900 755.700 ;
        RECT 541.800 755.100 558.900 756.600 ;
        RECT 556.800 754.500 558.900 755.100 ;
        RECT 563.100 756.000 565.200 757.050 ;
        RECT 563.100 755.100 568.200 756.000 ;
        RECT 571.800 755.400 573.600 757.200 ;
        RECT 590.100 755.400 591.300 771.600 ;
        RECT 602.100 760.050 603.900 761.850 ;
        RECT 605.100 760.050 606.300 773.400 ;
        RECT 607.950 765.450 610.050 769.050 ;
        RECT 617.100 768.300 618.900 779.400 ;
        RECT 620.100 769.200 621.900 780.000 ;
        RECT 623.100 768.300 624.900 779.400 ;
        RECT 617.100 767.400 624.900 768.300 ;
        RECT 626.100 767.400 627.900 779.400 ;
        RECT 638.100 773.400 639.900 780.000 ;
        RECT 641.100 773.400 642.900 779.400 ;
        RECT 644.100 773.400 645.900 780.000 ;
        RECT 622.950 765.450 625.050 766.050 ;
        RECT 607.950 765.000 625.050 765.450 ;
        RECT 608.550 764.550 625.050 765.000 ;
        RECT 622.950 763.950 625.050 764.550 ;
        RECT 612.000 762.450 616.050 763.050 ;
        RECT 611.550 760.950 616.050 762.450 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 563.100 754.950 565.200 755.100 ;
        RECT 539.400 750.600 540.900 753.900 ;
        RECT 557.100 752.700 558.900 754.500 ;
        RECT 566.400 754.200 568.200 755.100 ;
        RECT 572.700 752.400 573.600 755.400 ;
        RECT 574.500 754.200 591.300 755.400 ;
        RECT 574.500 753.300 576.600 754.200 ;
        RECT 585.300 752.700 587.100 753.300 ;
        RECT 545.100 750.600 551.700 752.400 ;
        RECT 566.400 751.200 573.600 752.400 ;
        RECT 578.700 751.500 587.100 752.700 ;
        RECT 566.400 750.600 567.300 751.200 ;
        RECT 569.400 750.600 571.200 751.200 ;
        RECT 578.700 750.600 580.200 751.500 ;
        RECT 590.100 750.600 591.300 754.200 ;
        RECT 531.300 744.600 533.100 750.600 ;
        RECT 536.700 744.000 538.500 750.600 ;
        RECT 539.400 749.400 543.600 750.600 ;
        RECT 541.800 744.600 543.600 749.400 ;
        RECT 545.700 747.600 547.800 749.700 ;
        RECT 548.700 747.600 550.800 749.700 ;
        RECT 551.700 747.600 553.800 749.700 ;
        RECT 554.700 747.600 556.800 749.700 ;
        RECT 560.100 748.500 562.800 750.600 ;
        RECT 564.600 749.400 567.300 750.600 ;
        RECT 564.600 748.500 566.400 749.400 ;
        RECT 546.000 744.600 547.800 747.600 ;
        RECT 549.000 744.600 550.800 747.600 ;
        RECT 552.000 744.600 553.800 747.600 ;
        RECT 555.000 744.600 556.800 747.600 ;
        RECT 558.000 744.000 559.800 747.600 ;
        RECT 561.000 744.600 562.800 748.500 ;
        RECT 568.200 747.600 570.300 749.700 ;
        RECT 571.200 747.600 573.300 749.700 ;
        RECT 574.200 747.600 576.300 749.700 ;
        RECT 565.500 744.000 567.300 747.600 ;
        RECT 568.500 744.600 570.300 747.600 ;
        RECT 571.500 744.600 573.300 747.600 ;
        RECT 574.500 744.600 576.300 747.600 ;
        RECT 578.700 744.600 580.500 750.600 ;
        RECT 584.100 744.000 585.900 750.600 ;
        RECT 589.500 744.600 591.300 750.600 ;
        RECT 605.100 747.600 606.300 757.950 ;
        RECT 611.550 757.050 612.450 760.950 ;
        RECT 620.250 760.050 622.050 761.850 ;
        RECT 626.700 760.050 627.600 767.400 ;
        RECT 633.000 762.450 637.050 763.050 ;
        RECT 632.550 760.950 637.050 762.450 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 611.550 755.550 616.050 757.050 ;
        RECT 617.100 756.150 618.900 757.950 ;
        RECT 623.250 756.150 625.050 757.950 ;
        RECT 612.000 754.950 616.050 755.550 ;
        RECT 626.700 750.600 627.600 757.950 ;
        RECT 632.550 757.050 633.450 760.950 ;
        RECT 641.100 760.050 642.300 773.400 ;
        RECT 659.400 767.400 661.200 780.000 ;
        RECT 664.500 768.900 666.300 779.400 ;
        RECT 667.500 773.400 669.300 780.000 ;
        RECT 667.200 770.100 669.000 771.900 ;
        RECT 664.500 767.400 666.900 768.900 ;
        RECT 683.100 767.400 684.900 780.000 ;
        RECT 659.100 760.050 660.900 761.850 ;
        RECT 665.700 760.050 666.900 767.400 ;
        RECT 686.100 766.500 687.900 779.400 ;
        RECT 689.100 767.400 690.900 780.000 ;
        RECT 692.100 766.500 693.900 779.400 ;
        RECT 695.100 767.400 696.900 780.000 ;
        RECT 698.100 766.500 699.900 779.400 ;
        RECT 701.100 767.400 702.900 780.000 ;
        RECT 704.100 766.500 705.900 779.400 ;
        RECT 707.100 767.400 708.900 780.000 ;
        RECT 722.100 767.400 723.900 779.400 ;
        RECT 725.100 767.400 726.900 780.000 ;
        RECT 737.100 767.400 738.900 780.000 ;
        RECT 742.200 768.600 744.000 779.400 ;
        RECT 740.400 767.400 744.000 768.600 ;
        RECT 758.100 767.400 759.900 779.400 ;
        RECT 761.100 769.200 762.900 780.000 ;
        RECT 764.100 773.400 765.900 779.400 ;
        RECT 686.100 765.300 690.000 766.500 ;
        RECT 692.100 765.300 696.000 766.500 ;
        RECT 698.100 765.300 702.000 766.500 ;
        RECT 704.100 765.300 706.950 766.500 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 685.800 757.950 687.900 760.050 ;
        RECT 632.550 755.550 637.050 757.050 ;
        RECT 638.250 756.150 640.050 757.950 ;
        RECT 633.000 754.950 637.050 755.550 ;
        RECT 641.100 752.700 642.300 757.950 ;
        RECT 644.100 756.150 645.900 757.950 ;
        RECT 662.100 756.150 663.900 757.950 ;
        RECT 665.700 753.600 666.900 757.950 ;
        RECT 668.100 756.150 669.900 757.950 ;
        RECT 685.800 756.150 687.600 757.950 ;
        RECT 688.800 754.800 690.000 765.300 ;
        RECT 691.200 754.800 693.000 755.400 ;
        RECT 688.800 753.600 693.000 754.800 ;
        RECT 694.800 754.800 696.000 765.300 ;
        RECT 697.200 754.800 699.000 755.400 ;
        RECT 694.800 753.600 699.000 754.800 ;
        RECT 700.800 754.800 702.000 765.300 ;
        RECT 705.900 760.050 706.950 765.300 ;
        RECT 722.700 760.050 723.900 767.400 ;
        RECT 737.250 760.050 739.050 761.850 ;
        RECT 740.400 760.050 741.300 767.400 ;
        RECT 743.100 760.050 744.900 761.850 ;
        RECT 758.100 760.050 759.300 767.400 ;
        RECT 764.700 766.500 765.900 773.400 ;
        RECT 779.400 767.400 781.200 780.000 ;
        RECT 784.500 768.900 786.300 779.400 ;
        RECT 787.500 773.400 789.300 780.000 ;
        RECT 787.200 770.100 789.000 771.900 ;
        RECT 784.500 767.400 786.900 768.900 ;
        RECT 803.100 768.600 804.900 779.400 ;
        RECT 806.100 769.500 807.900 780.000 ;
        RECT 809.100 778.500 816.900 779.400 ;
        RECT 809.100 768.600 810.900 778.500 ;
        RECT 803.100 767.700 810.900 768.600 ;
        RECT 760.200 765.600 765.900 766.500 ;
        RECT 760.200 764.700 762.000 765.600 ;
        RECT 703.800 757.950 706.950 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 736.950 757.950 739.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 758.100 757.950 760.200 760.050 ;
        RECT 703.200 754.800 705.000 755.400 ;
        RECT 700.800 753.600 705.000 754.800 ;
        RECT 665.700 752.700 669.300 753.600 ;
        RECT 688.800 752.700 690.000 753.600 ;
        RECT 694.800 752.700 696.000 753.600 ;
        RECT 700.800 752.700 702.000 753.600 ;
        RECT 705.900 752.700 706.950 757.950 ;
        RECT 641.100 751.800 645.300 752.700 ;
        RECT 602.100 744.000 603.900 747.600 ;
        RECT 605.100 744.600 606.900 747.600 ;
        RECT 618.000 744.000 619.800 750.600 ;
        RECT 622.500 749.400 627.600 750.600 ;
        RECT 622.500 744.600 624.300 749.400 ;
        RECT 625.500 744.000 627.300 747.600 ;
        RECT 638.400 744.000 640.200 750.600 ;
        RECT 643.500 744.600 645.300 751.800 ;
        RECT 659.100 749.700 666.900 751.050 ;
        RECT 659.100 744.600 660.900 749.700 ;
        RECT 662.100 744.000 663.900 748.800 ;
        RECT 665.100 744.600 666.900 749.700 ;
        RECT 668.100 750.600 669.300 752.700 ;
        RECT 686.100 751.500 690.000 752.700 ;
        RECT 692.100 751.500 696.000 752.700 ;
        RECT 698.100 751.500 702.000 752.700 ;
        RECT 704.100 751.500 706.950 752.700 ;
        RECT 668.100 744.600 669.900 750.600 ;
        RECT 683.100 744.000 684.900 750.600 ;
        RECT 686.100 744.600 687.900 751.500 ;
        RECT 689.100 744.000 690.900 750.600 ;
        RECT 692.100 744.600 693.900 751.500 ;
        RECT 695.100 744.000 696.900 750.600 ;
        RECT 698.100 744.600 699.900 751.500 ;
        RECT 701.100 744.000 702.900 750.600 ;
        RECT 704.100 744.600 705.900 751.500 ;
        RECT 722.700 750.600 723.900 757.950 ;
        RECT 725.100 756.150 726.900 757.950 ;
        RECT 707.100 744.000 708.900 750.600 ;
        RECT 722.100 744.600 723.900 750.600 ;
        RECT 725.100 744.000 726.900 750.600 ;
        RECT 740.400 747.600 741.300 757.950 ;
        RECT 758.100 750.600 759.300 757.950 ;
        RECT 761.100 753.300 762.000 764.700 ;
        RECT 772.950 765.450 775.050 766.050 ;
        RECT 781.950 765.450 784.050 766.200 ;
        RECT 772.950 764.550 784.050 765.450 ;
        RECT 772.950 763.950 775.050 764.550 ;
        RECT 781.950 764.100 784.050 764.550 ;
        RECT 763.800 760.050 765.600 761.850 ;
        RECT 779.100 760.050 780.900 761.850 ;
        RECT 785.700 760.050 786.900 767.400 ;
        RECT 812.100 766.500 813.900 777.600 ;
        RECT 815.100 767.400 816.900 778.500 ;
        RECT 830.400 767.400 832.200 780.000 ;
        RECT 835.500 768.900 837.300 779.400 ;
        RECT 838.500 773.400 840.300 780.000 ;
        RECT 854.700 773.400 856.500 780.000 ;
        RECT 838.200 770.100 840.000 771.900 ;
        RECT 855.000 770.100 856.800 771.900 ;
        RECT 857.700 768.900 859.500 779.400 ;
        RECT 835.500 767.400 837.900 768.900 ;
        RECT 793.950 765.450 796.050 766.050 ;
        RECT 805.950 765.450 808.050 766.050 ;
        RECT 793.950 764.550 808.050 765.450 ;
        RECT 793.950 763.950 796.050 764.550 ;
        RECT 805.950 763.950 808.050 764.550 ;
        RECT 809.100 765.600 813.900 766.500 ;
        RECT 806.250 760.050 808.050 761.850 ;
        RECT 809.100 760.050 810.000 765.600 ;
        RECT 812.100 760.050 813.900 761.850 ;
        RECT 830.100 760.050 831.900 761.850 ;
        RECT 836.700 760.050 837.900 767.400 ;
        RECT 857.100 767.400 859.500 768.900 ;
        RECT 862.800 767.400 864.600 780.000 ;
        RECT 875.100 778.500 882.900 779.400 ;
        RECT 875.100 767.400 876.900 778.500 ;
        RECT 857.100 760.050 858.300 767.400 ;
        RECT 878.100 766.500 879.900 777.600 ;
        RECT 881.100 768.600 882.900 778.500 ;
        RECT 884.100 769.500 885.900 780.000 ;
        RECT 887.100 768.600 888.900 779.400 ;
        RECT 902.700 773.400 904.500 780.000 ;
        RECT 903.000 770.100 904.800 771.900 ;
        RECT 905.700 768.900 907.500 779.400 ;
        RECT 881.100 767.700 888.900 768.600 ;
        RECT 905.100 767.400 907.500 768.900 ;
        RECT 910.800 767.400 912.600 780.000 ;
        RECT 926.100 773.400 927.900 779.400 ;
        RECT 929.100 773.400 930.900 780.000 ;
        RECT 878.100 765.600 882.900 766.500 ;
        RECT 863.100 760.050 864.900 761.850 ;
        RECT 878.100 760.050 879.900 761.850 ;
        RECT 882.000 760.050 882.900 765.600 ;
        RECT 883.950 760.050 885.750 761.850 ;
        RECT 905.100 760.050 906.300 767.400 ;
        RECT 911.100 760.050 912.900 761.850 ;
        RECT 926.700 760.050 927.900 773.400 ;
        RECT 929.100 760.050 930.900 761.850 ;
        RECT 763.500 757.950 765.600 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 856.950 757.950 859.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 880.950 757.950 883.050 760.050 ;
        RECT 883.950 757.950 886.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 901.950 757.950 904.050 760.050 ;
        RECT 904.950 757.950 907.050 760.050 ;
        RECT 907.950 757.950 910.050 760.050 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 925.950 757.950 928.050 760.050 ;
        RECT 928.950 757.950 931.050 760.050 ;
        RECT 766.950 756.450 769.050 757.050 ;
        RECT 775.950 756.450 778.050 757.050 ;
        RECT 766.950 755.550 778.050 756.450 ;
        RECT 782.100 756.150 783.900 757.950 ;
        RECT 766.950 754.950 769.050 755.550 ;
        RECT 775.950 754.950 778.050 755.550 ;
        RECT 760.200 752.400 762.000 753.300 ;
        RECT 785.700 753.600 786.900 757.950 ;
        RECT 788.100 756.150 789.900 757.950 ;
        RECT 803.250 756.150 805.050 757.950 ;
        RECT 785.700 752.700 789.300 753.600 ;
        RECT 760.200 751.500 765.900 752.400 ;
        RECT 737.100 744.000 738.900 747.600 ;
        RECT 740.100 744.600 741.900 747.600 ;
        RECT 743.100 744.000 744.900 747.600 ;
        RECT 758.100 744.600 759.900 750.600 ;
        RECT 761.100 744.000 762.900 750.600 ;
        RECT 764.700 747.600 765.900 751.500 ;
        RECT 764.100 744.600 765.900 747.600 ;
        RECT 779.100 749.700 786.900 751.050 ;
        RECT 779.100 744.600 780.900 749.700 ;
        RECT 782.100 744.000 783.900 748.800 ;
        RECT 785.100 744.600 786.900 749.700 ;
        RECT 788.100 750.600 789.300 752.700 ;
        RECT 790.950 753.450 793.050 754.050 ;
        RECT 805.950 753.450 808.050 754.050 ;
        RECT 790.950 752.550 808.050 753.450 ;
        RECT 790.950 751.950 793.050 752.550 ;
        RECT 805.950 751.950 808.050 752.550 ;
        RECT 809.100 750.600 810.300 757.950 ;
        RECT 815.100 756.150 816.900 757.950 ;
        RECT 833.100 756.150 834.900 757.950 ;
        RECT 836.700 753.600 837.900 757.950 ;
        RECT 839.100 756.150 840.900 757.950 ;
        RECT 854.100 756.150 855.900 757.950 ;
        RECT 857.100 753.600 858.300 757.950 ;
        RECT 860.100 756.150 861.900 757.950 ;
        RECT 875.100 756.150 876.900 757.950 ;
        RECT 836.700 752.700 840.300 753.600 ;
        RECT 788.100 744.600 789.900 750.600 ;
        RECT 803.700 744.000 805.500 750.600 ;
        RECT 808.200 744.600 810.000 750.600 ;
        RECT 812.700 744.000 814.500 750.600 ;
        RECT 830.100 749.700 837.900 751.050 ;
        RECT 830.100 744.600 831.900 749.700 ;
        RECT 833.100 744.000 834.900 748.800 ;
        RECT 836.100 744.600 837.900 749.700 ;
        RECT 839.100 750.600 840.300 752.700 ;
        RECT 854.700 752.700 858.300 753.600 ;
        RECT 868.950 753.450 871.050 754.050 ;
        RECT 877.950 753.450 880.050 754.050 ;
        RECT 854.700 750.600 855.900 752.700 ;
        RECT 868.950 752.550 880.050 753.450 ;
        RECT 868.950 751.950 871.050 752.550 ;
        RECT 877.950 751.950 880.050 752.550 ;
        RECT 839.100 744.600 840.900 750.600 ;
        RECT 854.100 744.600 855.900 750.600 ;
        RECT 857.100 749.700 864.900 751.050 ;
        RECT 881.700 750.600 882.900 757.950 ;
        RECT 886.950 756.150 888.750 757.950 ;
        RECT 902.100 756.150 903.900 757.950 ;
        RECT 905.100 753.600 906.300 757.950 ;
        RECT 908.100 756.150 909.900 757.950 ;
        RECT 902.700 752.700 906.300 753.600 ;
        RECT 902.700 750.600 903.900 752.700 ;
        RECT 857.100 744.600 858.900 749.700 ;
        RECT 860.100 744.000 861.900 748.800 ;
        RECT 863.100 744.600 864.900 749.700 ;
        RECT 877.500 744.000 879.300 750.600 ;
        RECT 882.000 744.600 883.800 750.600 ;
        RECT 886.500 744.000 888.300 750.600 ;
        RECT 902.100 744.600 903.900 750.600 ;
        RECT 905.100 749.700 912.900 751.050 ;
        RECT 905.100 744.600 906.900 749.700 ;
        RECT 908.100 744.000 909.900 748.800 ;
        RECT 911.100 744.600 912.900 749.700 ;
        RECT 926.700 747.600 927.900 757.950 ;
        RECT 926.100 744.600 927.900 747.600 ;
        RECT 929.100 744.000 930.900 747.600 ;
        RECT 14.100 734.400 15.900 740.400 ;
        RECT 14.700 732.300 15.900 734.400 ;
        RECT 17.100 735.300 18.900 740.400 ;
        RECT 20.100 736.200 21.900 741.000 ;
        RECT 23.100 735.300 24.900 740.400 ;
        RECT 17.100 733.950 24.900 735.300 ;
        RECT 38.100 734.400 39.900 740.400 ;
        RECT 41.100 734.400 42.900 741.000 ;
        RECT 44.100 737.400 45.900 740.400 ;
        RECT 59.100 737.400 60.900 741.000 ;
        RECT 62.100 737.400 63.900 740.400 ;
        RECT 65.100 737.400 66.900 741.000 ;
        RECT 14.700 731.400 18.300 732.300 ;
        RECT 14.100 727.050 15.900 728.850 ;
        RECT 17.100 727.050 18.300 731.400 ;
        RECT 20.100 727.050 21.900 728.850 ;
        RECT 38.100 727.050 39.300 734.400 ;
        RECT 44.700 733.500 45.900 737.400 ;
        RECT 40.200 732.600 45.900 733.500 ;
        RECT 40.200 731.700 42.000 732.600 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 22.950 724.950 25.050 727.050 ;
        RECT 38.100 724.950 40.200 727.050 ;
        RECT 17.100 717.600 18.300 724.950 ;
        RECT 23.100 723.150 24.900 724.950 ;
        RECT 38.100 717.600 39.300 724.950 ;
        RECT 41.100 720.300 42.000 731.700 ;
        RECT 62.400 727.050 63.300 737.400 ;
        RECT 77.100 735.000 78.900 740.400 ;
        RECT 80.100 735.900 81.900 741.000 ;
        RECT 83.100 739.500 90.900 740.400 ;
        RECT 83.100 735.000 84.900 739.500 ;
        RECT 77.100 734.100 84.900 735.000 ;
        RECT 86.100 734.400 87.900 738.600 ;
        RECT 89.100 734.400 90.900 739.500 ;
        RECT 104.100 734.400 105.900 740.400 ;
        RECT 86.400 732.900 87.300 734.400 ;
        RECT 82.950 731.700 87.300 732.900 ;
        RECT 104.700 732.300 105.900 734.400 ;
        RECT 107.100 735.300 108.900 740.400 ;
        RECT 110.100 736.200 111.900 741.000 ;
        RECT 113.100 735.300 114.900 740.400 ;
        RECT 129.600 736.200 131.400 740.400 ;
        RECT 107.100 733.950 114.900 735.300 ;
        RECT 128.700 734.400 131.400 736.200 ;
        RECT 132.600 734.400 134.400 741.000 ;
        RECT 80.250 727.050 82.050 728.850 ;
        RECT 43.500 724.950 45.600 727.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 61.950 724.950 64.050 727.050 ;
        RECT 64.950 724.950 67.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 82.950 727.050 84.000 731.700 ;
        RECT 104.700 731.400 108.300 732.300 ;
        RECT 85.950 727.050 87.750 728.850 ;
        RECT 104.100 727.050 105.900 728.850 ;
        RECT 107.100 727.050 108.300 731.400 ;
        RECT 115.950 729.450 118.050 730.050 ;
        RECT 121.950 729.450 124.050 730.050 ;
        RECT 110.100 727.050 111.900 728.850 ;
        RECT 115.950 728.550 124.050 729.450 ;
        RECT 115.950 727.950 118.050 728.550 ;
        RECT 121.950 727.950 124.050 728.550 ;
        RECT 128.700 727.050 129.600 734.400 ;
        RECT 130.500 732.600 132.300 733.500 ;
        RECT 137.100 732.600 138.900 740.400 ;
        RECT 130.500 731.700 138.900 732.600 ;
        RECT 149.100 734.400 150.900 740.400 ;
        RECT 152.100 734.400 153.900 741.000 ;
        RECT 155.100 737.400 156.900 740.400 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 128.100 724.950 130.200 727.050 ;
        RECT 131.400 724.950 133.500 727.050 ;
        RECT 43.800 723.150 45.600 724.950 ;
        RECT 59.250 723.150 61.050 724.950 ;
        RECT 40.200 719.400 42.000 720.300 ;
        RECT 40.200 718.500 45.900 719.400 ;
        RECT 17.100 716.100 19.500 717.600 ;
        RECT 15.000 713.100 16.800 714.900 ;
        RECT 14.700 705.000 16.500 711.600 ;
        RECT 17.700 705.600 19.500 716.100 ;
        RECT 22.800 705.000 24.600 717.600 ;
        RECT 38.100 705.600 39.900 717.600 ;
        RECT 41.100 705.000 42.900 715.800 ;
        RECT 44.700 711.600 45.900 718.500 ;
        RECT 62.400 717.600 63.300 724.950 ;
        RECT 65.100 723.150 66.900 724.950 ;
        RECT 77.100 723.150 78.900 724.950 ;
        RECT 82.950 717.600 84.000 724.950 ;
        RECT 88.950 723.150 90.750 724.950 ;
        RECT 107.100 717.600 108.300 724.950 ;
        RECT 113.100 723.150 114.900 724.950 ;
        RECT 109.950 720.450 112.050 720.750 ;
        RECT 121.950 720.450 124.050 721.050 ;
        RECT 109.950 719.550 124.050 720.450 ;
        RECT 109.950 718.650 112.050 719.550 ;
        RECT 121.950 718.950 124.050 719.550 ;
        RECT 128.700 717.600 129.600 724.950 ;
        RECT 132.000 723.150 133.800 724.950 ;
        RECT 44.100 705.600 45.900 711.600 ;
        RECT 59.100 705.000 60.900 717.600 ;
        RECT 62.400 716.400 66.000 717.600 ;
        RECT 64.200 705.600 66.000 716.400 ;
        RECT 77.100 705.000 78.900 717.600 ;
        RECT 81.600 705.600 84.900 717.600 ;
        RECT 87.600 705.000 89.400 717.600 ;
        RECT 107.100 716.100 109.500 717.600 ;
        RECT 105.000 713.100 106.800 714.900 ;
        RECT 104.700 705.000 106.500 711.600 ;
        RECT 107.700 705.600 109.500 716.100 ;
        RECT 112.800 705.000 114.600 717.600 ;
        RECT 128.100 705.600 129.900 717.600 ;
        RECT 131.100 705.000 132.900 717.000 ;
        RECT 135.000 711.600 135.900 731.700 ;
        RECT 136.950 727.050 138.750 728.850 ;
        RECT 149.100 727.050 150.300 734.400 ;
        RECT 155.700 733.500 156.900 737.400 ;
        RECT 170.100 734.400 171.900 740.400 ;
        RECT 151.200 732.600 156.900 733.500 ;
        RECT 151.200 731.700 153.000 732.600 ;
        RECT 136.800 724.950 138.900 727.050 ;
        RECT 149.100 724.950 151.200 727.050 ;
        RECT 149.100 717.600 150.300 724.950 ;
        RECT 152.100 720.300 153.000 731.700 ;
        RECT 170.700 732.300 171.900 734.400 ;
        RECT 173.100 735.300 174.900 740.400 ;
        RECT 176.100 736.200 177.900 741.000 ;
        RECT 179.100 735.300 180.900 740.400 ;
        RECT 191.700 737.400 193.500 741.000 ;
        RECT 194.700 735.600 196.500 740.400 ;
        RECT 173.100 733.950 180.900 735.300 ;
        RECT 191.400 734.400 196.500 735.600 ;
        RECT 199.200 734.400 201.000 741.000 ;
        RECT 215.100 735.300 216.900 740.400 ;
        RECT 218.100 736.200 219.900 741.000 ;
        RECT 221.100 735.300 222.900 740.400 ;
        RECT 170.700 731.400 174.300 732.300 ;
        RECT 170.100 727.050 171.900 728.850 ;
        RECT 173.100 727.050 174.300 731.400 ;
        RECT 176.100 727.050 177.900 728.850 ;
        RECT 191.400 727.050 192.300 734.400 ;
        RECT 215.100 733.950 222.900 735.300 ;
        RECT 224.100 734.400 225.900 740.400 ;
        RECT 236.100 734.400 237.900 740.400 ;
        RECT 224.100 732.300 225.300 734.400 ;
        RECT 221.700 731.400 225.300 732.300 ;
        RECT 236.700 732.300 237.900 734.400 ;
        RECT 239.100 735.300 240.900 740.400 ;
        RECT 242.100 736.200 243.900 741.000 ;
        RECT 245.100 735.300 246.900 740.400 ;
        RECT 239.100 733.950 246.900 735.300 ;
        RECT 257.100 734.400 258.900 740.400 ;
        RECT 260.100 735.300 261.900 741.000 ;
        RECT 264.600 734.400 266.400 740.400 ;
        RECT 269.100 735.300 270.900 741.000 ;
        RECT 272.100 734.400 273.900 740.400 ;
        RECT 284.100 737.400 285.900 741.000 ;
        RECT 287.100 737.400 288.900 740.400 ;
        RECT 290.100 737.400 291.900 741.000 ;
        RECT 257.700 732.600 258.900 734.400 ;
        RECT 264.900 732.900 266.100 734.400 ;
        RECT 269.100 733.500 273.900 734.400 ;
        RECT 236.700 731.400 240.300 732.300 ;
        RECT 257.700 731.700 264.000 732.600 ;
        RECT 193.950 727.050 195.750 728.850 ;
        RECT 200.100 727.050 201.900 728.850 ;
        RECT 218.100 727.050 219.900 728.850 ;
        RECT 221.700 727.050 222.900 731.400 ;
        RECT 224.100 727.050 225.900 728.850 ;
        RECT 236.100 727.050 237.900 728.850 ;
        RECT 239.100 727.050 240.300 731.400 ;
        RECT 261.900 729.600 264.000 731.700 ;
        RECT 242.100 727.050 243.900 728.850 ;
        RECT 257.400 727.050 259.200 728.850 ;
        RECT 262.200 727.800 264.000 729.600 ;
        RECT 264.900 730.800 267.900 732.900 ;
        RECT 269.100 732.300 271.200 733.500 ;
        RECT 283.950 732.450 286.050 736.050 ;
        RECT 281.550 732.000 286.050 732.450 ;
        RECT 281.550 731.550 285.450 732.000 ;
        RECT 154.500 724.950 156.600 727.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 220.950 724.950 223.050 727.050 ;
        RECT 223.950 724.950 226.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 257.100 726.300 259.200 727.050 ;
        RECT 257.100 724.950 264.000 726.300 ;
        RECT 154.800 723.150 156.600 724.950 ;
        RECT 151.200 719.400 153.000 720.300 ;
        RECT 160.950 720.450 163.050 721.050 ;
        RECT 169.950 720.450 172.050 721.050 ;
        RECT 160.950 719.550 172.050 720.450 ;
        RECT 151.200 718.500 156.900 719.400 ;
        RECT 160.950 718.950 163.050 719.550 ;
        RECT 169.950 718.950 172.050 719.550 ;
        RECT 134.100 705.600 135.900 711.600 ;
        RECT 137.100 705.000 138.900 711.600 ;
        RECT 149.100 705.600 150.900 717.600 ;
        RECT 152.100 705.000 153.900 715.800 ;
        RECT 155.700 711.600 156.900 718.500 ;
        RECT 173.100 717.600 174.300 724.950 ;
        RECT 179.100 723.150 180.900 724.950 ;
        RECT 191.400 717.600 192.300 724.950 ;
        RECT 196.950 723.150 198.750 724.950 ;
        RECT 215.100 723.150 216.900 724.950 ;
        RECT 193.950 720.450 196.050 721.050 ;
        RECT 205.950 720.450 208.050 721.050 ;
        RECT 193.950 719.550 208.050 720.450 ;
        RECT 193.950 718.950 196.050 719.550 ;
        RECT 205.950 718.950 208.050 719.550 ;
        RECT 221.700 717.600 222.900 724.950 ;
        RECT 173.100 716.100 175.500 717.600 ;
        RECT 171.000 713.100 172.800 714.900 ;
        RECT 155.100 705.600 156.900 711.600 ;
        RECT 170.700 705.000 172.500 711.600 ;
        RECT 173.700 705.600 175.500 716.100 ;
        RECT 178.800 705.000 180.600 717.600 ;
        RECT 191.100 705.600 192.900 717.600 ;
        RECT 194.100 716.700 201.900 717.600 ;
        RECT 194.100 705.600 195.900 716.700 ;
        RECT 197.100 705.000 198.900 715.800 ;
        RECT 200.100 705.600 201.900 716.700 ;
        RECT 215.400 705.000 217.200 717.600 ;
        RECT 220.500 716.100 222.900 717.600 ;
        RECT 239.100 717.600 240.300 724.950 ;
        RECT 245.100 723.150 246.900 724.950 ;
        RECT 262.200 724.500 264.000 724.950 ;
        RECT 264.900 725.100 266.100 730.800 ;
        RECT 267.000 727.800 269.100 729.900 ;
        RECT 281.550 729.450 282.450 731.550 ;
        RECT 267.300 726.000 269.100 727.800 ;
        RECT 278.550 728.550 282.450 729.450 ;
        RECT 264.900 724.200 267.300 725.100 ;
        RECT 265.800 724.050 267.300 724.200 ;
        RECT 271.800 724.950 273.900 727.050 ;
        RECT 261.000 721.500 264.900 723.300 ;
        RECT 262.800 721.200 264.900 721.500 ;
        RECT 265.800 721.950 267.900 724.050 ;
        RECT 271.800 723.150 273.600 724.950 ;
        RECT 265.800 720.000 266.700 721.950 ;
        RECT 259.500 717.600 261.600 719.700 ;
        RECT 265.200 718.950 266.700 720.000 ;
        RECT 278.550 720.450 279.450 728.550 ;
        RECT 287.400 727.050 288.300 737.400 ;
        RECT 305.400 734.400 307.200 741.000 ;
        RECT 310.500 733.200 312.300 740.400 ;
        RECT 326.400 734.400 328.200 741.000 ;
        RECT 331.500 733.200 333.300 740.400 ;
        RECT 344.100 734.400 345.900 740.400 ;
        RECT 289.950 732.450 292.050 733.050 ;
        RECT 298.950 732.450 301.050 733.050 ;
        RECT 303.000 732.450 307.050 733.050 ;
        RECT 289.950 731.550 301.050 732.450 ;
        RECT 289.950 730.950 292.050 731.550 ;
        RECT 298.950 730.950 301.050 731.550 ;
        RECT 302.550 730.950 307.050 732.450 ;
        RECT 308.100 732.300 312.300 733.200 ;
        RECT 302.550 729.450 303.450 730.950 ;
        RECT 296.550 728.550 303.450 729.450 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 286.950 724.950 289.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 284.250 723.150 286.050 724.950 ;
        RECT 283.950 720.450 286.050 721.050 ;
        RECT 278.550 719.550 286.050 720.450 ;
        RECT 283.950 718.950 286.050 719.550 ;
        RECT 265.200 717.600 266.400 718.950 ;
        RECT 239.100 716.100 241.500 717.600 ;
        RECT 220.500 705.600 222.300 716.100 ;
        RECT 223.200 713.100 225.000 714.900 ;
        RECT 237.000 713.100 238.800 714.900 ;
        RECT 223.500 705.000 225.300 711.600 ;
        RECT 236.700 705.000 238.500 711.600 ;
        RECT 239.700 705.600 241.500 716.100 ;
        RECT 244.800 705.000 246.600 717.600 ;
        RECT 257.100 716.700 261.600 717.600 ;
        RECT 257.100 705.600 258.900 716.700 ;
        RECT 260.100 705.000 261.900 715.500 ;
        RECT 264.600 705.600 266.400 717.600 ;
        RECT 269.100 717.600 271.200 718.500 ;
        RECT 287.400 717.600 288.300 724.950 ;
        RECT 290.100 723.150 291.900 724.950 ;
        RECT 296.550 724.050 297.450 728.550 ;
        RECT 305.250 727.050 307.050 728.850 ;
        RECT 308.100 727.050 309.300 732.300 ;
        RECT 313.950 729.450 316.050 733.050 ;
        RECT 329.100 732.300 333.300 733.200 ;
        RECT 344.700 732.300 345.900 734.400 ;
        RECT 347.100 735.300 348.900 740.400 ;
        RECT 350.100 736.200 351.900 741.000 ;
        RECT 353.100 735.300 354.900 740.400 ;
        RECT 347.100 733.950 354.900 735.300 ;
        RECT 365.100 735.300 366.900 740.400 ;
        RECT 368.100 736.200 369.900 741.000 ;
        RECT 371.100 735.300 372.900 740.400 ;
        RECT 365.100 733.950 372.900 735.300 ;
        RECT 374.100 734.400 375.900 740.400 ;
        RECT 389.100 735.300 390.900 740.400 ;
        RECT 392.100 736.200 393.900 741.000 ;
        RECT 395.100 735.300 396.900 740.400 ;
        RECT 374.100 732.300 375.300 734.400 ;
        RECT 389.100 733.950 396.900 735.300 ;
        RECT 398.100 734.400 399.900 740.400 ;
        RECT 413.100 734.400 414.900 740.400 ;
        RECT 398.100 732.300 399.300 734.400 ;
        RECT 319.950 729.450 322.050 729.900 ;
        RECT 313.950 729.000 322.050 729.450 ;
        RECT 311.100 727.050 312.900 728.850 ;
        RECT 314.550 728.550 322.050 729.000 ;
        RECT 319.950 727.800 322.050 728.550 ;
        RECT 326.250 727.050 328.050 728.850 ;
        RECT 329.100 727.050 330.300 732.300 ;
        RECT 344.700 731.400 348.300 732.300 ;
        RECT 334.950 729.450 339.000 730.050 ;
        RECT 332.100 727.050 333.900 728.850 ;
        RECT 334.950 727.950 339.450 729.450 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 331.950 724.950 334.050 727.050 ;
        RECT 292.950 722.550 297.450 724.050 ;
        RECT 292.950 721.950 297.000 722.550 ;
        RECT 269.100 716.400 273.900 717.600 ;
        RECT 269.100 705.000 270.900 715.500 ;
        RECT 272.100 705.600 273.900 716.400 ;
        RECT 284.100 705.000 285.900 717.600 ;
        RECT 287.400 716.400 291.000 717.600 ;
        RECT 289.200 705.600 291.000 716.400 ;
        RECT 308.100 711.600 309.300 724.950 ;
        RECT 310.950 717.450 313.050 718.050 ;
        RECT 325.950 717.450 328.050 718.050 ;
        RECT 310.950 716.550 328.050 717.450 ;
        RECT 310.950 715.950 313.050 716.550 ;
        RECT 325.950 715.950 328.050 716.550 ;
        RECT 329.100 711.600 330.300 724.950 ;
        RECT 338.550 724.050 339.450 727.950 ;
        RECT 344.100 727.050 345.900 728.850 ;
        RECT 347.100 727.050 348.300 731.400 ;
        RECT 371.700 731.400 375.300 732.300 ;
        RECT 395.700 731.400 399.300 732.300 ;
        RECT 413.700 732.300 414.900 734.400 ;
        RECT 416.100 735.300 417.900 740.400 ;
        RECT 419.100 736.200 420.900 741.000 ;
        RECT 422.100 735.300 423.900 740.400 ;
        RECT 416.100 733.950 423.900 735.300 ;
        RECT 437.100 737.400 438.900 740.400 ;
        RECT 437.100 733.500 438.300 737.400 ;
        RECT 440.100 734.400 441.900 741.000 ;
        RECT 443.100 734.400 444.900 740.400 ;
        RECT 458.100 734.400 459.900 740.400 ;
        RECT 437.100 732.600 442.800 733.500 ;
        RECT 413.700 731.400 417.300 732.300 ;
        RECT 350.100 727.050 351.900 728.850 ;
        RECT 368.100 727.050 369.900 728.850 ;
        RECT 371.700 727.050 372.900 731.400 ;
        RECT 374.100 727.050 375.900 728.850 ;
        RECT 392.100 727.050 393.900 728.850 ;
        RECT 395.700 727.050 396.900 731.400 ;
        RECT 400.950 729.450 403.050 730.050 ;
        RECT 398.100 727.050 399.900 728.850 ;
        RECT 400.950 728.550 408.450 729.450 ;
        RECT 400.950 727.950 403.050 728.550 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 338.550 722.550 343.050 724.050 ;
        RECT 339.000 721.950 343.050 722.550 ;
        RECT 347.100 717.600 348.300 724.950 ;
        RECT 353.100 723.150 354.900 724.950 ;
        RECT 365.100 723.150 366.900 724.950 ;
        RECT 371.700 717.600 372.900 724.950 ;
        RECT 389.100 723.150 390.900 724.950 ;
        RECT 395.700 717.600 396.900 724.950 ;
        RECT 407.550 724.050 408.450 728.550 ;
        RECT 413.100 727.050 414.900 728.850 ;
        RECT 416.100 727.050 417.300 731.400 ;
        RECT 441.000 731.700 442.800 732.600 ;
        RECT 419.100 727.050 420.900 728.850 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 437.400 724.950 439.500 727.050 ;
        RECT 407.550 722.550 412.050 724.050 ;
        RECT 408.000 721.950 412.050 722.550 ;
        RECT 347.100 716.100 349.500 717.600 ;
        RECT 345.000 713.100 346.800 714.900 ;
        RECT 305.100 705.000 306.900 711.600 ;
        RECT 308.100 705.600 309.900 711.600 ;
        RECT 311.100 705.000 312.900 711.600 ;
        RECT 326.100 705.000 327.900 711.600 ;
        RECT 329.100 705.600 330.900 711.600 ;
        RECT 332.100 705.000 333.900 711.600 ;
        RECT 344.700 705.000 346.500 711.600 ;
        RECT 347.700 705.600 349.500 716.100 ;
        RECT 352.800 705.000 354.600 717.600 ;
        RECT 365.400 705.000 367.200 717.600 ;
        RECT 370.500 716.100 372.900 717.600 ;
        RECT 370.500 705.600 372.300 716.100 ;
        RECT 373.200 713.100 375.000 714.900 ;
        RECT 373.500 705.000 375.300 711.600 ;
        RECT 389.400 705.000 391.200 717.600 ;
        RECT 394.500 716.100 396.900 717.600 ;
        RECT 416.100 717.600 417.300 724.950 ;
        RECT 422.100 723.150 423.900 724.950 ;
        RECT 437.400 723.150 439.200 724.950 ;
        RECT 441.000 720.300 441.900 731.700 ;
        RECT 443.700 727.050 444.900 734.400 ;
        RECT 458.700 732.300 459.900 734.400 ;
        RECT 461.100 735.300 462.900 740.400 ;
        RECT 464.100 736.200 465.900 741.000 ;
        RECT 467.100 735.300 468.900 740.400 ;
        RECT 461.100 733.950 468.900 735.300 ;
        RECT 482.100 737.400 483.900 740.400 ;
        RECT 482.100 733.500 483.300 737.400 ;
        RECT 485.100 734.400 486.900 741.000 ;
        RECT 488.100 734.400 489.900 740.400 ;
        RECT 482.100 732.600 487.800 733.500 ;
        RECT 458.700 731.400 462.300 732.300 ;
        RECT 458.100 727.050 459.900 728.850 ;
        RECT 461.100 727.050 462.300 731.400 ;
        RECT 486.000 731.700 487.800 732.600 ;
        RECT 464.100 727.050 465.900 728.850 ;
        RECT 442.800 724.950 444.900 727.050 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 482.400 724.950 484.500 727.050 ;
        RECT 441.000 719.400 442.800 720.300 ;
        RECT 437.100 718.500 442.800 719.400 ;
        RECT 416.100 716.100 418.500 717.600 ;
        RECT 394.500 705.600 396.300 716.100 ;
        RECT 397.200 713.100 399.000 714.900 ;
        RECT 400.950 714.450 403.050 715.050 ;
        RECT 406.950 714.450 409.050 714.900 ;
        RECT 400.950 713.550 409.050 714.450 ;
        RECT 400.950 712.950 403.050 713.550 ;
        RECT 406.950 712.800 409.050 713.550 ;
        RECT 414.000 713.100 415.800 714.900 ;
        RECT 397.500 705.000 399.300 711.600 ;
        RECT 413.700 705.000 415.500 711.600 ;
        RECT 416.700 705.600 418.500 716.100 ;
        RECT 421.800 705.000 423.600 717.600 ;
        RECT 424.950 708.450 427.050 712.050 ;
        RECT 437.100 711.600 438.300 718.500 ;
        RECT 443.700 717.600 444.900 724.950 ;
        RECT 433.950 708.450 436.050 709.050 ;
        RECT 424.950 708.000 436.050 708.450 ;
        RECT 425.550 707.550 436.050 708.000 ;
        RECT 433.950 706.950 436.050 707.550 ;
        RECT 437.100 705.600 438.900 711.600 ;
        RECT 440.100 705.000 441.900 715.800 ;
        RECT 443.100 705.600 444.900 717.600 ;
        RECT 461.100 717.600 462.300 724.950 ;
        RECT 467.100 723.150 468.900 724.950 ;
        RECT 482.400 723.150 484.200 724.950 ;
        RECT 486.000 720.300 486.900 731.700 ;
        RECT 488.700 727.050 489.900 734.400 ;
        RECT 500.700 733.200 502.500 740.400 ;
        RECT 505.800 734.400 507.600 741.000 ;
        RECT 522.000 734.400 523.800 741.000 ;
        RECT 526.500 735.600 528.300 740.400 ;
        RECT 529.500 737.400 531.300 741.000 ;
        RECT 526.500 734.400 531.600 735.600 ;
        RECT 545.100 734.400 546.900 740.400 ;
        RECT 500.700 732.300 504.900 733.200 ;
        RECT 500.100 727.050 501.900 728.850 ;
        RECT 503.700 727.050 504.900 732.300 ;
        RECT 505.950 727.050 507.750 728.850 ;
        RECT 521.100 727.050 522.900 728.850 ;
        RECT 527.250 727.050 529.050 728.850 ;
        RECT 530.700 727.050 531.600 734.400 ;
        RECT 535.950 730.950 538.050 733.050 ;
        RECT 545.700 732.300 546.900 734.400 ;
        RECT 548.100 735.300 549.900 740.400 ;
        RECT 551.100 736.200 552.900 741.000 ;
        RECT 554.100 735.300 555.900 740.400 ;
        RECT 548.100 733.950 555.900 735.300 ;
        RECT 566.100 737.400 567.900 740.400 ;
        RECT 566.100 733.500 567.300 737.400 ;
        RECT 569.100 734.400 570.900 741.000 ;
        RECT 572.100 734.400 573.900 740.400 ;
        RECT 587.100 734.400 588.900 741.000 ;
        RECT 590.100 734.400 591.900 740.400 ;
        RECT 593.100 734.400 594.900 741.000 ;
        RECT 608.100 737.400 609.900 740.400 ;
        RECT 566.100 732.600 571.800 733.500 ;
        RECT 545.700 731.400 549.300 732.300 ;
        RECT 487.800 724.950 489.900 727.050 ;
        RECT 499.950 724.950 502.050 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 523.950 724.950 526.050 727.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 486.000 719.400 487.800 720.300 ;
        RECT 482.100 718.500 487.800 719.400 ;
        RECT 461.100 716.100 463.500 717.600 ;
        RECT 459.000 713.100 460.800 714.900 ;
        RECT 458.700 705.000 460.500 711.600 ;
        RECT 461.700 705.600 463.500 716.100 ;
        RECT 466.800 705.000 468.600 717.600 ;
        RECT 482.100 711.600 483.300 718.500 ;
        RECT 488.700 717.600 489.900 724.950 ;
        RECT 482.100 705.600 483.900 711.600 ;
        RECT 485.100 705.000 486.900 715.800 ;
        RECT 488.100 705.600 489.900 717.600 ;
        RECT 503.700 711.600 504.900 724.950 ;
        RECT 524.250 723.150 526.050 724.950 ;
        RECT 530.700 717.600 531.600 724.950 ;
        RECT 536.550 723.450 537.450 730.950 ;
        RECT 545.100 727.050 546.900 728.850 ;
        RECT 548.100 727.050 549.300 731.400 ;
        RECT 570.000 731.700 571.800 732.600 ;
        RECT 551.100 727.050 552.900 728.850 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 566.400 724.950 568.500 727.050 ;
        RECT 541.950 723.450 544.050 724.050 ;
        RECT 536.550 722.550 544.050 723.450 ;
        RECT 541.950 721.950 544.050 722.550 ;
        RECT 548.100 717.600 549.300 724.950 ;
        RECT 554.100 723.150 555.900 724.950 ;
        RECT 566.400 723.150 568.200 724.950 ;
        RECT 570.000 720.300 570.900 731.700 ;
        RECT 572.700 727.050 573.900 734.400 ;
        RECT 571.800 724.950 573.900 727.050 ;
        RECT 587.400 727.050 589.200 728.850 ;
        RECT 590.400 727.050 591.450 734.400 ;
        RECT 608.100 733.500 609.300 737.400 ;
        RECT 611.100 734.400 612.900 741.000 ;
        RECT 614.100 734.400 615.900 740.400 ;
        RECT 617.700 737.400 619.500 741.000 ;
        RECT 620.700 737.400 622.500 740.400 ;
        RECT 608.100 732.600 613.800 733.500 ;
        RECT 612.000 731.700 613.800 732.600 ;
        RECT 587.400 724.950 589.500 727.050 ;
        RECT 590.400 724.950 594.600 727.050 ;
        RECT 608.400 724.950 610.500 727.050 ;
        RECT 570.000 719.400 571.800 720.300 ;
        RECT 566.100 718.500 571.800 719.400 ;
        RECT 521.100 716.700 528.900 717.600 ;
        RECT 500.100 705.000 501.900 711.600 ;
        RECT 503.100 705.600 504.900 711.600 ;
        RECT 506.100 705.000 507.900 711.600 ;
        RECT 521.100 705.600 522.900 716.700 ;
        RECT 524.100 705.000 525.900 715.800 ;
        RECT 527.100 705.600 528.900 716.700 ;
        RECT 530.100 705.600 531.900 717.600 ;
        RECT 548.100 716.100 550.500 717.600 ;
        RECT 546.000 713.100 547.800 714.900 ;
        RECT 545.700 705.000 547.500 711.600 ;
        RECT 548.700 705.600 550.500 716.100 ;
        RECT 553.800 705.000 555.600 717.600 ;
        RECT 566.100 711.600 567.300 718.500 ;
        RECT 572.700 717.600 573.900 724.950 ;
        RECT 590.400 717.600 591.450 724.950 ;
        RECT 608.400 723.150 610.200 724.950 ;
        RECT 612.000 720.300 612.900 731.700 ;
        RECT 614.700 727.050 615.900 734.400 ;
        RECT 613.800 724.950 615.900 727.050 ;
        RECT 612.000 719.400 613.800 720.300 ;
        RECT 608.100 718.500 613.800 719.400 ;
        RECT 566.100 705.600 567.900 711.600 ;
        RECT 569.100 705.000 570.900 715.800 ;
        RECT 572.100 705.600 573.900 717.600 ;
        RECT 587.100 705.000 588.900 717.600 ;
        RECT 590.100 705.600 591.900 717.600 ;
        RECT 593.100 705.000 594.900 717.600 ;
        RECT 608.100 711.600 609.300 718.500 ;
        RECT 614.700 717.600 615.900 724.950 ;
        RECT 621.000 724.050 622.500 737.400 ;
        RECT 620.100 721.950 622.500 724.050 ;
        RECT 608.100 705.600 609.900 711.600 ;
        RECT 611.100 705.000 612.900 715.800 ;
        RECT 614.100 705.600 615.900 717.600 ;
        RECT 621.000 711.600 622.500 721.950 ;
        RECT 624.300 734.400 626.100 740.400 ;
        RECT 629.700 734.400 631.500 741.000 ;
        RECT 634.800 735.600 636.600 740.400 ;
        RECT 639.000 737.400 640.800 740.400 ;
        RECT 642.000 737.400 643.800 740.400 ;
        RECT 645.000 737.400 646.800 740.400 ;
        RECT 648.000 737.400 649.800 740.400 ;
        RECT 651.000 737.400 652.800 741.000 ;
        RECT 632.400 734.400 636.600 735.600 ;
        RECT 638.700 735.300 640.800 737.400 ;
        RECT 641.700 735.300 643.800 737.400 ;
        RECT 644.700 735.300 646.800 737.400 ;
        RECT 647.700 735.300 649.800 737.400 ;
        RECT 654.000 736.500 655.800 740.400 ;
        RECT 658.500 737.400 660.300 741.000 ;
        RECT 661.500 737.400 663.300 740.400 ;
        RECT 664.500 737.400 666.300 740.400 ;
        RECT 667.500 737.400 669.300 740.400 ;
        RECT 653.100 734.400 655.800 736.500 ;
        RECT 657.600 735.600 659.400 736.500 ;
        RECT 657.600 734.400 660.300 735.600 ;
        RECT 661.200 735.300 663.300 737.400 ;
        RECT 664.200 735.300 666.300 737.400 ;
        RECT 667.200 735.300 669.300 737.400 ;
        RECT 671.700 734.400 673.500 740.400 ;
        RECT 677.100 734.400 678.900 741.000 ;
        RECT 682.500 734.400 684.300 740.400 ;
        RECT 699.000 734.400 700.800 741.000 ;
        RECT 703.500 735.600 705.300 740.400 ;
        RECT 706.500 737.400 708.300 741.000 ;
        RECT 703.500 734.400 708.600 735.600 ;
        RECT 721.500 734.400 723.300 741.000 ;
        RECT 726.000 734.400 727.800 740.400 ;
        RECT 730.500 734.400 732.300 741.000 ;
        RECT 733.950 735.450 736.050 739.050 ;
        RECT 746.100 737.400 747.900 741.000 ;
        RECT 749.100 737.400 750.900 740.400 ;
        RECT 745.950 735.450 748.050 736.050 ;
        RECT 733.950 735.000 748.050 735.450 ;
        RECT 734.550 734.550 748.050 735.000 ;
        RECT 624.300 717.600 625.200 734.400 ;
        RECT 632.400 731.100 633.900 734.400 ;
        RECT 638.100 732.600 644.700 734.400 ;
        RECT 659.400 733.800 660.300 734.400 ;
        RECT 662.400 733.800 664.200 734.400 ;
        RECT 659.400 732.600 666.600 733.800 ;
        RECT 626.100 729.300 633.900 731.100 ;
        RECT 650.100 730.500 651.900 732.300 ;
        RECT 649.800 729.900 651.900 730.500 ;
        RECT 634.800 728.400 651.900 729.900 ;
        RECT 656.100 729.900 658.200 730.050 ;
        RECT 659.400 729.900 661.200 730.800 ;
        RECT 656.100 729.000 661.200 729.900 ;
        RECT 665.700 729.600 666.600 732.600 ;
        RECT 671.700 733.500 673.200 734.400 ;
        RECT 671.700 732.300 680.100 733.500 ;
        RECT 678.300 731.700 680.100 732.300 ;
        RECT 667.500 730.800 669.600 731.700 ;
        RECT 683.100 730.800 684.300 734.400 ;
        RECT 667.500 729.600 684.300 730.800 ;
        RECT 629.700 726.900 636.300 728.400 ;
        RECT 656.100 727.950 658.200 729.000 ;
        RECT 664.800 727.800 666.600 729.600 ;
        RECT 629.700 724.050 631.200 726.900 ;
        RECT 637.500 725.700 681.900 726.900 ;
        RECT 637.500 724.200 638.400 725.700 ;
        RECT 629.100 721.950 631.200 724.050 ;
        RECT 633.300 722.400 638.400 724.200 ;
        RECT 641.100 723.900 654.600 724.800 ;
        RECT 661.800 723.900 663.600 724.500 ;
        RECT 680.100 724.050 681.900 725.700 ;
        RECT 641.100 722.700 642.000 723.900 ;
        RECT 641.100 720.900 642.900 722.700 ;
        RECT 647.100 721.200 651.000 723.000 ;
        RECT 652.500 722.700 663.600 723.900 ;
        RECT 674.100 723.750 676.200 724.050 ;
        RECT 652.500 721.800 654.600 722.700 ;
        RECT 672.300 721.950 676.200 723.750 ;
        RECT 680.100 721.950 682.200 724.050 ;
        RECT 672.300 721.200 674.100 721.950 ;
        RECT 647.100 720.900 649.200 721.200 ;
        RECT 660.600 720.300 674.100 721.200 ;
        RECT 626.100 719.700 627.900 720.300 ;
        RECT 660.600 719.700 661.800 720.300 ;
        RECT 626.100 718.500 661.800 719.700 ;
        RECT 664.500 718.500 666.600 718.800 ;
        RECT 624.300 716.700 640.800 717.600 ;
        RECT 624.300 713.400 625.200 716.700 ;
        RECT 629.100 714.600 634.800 715.800 ;
        RECT 638.700 715.500 640.800 716.700 ;
        RECT 644.100 716.400 661.800 717.600 ;
        RECT 664.500 717.300 676.500 718.500 ;
        RECT 664.500 716.700 666.600 717.300 ;
        RECT 674.700 716.700 676.500 717.300 ;
        RECT 644.100 715.500 646.200 716.400 ;
        RECT 660.600 715.800 661.800 716.400 ;
        RECT 678.000 715.800 679.800 716.100 ;
        RECT 629.100 714.000 630.900 714.600 ;
        RECT 624.300 712.500 628.200 713.400 ;
        RECT 627.000 711.600 628.200 712.500 ;
        RECT 633.600 711.600 634.800 714.600 ;
        RECT 635.700 713.700 637.500 714.300 ;
        RECT 635.700 712.500 643.800 713.700 ;
        RECT 641.700 711.600 643.800 712.500 ;
        RECT 647.100 711.600 649.800 715.500 ;
        RECT 652.500 713.100 655.800 715.200 ;
        RECT 660.600 714.600 679.800 715.800 ;
        RECT 617.700 705.000 619.500 711.600 ;
        RECT 620.700 705.600 622.500 711.600 ;
        RECT 624.000 705.000 625.800 711.600 ;
        RECT 627.000 705.600 628.800 711.600 ;
        RECT 630.000 705.000 631.800 711.600 ;
        RECT 633.000 705.600 634.800 711.600 ;
        RECT 636.000 705.000 637.800 711.600 ;
        RECT 638.700 708.600 640.800 710.700 ;
        RECT 641.700 708.600 643.800 710.700 ;
        RECT 644.700 708.600 646.800 710.700 ;
        RECT 639.000 705.600 640.800 708.600 ;
        RECT 642.000 705.600 643.800 708.600 ;
        RECT 645.000 705.600 646.800 708.600 ;
        RECT 648.000 705.600 649.800 711.600 ;
        RECT 651.000 705.000 652.800 711.600 ;
        RECT 654.000 705.600 655.800 713.100 ;
        RECT 661.200 711.600 663.300 713.700 ;
        RECT 657.900 705.000 659.700 711.600 ;
        RECT 660.900 705.600 662.700 711.600 ;
        RECT 663.600 708.600 665.700 710.700 ;
        RECT 666.600 708.600 668.700 710.700 ;
        RECT 663.900 705.600 665.700 708.600 ;
        RECT 666.900 705.600 668.700 708.600 ;
        RECT 670.500 705.000 672.300 711.600 ;
        RECT 673.500 705.600 675.300 714.600 ;
        RECT 678.000 714.300 679.800 714.600 ;
        RECT 683.100 713.400 684.300 729.600 ;
        RECT 698.100 727.050 699.900 728.850 ;
        RECT 704.250 727.050 706.050 728.850 ;
        RECT 707.700 727.050 708.600 734.400 ;
        RECT 719.100 727.050 720.900 728.850 ;
        RECT 725.700 727.050 726.900 734.400 ;
        RECT 745.950 733.950 748.050 734.550 ;
        RECT 727.950 732.450 730.050 733.050 ;
        RECT 742.950 732.450 745.050 733.050 ;
        RECT 727.950 731.550 745.050 732.450 ;
        RECT 727.950 730.950 730.050 731.550 ;
        RECT 742.950 730.950 745.050 731.550 ;
        RECT 730.950 727.050 732.750 728.850 ;
        RECT 749.100 727.050 750.300 737.400 ;
        RECT 751.950 735.450 754.050 736.050 ;
        RECT 757.950 735.450 760.050 736.050 ;
        RECT 751.950 734.550 760.050 735.450 ;
        RECT 751.950 733.950 754.050 734.550 ;
        RECT 757.950 733.950 760.050 734.550 ;
        RECT 761.100 735.300 762.900 740.400 ;
        RECT 764.100 736.200 765.900 741.000 ;
        RECT 767.100 735.300 768.900 740.400 ;
        RECT 761.100 733.950 768.900 735.300 ;
        RECT 770.100 734.400 771.900 740.400 ;
        RECT 770.100 732.300 771.300 734.400 ;
        RECT 767.700 731.400 771.300 732.300 ;
        RECT 784.500 732.000 786.300 740.400 ;
        RECT 764.100 727.050 765.900 728.850 ;
        RECT 767.700 727.050 768.900 731.400 ;
        RECT 783.000 730.800 786.300 732.000 ;
        RECT 791.100 731.400 792.900 741.000 ;
        RECT 806.100 737.400 807.900 741.000 ;
        RECT 809.100 737.400 810.900 740.400 ;
        RECT 770.100 727.050 771.900 728.850 ;
        RECT 783.000 727.050 783.900 730.800 ;
        RECT 785.100 727.050 786.900 728.850 ;
        RECT 791.100 727.050 792.900 728.850 ;
        RECT 809.100 727.050 810.300 737.400 ;
        RECT 824.100 735.300 825.900 740.400 ;
        RECT 827.100 736.200 828.900 741.000 ;
        RECT 830.100 735.300 831.900 740.400 ;
        RECT 824.100 733.950 831.900 735.300 ;
        RECT 833.100 734.400 834.900 740.400 ;
        RECT 833.100 732.300 834.300 734.400 ;
        RECT 830.700 731.400 834.300 732.300 ;
        RECT 848.100 731.400 849.900 741.000 ;
        RECT 854.700 732.000 856.500 740.400 ;
        RECT 872.100 734.400 873.900 740.400 ;
        RECT 872.700 732.300 873.900 734.400 ;
        RECT 875.100 735.300 876.900 740.400 ;
        RECT 878.100 736.200 879.900 741.000 ;
        RECT 881.100 735.300 882.900 740.400 ;
        RECT 875.100 733.950 882.900 735.300 ;
        RECT 893.100 735.300 894.900 740.400 ;
        RECT 896.100 736.200 897.900 741.000 ;
        RECT 899.100 735.300 900.900 740.400 ;
        RECT 893.100 733.950 900.900 735.300 ;
        RECT 902.100 734.400 903.900 740.400 ;
        RECT 914.100 737.400 915.900 741.000 ;
        RECT 917.100 737.400 918.900 740.400 ;
        RECT 920.100 737.400 921.900 741.000 ;
        RECT 902.100 732.300 903.300 734.400 ;
        RECT 827.100 727.050 828.900 728.850 ;
        RECT 830.700 727.050 831.900 731.400 ;
        RECT 854.700 730.800 858.000 732.000 ;
        RECT 872.700 731.400 876.300 732.300 ;
        RECT 833.100 727.050 834.900 728.850 ;
        RECT 848.100 727.050 849.900 728.850 ;
        RECT 854.100 727.050 855.900 728.850 ;
        RECT 857.100 727.050 858.000 730.800 ;
        RECT 872.100 727.050 873.900 728.850 ;
        RECT 875.100 727.050 876.300 731.400 ;
        RECT 899.700 731.400 903.300 732.300 ;
        RECT 907.950 732.450 910.050 733.050 ;
        RECT 913.950 732.450 916.050 733.050 ;
        RECT 907.950 731.550 916.050 732.450 ;
        RECT 878.100 727.050 879.900 728.850 ;
        RECT 896.100 727.050 897.900 728.850 ;
        RECT 899.700 727.050 900.900 731.400 ;
        RECT 907.950 730.950 910.050 731.550 ;
        RECT 913.950 730.950 916.050 731.550 ;
        RECT 902.100 727.050 903.900 728.850 ;
        RECT 917.700 727.050 918.600 737.400 ;
        RECT 935.100 734.400 936.900 740.400 ;
        RECT 935.700 732.300 936.900 734.400 ;
        RECT 938.100 735.300 939.900 740.400 ;
        RECT 941.100 736.200 942.900 741.000 ;
        RECT 944.100 735.300 945.900 740.400 ;
        RECT 938.100 733.950 945.900 735.300 ;
        RECT 935.700 731.400 939.300 732.300 ;
        RECT 935.100 727.050 936.900 728.850 ;
        RECT 938.100 727.050 939.300 731.400 ;
        RECT 941.100 727.050 942.900 728.850 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 760.950 724.950 763.050 727.050 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 787.950 724.950 790.050 727.050 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 832.950 724.950 835.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 856.950 724.950 859.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 877.950 724.950 880.050 727.050 ;
        RECT 880.950 724.950 883.050 727.050 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 898.950 724.950 901.050 727.050 ;
        RECT 901.950 724.950 904.050 727.050 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 916.950 724.950 919.050 727.050 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 934.950 724.950 937.050 727.050 ;
        RECT 937.950 724.950 940.050 727.050 ;
        RECT 940.950 724.950 943.050 727.050 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 701.250 723.150 703.050 724.950 ;
        RECT 707.700 717.600 708.600 724.950 ;
        RECT 722.100 723.150 723.900 724.950 ;
        RECT 726.000 719.400 726.900 724.950 ;
        RECT 727.950 723.150 729.750 724.950 ;
        RECT 746.100 723.150 747.900 724.950 ;
        RECT 722.100 718.500 726.900 719.400 ;
        RECT 680.700 712.500 684.300 713.400 ;
        RECT 698.100 716.700 705.900 717.600 ;
        RECT 680.700 711.600 681.600 712.500 ;
        RECT 676.500 705.000 678.300 711.600 ;
        RECT 679.500 710.700 681.600 711.600 ;
        RECT 679.500 705.600 681.300 710.700 ;
        RECT 682.500 705.000 684.300 711.600 ;
        RECT 698.100 705.600 699.900 716.700 ;
        RECT 701.100 705.000 702.900 715.800 ;
        RECT 704.100 705.600 705.900 716.700 ;
        RECT 707.100 705.600 708.900 717.600 ;
        RECT 719.100 706.500 720.900 717.600 ;
        RECT 722.100 707.400 723.900 718.500 ;
        RECT 725.100 716.400 732.900 717.300 ;
        RECT 725.100 706.500 726.900 716.400 ;
        RECT 719.100 705.600 726.900 706.500 ;
        RECT 728.100 705.000 729.900 715.500 ;
        RECT 731.100 705.600 732.900 716.400 ;
        RECT 749.100 711.600 750.300 724.950 ;
        RECT 761.100 723.150 762.900 724.950 ;
        RECT 767.700 717.600 768.900 724.950 ;
        RECT 746.100 705.000 747.900 711.600 ;
        RECT 749.100 705.600 750.900 711.600 ;
        RECT 761.400 705.000 763.200 717.600 ;
        RECT 766.500 716.100 768.900 717.600 ;
        RECT 766.500 705.600 768.300 716.100 ;
        RECT 769.200 713.100 771.000 714.900 ;
        RECT 783.000 712.800 783.900 724.950 ;
        RECT 788.100 723.150 789.900 724.950 ;
        RECT 806.100 723.150 807.900 724.950 ;
        RECT 784.950 720.450 787.050 720.750 ;
        RECT 790.950 720.450 793.050 721.050 ;
        RECT 805.950 720.450 808.050 721.050 ;
        RECT 784.950 719.550 808.050 720.450 ;
        RECT 784.950 718.650 787.050 719.550 ;
        RECT 790.950 718.950 793.050 719.550 ;
        RECT 805.950 718.950 808.050 719.550 ;
        RECT 783.000 711.900 789.600 712.800 ;
        RECT 783.000 711.600 783.900 711.900 ;
        RECT 769.500 705.000 771.300 711.600 ;
        RECT 782.100 705.600 783.900 711.600 ;
        RECT 788.100 711.600 789.600 711.900 ;
        RECT 809.100 711.600 810.300 724.950 ;
        RECT 824.100 723.150 825.900 724.950 ;
        RECT 814.950 720.450 817.050 721.050 ;
        RECT 826.950 720.450 829.050 720.750 ;
        RECT 814.950 719.550 829.050 720.450 ;
        RECT 814.950 718.950 817.050 719.550 ;
        RECT 826.950 718.650 829.050 719.550 ;
        RECT 830.700 717.600 831.900 724.950 ;
        RECT 851.100 723.150 852.900 724.950 ;
        RECT 785.100 705.000 786.900 711.000 ;
        RECT 788.100 705.600 789.900 711.600 ;
        RECT 791.100 705.000 792.900 711.600 ;
        RECT 806.100 705.000 807.900 711.600 ;
        RECT 809.100 705.600 810.900 711.600 ;
        RECT 824.400 705.000 826.200 717.600 ;
        RECT 829.500 716.100 831.900 717.600 ;
        RECT 832.950 717.450 835.050 718.050 ;
        RECT 841.950 717.450 844.050 718.050 ;
        RECT 832.950 716.550 844.050 717.450 ;
        RECT 829.500 705.600 831.300 716.100 ;
        RECT 832.950 715.950 835.050 716.550 ;
        RECT 841.950 715.950 844.050 716.550 ;
        RECT 832.200 713.100 834.000 714.900 ;
        RECT 857.100 712.800 858.000 724.950 ;
        RECT 875.100 717.600 876.300 724.950 ;
        RECT 881.100 723.150 882.900 724.950 ;
        RECT 893.100 723.150 894.900 724.950 ;
        RECT 899.700 717.600 900.900 724.950 ;
        RECT 914.100 723.150 915.900 724.950 ;
        RECT 917.700 717.600 918.600 724.950 ;
        RECT 919.950 723.150 921.750 724.950 ;
        RECT 938.100 717.600 939.300 724.950 ;
        RECT 944.100 723.150 945.900 724.950 ;
        RECT 875.100 716.100 877.500 717.600 ;
        RECT 873.000 713.100 874.800 714.900 ;
        RECT 851.400 711.900 858.000 712.800 ;
        RECT 851.400 711.600 852.900 711.900 ;
        RECT 832.500 705.000 834.300 711.600 ;
        RECT 848.100 705.000 849.900 711.600 ;
        RECT 851.100 705.600 852.900 711.600 ;
        RECT 857.100 711.600 858.000 711.900 ;
        RECT 854.100 705.000 855.900 711.000 ;
        RECT 857.100 705.600 858.900 711.600 ;
        RECT 872.700 705.000 874.500 711.600 ;
        RECT 875.700 705.600 877.500 716.100 ;
        RECT 880.800 705.000 882.600 717.600 ;
        RECT 893.400 705.000 895.200 717.600 ;
        RECT 898.500 716.100 900.900 717.600 ;
        RECT 915.000 716.400 918.600 717.600 ;
        RECT 898.500 705.600 900.300 716.100 ;
        RECT 901.200 713.100 903.000 714.900 ;
        RECT 901.500 705.000 903.300 711.600 ;
        RECT 915.000 705.600 916.800 716.400 ;
        RECT 920.100 705.000 921.900 717.600 ;
        RECT 938.100 716.100 940.500 717.600 ;
        RECT 936.000 713.100 937.800 714.900 ;
        RECT 935.700 705.000 937.500 711.600 ;
        RECT 938.700 705.600 940.500 716.100 ;
        RECT 943.800 705.000 945.600 717.600 ;
        RECT 11.100 689.400 12.900 702.000 ;
        RECT 14.100 689.400 15.900 701.400 ;
        RECT 17.100 689.400 18.900 702.000 ;
        RECT 32.100 689.400 33.900 702.000 ;
        RECT 35.100 689.400 36.900 701.400 ;
        RECT 51.000 690.600 52.800 701.400 ;
        RECT 51.000 689.400 54.600 690.600 ;
        RECT 56.100 689.400 57.900 702.000 ;
        RECT 71.100 700.500 78.900 701.400 ;
        RECT 71.100 689.400 72.900 700.500 ;
        RECT 14.400 682.050 15.450 689.400 ;
        RECT 35.100 682.050 36.300 689.400 ;
        RECT 50.100 682.050 51.900 683.850 ;
        RECT 53.700 682.050 54.600 689.400 ;
        RECT 74.100 688.500 75.900 699.600 ;
        RECT 77.100 690.600 78.900 700.500 ;
        RECT 80.100 691.500 81.900 702.000 ;
        RECT 83.100 690.600 84.900 701.400 ;
        RECT 95.100 695.400 96.900 702.000 ;
        RECT 98.100 695.400 99.900 701.400 ;
        RECT 101.100 695.400 102.900 702.000 ;
        RECT 116.700 695.400 118.500 702.000 ;
        RECT 77.100 689.700 84.900 690.600 ;
        RECT 74.100 687.600 78.900 688.500 ;
        RECT 55.950 682.050 57.750 683.850 ;
        RECT 74.100 682.050 75.900 683.850 ;
        RECT 78.000 682.050 78.900 687.600 ;
        RECT 79.950 682.050 81.750 683.850 ;
        RECT 98.100 682.050 99.300 695.400 ;
        RECT 117.000 692.100 118.800 693.900 ;
        RECT 119.700 690.900 121.500 701.400 ;
        RECT 119.100 689.400 121.500 690.900 ;
        RECT 124.800 689.400 126.600 702.000 ;
        RECT 140.100 689.400 141.900 701.400 ;
        RECT 143.100 690.000 144.900 702.000 ;
        RECT 146.100 695.400 147.900 701.400 ;
        RECT 149.100 695.400 150.900 702.000 ;
        RECT 161.100 695.400 162.900 702.000 ;
        RECT 164.100 695.400 165.900 701.400 ;
        RECT 179.100 695.400 180.900 702.000 ;
        RECT 182.100 695.400 183.900 701.400 ;
        RECT 185.100 695.400 186.900 702.000 ;
        RECT 190.950 696.450 193.050 696.900 ;
        RECT 196.950 696.450 199.050 697.050 ;
        RECT 190.950 695.550 199.050 696.450 ;
        RECT 119.100 682.050 120.300 689.400 ;
        RECT 121.950 687.450 124.050 688.050 ;
        RECT 133.950 687.450 136.050 688.050 ;
        RECT 121.950 686.550 136.050 687.450 ;
        RECT 121.950 685.950 124.050 686.550 ;
        RECT 133.950 685.950 136.050 686.550 ;
        RECT 125.100 682.050 126.900 683.850 ;
        RECT 140.700 682.050 141.600 689.400 ;
        RECT 144.000 682.050 145.800 683.850 ;
        RECT 11.400 679.950 13.500 682.050 ;
        RECT 14.400 679.950 18.600 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 73.950 679.950 76.050 682.050 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 94.950 679.950 97.050 682.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 121.950 679.950 124.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 140.100 679.950 142.200 682.050 ;
        RECT 143.400 679.950 145.500 682.050 ;
        RECT 11.400 678.150 13.200 679.950 ;
        RECT 14.400 672.600 15.450 679.950 ;
        RECT 32.100 678.150 33.900 679.950 ;
        RECT 35.100 672.600 36.300 679.950 ;
        RECT 11.100 666.000 12.900 672.600 ;
        RECT 14.100 666.600 15.900 672.600 ;
        RECT 17.100 666.000 18.900 672.600 ;
        RECT 32.100 666.000 33.900 672.600 ;
        RECT 35.100 666.600 36.900 672.600 ;
        RECT 53.700 669.600 54.600 679.950 ;
        RECT 71.100 678.150 72.900 679.950 ;
        RECT 77.700 672.600 78.900 679.950 ;
        RECT 82.950 678.150 84.750 679.950 ;
        RECT 95.250 678.150 97.050 679.950 ;
        RECT 98.100 674.700 99.300 679.950 ;
        RECT 101.100 678.150 102.900 679.950 ;
        RECT 116.100 678.150 117.900 679.950 ;
        RECT 119.100 675.600 120.300 679.950 ;
        RECT 122.100 678.150 123.900 679.950 ;
        RECT 116.700 674.700 120.300 675.600 ;
        RECT 98.100 673.800 102.300 674.700 ;
        RECT 50.100 666.000 51.900 669.600 ;
        RECT 53.100 666.600 54.900 669.600 ;
        RECT 56.100 666.000 57.900 669.600 ;
        RECT 73.500 666.000 75.300 672.600 ;
        RECT 78.000 666.600 79.800 672.600 ;
        RECT 82.500 666.000 84.300 672.600 ;
        RECT 95.400 666.000 97.200 672.600 ;
        RECT 100.500 666.600 102.300 673.800 ;
        RECT 116.700 672.600 117.900 674.700 ;
        RECT 116.100 666.600 117.900 672.600 ;
        RECT 119.100 671.700 126.900 673.050 ;
        RECT 119.100 666.600 120.900 671.700 ;
        RECT 122.100 666.000 123.900 670.800 ;
        RECT 125.100 666.600 126.900 671.700 ;
        RECT 140.700 672.600 141.600 679.950 ;
        RECT 147.000 675.300 147.900 695.400 ;
        RECT 161.100 682.050 162.900 683.850 ;
        RECT 164.100 682.050 165.300 695.400 ;
        RECT 182.700 682.050 183.900 695.400 ;
        RECT 190.950 694.800 193.050 695.550 ;
        RECT 196.950 694.950 199.050 695.550 ;
        RECT 200.100 690.600 201.900 701.400 ;
        RECT 203.100 691.500 204.900 702.000 ;
        RECT 206.100 700.500 213.900 701.400 ;
        RECT 206.100 690.600 207.900 700.500 ;
        RECT 200.100 689.700 207.900 690.600 ;
        RECT 209.100 688.500 210.900 699.600 ;
        RECT 212.100 689.400 213.900 700.500 ;
        RECT 227.100 695.400 228.900 702.000 ;
        RECT 230.100 695.400 231.900 701.400 ;
        RECT 233.100 695.400 234.900 702.000 ;
        RECT 245.100 695.400 246.900 702.000 ;
        RECT 248.100 695.400 249.900 701.400 ;
        RECT 251.100 695.400 252.900 702.000 ;
        RECT 193.950 687.450 196.050 688.050 ;
        RECT 202.950 687.450 205.050 688.050 ;
        RECT 193.950 686.550 205.050 687.450 ;
        RECT 193.950 685.950 196.050 686.550 ;
        RECT 202.950 685.950 205.050 686.550 ;
        RECT 206.100 687.600 210.900 688.500 ;
        RECT 195.000 684.450 199.050 685.050 ;
        RECT 194.550 682.950 199.050 684.450 ;
        RECT 148.800 679.950 150.900 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 148.950 678.150 150.750 679.950 ;
        RECT 142.500 674.400 150.900 675.300 ;
        RECT 142.500 673.500 144.300 674.400 ;
        RECT 140.700 670.800 143.400 672.600 ;
        RECT 141.600 666.600 143.400 670.800 ;
        RECT 144.600 666.000 146.400 672.600 ;
        RECT 149.100 666.600 150.900 674.400 ;
        RECT 164.100 669.600 165.300 679.950 ;
        RECT 179.100 678.150 180.900 679.950 ;
        RECT 182.700 674.700 183.900 679.950 ;
        RECT 184.950 678.150 186.750 679.950 ;
        RECT 179.700 673.800 183.900 674.700 ;
        RECT 184.950 675.450 187.050 676.050 ;
        RECT 194.550 675.450 195.450 682.950 ;
        RECT 203.250 682.050 205.050 683.850 ;
        RECT 206.100 682.050 207.000 687.600 ;
        RECT 214.950 684.450 219.000 685.050 ;
        RECT 209.100 682.050 210.900 683.850 ;
        RECT 214.950 682.950 219.450 684.450 ;
        RECT 199.950 679.950 202.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 200.250 678.150 202.050 679.950 ;
        RECT 184.950 674.550 195.450 675.450 ;
        RECT 184.950 673.950 187.050 674.550 ;
        RECT 161.100 666.000 162.900 669.600 ;
        RECT 164.100 666.600 165.900 669.600 ;
        RECT 179.700 666.600 181.500 673.800 ;
        RECT 206.100 672.600 207.300 679.950 ;
        RECT 212.100 678.150 213.900 679.950 ;
        RECT 211.950 675.450 214.050 676.050 ;
        RECT 218.550 675.450 219.450 682.950 ;
        RECT 230.700 682.050 231.900 695.400 ;
        RECT 248.700 682.050 249.900 695.400 ;
        RECT 266.100 689.400 267.900 701.400 ;
        RECT 269.100 690.000 270.900 702.000 ;
        RECT 272.100 695.400 273.900 701.400 ;
        RECT 275.100 695.400 276.900 702.000 ;
        RECT 266.700 682.050 267.600 689.400 ;
        RECT 270.000 682.050 271.800 683.850 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 244.950 679.950 247.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 266.100 679.950 268.200 682.050 ;
        RECT 269.400 679.950 271.500 682.050 ;
        RECT 227.100 678.150 228.900 679.950 ;
        RECT 211.950 674.550 219.450 675.450 ;
        RECT 230.700 674.700 231.900 679.950 ;
        RECT 232.950 678.150 234.750 679.950 ;
        RECT 245.100 678.150 246.900 679.950 ;
        RECT 248.700 674.700 249.900 679.950 ;
        RECT 250.950 678.150 252.750 679.950 ;
        RECT 211.950 673.950 214.050 674.550 ;
        RECT 227.700 673.800 231.900 674.700 ;
        RECT 245.700 673.800 249.900 674.700 ;
        RECT 184.800 666.000 186.600 672.600 ;
        RECT 200.700 666.000 202.500 672.600 ;
        RECT 205.200 666.600 207.000 672.600 ;
        RECT 209.700 666.000 211.500 672.600 ;
        RECT 227.700 666.600 229.500 673.800 ;
        RECT 232.800 666.000 234.600 672.600 ;
        RECT 245.700 666.600 247.500 673.800 ;
        RECT 266.700 672.600 267.600 679.950 ;
        RECT 273.000 675.300 273.900 695.400 ;
        RECT 290.100 689.400 291.900 701.400 ;
        RECT 293.100 691.200 294.900 702.000 ;
        RECT 296.100 695.400 297.900 701.400 ;
        RECT 308.700 695.400 310.500 702.000 ;
        RECT 274.950 688.050 277.050 688.200 ;
        RECT 274.950 687.450 279.000 688.050 ;
        RECT 274.950 686.100 279.450 687.450 ;
        RECT 276.000 685.950 279.450 686.100 ;
        RECT 274.800 679.950 276.900 682.050 ;
        RECT 274.950 678.150 276.750 679.950 ;
        RECT 278.550 675.900 279.450 685.950 ;
        RECT 280.950 684.450 283.050 685.050 ;
        RECT 286.950 684.450 289.050 685.050 ;
        RECT 280.950 683.550 289.050 684.450 ;
        RECT 280.950 682.950 283.050 683.550 ;
        RECT 286.950 682.950 289.050 683.550 ;
        RECT 290.100 682.050 291.300 689.400 ;
        RECT 296.700 688.500 297.900 695.400 ;
        RECT 309.000 692.100 310.800 693.900 ;
        RECT 311.700 690.900 313.500 701.400 ;
        RECT 292.200 687.600 297.900 688.500 ;
        RECT 311.100 689.400 313.500 690.900 ;
        RECT 316.800 689.400 318.600 702.000 ;
        RECT 320.700 695.400 322.500 702.000 ;
        RECT 323.700 695.400 325.500 701.400 ;
        RECT 327.000 695.400 328.800 702.000 ;
        RECT 330.000 695.400 331.800 701.400 ;
        RECT 333.000 695.400 334.800 702.000 ;
        RECT 336.000 695.400 337.800 701.400 ;
        RECT 339.000 695.400 340.800 702.000 ;
        RECT 342.000 698.400 343.800 701.400 ;
        RECT 345.000 698.400 346.800 701.400 ;
        RECT 348.000 698.400 349.800 701.400 ;
        RECT 341.700 696.300 343.800 698.400 ;
        RECT 344.700 696.300 346.800 698.400 ;
        RECT 347.700 696.300 349.800 698.400 ;
        RECT 351.000 695.400 352.800 701.400 ;
        RECT 354.000 695.400 355.800 702.000 ;
        RECT 292.200 686.700 294.000 687.600 ;
        RECT 290.100 679.950 292.200 682.050 ;
        RECT 268.500 674.400 276.900 675.300 ;
        RECT 268.500 673.500 270.300 674.400 ;
        RECT 250.800 666.000 252.600 672.600 ;
        RECT 266.700 670.800 269.400 672.600 ;
        RECT 267.600 666.600 269.400 670.800 ;
        RECT 270.600 666.000 272.400 672.600 ;
        RECT 275.100 666.600 276.900 674.400 ;
        RECT 277.950 673.800 280.050 675.900 ;
        RECT 290.100 672.600 291.300 679.950 ;
        RECT 293.100 675.300 294.000 686.700 ;
        RECT 303.000 684.450 307.050 685.050 ;
        RECT 295.800 682.050 297.600 683.850 ;
        RECT 295.500 679.950 297.600 682.050 ;
        RECT 302.550 682.950 307.050 684.450 ;
        RECT 302.550 678.450 303.450 682.950 ;
        RECT 311.100 682.050 312.300 689.400 ;
        RECT 324.000 685.050 325.500 695.400 ;
        RECT 330.000 694.500 331.200 695.400 ;
        RECT 317.100 682.050 318.900 683.850 ;
        RECT 323.100 682.950 325.500 685.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 302.550 678.000 306.450 678.450 ;
        RECT 308.100 678.150 309.900 679.950 ;
        RECT 302.550 677.550 307.050 678.000 ;
        RECT 292.200 674.400 294.000 675.300 ;
        RECT 292.200 673.500 297.900 674.400 ;
        RECT 304.950 673.950 307.050 677.550 ;
        RECT 311.100 675.600 312.300 679.950 ;
        RECT 314.100 678.150 315.900 679.950 ;
        RECT 308.700 674.700 312.300 675.600 ;
        RECT 290.100 666.600 291.900 672.600 ;
        RECT 293.100 666.000 294.900 672.600 ;
        RECT 296.700 669.600 297.900 673.500 ;
        RECT 308.700 672.600 309.900 674.700 ;
        RECT 296.100 666.600 297.900 669.600 ;
        RECT 308.100 666.600 309.900 672.600 ;
        RECT 311.100 671.700 318.900 673.050 ;
        RECT 311.100 666.600 312.900 671.700 ;
        RECT 314.100 666.000 315.900 670.800 ;
        RECT 317.100 666.600 318.900 671.700 ;
        RECT 324.000 669.600 325.500 682.950 ;
        RECT 320.700 666.000 322.500 669.600 ;
        RECT 323.700 666.600 325.500 669.600 ;
        RECT 327.300 693.600 331.200 694.500 ;
        RECT 327.300 690.300 328.200 693.600 ;
        RECT 332.100 692.400 333.900 693.000 ;
        RECT 336.600 692.400 337.800 695.400 ;
        RECT 344.700 694.500 346.800 695.400 ;
        RECT 338.700 693.300 346.800 694.500 ;
        RECT 338.700 692.700 340.500 693.300 ;
        RECT 332.100 691.200 337.800 692.400 ;
        RECT 350.100 691.500 352.800 695.400 ;
        RECT 357.000 693.900 358.800 701.400 ;
        RECT 360.900 695.400 362.700 702.000 ;
        RECT 363.900 695.400 365.700 701.400 ;
        RECT 366.900 698.400 368.700 701.400 ;
        RECT 369.900 698.400 371.700 701.400 ;
        RECT 366.600 696.300 368.700 698.400 ;
        RECT 369.600 696.300 371.700 698.400 ;
        RECT 373.500 695.400 375.300 702.000 ;
        RECT 355.500 691.800 358.800 693.900 ;
        RECT 364.200 693.300 366.300 695.400 ;
        RECT 376.500 692.400 378.300 701.400 ;
        RECT 379.500 695.400 381.300 702.000 ;
        RECT 382.500 696.300 384.300 701.400 ;
        RECT 382.500 695.400 384.600 696.300 ;
        RECT 385.500 695.400 387.300 702.000 ;
        RECT 383.700 694.500 384.600 695.400 ;
        RECT 383.700 693.600 387.300 694.500 ;
        RECT 381.000 692.400 382.800 692.700 ;
        RECT 341.700 690.300 343.800 691.500 ;
        RECT 327.300 689.400 343.800 690.300 ;
        RECT 347.100 690.600 349.200 691.500 ;
        RECT 363.600 691.200 382.800 692.400 ;
        RECT 363.600 690.600 364.800 691.200 ;
        RECT 381.000 690.900 382.800 691.200 ;
        RECT 347.100 689.400 364.800 690.600 ;
        RECT 367.500 689.700 369.600 690.300 ;
        RECT 377.700 689.700 379.500 690.300 ;
        RECT 327.300 672.600 328.200 689.400 ;
        RECT 367.500 688.500 379.500 689.700 ;
        RECT 329.100 687.300 364.800 688.500 ;
        RECT 367.500 688.200 369.600 688.500 ;
        RECT 329.100 686.700 330.900 687.300 ;
        RECT 363.600 686.700 364.800 687.300 ;
        RECT 332.100 682.950 334.200 685.050 ;
        RECT 332.700 680.100 334.200 682.950 ;
        RECT 336.300 682.800 341.400 684.600 ;
        RECT 340.500 681.300 341.400 682.800 ;
        RECT 344.100 684.300 345.900 686.100 ;
        RECT 350.100 685.800 352.200 686.100 ;
        RECT 363.600 685.800 377.100 686.700 ;
        RECT 344.100 683.100 345.000 684.300 ;
        RECT 350.100 684.000 354.000 685.800 ;
        RECT 355.500 684.300 357.600 685.200 ;
        RECT 375.300 685.050 377.100 685.800 ;
        RECT 355.500 683.100 366.600 684.300 ;
        RECT 375.300 683.250 379.200 685.050 ;
        RECT 344.100 682.200 357.600 683.100 ;
        RECT 364.800 682.500 366.600 683.100 ;
        RECT 377.100 682.950 379.200 683.250 ;
        RECT 383.100 682.950 385.200 685.050 ;
        RECT 383.100 681.300 384.900 682.950 ;
        RECT 340.500 680.100 384.900 681.300 ;
        RECT 332.700 678.600 339.300 680.100 ;
        RECT 329.100 675.900 336.900 677.700 ;
        RECT 337.800 677.100 354.900 678.600 ;
        RECT 352.800 676.500 354.900 677.100 ;
        RECT 359.100 678.000 361.200 679.050 ;
        RECT 359.100 677.100 364.200 678.000 ;
        RECT 367.800 677.400 369.600 679.200 ;
        RECT 386.100 677.400 387.300 693.600 ;
        RECT 401.400 689.400 403.200 702.000 ;
        RECT 406.500 690.900 408.300 701.400 ;
        RECT 409.500 695.400 411.300 702.000 ;
        RECT 418.950 696.450 421.050 697.050 ;
        RECT 413.550 695.550 421.050 696.450 ;
        RECT 409.200 692.100 411.000 693.900 ;
        RECT 413.550 691.050 414.450 695.550 ;
        RECT 418.950 694.950 421.050 695.550 ;
        RECT 422.100 695.400 423.900 702.000 ;
        RECT 425.100 695.400 426.900 701.400 ;
        RECT 428.100 695.400 429.900 702.000 ;
        RECT 431.700 695.400 433.500 702.000 ;
        RECT 434.700 696.300 436.500 701.400 ;
        RECT 434.400 695.400 436.500 696.300 ;
        RECT 437.700 695.400 439.500 702.000 ;
        RECT 406.500 689.400 408.900 690.900 ;
        RECT 401.100 682.050 402.900 683.850 ;
        RECT 407.700 682.050 408.900 689.400 ;
        RECT 409.950 689.550 414.450 691.050 ;
        RECT 409.950 688.950 414.000 689.550 ;
        RECT 420.000 687.450 424.050 688.050 ;
        RECT 419.550 685.950 424.050 687.450 ;
        RECT 419.550 684.450 420.450 685.950 ;
        RECT 416.550 683.550 420.450 684.450 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 404.100 678.150 405.900 679.950 ;
        RECT 359.100 676.950 361.200 677.100 ;
        RECT 335.400 672.600 336.900 675.900 ;
        RECT 353.100 674.700 354.900 676.500 ;
        RECT 362.400 676.200 364.200 677.100 ;
        RECT 368.700 674.400 369.600 677.400 ;
        RECT 370.500 676.200 387.300 677.400 ;
        RECT 370.500 675.300 372.600 676.200 ;
        RECT 381.300 674.700 383.100 675.300 ;
        RECT 341.100 672.600 347.700 674.400 ;
        RECT 362.400 673.200 369.600 674.400 ;
        RECT 374.700 673.500 383.100 674.700 ;
        RECT 362.400 672.600 363.300 673.200 ;
        RECT 365.400 672.600 367.200 673.200 ;
        RECT 374.700 672.600 376.200 673.500 ;
        RECT 386.100 672.600 387.300 676.200 ;
        RECT 407.700 675.600 408.900 679.950 ;
        RECT 410.100 678.150 411.900 679.950 ;
        RECT 416.550 679.050 417.450 683.550 ;
        RECT 425.700 682.050 426.900 695.400 ;
        RECT 434.400 694.500 435.300 695.400 ;
        RECT 431.700 693.600 435.300 694.500 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 416.550 677.550 421.050 679.050 ;
        RECT 422.100 678.150 423.900 679.950 ;
        RECT 417.000 676.950 421.050 677.550 ;
        RECT 407.700 674.700 411.300 675.600 ;
        RECT 425.700 674.700 426.900 679.950 ;
        RECT 427.950 678.150 429.750 679.950 ;
        RECT 327.300 666.600 329.100 672.600 ;
        RECT 332.700 666.000 334.500 672.600 ;
        RECT 335.400 671.400 339.600 672.600 ;
        RECT 337.800 666.600 339.600 671.400 ;
        RECT 341.700 669.600 343.800 671.700 ;
        RECT 344.700 669.600 346.800 671.700 ;
        RECT 347.700 669.600 349.800 671.700 ;
        RECT 350.700 669.600 352.800 671.700 ;
        RECT 356.100 670.500 358.800 672.600 ;
        RECT 360.600 671.400 363.300 672.600 ;
        RECT 360.600 670.500 362.400 671.400 ;
        RECT 342.000 666.600 343.800 669.600 ;
        RECT 345.000 666.600 346.800 669.600 ;
        RECT 348.000 666.600 349.800 669.600 ;
        RECT 351.000 666.600 352.800 669.600 ;
        RECT 354.000 666.000 355.800 669.600 ;
        RECT 357.000 666.600 358.800 670.500 ;
        RECT 364.200 669.600 366.300 671.700 ;
        RECT 367.200 669.600 369.300 671.700 ;
        RECT 370.200 669.600 372.300 671.700 ;
        RECT 361.500 666.000 363.300 669.600 ;
        RECT 364.500 666.600 366.300 669.600 ;
        RECT 367.500 666.600 369.300 669.600 ;
        RECT 370.500 666.600 372.300 669.600 ;
        RECT 374.700 666.600 376.500 672.600 ;
        RECT 380.100 666.000 381.900 672.600 ;
        RECT 385.500 666.600 387.300 672.600 ;
        RECT 401.100 671.700 408.900 673.050 ;
        RECT 401.100 666.600 402.900 671.700 ;
        RECT 404.100 666.000 405.900 670.800 ;
        RECT 407.100 666.600 408.900 671.700 ;
        RECT 410.100 672.600 411.300 674.700 ;
        RECT 422.700 673.800 426.900 674.700 ;
        RECT 431.700 677.400 432.900 693.600 ;
        RECT 436.200 692.400 438.000 692.700 ;
        RECT 440.700 692.400 442.500 701.400 ;
        RECT 443.700 695.400 445.500 702.000 ;
        RECT 447.300 698.400 449.100 701.400 ;
        RECT 450.300 698.400 452.100 701.400 ;
        RECT 447.300 696.300 449.400 698.400 ;
        RECT 450.300 696.300 452.400 698.400 ;
        RECT 453.300 695.400 455.100 701.400 ;
        RECT 456.300 695.400 458.100 702.000 ;
        RECT 452.700 693.300 454.800 695.400 ;
        RECT 460.200 693.900 462.000 701.400 ;
        RECT 463.200 695.400 465.000 702.000 ;
        RECT 466.200 695.400 468.000 701.400 ;
        RECT 469.200 698.400 471.000 701.400 ;
        RECT 472.200 698.400 474.000 701.400 ;
        RECT 475.200 698.400 477.000 701.400 ;
        RECT 469.200 696.300 471.300 698.400 ;
        RECT 472.200 696.300 474.300 698.400 ;
        RECT 475.200 696.300 477.300 698.400 ;
        RECT 478.200 695.400 480.000 702.000 ;
        RECT 481.200 695.400 483.000 701.400 ;
        RECT 484.200 695.400 486.000 702.000 ;
        RECT 487.200 695.400 489.000 701.400 ;
        RECT 490.200 695.400 492.000 702.000 ;
        RECT 493.500 695.400 495.300 701.400 ;
        RECT 496.500 695.400 498.300 702.000 ;
        RECT 436.200 691.200 455.400 692.400 ;
        RECT 460.200 691.800 463.500 693.900 ;
        RECT 466.200 691.500 468.900 695.400 ;
        RECT 472.200 694.500 474.300 695.400 ;
        RECT 472.200 693.300 480.300 694.500 ;
        RECT 478.500 692.700 480.300 693.300 ;
        RECT 481.200 692.400 482.400 695.400 ;
        RECT 487.800 694.500 489.000 695.400 ;
        RECT 487.800 693.600 491.700 694.500 ;
        RECT 485.100 692.400 486.900 693.000 ;
        RECT 436.200 690.900 438.000 691.200 ;
        RECT 454.200 690.600 455.400 691.200 ;
        RECT 469.800 690.600 471.900 691.500 ;
        RECT 439.500 689.700 441.300 690.300 ;
        RECT 449.400 689.700 451.500 690.300 ;
        RECT 439.500 688.500 451.500 689.700 ;
        RECT 454.200 689.400 471.900 690.600 ;
        RECT 475.200 690.300 477.300 691.500 ;
        RECT 481.200 691.200 486.900 692.400 ;
        RECT 490.800 690.300 491.700 693.600 ;
        RECT 475.200 689.400 491.700 690.300 ;
        RECT 449.400 688.200 451.500 688.500 ;
        RECT 454.200 687.300 489.900 688.500 ;
        RECT 454.200 686.700 455.400 687.300 ;
        RECT 488.100 686.700 489.900 687.300 ;
        RECT 441.900 685.800 455.400 686.700 ;
        RECT 466.800 685.800 468.900 686.100 ;
        RECT 441.900 685.050 443.700 685.800 ;
        RECT 433.800 682.950 435.900 685.050 ;
        RECT 439.800 683.250 443.700 685.050 ;
        RECT 461.400 684.300 463.500 685.200 ;
        RECT 439.800 682.950 441.900 683.250 ;
        RECT 452.400 683.100 463.500 684.300 ;
        RECT 465.000 684.000 468.900 685.800 ;
        RECT 473.100 684.300 474.900 686.100 ;
        RECT 474.000 683.100 474.900 684.300 ;
        RECT 434.100 681.300 435.900 682.950 ;
        RECT 452.400 682.500 454.200 683.100 ;
        RECT 461.400 682.200 474.900 683.100 ;
        RECT 477.600 682.800 482.700 684.600 ;
        RECT 484.800 682.950 486.900 685.050 ;
        RECT 477.600 681.300 478.500 682.800 ;
        RECT 434.100 680.100 478.500 681.300 ;
        RECT 484.800 680.100 486.300 682.950 ;
        RECT 449.400 677.400 451.200 679.200 ;
        RECT 457.800 678.000 459.900 679.050 ;
        RECT 479.700 678.600 486.300 680.100 ;
        RECT 431.700 676.200 448.500 677.400 ;
        RECT 410.100 666.600 411.900 672.600 ;
        RECT 422.700 666.600 424.500 673.800 ;
        RECT 431.700 672.600 432.900 676.200 ;
        RECT 446.400 675.300 448.500 676.200 ;
        RECT 435.900 674.700 437.700 675.300 ;
        RECT 435.900 673.500 444.300 674.700 ;
        RECT 442.800 672.600 444.300 673.500 ;
        RECT 449.400 674.400 450.300 677.400 ;
        RECT 454.800 677.100 459.900 678.000 ;
        RECT 454.800 676.200 456.600 677.100 ;
        RECT 457.800 676.950 459.900 677.100 ;
        RECT 464.100 677.100 481.200 678.600 ;
        RECT 464.100 676.500 466.200 677.100 ;
        RECT 464.100 674.700 465.900 676.500 ;
        RECT 482.100 675.900 489.900 677.700 ;
        RECT 449.400 673.200 456.600 674.400 ;
        RECT 451.800 672.600 453.600 673.200 ;
        RECT 455.700 672.600 456.600 673.200 ;
        RECT 471.300 672.600 477.900 674.400 ;
        RECT 482.100 672.600 483.600 675.900 ;
        RECT 490.800 672.600 491.700 689.400 ;
        RECT 427.800 666.000 429.600 672.600 ;
        RECT 431.700 666.600 433.500 672.600 ;
        RECT 437.100 666.000 438.900 672.600 ;
        RECT 442.500 666.600 444.300 672.600 ;
        RECT 446.700 669.600 448.800 671.700 ;
        RECT 449.700 669.600 451.800 671.700 ;
        RECT 452.700 669.600 454.800 671.700 ;
        RECT 455.700 671.400 458.400 672.600 ;
        RECT 456.600 670.500 458.400 671.400 ;
        RECT 460.200 670.500 462.900 672.600 ;
        RECT 446.700 666.600 448.500 669.600 ;
        RECT 449.700 666.600 451.500 669.600 ;
        RECT 452.700 666.600 454.500 669.600 ;
        RECT 455.700 666.000 457.500 669.600 ;
        RECT 460.200 666.600 462.000 670.500 ;
        RECT 466.200 669.600 468.300 671.700 ;
        RECT 469.200 669.600 471.300 671.700 ;
        RECT 472.200 669.600 474.300 671.700 ;
        RECT 475.200 669.600 477.300 671.700 ;
        RECT 479.400 671.400 483.600 672.600 ;
        RECT 463.200 666.000 465.000 669.600 ;
        RECT 466.200 666.600 468.000 669.600 ;
        RECT 469.200 666.600 471.000 669.600 ;
        RECT 472.200 666.600 474.000 669.600 ;
        RECT 475.200 666.600 477.000 669.600 ;
        RECT 479.400 666.600 481.200 671.400 ;
        RECT 484.500 666.000 486.300 672.600 ;
        RECT 489.900 666.600 491.700 672.600 ;
        RECT 493.500 685.050 495.000 695.400 ;
        RECT 512.100 689.400 513.900 702.000 ;
        RECT 515.100 688.500 516.900 701.400 ;
        RECT 518.100 689.400 519.900 702.000 ;
        RECT 521.100 688.500 522.900 701.400 ;
        RECT 524.100 689.400 525.900 702.000 ;
        RECT 527.100 688.500 528.900 701.400 ;
        RECT 530.100 689.400 531.900 702.000 ;
        RECT 533.100 688.500 534.900 701.400 ;
        RECT 536.100 689.400 537.900 702.000 ;
        RECT 551.100 689.400 552.900 702.000 ;
        RECT 554.100 688.500 555.900 701.400 ;
        RECT 557.100 689.400 558.900 702.000 ;
        RECT 560.100 688.500 561.900 701.400 ;
        RECT 563.100 689.400 564.900 702.000 ;
        RECT 566.100 688.500 567.900 701.400 ;
        RECT 569.100 689.400 570.900 702.000 ;
        RECT 572.100 688.500 573.900 701.400 ;
        RECT 575.100 689.400 576.900 702.000 ;
        RECT 587.100 695.400 588.900 702.000 ;
        RECT 590.100 695.400 591.900 701.400 ;
        RECT 514.050 687.300 516.900 688.500 ;
        RECT 519.000 687.300 522.900 688.500 ;
        RECT 525.000 687.300 528.900 688.500 ;
        RECT 531.000 687.300 534.900 688.500 ;
        RECT 553.050 687.300 555.900 688.500 ;
        RECT 558.000 687.300 561.900 688.500 ;
        RECT 564.000 687.300 567.900 688.500 ;
        RECT 570.000 687.300 573.900 688.500 ;
        RECT 493.500 682.950 495.900 685.050 ;
        RECT 493.500 669.600 495.000 682.950 ;
        RECT 514.050 682.050 515.100 687.300 ;
        RECT 514.050 679.950 517.200 682.050 ;
        RECT 514.050 674.700 515.100 679.950 ;
        RECT 516.000 676.800 517.800 677.400 ;
        RECT 519.000 676.800 520.200 687.300 ;
        RECT 516.000 675.600 520.200 676.800 ;
        RECT 522.000 676.800 523.800 677.400 ;
        RECT 525.000 676.800 526.200 687.300 ;
        RECT 522.000 675.600 526.200 676.800 ;
        RECT 528.000 676.800 529.800 677.400 ;
        RECT 531.000 676.800 532.200 687.300 ;
        RECT 553.050 682.050 554.100 687.300 ;
        RECT 533.100 679.950 535.200 682.050 ;
        RECT 533.400 678.150 535.200 679.950 ;
        RECT 553.050 679.950 556.200 682.050 ;
        RECT 528.000 675.600 532.200 676.800 ;
        RECT 519.000 674.700 520.200 675.600 ;
        RECT 525.000 674.700 526.200 675.600 ;
        RECT 531.000 674.700 532.200 675.600 ;
        RECT 553.050 674.700 554.100 679.950 ;
        RECT 555.000 676.800 556.800 677.400 ;
        RECT 558.000 676.800 559.200 687.300 ;
        RECT 555.000 675.600 559.200 676.800 ;
        RECT 561.000 676.800 562.800 677.400 ;
        RECT 564.000 676.800 565.200 687.300 ;
        RECT 561.000 675.600 565.200 676.800 ;
        RECT 567.000 676.800 568.800 677.400 ;
        RECT 570.000 676.800 571.200 687.300 ;
        RECT 587.100 682.050 588.900 683.850 ;
        RECT 590.100 682.050 591.300 695.400 ;
        RECT 605.400 689.400 607.200 702.000 ;
        RECT 610.500 690.900 612.300 701.400 ;
        RECT 613.500 695.400 615.300 702.000 ;
        RECT 617.700 695.400 619.500 702.000 ;
        RECT 620.700 695.400 622.500 701.400 ;
        RECT 624.000 695.400 625.800 702.000 ;
        RECT 627.000 695.400 628.800 701.400 ;
        RECT 630.000 695.400 631.800 702.000 ;
        RECT 633.000 695.400 634.800 701.400 ;
        RECT 636.000 695.400 637.800 702.000 ;
        RECT 639.000 698.400 640.800 701.400 ;
        RECT 642.000 698.400 643.800 701.400 ;
        RECT 645.000 698.400 646.800 701.400 ;
        RECT 638.700 696.300 640.800 698.400 ;
        RECT 641.700 696.300 643.800 698.400 ;
        RECT 644.700 696.300 646.800 698.400 ;
        RECT 648.000 695.400 649.800 701.400 ;
        RECT 651.000 695.400 652.800 702.000 ;
        RECT 613.200 692.100 615.000 693.900 ;
        RECT 610.500 689.400 612.900 690.900 ;
        RECT 604.950 687.450 607.050 688.050 ;
        RECT 596.550 686.550 607.050 687.450 ;
        RECT 572.100 679.950 574.200 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 572.400 678.150 574.200 679.950 ;
        RECT 567.000 675.600 571.200 676.800 ;
        RECT 558.000 674.700 559.200 675.600 ;
        RECT 564.000 674.700 565.200 675.600 ;
        RECT 570.000 674.700 571.200 675.600 ;
        RECT 514.050 673.500 516.900 674.700 ;
        RECT 519.000 673.500 522.900 674.700 ;
        RECT 525.000 673.500 528.900 674.700 ;
        RECT 531.000 673.500 534.900 674.700 ;
        RECT 553.050 673.500 555.900 674.700 ;
        RECT 558.000 673.500 561.900 674.700 ;
        RECT 564.000 673.500 567.900 674.700 ;
        RECT 570.000 673.500 573.900 674.700 ;
        RECT 493.500 666.600 495.300 669.600 ;
        RECT 496.500 666.000 498.300 669.600 ;
        RECT 512.100 666.000 513.900 672.600 ;
        RECT 515.100 666.600 516.900 673.500 ;
        RECT 518.100 666.000 519.900 672.600 ;
        RECT 521.100 666.600 522.900 673.500 ;
        RECT 524.100 666.000 525.900 672.600 ;
        RECT 527.100 666.600 528.900 673.500 ;
        RECT 530.100 666.000 531.900 672.600 ;
        RECT 533.100 666.600 534.900 673.500 ;
        RECT 536.100 666.000 537.900 672.600 ;
        RECT 551.100 666.000 552.900 672.600 ;
        RECT 554.100 666.600 555.900 673.500 ;
        RECT 557.100 666.000 558.900 672.600 ;
        RECT 560.100 666.600 561.900 673.500 ;
        RECT 563.100 666.000 564.900 672.600 ;
        RECT 566.100 666.600 567.900 673.500 ;
        RECT 569.100 666.000 570.900 672.600 ;
        RECT 572.100 666.600 573.900 673.500 ;
        RECT 575.100 666.000 576.900 672.600 ;
        RECT 577.950 672.450 580.050 673.050 ;
        RECT 586.950 672.450 589.050 673.050 ;
        RECT 577.950 671.550 589.050 672.450 ;
        RECT 577.950 670.950 580.050 671.550 ;
        RECT 586.950 670.950 589.050 671.550 ;
        RECT 590.100 669.600 591.300 679.950 ;
        RECT 596.550 675.900 597.450 686.550 ;
        RECT 604.950 685.950 607.050 686.550 ;
        RECT 600.000 684.450 604.050 685.050 ;
        RECT 599.550 682.950 604.050 684.450 ;
        RECT 599.550 679.050 600.450 682.950 ;
        RECT 605.100 682.050 606.900 683.850 ;
        RECT 611.700 682.050 612.900 689.400 ;
        RECT 621.000 685.050 622.500 695.400 ;
        RECT 627.000 694.500 628.200 695.400 ;
        RECT 620.100 682.950 622.500 685.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 607.950 679.950 610.050 682.050 ;
        RECT 610.950 679.950 613.050 682.050 ;
        RECT 613.950 679.950 616.050 682.050 ;
        RECT 599.550 677.550 604.050 679.050 ;
        RECT 608.100 678.150 609.900 679.950 ;
        RECT 600.000 676.950 604.050 677.550 ;
        RECT 595.950 673.800 598.050 675.900 ;
        RECT 611.700 675.600 612.900 679.950 ;
        RECT 614.100 678.150 615.900 679.950 ;
        RECT 611.700 674.700 615.300 675.600 ;
        RECT 605.100 671.700 612.900 673.050 ;
        RECT 587.100 666.000 588.900 669.600 ;
        RECT 590.100 666.600 591.900 669.600 ;
        RECT 605.100 666.600 606.900 671.700 ;
        RECT 608.100 666.000 609.900 670.800 ;
        RECT 611.100 666.600 612.900 671.700 ;
        RECT 614.100 672.600 615.300 674.700 ;
        RECT 614.100 666.600 615.900 672.600 ;
        RECT 621.000 669.600 622.500 682.950 ;
        RECT 617.700 666.000 619.500 669.600 ;
        RECT 620.700 666.600 622.500 669.600 ;
        RECT 624.300 693.600 628.200 694.500 ;
        RECT 624.300 690.300 625.200 693.600 ;
        RECT 629.100 692.400 630.900 693.000 ;
        RECT 633.600 692.400 634.800 695.400 ;
        RECT 641.700 694.500 643.800 695.400 ;
        RECT 635.700 693.300 643.800 694.500 ;
        RECT 635.700 692.700 637.500 693.300 ;
        RECT 629.100 691.200 634.800 692.400 ;
        RECT 647.100 691.500 649.800 695.400 ;
        RECT 654.000 693.900 655.800 701.400 ;
        RECT 657.900 695.400 659.700 702.000 ;
        RECT 660.900 695.400 662.700 701.400 ;
        RECT 663.900 698.400 665.700 701.400 ;
        RECT 666.900 698.400 668.700 701.400 ;
        RECT 663.600 696.300 665.700 698.400 ;
        RECT 666.600 696.300 668.700 698.400 ;
        RECT 670.500 695.400 672.300 702.000 ;
        RECT 652.500 691.800 655.800 693.900 ;
        RECT 661.200 693.300 663.300 695.400 ;
        RECT 673.500 692.400 675.300 701.400 ;
        RECT 676.500 695.400 678.300 702.000 ;
        RECT 679.500 696.300 681.300 701.400 ;
        RECT 679.500 695.400 681.600 696.300 ;
        RECT 682.500 695.400 684.300 702.000 ;
        RECT 686.700 695.400 688.500 702.000 ;
        RECT 689.700 696.300 691.500 701.400 ;
        RECT 689.400 695.400 691.500 696.300 ;
        RECT 692.700 695.400 694.500 702.000 ;
        RECT 680.700 694.500 681.600 695.400 ;
        RECT 689.400 694.500 690.300 695.400 ;
        RECT 680.700 693.600 684.300 694.500 ;
        RECT 678.000 692.400 679.800 692.700 ;
        RECT 638.700 690.300 640.800 691.500 ;
        RECT 624.300 689.400 640.800 690.300 ;
        RECT 644.100 690.600 646.200 691.500 ;
        RECT 660.600 691.200 679.800 692.400 ;
        RECT 660.600 690.600 661.800 691.200 ;
        RECT 678.000 690.900 679.800 691.200 ;
        RECT 644.100 689.400 661.800 690.600 ;
        RECT 664.500 689.700 666.600 690.300 ;
        RECT 674.700 689.700 676.500 690.300 ;
        RECT 624.300 672.600 625.200 689.400 ;
        RECT 664.500 688.500 676.500 689.700 ;
        RECT 626.100 687.300 661.800 688.500 ;
        RECT 664.500 688.200 666.600 688.500 ;
        RECT 626.100 686.700 627.900 687.300 ;
        RECT 660.600 686.700 661.800 687.300 ;
        RECT 629.100 682.950 631.200 685.050 ;
        RECT 629.700 680.100 631.200 682.950 ;
        RECT 633.300 682.800 638.400 684.600 ;
        RECT 637.500 681.300 638.400 682.800 ;
        RECT 641.100 684.300 642.900 686.100 ;
        RECT 647.100 685.800 649.200 686.100 ;
        RECT 660.600 685.800 674.100 686.700 ;
        RECT 641.100 683.100 642.000 684.300 ;
        RECT 647.100 684.000 651.000 685.800 ;
        RECT 652.500 684.300 654.600 685.200 ;
        RECT 672.300 685.050 674.100 685.800 ;
        RECT 652.500 683.100 663.600 684.300 ;
        RECT 672.300 683.250 676.200 685.050 ;
        RECT 641.100 682.200 654.600 683.100 ;
        RECT 661.800 682.500 663.600 683.100 ;
        RECT 674.100 682.950 676.200 683.250 ;
        RECT 680.100 682.950 682.200 685.050 ;
        RECT 680.100 681.300 681.900 682.950 ;
        RECT 637.500 680.100 681.900 681.300 ;
        RECT 629.700 678.600 636.300 680.100 ;
        RECT 626.100 675.900 633.900 677.700 ;
        RECT 634.800 677.100 651.900 678.600 ;
        RECT 649.800 676.500 651.900 677.100 ;
        RECT 656.100 678.000 658.200 679.050 ;
        RECT 656.100 677.100 661.200 678.000 ;
        RECT 664.800 677.400 666.600 679.200 ;
        RECT 683.100 677.400 684.300 693.600 ;
        RECT 656.100 676.950 658.200 677.100 ;
        RECT 632.400 672.600 633.900 675.900 ;
        RECT 650.100 674.700 651.900 676.500 ;
        RECT 659.400 676.200 661.200 677.100 ;
        RECT 665.700 674.400 666.600 677.400 ;
        RECT 667.500 676.200 684.300 677.400 ;
        RECT 667.500 675.300 669.600 676.200 ;
        RECT 678.300 674.700 680.100 675.300 ;
        RECT 638.100 672.600 644.700 674.400 ;
        RECT 659.400 673.200 666.600 674.400 ;
        RECT 671.700 673.500 680.100 674.700 ;
        RECT 659.400 672.600 660.300 673.200 ;
        RECT 662.400 672.600 664.200 673.200 ;
        RECT 671.700 672.600 673.200 673.500 ;
        RECT 683.100 672.600 684.300 676.200 ;
        RECT 624.300 666.600 626.100 672.600 ;
        RECT 629.700 666.000 631.500 672.600 ;
        RECT 632.400 671.400 636.600 672.600 ;
        RECT 634.800 666.600 636.600 671.400 ;
        RECT 638.700 669.600 640.800 671.700 ;
        RECT 641.700 669.600 643.800 671.700 ;
        RECT 644.700 669.600 646.800 671.700 ;
        RECT 647.700 669.600 649.800 671.700 ;
        RECT 653.100 670.500 655.800 672.600 ;
        RECT 657.600 671.400 660.300 672.600 ;
        RECT 657.600 670.500 659.400 671.400 ;
        RECT 639.000 666.600 640.800 669.600 ;
        RECT 642.000 666.600 643.800 669.600 ;
        RECT 645.000 666.600 646.800 669.600 ;
        RECT 648.000 666.600 649.800 669.600 ;
        RECT 651.000 666.000 652.800 669.600 ;
        RECT 654.000 666.600 655.800 670.500 ;
        RECT 661.200 669.600 663.300 671.700 ;
        RECT 664.200 669.600 666.300 671.700 ;
        RECT 667.200 669.600 669.300 671.700 ;
        RECT 658.500 666.000 660.300 669.600 ;
        RECT 661.500 666.600 663.300 669.600 ;
        RECT 664.500 666.600 666.300 669.600 ;
        RECT 667.500 666.600 669.300 669.600 ;
        RECT 671.700 666.600 673.500 672.600 ;
        RECT 677.100 666.000 678.900 672.600 ;
        RECT 682.500 666.600 684.300 672.600 ;
        RECT 686.700 693.600 690.300 694.500 ;
        RECT 686.700 677.400 687.900 693.600 ;
        RECT 691.200 692.400 693.000 692.700 ;
        RECT 695.700 692.400 697.500 701.400 ;
        RECT 698.700 695.400 700.500 702.000 ;
        RECT 702.300 698.400 704.100 701.400 ;
        RECT 705.300 698.400 707.100 701.400 ;
        RECT 702.300 696.300 704.400 698.400 ;
        RECT 705.300 696.300 707.400 698.400 ;
        RECT 708.300 695.400 710.100 701.400 ;
        RECT 711.300 695.400 713.100 702.000 ;
        RECT 707.700 693.300 709.800 695.400 ;
        RECT 715.200 693.900 717.000 701.400 ;
        RECT 718.200 695.400 720.000 702.000 ;
        RECT 721.200 695.400 723.000 701.400 ;
        RECT 724.200 698.400 726.000 701.400 ;
        RECT 727.200 698.400 729.000 701.400 ;
        RECT 730.200 698.400 732.000 701.400 ;
        RECT 724.200 696.300 726.300 698.400 ;
        RECT 727.200 696.300 729.300 698.400 ;
        RECT 730.200 696.300 732.300 698.400 ;
        RECT 733.200 695.400 735.000 702.000 ;
        RECT 736.200 695.400 738.000 701.400 ;
        RECT 739.200 695.400 741.000 702.000 ;
        RECT 742.200 695.400 744.000 701.400 ;
        RECT 745.200 695.400 747.000 702.000 ;
        RECT 748.500 695.400 750.300 701.400 ;
        RECT 751.500 695.400 753.300 702.000 ;
        RECT 691.200 691.200 710.400 692.400 ;
        RECT 715.200 691.800 718.500 693.900 ;
        RECT 721.200 691.500 723.900 695.400 ;
        RECT 727.200 694.500 729.300 695.400 ;
        RECT 727.200 693.300 735.300 694.500 ;
        RECT 733.500 692.700 735.300 693.300 ;
        RECT 736.200 692.400 737.400 695.400 ;
        RECT 742.800 694.500 744.000 695.400 ;
        RECT 742.800 693.600 746.700 694.500 ;
        RECT 740.100 692.400 741.900 693.000 ;
        RECT 691.200 690.900 693.000 691.200 ;
        RECT 709.200 690.600 710.400 691.200 ;
        RECT 724.800 690.600 726.900 691.500 ;
        RECT 694.500 689.700 696.300 690.300 ;
        RECT 704.400 689.700 706.500 690.300 ;
        RECT 694.500 688.500 706.500 689.700 ;
        RECT 709.200 689.400 726.900 690.600 ;
        RECT 730.200 690.300 732.300 691.500 ;
        RECT 736.200 691.200 741.900 692.400 ;
        RECT 745.800 690.300 746.700 693.600 ;
        RECT 730.200 689.400 746.700 690.300 ;
        RECT 704.400 688.200 706.500 688.500 ;
        RECT 709.200 687.300 744.900 688.500 ;
        RECT 709.200 686.700 710.400 687.300 ;
        RECT 743.100 686.700 744.900 687.300 ;
        RECT 696.900 685.800 710.400 686.700 ;
        RECT 721.800 685.800 723.900 686.100 ;
        RECT 696.900 685.050 698.700 685.800 ;
        RECT 688.800 682.950 690.900 685.050 ;
        RECT 694.800 683.250 698.700 685.050 ;
        RECT 716.400 684.300 718.500 685.200 ;
        RECT 694.800 682.950 696.900 683.250 ;
        RECT 707.400 683.100 718.500 684.300 ;
        RECT 720.000 684.000 723.900 685.800 ;
        RECT 728.100 684.300 729.900 686.100 ;
        RECT 729.000 683.100 729.900 684.300 ;
        RECT 689.100 681.300 690.900 682.950 ;
        RECT 707.400 682.500 709.200 683.100 ;
        RECT 716.400 682.200 729.900 683.100 ;
        RECT 732.600 682.800 737.700 684.600 ;
        RECT 739.800 682.950 741.900 685.050 ;
        RECT 732.600 681.300 733.500 682.800 ;
        RECT 689.100 680.100 733.500 681.300 ;
        RECT 739.800 680.100 741.300 682.950 ;
        RECT 704.400 677.400 706.200 679.200 ;
        RECT 712.800 678.000 714.900 679.050 ;
        RECT 734.700 678.600 741.300 680.100 ;
        RECT 686.700 676.200 703.500 677.400 ;
        RECT 686.700 672.600 687.900 676.200 ;
        RECT 701.400 675.300 703.500 676.200 ;
        RECT 690.900 674.700 692.700 675.300 ;
        RECT 690.900 673.500 699.300 674.700 ;
        RECT 697.800 672.600 699.300 673.500 ;
        RECT 704.400 674.400 705.300 677.400 ;
        RECT 709.800 677.100 714.900 678.000 ;
        RECT 709.800 676.200 711.600 677.100 ;
        RECT 712.800 676.950 714.900 677.100 ;
        RECT 719.100 677.100 736.200 678.600 ;
        RECT 719.100 676.500 721.200 677.100 ;
        RECT 719.100 674.700 720.900 676.500 ;
        RECT 737.100 675.900 744.900 677.700 ;
        RECT 704.400 673.200 711.600 674.400 ;
        RECT 706.800 672.600 708.600 673.200 ;
        RECT 710.700 672.600 711.600 673.200 ;
        RECT 726.300 672.600 732.900 674.400 ;
        RECT 737.100 672.600 738.600 675.900 ;
        RECT 745.800 672.600 746.700 689.400 ;
        RECT 686.700 666.600 688.500 672.600 ;
        RECT 692.100 666.000 693.900 672.600 ;
        RECT 697.500 666.600 699.300 672.600 ;
        RECT 701.700 669.600 703.800 671.700 ;
        RECT 704.700 669.600 706.800 671.700 ;
        RECT 707.700 669.600 709.800 671.700 ;
        RECT 710.700 671.400 713.400 672.600 ;
        RECT 711.600 670.500 713.400 671.400 ;
        RECT 715.200 670.500 717.900 672.600 ;
        RECT 701.700 666.600 703.500 669.600 ;
        RECT 704.700 666.600 706.500 669.600 ;
        RECT 707.700 666.600 709.500 669.600 ;
        RECT 710.700 666.000 712.500 669.600 ;
        RECT 715.200 666.600 717.000 670.500 ;
        RECT 721.200 669.600 723.300 671.700 ;
        RECT 724.200 669.600 726.300 671.700 ;
        RECT 727.200 669.600 729.300 671.700 ;
        RECT 730.200 669.600 732.300 671.700 ;
        RECT 734.400 671.400 738.600 672.600 ;
        RECT 718.200 666.000 720.000 669.600 ;
        RECT 721.200 666.600 723.000 669.600 ;
        RECT 724.200 666.600 726.000 669.600 ;
        RECT 727.200 666.600 729.000 669.600 ;
        RECT 730.200 666.600 732.000 669.600 ;
        RECT 734.400 666.600 736.200 671.400 ;
        RECT 739.500 666.000 741.300 672.600 ;
        RECT 744.900 666.600 746.700 672.600 ;
        RECT 748.500 685.050 750.000 695.400 ;
        RECT 767.100 689.400 768.900 701.400 ;
        RECT 770.100 690.300 771.900 701.400 ;
        RECT 773.100 691.200 774.900 702.000 ;
        RECT 776.100 690.300 777.900 701.400 ;
        RECT 791.100 695.400 792.900 701.400 ;
        RECT 794.100 696.000 795.900 702.000 ;
        RECT 770.100 689.400 777.900 690.300 ;
        RECT 792.000 695.100 792.900 695.400 ;
        RECT 797.100 695.400 798.900 701.400 ;
        RECT 800.100 695.400 801.900 702.000 ;
        RECT 812.100 695.400 813.900 701.400 ;
        RECT 815.100 695.400 816.900 702.000 ;
        RECT 797.100 695.100 798.600 695.400 ;
        RECT 792.000 694.200 798.600 695.100 ;
        RECT 748.500 682.950 750.900 685.050 ;
        RECT 748.500 669.600 750.000 682.950 ;
        RECT 767.400 682.050 768.300 689.400 ;
        RECT 772.950 682.050 774.750 683.850 ;
        RECT 792.000 682.050 792.900 694.200 ;
        RECT 797.100 682.050 798.900 683.850 ;
        RECT 812.700 682.050 813.900 695.400 ;
        RECT 830.400 689.400 832.200 702.000 ;
        RECT 835.500 690.900 837.300 701.400 ;
        RECT 838.500 695.400 840.300 702.000 ;
        RECT 854.100 695.400 855.900 702.000 ;
        RECT 857.100 695.400 858.900 701.400 ;
        RECT 860.100 695.400 861.900 702.000 ;
        RECT 838.200 692.100 840.000 693.900 ;
        RECT 835.500 689.400 837.900 690.900 ;
        RECT 815.100 682.050 816.900 683.850 ;
        RECT 830.100 682.050 831.900 683.850 ;
        RECT 836.700 682.050 837.900 689.400 ;
        RECT 857.700 682.050 858.900 695.400 ;
        RECT 872.100 690.300 873.900 701.400 ;
        RECT 875.100 691.200 876.900 702.000 ;
        RECT 878.100 690.300 879.900 701.400 ;
        RECT 872.100 689.400 879.900 690.300 ;
        RECT 881.100 689.400 882.900 701.400 ;
        RECT 896.100 695.400 897.900 702.000 ;
        RECT 899.100 695.400 900.900 701.400 ;
        RECT 902.100 695.400 903.900 702.000 ;
        RECT 875.250 682.050 877.050 683.850 ;
        RECT 881.700 682.050 882.600 689.400 ;
        RECT 891.000 684.450 895.050 685.050 ;
        RECT 890.550 682.950 895.050 684.450 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 767.400 672.600 768.300 679.950 ;
        RECT 769.950 678.150 771.750 679.950 ;
        RECT 776.100 678.150 777.900 679.950 ;
        RECT 792.000 676.200 792.900 679.950 ;
        RECT 794.100 678.150 795.900 679.950 ;
        RECT 800.100 678.150 801.900 679.950 ;
        RECT 792.000 675.000 795.300 676.200 ;
        RECT 767.400 671.400 772.500 672.600 ;
        RECT 748.500 666.600 750.300 669.600 ;
        RECT 751.500 666.000 753.300 669.600 ;
        RECT 767.700 666.000 769.500 669.600 ;
        RECT 770.700 666.600 772.500 671.400 ;
        RECT 775.200 666.000 777.000 672.600 ;
        RECT 793.500 666.600 795.300 675.000 ;
        RECT 800.100 666.000 801.900 675.600 ;
        RECT 812.700 669.600 813.900 679.950 ;
        RECT 833.100 678.150 834.900 679.950 ;
        RECT 836.700 675.600 837.900 679.950 ;
        RECT 839.100 678.150 840.900 679.950 ;
        RECT 844.950 678.450 847.050 679.050 ;
        RECT 850.950 678.450 853.050 679.050 ;
        RECT 844.950 677.550 853.050 678.450 ;
        RECT 854.100 678.150 855.900 679.950 ;
        RECT 844.950 676.950 847.050 677.550 ;
        RECT 850.950 676.950 853.050 677.550 ;
        RECT 836.700 674.700 840.300 675.600 ;
        RECT 857.700 674.700 858.900 679.950 ;
        RECT 859.950 678.150 861.750 679.950 ;
        RECT 872.100 678.150 873.900 679.950 ;
        RECT 878.250 678.150 880.050 679.950 ;
        RECT 830.100 671.700 837.900 673.050 ;
        RECT 812.100 666.600 813.900 669.600 ;
        RECT 815.100 666.000 816.900 669.600 ;
        RECT 830.100 666.600 831.900 671.700 ;
        RECT 833.100 666.000 834.900 670.800 ;
        RECT 836.100 666.600 837.900 671.700 ;
        RECT 839.100 672.600 840.300 674.700 ;
        RECT 854.700 673.800 858.900 674.700 ;
        RECT 839.100 666.600 840.900 672.600 ;
        RECT 854.700 666.600 856.500 673.800 ;
        RECT 881.700 672.600 882.600 679.950 ;
        RECT 883.950 678.450 886.050 679.050 ;
        RECT 890.550 678.450 891.450 682.950 ;
        RECT 899.700 682.050 900.900 695.400 ;
        RECT 914.100 690.600 915.900 701.400 ;
        RECT 917.100 691.500 918.900 702.000 ;
        RECT 920.100 700.500 927.900 701.400 ;
        RECT 920.100 690.600 921.900 700.500 ;
        RECT 914.100 689.700 921.900 690.600 ;
        RECT 923.100 688.500 924.900 699.600 ;
        RECT 926.100 689.400 927.900 700.500 ;
        RECT 938.100 695.400 939.900 702.000 ;
        RECT 941.100 695.400 942.900 701.400 ;
        RECT 944.100 695.400 945.900 702.000 ;
        RECT 920.100 687.600 924.900 688.500 ;
        RECT 904.950 684.450 909.000 685.050 ;
        RECT 904.950 682.950 909.450 684.450 ;
        RECT 895.950 679.950 898.050 682.050 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 883.950 677.550 891.450 678.450 ;
        RECT 896.100 678.150 897.900 679.950 ;
        RECT 883.950 676.950 886.050 677.550 ;
        RECT 899.700 674.700 900.900 679.950 ;
        RECT 901.950 678.150 903.750 679.950 ;
        RECT 859.800 666.000 861.600 672.600 ;
        RECT 873.000 666.000 874.800 672.600 ;
        RECT 877.500 671.400 882.600 672.600 ;
        RECT 896.700 673.800 900.900 674.700 ;
        RECT 901.950 675.450 904.050 676.050 ;
        RECT 908.550 675.450 909.450 682.950 ;
        RECT 917.250 682.050 919.050 683.850 ;
        RECT 920.100 682.050 921.000 687.600 ;
        RECT 923.100 682.050 924.900 683.850 ;
        RECT 941.700 682.050 942.900 695.400 ;
        RECT 913.950 679.950 916.050 682.050 ;
        RECT 916.950 679.950 919.050 682.050 ;
        RECT 919.950 679.950 922.050 682.050 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 925.950 679.950 928.050 682.050 ;
        RECT 937.950 679.950 940.050 682.050 ;
        RECT 940.950 679.950 943.050 682.050 ;
        RECT 943.950 679.950 946.050 682.050 ;
        RECT 914.250 678.150 916.050 679.950 ;
        RECT 901.950 674.550 909.450 675.450 ;
        RECT 901.950 673.950 904.050 674.550 ;
        RECT 877.500 666.600 879.300 671.400 ;
        RECT 880.500 666.000 882.300 669.600 ;
        RECT 896.700 666.600 898.500 673.800 ;
        RECT 920.100 672.600 921.300 679.950 ;
        RECT 926.100 678.150 927.900 679.950 ;
        RECT 938.100 678.150 939.900 679.950 ;
        RECT 941.700 674.700 942.900 679.950 ;
        RECT 943.950 678.150 945.750 679.950 ;
        RECT 938.700 673.800 942.900 674.700 ;
        RECT 901.800 666.000 903.600 672.600 ;
        RECT 914.700 666.000 916.500 672.600 ;
        RECT 919.200 666.600 921.000 672.600 ;
        RECT 923.700 666.000 925.500 672.600 ;
        RECT 938.700 666.600 940.500 673.800 ;
        RECT 943.800 666.000 945.600 672.600 ;
        RECT 14.100 659.400 15.900 662.400 ;
        RECT 14.100 655.500 15.300 659.400 ;
        RECT 17.100 656.400 18.900 663.000 ;
        RECT 20.100 656.400 21.900 662.400 ;
        RECT 36.600 658.200 38.400 662.400 ;
        RECT 14.100 654.600 19.800 655.500 ;
        RECT 18.000 653.700 19.800 654.600 ;
        RECT 14.400 646.950 16.500 649.050 ;
        RECT 14.400 645.150 16.200 646.950 ;
        RECT 18.000 642.300 18.900 653.700 ;
        RECT 20.700 649.050 21.900 656.400 ;
        RECT 35.700 656.400 38.400 658.200 ;
        RECT 39.600 656.400 41.400 663.000 ;
        RECT 35.700 649.050 36.600 656.400 ;
        RECT 37.500 654.600 39.300 655.500 ;
        RECT 44.100 654.600 45.900 662.400 ;
        RECT 56.400 656.400 58.200 663.000 ;
        RECT 61.500 655.200 63.300 662.400 ;
        RECT 76.500 656.400 78.300 663.000 ;
        RECT 81.000 656.400 82.800 662.400 ;
        RECT 85.500 656.400 87.300 663.000 ;
        RECT 101.100 656.400 102.900 662.400 ;
        RECT 37.500 653.700 45.900 654.600 ;
        RECT 59.100 654.300 63.300 655.200 ;
        RECT 19.800 646.950 21.900 649.050 ;
        RECT 35.100 646.950 37.200 649.050 ;
        RECT 38.400 646.950 40.500 649.050 ;
        RECT 18.000 641.400 19.800 642.300 ;
        RECT 14.100 640.500 19.800 641.400 ;
        RECT 14.100 633.600 15.300 640.500 ;
        RECT 20.700 639.600 21.900 646.950 ;
        RECT 35.700 639.600 36.600 646.950 ;
        RECT 39.000 645.150 40.800 646.950 ;
        RECT 14.100 627.600 15.900 633.600 ;
        RECT 17.100 627.000 18.900 637.800 ;
        RECT 20.100 627.600 21.900 639.600 ;
        RECT 35.100 627.600 36.900 639.600 ;
        RECT 38.100 627.000 39.900 639.000 ;
        RECT 42.000 633.600 42.900 653.700 ;
        RECT 43.950 649.050 45.750 650.850 ;
        RECT 56.250 649.050 58.050 650.850 ;
        RECT 59.100 649.050 60.300 654.300 ;
        RECT 62.100 649.050 63.900 650.850 ;
        RECT 74.100 649.050 75.900 650.850 ;
        RECT 80.700 649.050 81.900 656.400 ;
        RECT 101.700 654.300 102.900 656.400 ;
        RECT 104.100 657.300 105.900 662.400 ;
        RECT 107.100 658.200 108.900 663.000 ;
        RECT 110.100 657.300 111.900 662.400 ;
        RECT 104.100 655.950 111.900 657.300 ;
        RECT 112.950 657.450 115.050 658.050 ;
        RECT 118.950 657.450 121.050 658.050 ;
        RECT 112.950 656.550 121.050 657.450 ;
        RECT 112.950 655.950 115.050 656.550 ;
        RECT 118.950 655.950 121.050 656.550 ;
        RECT 125.400 656.400 127.200 663.000 ;
        RECT 130.500 655.200 132.300 662.400 ;
        RECT 115.950 654.450 118.050 655.050 ;
        RECT 124.950 654.450 127.050 655.050 ;
        RECT 101.700 653.400 105.300 654.300 ;
        RECT 85.950 649.050 87.750 650.850 ;
        RECT 101.100 649.050 102.900 650.850 ;
        RECT 104.100 649.050 105.300 653.400 ;
        RECT 115.950 653.550 127.050 654.450 ;
        RECT 115.950 652.950 118.050 653.550 ;
        RECT 124.950 652.950 127.050 653.550 ;
        RECT 128.100 654.300 132.300 655.200 ;
        RECT 146.100 656.400 147.900 662.400 ;
        RECT 149.100 656.400 150.900 663.000 ;
        RECT 152.100 659.400 153.900 662.400 ;
        RECT 107.100 649.050 108.900 650.850 ;
        RECT 125.250 649.050 127.050 650.850 ;
        RECT 128.100 649.050 129.300 654.300 ;
        RECT 133.950 651.450 136.050 652.050 ;
        RECT 142.950 651.450 145.050 652.050 ;
        RECT 131.100 649.050 132.900 650.850 ;
        RECT 133.950 650.550 145.050 651.450 ;
        RECT 133.950 649.950 136.050 650.550 ;
        RECT 142.950 649.950 145.050 650.550 ;
        RECT 146.100 649.050 147.300 656.400 ;
        RECT 152.700 655.500 153.900 659.400 ;
        RECT 167.700 656.400 169.500 663.000 ;
        RECT 172.200 656.400 174.000 662.400 ;
        RECT 176.700 656.400 178.500 663.000 ;
        RECT 194.100 656.400 195.900 662.400 ;
        RECT 148.200 654.600 153.900 655.500 ;
        RECT 148.200 653.700 150.000 654.600 ;
        RECT 43.800 646.950 45.900 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 130.950 646.950 133.050 649.050 ;
        RECT 146.100 646.950 148.200 649.050 ;
        RECT 59.100 633.600 60.300 646.950 ;
        RECT 77.100 645.150 78.900 646.950 ;
        RECT 61.950 642.450 64.050 643.050 ;
        RECT 70.950 642.450 73.050 643.050 ;
        RECT 61.950 641.550 73.050 642.450 ;
        RECT 61.950 640.950 64.050 641.550 ;
        RECT 70.950 640.950 73.050 641.550 ;
        RECT 81.000 641.400 81.900 646.950 ;
        RECT 82.950 645.150 84.750 646.950 ;
        RECT 77.100 640.500 81.900 641.400 ;
        RECT 41.100 627.600 42.900 633.600 ;
        RECT 44.100 627.000 45.900 633.600 ;
        RECT 56.100 627.000 57.900 633.600 ;
        RECT 59.100 627.600 60.900 633.600 ;
        RECT 62.100 627.000 63.900 633.600 ;
        RECT 74.100 628.500 75.900 639.600 ;
        RECT 77.100 629.400 78.900 640.500 ;
        RECT 104.100 639.600 105.300 646.950 ;
        RECT 110.100 645.150 111.900 646.950 ;
        RECT 80.100 638.400 87.900 639.300 ;
        RECT 80.100 628.500 81.900 638.400 ;
        RECT 74.100 627.600 81.900 628.500 ;
        RECT 83.100 627.000 84.900 637.500 ;
        RECT 86.100 627.600 87.900 638.400 ;
        RECT 104.100 638.100 106.500 639.600 ;
        RECT 102.000 635.100 103.800 636.900 ;
        RECT 101.700 627.000 103.500 633.600 ;
        RECT 104.700 627.600 106.500 638.100 ;
        RECT 109.800 627.000 111.600 639.600 ;
        RECT 128.100 633.600 129.300 646.950 ;
        RECT 146.100 639.600 147.300 646.950 ;
        RECT 149.100 642.300 150.000 653.700 ;
        RECT 162.000 651.450 166.050 652.050 ;
        RECT 161.550 649.950 166.050 651.450 ;
        RECT 151.500 646.950 153.600 649.050 ;
        RECT 151.800 645.150 153.600 646.950 ;
        RECT 161.550 646.050 162.450 649.950 ;
        RECT 167.250 649.050 169.050 650.850 ;
        RECT 173.100 649.050 174.300 656.400 ;
        RECT 194.700 654.300 195.900 656.400 ;
        RECT 197.100 657.300 198.900 662.400 ;
        RECT 200.100 658.200 201.900 663.000 ;
        RECT 203.100 657.300 204.900 662.400 ;
        RECT 197.100 655.950 204.900 657.300 ;
        RECT 218.400 656.400 220.200 663.000 ;
        RECT 223.500 655.200 225.300 662.400 ;
        RECT 236.100 656.400 237.900 662.400 ;
        RECT 221.100 654.300 225.300 655.200 ;
        RECT 236.700 654.300 237.900 656.400 ;
        RECT 239.100 657.300 240.900 662.400 ;
        RECT 242.100 658.200 243.900 663.000 ;
        RECT 245.100 657.300 246.900 662.400 ;
        RECT 258.600 658.200 260.400 662.400 ;
        RECT 239.100 655.950 246.900 657.300 ;
        RECT 257.700 656.400 260.400 658.200 ;
        RECT 261.600 656.400 263.400 663.000 ;
        RECT 194.700 653.400 198.300 654.300 ;
        RECT 179.100 649.050 180.900 650.850 ;
        RECT 194.100 649.050 195.900 650.850 ;
        RECT 197.100 649.050 198.300 653.400 ;
        RECT 200.100 649.050 201.900 650.850 ;
        RECT 218.250 649.050 220.050 650.850 ;
        RECT 221.100 649.050 222.300 654.300 ;
        RECT 236.700 653.400 240.300 654.300 ;
        RECT 224.100 649.050 225.900 650.850 ;
        RECT 236.100 649.050 237.900 650.850 ;
        RECT 239.100 649.050 240.300 653.400 ;
        RECT 242.100 649.050 243.900 650.850 ;
        RECT 257.700 649.050 258.600 656.400 ;
        RECT 259.500 654.600 261.300 655.500 ;
        RECT 266.100 654.600 267.900 662.400 ;
        RECT 259.500 653.700 267.900 654.600 ;
        RECT 283.500 654.000 285.300 662.400 ;
        RECT 166.950 646.950 169.050 649.050 ;
        RECT 169.950 646.950 172.050 649.050 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 193.950 646.950 196.050 649.050 ;
        RECT 196.950 646.950 199.050 649.050 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 217.950 646.950 220.050 649.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 241.950 646.950 244.050 649.050 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 257.100 646.950 259.200 649.050 ;
        RECT 260.400 646.950 262.500 649.050 ;
        RECT 161.550 644.550 166.050 646.050 ;
        RECT 170.250 645.150 172.050 646.950 ;
        RECT 162.000 643.950 166.050 644.550 ;
        RECT 148.200 641.400 150.000 642.300 ;
        RECT 173.100 641.400 174.000 646.950 ;
        RECT 176.100 645.150 177.900 646.950 ;
        RECT 148.200 640.500 153.900 641.400 ;
        RECT 173.100 640.500 177.900 641.400 ;
        RECT 125.100 627.000 126.900 633.600 ;
        RECT 128.100 627.600 129.900 633.600 ;
        RECT 131.100 627.000 132.900 633.600 ;
        RECT 146.100 627.600 147.900 639.600 ;
        RECT 149.100 627.000 150.900 637.800 ;
        RECT 152.700 633.600 153.900 640.500 ;
        RECT 152.100 627.600 153.900 633.600 ;
        RECT 167.100 638.400 174.900 639.300 ;
        RECT 167.100 627.600 168.900 638.400 ;
        RECT 170.100 627.000 171.900 637.500 ;
        RECT 173.100 628.500 174.900 638.400 ;
        RECT 176.100 629.400 177.900 640.500 ;
        RECT 197.100 639.600 198.300 646.950 ;
        RECT 203.100 645.150 204.900 646.950 ;
        RECT 179.100 628.500 180.900 639.600 ;
        RECT 197.100 638.100 199.500 639.600 ;
        RECT 195.000 635.100 196.800 636.900 ;
        RECT 173.100 627.600 180.900 628.500 ;
        RECT 194.700 627.000 196.500 633.600 ;
        RECT 197.700 627.600 199.500 638.100 ;
        RECT 202.800 627.000 204.600 639.600 ;
        RECT 221.100 633.600 222.300 646.950 ;
        RECT 239.100 639.600 240.300 646.950 ;
        RECT 245.100 645.150 246.900 646.950 ;
        RECT 257.700 639.600 258.600 646.950 ;
        RECT 261.000 645.150 262.800 646.950 ;
        RECT 239.100 638.100 241.500 639.600 ;
        RECT 237.000 635.100 238.800 636.900 ;
        RECT 218.100 627.000 219.900 633.600 ;
        RECT 221.100 627.600 222.900 633.600 ;
        RECT 224.100 627.000 225.900 633.600 ;
        RECT 236.700 627.000 238.500 633.600 ;
        RECT 239.700 627.600 241.500 638.100 ;
        RECT 244.800 627.000 246.600 639.600 ;
        RECT 257.100 627.600 258.900 639.600 ;
        RECT 260.100 627.000 261.900 639.000 ;
        RECT 264.000 633.600 264.900 653.700 ;
        RECT 282.000 652.800 285.300 654.000 ;
        RECT 290.100 653.400 291.900 663.000 ;
        RECT 305.100 659.400 306.900 663.000 ;
        RECT 308.100 659.400 309.900 662.400 ;
        RECT 265.950 649.050 267.750 650.850 ;
        RECT 282.000 649.050 282.900 652.800 ;
        RECT 284.100 649.050 285.900 650.850 ;
        RECT 290.100 649.050 291.900 650.850 ;
        RECT 308.100 649.050 309.300 659.400 ;
        RECT 320.400 656.400 322.200 663.000 ;
        RECT 325.500 655.200 327.300 662.400 ;
        RECT 338.100 656.400 339.900 662.400 ;
        RECT 341.100 657.300 342.900 663.000 ;
        RECT 345.600 656.400 347.400 662.400 ;
        RECT 350.100 657.300 351.900 663.000 ;
        RECT 353.100 656.400 354.900 662.400 ;
        RECT 356.700 659.400 358.500 663.000 ;
        RECT 359.700 659.400 361.500 662.400 ;
        RECT 338.100 655.500 342.900 656.400 ;
        RECT 323.100 654.300 327.300 655.200 ;
        RECT 340.800 654.300 342.900 655.500 ;
        RECT 345.900 654.900 347.100 656.400 ;
        RECT 320.250 649.050 322.050 650.850 ;
        RECT 323.100 649.050 324.300 654.300 ;
        RECT 344.100 652.800 347.100 654.900 ;
        RECT 353.100 654.600 354.300 656.400 ;
        RECT 326.100 649.050 327.900 650.850 ;
        RECT 342.900 649.800 345.000 651.900 ;
        RECT 265.800 646.950 267.900 649.050 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 307.950 646.950 310.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 325.950 646.950 328.050 649.050 ;
        RECT 338.100 646.950 340.200 649.050 ;
        RECT 342.900 648.000 344.700 649.800 ;
        RECT 345.900 647.100 347.100 652.800 ;
        RECT 348.000 653.700 354.300 654.600 ;
        RECT 348.000 651.600 350.100 653.700 ;
        RECT 348.000 649.800 349.800 651.600 ;
        RECT 352.800 649.050 354.600 650.850 ;
        RECT 352.800 648.300 354.900 649.050 ;
        RECT 282.000 634.800 282.900 646.950 ;
        RECT 287.100 645.150 288.900 646.950 ;
        RECT 305.100 645.150 306.900 646.950 ;
        RECT 282.000 633.900 288.600 634.800 ;
        RECT 282.000 633.600 282.900 633.900 ;
        RECT 263.100 627.600 264.900 633.600 ;
        RECT 266.100 627.000 267.900 633.600 ;
        RECT 281.100 627.600 282.900 633.600 ;
        RECT 287.100 633.600 288.600 633.900 ;
        RECT 308.100 633.600 309.300 646.950 ;
        RECT 323.100 633.600 324.300 646.950 ;
        RECT 338.400 645.150 340.200 646.950 ;
        RECT 344.700 646.200 347.100 647.100 ;
        RECT 348.000 646.950 354.900 648.300 ;
        RECT 348.000 646.500 349.800 646.950 ;
        RECT 344.700 646.050 346.200 646.200 ;
        RECT 360.000 646.050 361.500 659.400 ;
        RECT 344.100 643.950 346.200 646.050 ;
        RECT 345.300 642.000 346.200 643.950 ;
        RECT 347.100 643.500 351.000 645.300 ;
        RECT 359.100 643.950 361.500 646.050 ;
        RECT 347.100 643.200 349.200 643.500 ;
        RECT 345.300 640.950 346.800 642.000 ;
        RECT 340.800 639.600 342.900 640.500 ;
        RECT 338.100 638.400 342.900 639.600 ;
        RECT 345.600 639.600 346.800 640.950 ;
        RECT 350.400 639.600 352.500 641.700 ;
        RECT 284.100 627.000 285.900 633.000 ;
        RECT 287.100 627.600 288.900 633.600 ;
        RECT 290.100 627.000 291.900 633.600 ;
        RECT 305.100 627.000 306.900 633.600 ;
        RECT 308.100 627.600 309.900 633.600 ;
        RECT 320.100 627.000 321.900 633.600 ;
        RECT 323.100 627.600 324.900 633.600 ;
        RECT 326.100 627.000 327.900 633.600 ;
        RECT 338.100 627.600 339.900 638.400 ;
        RECT 341.100 627.000 342.900 637.500 ;
        RECT 345.600 627.600 347.400 639.600 ;
        RECT 350.400 638.700 354.900 639.600 ;
        RECT 350.100 627.000 351.900 637.500 ;
        RECT 353.100 627.600 354.900 638.700 ;
        RECT 360.000 633.600 361.500 643.950 ;
        RECT 363.300 656.400 365.100 662.400 ;
        RECT 368.700 656.400 370.500 663.000 ;
        RECT 373.800 657.600 375.600 662.400 ;
        RECT 378.000 659.400 379.800 662.400 ;
        RECT 381.000 659.400 382.800 662.400 ;
        RECT 384.000 659.400 385.800 662.400 ;
        RECT 387.000 659.400 388.800 662.400 ;
        RECT 390.000 659.400 391.800 663.000 ;
        RECT 371.400 656.400 375.600 657.600 ;
        RECT 377.700 657.300 379.800 659.400 ;
        RECT 380.700 657.300 382.800 659.400 ;
        RECT 383.700 657.300 385.800 659.400 ;
        RECT 386.700 657.300 388.800 659.400 ;
        RECT 393.000 658.500 394.800 662.400 ;
        RECT 397.500 659.400 399.300 663.000 ;
        RECT 400.500 659.400 402.300 662.400 ;
        RECT 403.500 659.400 405.300 662.400 ;
        RECT 406.500 659.400 408.300 662.400 ;
        RECT 392.100 656.400 394.800 658.500 ;
        RECT 396.600 657.600 398.400 658.500 ;
        RECT 396.600 656.400 399.300 657.600 ;
        RECT 400.200 657.300 402.300 659.400 ;
        RECT 403.200 657.300 405.300 659.400 ;
        RECT 406.200 657.300 408.300 659.400 ;
        RECT 410.700 656.400 412.500 662.400 ;
        RECT 416.100 656.400 417.900 663.000 ;
        RECT 421.500 656.400 423.300 662.400 ;
        RECT 437.400 656.400 439.200 663.000 ;
        RECT 363.300 639.600 364.200 656.400 ;
        RECT 371.400 653.100 372.900 656.400 ;
        RECT 377.100 654.600 383.700 656.400 ;
        RECT 398.400 655.800 399.300 656.400 ;
        RECT 401.400 655.800 403.200 656.400 ;
        RECT 398.400 654.600 405.600 655.800 ;
        RECT 365.100 651.300 372.900 653.100 ;
        RECT 389.100 652.500 390.900 654.300 ;
        RECT 388.800 651.900 390.900 652.500 ;
        RECT 373.800 650.400 390.900 651.900 ;
        RECT 395.100 651.900 397.200 652.050 ;
        RECT 398.400 651.900 400.200 652.800 ;
        RECT 395.100 651.000 400.200 651.900 ;
        RECT 404.700 651.600 405.600 654.600 ;
        RECT 410.700 655.500 412.200 656.400 ;
        RECT 410.700 654.300 419.100 655.500 ;
        RECT 417.300 653.700 419.100 654.300 ;
        RECT 406.500 652.800 408.600 653.700 ;
        RECT 422.100 652.800 423.300 656.400 ;
        RECT 442.500 655.200 444.300 662.400 ;
        RECT 406.500 651.600 423.300 652.800 ;
        RECT 368.700 648.900 375.300 650.400 ;
        RECT 395.100 649.950 397.200 651.000 ;
        RECT 403.800 649.800 405.600 651.600 ;
        RECT 368.700 646.050 370.200 648.900 ;
        RECT 376.500 647.700 420.900 648.900 ;
        RECT 376.500 646.200 377.400 647.700 ;
        RECT 368.100 643.950 370.200 646.050 ;
        RECT 372.300 644.400 377.400 646.200 ;
        RECT 380.100 645.900 393.600 646.800 ;
        RECT 400.800 645.900 402.600 646.500 ;
        RECT 419.100 646.050 420.900 647.700 ;
        RECT 380.100 644.700 381.000 645.900 ;
        RECT 380.100 642.900 381.900 644.700 ;
        RECT 386.100 643.200 390.000 645.000 ;
        RECT 391.500 644.700 402.600 645.900 ;
        RECT 413.100 645.750 415.200 646.050 ;
        RECT 391.500 643.800 393.600 644.700 ;
        RECT 411.300 643.950 415.200 645.750 ;
        RECT 419.100 643.950 421.200 646.050 ;
        RECT 411.300 643.200 413.100 643.950 ;
        RECT 386.100 642.900 388.200 643.200 ;
        RECT 399.600 642.300 413.100 643.200 ;
        RECT 365.100 641.700 366.900 642.300 ;
        RECT 399.600 641.700 400.800 642.300 ;
        RECT 365.100 640.500 400.800 641.700 ;
        RECT 403.500 640.500 405.600 640.800 ;
        RECT 363.300 638.700 379.800 639.600 ;
        RECT 363.300 635.400 364.200 638.700 ;
        RECT 368.100 636.600 373.800 637.800 ;
        RECT 377.700 637.500 379.800 638.700 ;
        RECT 383.100 638.400 400.800 639.600 ;
        RECT 403.500 639.300 415.500 640.500 ;
        RECT 403.500 638.700 405.600 639.300 ;
        RECT 413.700 638.700 415.500 639.300 ;
        RECT 383.100 637.500 385.200 638.400 ;
        RECT 399.600 637.800 400.800 638.400 ;
        RECT 417.000 637.800 418.800 638.100 ;
        RECT 368.100 636.000 369.900 636.600 ;
        RECT 363.300 634.500 367.200 635.400 ;
        RECT 366.000 633.600 367.200 634.500 ;
        RECT 372.600 633.600 373.800 636.600 ;
        RECT 374.700 635.700 376.500 636.300 ;
        RECT 374.700 634.500 382.800 635.700 ;
        RECT 380.700 633.600 382.800 634.500 ;
        RECT 386.100 633.600 388.800 637.500 ;
        RECT 391.500 635.100 394.800 637.200 ;
        RECT 399.600 636.600 418.800 637.800 ;
        RECT 356.700 627.000 358.500 633.600 ;
        RECT 359.700 627.600 361.500 633.600 ;
        RECT 363.000 627.000 364.800 633.600 ;
        RECT 366.000 627.600 367.800 633.600 ;
        RECT 369.000 627.000 370.800 633.600 ;
        RECT 372.000 627.600 373.800 633.600 ;
        RECT 375.000 627.000 376.800 633.600 ;
        RECT 377.700 630.600 379.800 632.700 ;
        RECT 380.700 630.600 382.800 632.700 ;
        RECT 383.700 630.600 385.800 632.700 ;
        RECT 378.000 627.600 379.800 630.600 ;
        RECT 381.000 627.600 382.800 630.600 ;
        RECT 384.000 627.600 385.800 630.600 ;
        RECT 387.000 627.600 388.800 633.600 ;
        RECT 390.000 627.000 391.800 633.600 ;
        RECT 393.000 627.600 394.800 635.100 ;
        RECT 400.200 633.600 402.300 635.700 ;
        RECT 396.900 627.000 398.700 633.600 ;
        RECT 399.900 627.600 401.700 633.600 ;
        RECT 402.600 630.600 404.700 632.700 ;
        RECT 405.600 630.600 407.700 632.700 ;
        RECT 402.900 627.600 404.700 630.600 ;
        RECT 405.900 627.600 407.700 630.600 ;
        RECT 409.500 627.000 411.300 633.600 ;
        RECT 412.500 627.600 414.300 636.600 ;
        RECT 417.000 636.300 418.800 636.600 ;
        RECT 422.100 635.400 423.300 651.600 ;
        RECT 440.100 654.300 444.300 655.200 ;
        RECT 455.100 656.400 456.900 662.400 ;
        RECT 458.100 656.400 459.900 663.000 ;
        RECT 461.100 659.400 462.900 662.400 ;
        RECT 437.250 649.050 439.050 650.850 ;
        RECT 440.100 649.050 441.300 654.300 ;
        RECT 443.100 649.050 444.900 650.850 ;
        RECT 455.100 649.050 456.300 656.400 ;
        RECT 461.700 655.500 462.900 659.400 ;
        RECT 457.200 654.600 462.900 655.500 ;
        RECT 476.100 656.400 477.900 662.400 ;
        RECT 479.100 656.400 480.900 663.000 ;
        RECT 482.100 659.400 483.900 662.400 ;
        RECT 457.200 653.700 459.000 654.600 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 455.100 646.950 457.200 649.050 ;
        RECT 419.700 634.500 423.300 635.400 ;
        RECT 419.700 633.600 420.600 634.500 ;
        RECT 440.100 633.600 441.300 646.950 ;
        RECT 455.100 639.600 456.300 646.950 ;
        RECT 458.100 642.300 459.000 653.700 ;
        RECT 476.100 649.050 477.300 656.400 ;
        RECT 482.700 655.500 483.900 659.400 ;
        RECT 497.400 656.400 499.200 663.000 ;
        RECT 478.200 654.600 483.900 655.500 ;
        RECT 502.500 655.200 504.300 662.400 ;
        RECT 515.100 656.400 516.900 662.400 ;
        RECT 478.200 653.700 480.000 654.600 ;
        RECT 460.500 646.950 462.600 649.050 ;
        RECT 460.800 645.150 462.600 646.950 ;
        RECT 476.100 646.950 478.200 649.050 ;
        RECT 457.200 641.400 459.000 642.300 ;
        RECT 457.200 640.500 462.900 641.400 ;
        RECT 415.500 627.000 417.300 633.600 ;
        RECT 418.500 632.700 420.600 633.600 ;
        RECT 418.500 627.600 420.300 632.700 ;
        RECT 421.500 627.000 423.300 633.600 ;
        RECT 437.100 627.000 438.900 633.600 ;
        RECT 440.100 627.600 441.900 633.600 ;
        RECT 443.100 627.000 444.900 633.600 ;
        RECT 455.100 627.600 456.900 639.600 ;
        RECT 458.100 627.000 459.900 637.800 ;
        RECT 461.700 633.600 462.900 640.500 ;
        RECT 461.100 627.600 462.900 633.600 ;
        RECT 476.100 639.600 477.300 646.950 ;
        RECT 479.100 642.300 480.000 653.700 ;
        RECT 500.100 654.300 504.300 655.200 ;
        RECT 515.700 654.300 516.900 656.400 ;
        RECT 518.100 657.300 519.900 662.400 ;
        RECT 521.100 658.200 522.900 663.000 ;
        RECT 524.100 657.300 525.900 662.400 ;
        RECT 527.700 659.400 529.500 663.000 ;
        RECT 530.700 659.400 532.500 662.400 ;
        RECT 518.100 655.950 525.900 657.300 ;
        RECT 497.250 649.050 499.050 650.850 ;
        RECT 500.100 649.050 501.300 654.300 ;
        RECT 515.700 653.400 519.300 654.300 ;
        RECT 503.100 649.050 504.900 650.850 ;
        RECT 515.100 649.050 516.900 650.850 ;
        RECT 518.100 649.050 519.300 653.400 ;
        RECT 521.100 649.050 522.900 650.850 ;
        RECT 481.500 646.950 483.600 649.050 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 514.950 646.950 517.050 649.050 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 481.800 645.150 483.600 646.950 ;
        RECT 484.950 645.450 487.050 646.050 ;
        RECT 493.950 645.450 496.050 646.050 ;
        RECT 484.950 644.550 496.050 645.450 ;
        RECT 484.950 643.950 487.050 644.550 ;
        RECT 493.950 643.950 496.050 644.550 ;
        RECT 478.200 641.400 480.000 642.300 ;
        RECT 478.200 640.500 483.900 641.400 ;
        RECT 476.100 627.600 477.900 639.600 ;
        RECT 479.100 627.000 480.900 637.800 ;
        RECT 482.700 633.600 483.900 640.500 ;
        RECT 500.100 633.600 501.300 646.950 ;
        RECT 518.100 639.600 519.300 646.950 ;
        RECT 524.100 645.150 525.900 646.950 ;
        RECT 531.000 646.050 532.500 659.400 ;
        RECT 530.100 643.950 532.500 646.050 ;
        RECT 518.100 638.100 520.500 639.600 ;
        RECT 516.000 635.100 517.800 636.900 ;
        RECT 482.100 627.600 483.900 633.600 ;
        RECT 497.100 627.000 498.900 633.600 ;
        RECT 500.100 627.600 501.900 633.600 ;
        RECT 503.100 627.000 504.900 633.600 ;
        RECT 515.700 627.000 517.500 633.600 ;
        RECT 518.700 627.600 520.500 638.100 ;
        RECT 523.800 627.000 525.600 639.600 ;
        RECT 531.000 633.600 532.500 643.950 ;
        RECT 534.300 656.400 536.100 662.400 ;
        RECT 539.700 656.400 541.500 663.000 ;
        RECT 544.800 657.600 546.600 662.400 ;
        RECT 549.000 659.400 550.800 662.400 ;
        RECT 552.000 659.400 553.800 662.400 ;
        RECT 555.000 659.400 556.800 662.400 ;
        RECT 558.000 659.400 559.800 662.400 ;
        RECT 561.000 659.400 562.800 663.000 ;
        RECT 542.400 656.400 546.600 657.600 ;
        RECT 548.700 657.300 550.800 659.400 ;
        RECT 551.700 657.300 553.800 659.400 ;
        RECT 554.700 657.300 556.800 659.400 ;
        RECT 557.700 657.300 559.800 659.400 ;
        RECT 564.000 658.500 565.800 662.400 ;
        RECT 568.500 659.400 570.300 663.000 ;
        RECT 571.500 659.400 573.300 662.400 ;
        RECT 574.500 659.400 576.300 662.400 ;
        RECT 577.500 659.400 579.300 662.400 ;
        RECT 563.100 656.400 565.800 658.500 ;
        RECT 567.600 657.600 569.400 658.500 ;
        RECT 567.600 656.400 570.300 657.600 ;
        RECT 571.200 657.300 573.300 659.400 ;
        RECT 574.200 657.300 576.300 659.400 ;
        RECT 577.200 657.300 579.300 659.400 ;
        RECT 581.700 656.400 583.500 662.400 ;
        RECT 587.100 656.400 588.900 663.000 ;
        RECT 592.500 656.400 594.300 662.400 ;
        RECT 534.300 639.600 535.200 656.400 ;
        RECT 542.400 653.100 543.900 656.400 ;
        RECT 548.100 654.600 554.700 656.400 ;
        RECT 569.400 655.800 570.300 656.400 ;
        RECT 572.400 655.800 574.200 656.400 ;
        RECT 569.400 654.600 576.600 655.800 ;
        RECT 536.100 651.300 543.900 653.100 ;
        RECT 560.100 652.500 561.900 654.300 ;
        RECT 559.800 651.900 561.900 652.500 ;
        RECT 544.800 650.400 561.900 651.900 ;
        RECT 566.100 651.900 568.200 652.050 ;
        RECT 569.400 651.900 571.200 652.800 ;
        RECT 566.100 651.000 571.200 651.900 ;
        RECT 575.700 651.600 576.600 654.600 ;
        RECT 581.700 655.500 583.200 656.400 ;
        RECT 581.700 654.300 590.100 655.500 ;
        RECT 588.300 653.700 590.100 654.300 ;
        RECT 577.500 652.800 579.600 653.700 ;
        RECT 593.100 652.800 594.300 656.400 ;
        RECT 608.100 657.300 609.900 662.400 ;
        RECT 611.100 658.200 612.900 663.000 ;
        RECT 614.100 657.300 615.900 662.400 ;
        RECT 608.100 655.950 615.900 657.300 ;
        RECT 617.100 656.400 618.900 662.400 ;
        RECT 617.100 654.300 618.300 656.400 ;
        RECT 629.700 655.200 631.500 662.400 ;
        RECT 634.800 656.400 636.600 663.000 ;
        RECT 650.400 656.400 652.200 663.000 ;
        RECT 655.500 655.200 657.300 662.400 ;
        RECT 629.700 654.300 633.900 655.200 ;
        RECT 577.500 651.600 594.300 652.800 ;
        RECT 539.700 648.900 546.300 650.400 ;
        RECT 566.100 649.950 568.200 651.000 ;
        RECT 574.800 649.800 576.600 651.600 ;
        RECT 539.700 646.050 541.200 648.900 ;
        RECT 547.500 647.700 591.900 648.900 ;
        RECT 547.500 646.200 548.400 647.700 ;
        RECT 539.100 643.950 541.200 646.050 ;
        RECT 543.300 644.400 548.400 646.200 ;
        RECT 551.100 645.900 564.600 646.800 ;
        RECT 571.800 645.900 573.600 646.500 ;
        RECT 590.100 646.050 591.900 647.700 ;
        RECT 551.100 644.700 552.000 645.900 ;
        RECT 551.100 642.900 552.900 644.700 ;
        RECT 557.100 643.200 561.000 645.000 ;
        RECT 562.500 644.700 573.600 645.900 ;
        RECT 584.100 645.750 586.200 646.050 ;
        RECT 562.500 643.800 564.600 644.700 ;
        RECT 582.300 643.950 586.200 645.750 ;
        RECT 590.100 643.950 592.200 646.050 ;
        RECT 582.300 643.200 584.100 643.950 ;
        RECT 557.100 642.900 559.200 643.200 ;
        RECT 570.600 642.300 584.100 643.200 ;
        RECT 536.100 641.700 537.900 642.300 ;
        RECT 570.600 641.700 571.800 642.300 ;
        RECT 536.100 640.500 571.800 641.700 ;
        RECT 574.500 640.500 576.600 640.800 ;
        RECT 534.300 638.700 550.800 639.600 ;
        RECT 534.300 635.400 535.200 638.700 ;
        RECT 539.100 636.600 544.800 637.800 ;
        RECT 548.700 637.500 550.800 638.700 ;
        RECT 554.100 638.400 571.800 639.600 ;
        RECT 574.500 639.300 586.500 640.500 ;
        RECT 574.500 638.700 576.600 639.300 ;
        RECT 584.700 638.700 586.500 639.300 ;
        RECT 554.100 637.500 556.200 638.400 ;
        RECT 570.600 637.800 571.800 638.400 ;
        RECT 588.000 637.800 589.800 638.100 ;
        RECT 539.100 636.000 540.900 636.600 ;
        RECT 534.300 634.500 538.200 635.400 ;
        RECT 537.000 633.600 538.200 634.500 ;
        RECT 543.600 633.600 544.800 636.600 ;
        RECT 545.700 635.700 547.500 636.300 ;
        RECT 545.700 634.500 553.800 635.700 ;
        RECT 551.700 633.600 553.800 634.500 ;
        RECT 557.100 633.600 559.800 637.500 ;
        RECT 562.500 635.100 565.800 637.200 ;
        RECT 570.600 636.600 589.800 637.800 ;
        RECT 527.700 627.000 529.500 633.600 ;
        RECT 530.700 627.600 532.500 633.600 ;
        RECT 534.000 627.000 535.800 633.600 ;
        RECT 537.000 627.600 538.800 633.600 ;
        RECT 540.000 627.000 541.800 633.600 ;
        RECT 543.000 627.600 544.800 633.600 ;
        RECT 546.000 627.000 547.800 633.600 ;
        RECT 548.700 630.600 550.800 632.700 ;
        RECT 551.700 630.600 553.800 632.700 ;
        RECT 554.700 630.600 556.800 632.700 ;
        RECT 549.000 627.600 550.800 630.600 ;
        RECT 552.000 627.600 553.800 630.600 ;
        RECT 555.000 627.600 556.800 630.600 ;
        RECT 558.000 627.600 559.800 633.600 ;
        RECT 561.000 627.000 562.800 633.600 ;
        RECT 564.000 627.600 565.800 635.100 ;
        RECT 571.200 633.600 573.300 635.700 ;
        RECT 567.900 627.000 569.700 633.600 ;
        RECT 570.900 627.600 572.700 633.600 ;
        RECT 573.600 630.600 575.700 632.700 ;
        RECT 576.600 630.600 578.700 632.700 ;
        RECT 573.900 627.600 575.700 630.600 ;
        RECT 576.900 627.600 578.700 630.600 ;
        RECT 580.500 627.000 582.300 633.600 ;
        RECT 583.500 627.600 585.300 636.600 ;
        RECT 588.000 636.300 589.800 636.600 ;
        RECT 593.100 635.400 594.300 651.600 ;
        RECT 614.700 653.400 618.300 654.300 ;
        RECT 611.100 649.050 612.900 650.850 ;
        RECT 614.700 649.050 615.900 653.400 ;
        RECT 617.100 649.050 618.900 650.850 ;
        RECT 629.100 649.050 630.900 650.850 ;
        RECT 632.700 649.050 633.900 654.300 ;
        RECT 653.100 654.300 657.300 655.200 ;
        RECT 634.950 649.050 636.750 650.850 ;
        RECT 650.250 649.050 652.050 650.850 ;
        RECT 653.100 649.050 654.300 654.300 ;
        RECT 671.100 653.400 672.900 663.000 ;
        RECT 677.700 654.000 679.500 662.400 ;
        RECT 677.700 652.800 681.000 654.000 ;
        RECT 692.100 653.400 693.900 663.000 ;
        RECT 698.700 654.000 700.500 662.400 ;
        RECT 716.700 655.200 718.500 662.400 ;
        RECT 721.800 656.400 723.600 663.000 ;
        RECT 734.100 656.400 735.900 662.400 ;
        RECT 737.100 657.300 738.900 663.000 ;
        RECT 741.600 656.400 743.400 662.400 ;
        RECT 746.100 657.300 747.900 663.000 ;
        RECT 749.100 656.400 750.900 662.400 ;
        RECT 764.100 656.400 765.900 662.400 ;
        RECT 767.100 657.300 768.900 663.000 ;
        RECT 771.600 656.400 773.400 662.400 ;
        RECT 776.100 657.300 777.900 663.000 ;
        RECT 779.100 656.400 780.900 662.400 ;
        RECT 791.100 659.400 792.900 663.000 ;
        RECT 794.100 659.400 795.900 662.400 ;
        RECT 716.700 654.300 720.900 655.200 ;
        RECT 698.700 652.800 702.000 654.000 ;
        RECT 656.100 649.050 657.900 650.850 ;
        RECT 671.100 649.050 672.900 650.850 ;
        RECT 677.100 649.050 678.900 650.850 ;
        RECT 680.100 649.050 681.000 652.800 ;
        RECT 687.000 651.450 691.050 652.050 ;
        RECT 686.550 649.950 691.050 651.450 ;
        RECT 598.950 645.450 601.050 649.050 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 634.950 646.950 637.050 649.050 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 604.950 645.450 607.050 646.050 ;
        RECT 598.950 645.000 607.050 645.450 ;
        RECT 608.100 645.150 609.900 646.950 ;
        RECT 599.550 644.550 607.050 645.000 ;
        RECT 604.950 643.950 607.050 644.550 ;
        RECT 595.950 642.450 598.050 643.050 ;
        RECT 601.950 642.450 604.050 642.900 ;
        RECT 595.950 641.550 604.050 642.450 ;
        RECT 595.950 640.950 598.050 641.550 ;
        RECT 601.950 640.800 604.050 641.550 ;
        RECT 614.700 639.600 615.900 646.950 ;
        RECT 590.700 634.500 594.300 635.400 ;
        RECT 590.700 633.600 591.600 634.500 ;
        RECT 586.500 627.000 588.300 633.600 ;
        RECT 589.500 632.700 591.600 633.600 ;
        RECT 589.500 627.600 591.300 632.700 ;
        RECT 592.500 627.000 594.300 633.600 ;
        RECT 608.400 627.000 610.200 639.600 ;
        RECT 613.500 638.100 615.900 639.600 ;
        RECT 613.500 627.600 615.300 638.100 ;
        RECT 616.200 635.100 618.000 636.900 ;
        RECT 632.700 633.600 633.900 646.950 ;
        RECT 653.100 633.600 654.300 646.950 ;
        RECT 674.100 645.150 675.900 646.950 ;
        RECT 661.950 642.450 664.050 643.050 ;
        RECT 670.950 642.450 673.050 643.050 ;
        RECT 661.950 641.550 673.050 642.450 ;
        RECT 661.950 640.950 664.050 641.550 ;
        RECT 670.950 640.950 673.050 641.550 ;
        RECT 680.100 634.800 681.000 646.950 ;
        RECT 686.550 646.050 687.450 649.950 ;
        RECT 692.100 649.050 693.900 650.850 ;
        RECT 698.100 649.050 699.900 650.850 ;
        RECT 701.100 649.050 702.000 652.800 ;
        RECT 716.100 649.050 717.900 650.850 ;
        RECT 719.700 649.050 720.900 654.300 ;
        RECT 734.700 654.600 735.900 656.400 ;
        RECT 741.900 654.900 743.100 656.400 ;
        RECT 746.100 655.500 750.900 656.400 ;
        RECT 734.700 653.700 741.000 654.600 ;
        RECT 738.900 651.600 741.000 653.700 ;
        RECT 721.950 649.050 723.750 650.850 ;
        RECT 734.400 649.050 736.200 650.850 ;
        RECT 739.200 649.800 741.000 651.600 ;
        RECT 741.900 652.800 744.900 654.900 ;
        RECT 746.100 654.300 748.200 655.500 ;
        RECT 764.700 654.600 765.900 656.400 ;
        RECT 771.900 654.900 773.100 656.400 ;
        RECT 776.100 655.500 780.900 656.400 ;
        RECT 764.700 653.700 771.000 654.600 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 734.100 648.300 736.200 649.050 ;
        RECT 734.100 646.950 741.000 648.300 ;
        RECT 682.950 644.550 687.450 646.050 ;
        RECT 695.100 645.150 696.900 646.950 ;
        RECT 682.950 643.950 687.000 644.550 ;
        RECT 701.100 634.800 702.000 646.950 ;
        RECT 674.400 633.900 681.000 634.800 ;
        RECT 674.400 633.600 675.900 633.900 ;
        RECT 616.500 627.000 618.300 633.600 ;
        RECT 629.100 627.000 630.900 633.600 ;
        RECT 632.100 627.600 633.900 633.600 ;
        RECT 635.100 627.000 636.900 633.600 ;
        RECT 650.100 627.000 651.900 633.600 ;
        RECT 653.100 627.600 654.900 633.600 ;
        RECT 656.100 627.000 657.900 633.600 ;
        RECT 671.100 627.000 672.900 633.600 ;
        RECT 674.100 627.600 675.900 633.600 ;
        RECT 680.100 633.600 681.000 633.900 ;
        RECT 695.400 633.900 702.000 634.800 ;
        RECT 695.400 633.600 696.900 633.900 ;
        RECT 677.100 627.000 678.900 633.000 ;
        RECT 680.100 627.600 681.900 633.600 ;
        RECT 692.100 627.000 693.900 633.600 ;
        RECT 695.100 627.600 696.900 633.600 ;
        RECT 701.100 633.600 702.000 633.900 ;
        RECT 719.700 633.600 720.900 646.950 ;
        RECT 739.200 646.500 741.000 646.950 ;
        RECT 741.900 647.100 743.100 652.800 ;
        RECT 744.000 649.800 746.100 651.900 ;
        RECT 768.900 651.600 771.000 653.700 ;
        RECT 744.300 648.000 746.100 649.800 ;
        RECT 764.400 649.050 766.200 650.850 ;
        RECT 769.200 649.800 771.000 651.600 ;
        RECT 771.900 652.800 774.900 654.900 ;
        RECT 776.100 654.300 778.200 655.500 ;
        RECT 741.900 646.200 744.300 647.100 ;
        RECT 742.800 646.050 744.300 646.200 ;
        RECT 748.800 646.950 750.900 649.050 ;
        RECT 764.100 648.300 766.200 649.050 ;
        RECT 764.100 646.950 771.000 648.300 ;
        RECT 738.000 643.500 741.900 645.300 ;
        RECT 739.800 643.200 741.900 643.500 ;
        RECT 742.800 643.950 744.900 646.050 ;
        RECT 748.800 645.150 750.600 646.950 ;
        RECT 769.200 646.500 771.000 646.950 ;
        RECT 771.900 647.100 773.100 652.800 ;
        RECT 774.000 649.800 776.100 651.900 ;
        RECT 774.300 648.000 776.100 649.800 ;
        RECT 794.100 649.050 795.300 659.400 ;
        RECT 809.100 656.400 810.900 662.400 ;
        RECT 809.700 654.300 810.900 656.400 ;
        RECT 812.100 657.300 813.900 662.400 ;
        RECT 815.100 658.200 816.900 663.000 ;
        RECT 818.100 657.300 819.900 662.400 ;
        RECT 812.100 655.950 819.900 657.300 ;
        RECT 833.100 656.400 834.900 662.400 ;
        RECT 836.100 657.300 837.900 663.000 ;
        RECT 840.600 656.400 842.400 662.400 ;
        RECT 845.100 657.300 846.900 663.000 ;
        RECT 848.100 656.400 849.900 662.400 ;
        RECT 863.700 659.400 865.500 663.000 ;
        RECT 866.700 657.600 868.500 662.400 ;
        RECT 833.700 654.600 834.900 656.400 ;
        RECT 840.900 654.900 842.100 656.400 ;
        RECT 845.100 655.500 849.900 656.400 ;
        RECT 863.400 656.400 868.500 657.600 ;
        RECT 871.200 656.400 873.000 663.000 ;
        RECT 809.700 653.400 813.300 654.300 ;
        RECT 833.700 653.700 840.000 654.600 ;
        RECT 809.100 649.050 810.900 650.850 ;
        RECT 812.100 649.050 813.300 653.400 ;
        RECT 837.900 651.600 840.000 653.700 ;
        RECT 815.100 649.050 816.900 650.850 ;
        RECT 833.400 649.050 835.200 650.850 ;
        RECT 838.200 649.800 840.000 651.600 ;
        RECT 840.900 652.800 843.900 654.900 ;
        RECT 845.100 654.300 847.200 655.500 ;
        RECT 771.900 646.200 774.300 647.100 ;
        RECT 772.800 646.050 774.300 646.200 ;
        RECT 778.800 646.950 780.900 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 833.100 648.300 835.200 649.050 ;
        RECT 833.100 646.950 840.000 648.300 ;
        RECT 742.800 642.000 743.700 643.950 ;
        RECT 768.000 643.500 771.900 645.300 ;
        RECT 769.800 643.200 771.900 643.500 ;
        RECT 772.800 643.950 774.900 646.050 ;
        RECT 778.800 645.150 780.600 646.950 ;
        RECT 791.100 645.150 792.900 646.950 ;
        RECT 772.800 642.000 773.700 643.950 ;
        RECT 736.500 639.600 738.600 641.700 ;
        RECT 742.200 640.950 743.700 642.000 ;
        RECT 742.200 639.600 743.400 640.950 ;
        RECT 734.100 638.700 738.600 639.600 ;
        RECT 698.100 627.000 699.900 633.000 ;
        RECT 701.100 627.600 702.900 633.600 ;
        RECT 716.100 627.000 717.900 633.600 ;
        RECT 719.100 627.600 720.900 633.600 ;
        RECT 722.100 627.000 723.900 633.600 ;
        RECT 734.100 627.600 735.900 638.700 ;
        RECT 737.100 627.000 738.900 637.500 ;
        RECT 741.600 627.600 743.400 639.600 ;
        RECT 746.100 639.600 748.200 640.500 ;
        RECT 766.500 639.600 768.600 641.700 ;
        RECT 772.200 640.950 773.700 642.000 ;
        RECT 772.200 639.600 773.400 640.950 ;
        RECT 746.100 638.400 750.900 639.600 ;
        RECT 746.100 627.000 747.900 637.500 ;
        RECT 749.100 627.600 750.900 638.400 ;
        RECT 764.100 638.700 768.600 639.600 ;
        RECT 764.100 627.600 765.900 638.700 ;
        RECT 767.100 627.000 768.900 637.500 ;
        RECT 771.600 627.600 773.400 639.600 ;
        RECT 776.100 639.600 778.200 640.500 ;
        RECT 776.100 638.400 780.900 639.600 ;
        RECT 776.100 627.000 777.900 637.500 ;
        RECT 779.100 627.600 780.900 638.400 ;
        RECT 794.100 633.600 795.300 646.950 ;
        RECT 796.950 645.450 799.050 646.050 ;
        RECT 805.950 645.450 808.050 646.050 ;
        RECT 796.950 644.550 808.050 645.450 ;
        RECT 796.950 643.950 799.050 644.550 ;
        RECT 805.950 643.950 808.050 644.550 ;
        RECT 812.100 639.600 813.300 646.950 ;
        RECT 818.100 645.150 819.900 646.950 ;
        RECT 838.200 646.500 840.000 646.950 ;
        RECT 840.900 647.100 842.100 652.800 ;
        RECT 843.000 649.800 845.100 651.900 ;
        RECT 843.300 648.000 845.100 649.800 ;
        RECT 863.400 649.050 864.300 656.400 ;
        RECT 887.100 653.400 888.900 663.000 ;
        RECT 893.700 654.000 895.500 662.400 ;
        RECT 911.100 659.400 912.900 663.000 ;
        RECT 914.100 659.400 915.900 662.400 ;
        RECT 893.700 652.800 897.000 654.000 ;
        RECT 865.950 649.050 867.750 650.850 ;
        RECT 872.100 649.050 873.900 650.850 ;
        RECT 887.100 649.050 888.900 650.850 ;
        RECT 893.100 649.050 894.900 650.850 ;
        RECT 896.100 649.050 897.000 652.800 ;
        RECT 914.100 649.050 915.300 659.400 ;
        RECT 928.500 654.000 930.300 662.400 ;
        RECT 927.000 652.800 930.300 654.000 ;
        RECT 935.100 653.400 936.900 663.000 ;
        RECT 927.000 649.050 927.900 652.800 ;
        RECT 929.100 649.050 930.900 650.850 ;
        RECT 935.100 649.050 936.900 650.850 ;
        RECT 840.900 646.200 843.300 647.100 ;
        RECT 841.800 646.050 843.300 646.200 ;
        RECT 847.800 646.950 849.900 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 925.950 646.950 928.050 649.050 ;
        RECT 928.950 646.950 931.050 649.050 ;
        RECT 931.950 646.950 934.050 649.050 ;
        RECT 934.950 646.950 937.050 649.050 ;
        RECT 837.000 643.500 840.900 645.300 ;
        RECT 838.800 643.200 840.900 643.500 ;
        RECT 841.800 643.950 843.900 646.050 ;
        RECT 847.800 645.150 849.600 646.950 ;
        RECT 841.800 642.000 842.700 643.950 ;
        RECT 835.500 639.600 837.600 641.700 ;
        RECT 841.200 640.950 842.700 642.000 ;
        RECT 841.200 639.600 842.400 640.950 ;
        RECT 812.100 638.100 814.500 639.600 ;
        RECT 810.000 635.100 811.800 636.900 ;
        RECT 791.100 627.000 792.900 633.600 ;
        RECT 794.100 627.600 795.900 633.600 ;
        RECT 809.700 627.000 811.500 633.600 ;
        RECT 812.700 627.600 814.500 638.100 ;
        RECT 817.800 627.000 819.600 639.600 ;
        RECT 833.100 638.700 837.600 639.600 ;
        RECT 833.100 627.600 834.900 638.700 ;
        RECT 836.100 627.000 837.900 637.500 ;
        RECT 840.600 627.600 842.400 639.600 ;
        RECT 845.100 639.600 847.200 640.500 ;
        RECT 863.400 639.600 864.300 646.950 ;
        RECT 868.950 645.150 870.750 646.950 ;
        RECT 890.100 645.150 891.900 646.950 ;
        RECT 880.950 642.450 883.050 643.050 ;
        RECT 892.950 642.450 895.050 643.050 ;
        RECT 880.950 641.550 895.050 642.450 ;
        RECT 880.950 640.950 883.050 641.550 ;
        RECT 892.950 640.950 895.050 641.550 ;
        RECT 845.100 638.400 849.900 639.600 ;
        RECT 845.100 627.000 846.900 637.500 ;
        RECT 848.100 627.600 849.900 638.400 ;
        RECT 863.100 627.600 864.900 639.600 ;
        RECT 866.100 638.700 873.900 639.600 ;
        RECT 866.100 627.600 867.900 638.700 ;
        RECT 869.100 627.000 870.900 637.800 ;
        RECT 872.100 627.600 873.900 638.700 ;
        RECT 896.100 634.800 897.000 646.950 ;
        RECT 911.100 645.150 912.900 646.950 ;
        RECT 890.400 633.900 897.000 634.800 ;
        RECT 890.400 633.600 891.900 633.900 ;
        RECT 887.100 627.000 888.900 633.600 ;
        RECT 890.100 627.600 891.900 633.600 ;
        RECT 896.100 633.600 897.000 633.900 ;
        RECT 914.100 633.600 915.300 646.950 ;
        RECT 927.000 634.800 927.900 646.950 ;
        RECT 932.100 645.150 933.900 646.950 ;
        RECT 928.950 642.450 931.050 643.050 ;
        RECT 937.950 642.450 940.050 643.050 ;
        RECT 928.950 641.550 940.050 642.450 ;
        RECT 928.950 640.950 931.050 641.550 ;
        RECT 937.950 640.950 940.050 641.550 ;
        RECT 927.000 633.900 933.600 634.800 ;
        RECT 927.000 633.600 927.900 633.900 ;
        RECT 893.100 627.000 894.900 633.000 ;
        RECT 896.100 627.600 897.900 633.600 ;
        RECT 911.100 627.000 912.900 633.600 ;
        RECT 914.100 627.600 915.900 633.600 ;
        RECT 926.100 627.600 927.900 633.600 ;
        RECT 932.100 633.600 933.600 633.900 ;
        RECT 929.100 627.000 930.900 633.000 ;
        RECT 932.100 627.600 933.900 633.600 ;
        RECT 935.100 627.000 936.900 633.600 ;
        RECT 14.100 617.400 15.900 624.000 ;
        RECT 17.100 617.400 18.900 623.400 ;
        RECT 20.100 617.400 21.900 624.000 ;
        RECT 32.700 617.400 34.500 624.000 ;
        RECT 9.000 606.450 13.050 607.050 ;
        RECT 8.550 604.950 13.050 606.450 ;
        RECT 8.550 601.050 9.450 604.950 ;
        RECT 17.700 604.050 18.900 617.400 ;
        RECT 33.000 614.100 34.800 615.900 ;
        RECT 22.950 612.450 25.050 613.050 ;
        RECT 31.950 612.450 34.050 613.050 ;
        RECT 35.700 612.900 37.500 623.400 ;
        RECT 22.950 611.550 34.050 612.450 ;
        RECT 22.950 610.950 25.050 611.550 ;
        RECT 31.950 610.950 34.050 611.550 ;
        RECT 35.100 611.400 37.500 612.900 ;
        RECT 40.800 611.400 42.600 624.000 ;
        RECT 56.400 611.400 58.200 624.000 ;
        RECT 61.500 612.900 63.300 623.400 ;
        RECT 64.500 617.400 66.300 624.000 ;
        RECT 80.100 617.400 81.900 623.400 ;
        RECT 83.100 617.400 84.900 624.000 ;
        RECT 64.200 614.100 66.000 615.900 ;
        RECT 61.500 611.400 63.900 612.900 ;
        RECT 35.100 604.050 36.300 611.400 ;
        RECT 37.950 609.450 40.050 610.200 ;
        RECT 49.950 609.450 52.050 610.050 ;
        RECT 58.950 609.450 61.050 609.900 ;
        RECT 37.950 608.550 61.050 609.450 ;
        RECT 37.950 608.100 40.050 608.550 ;
        RECT 49.950 607.950 52.050 608.550 ;
        RECT 58.950 607.800 61.050 608.550 ;
        RECT 41.100 604.050 42.900 605.850 ;
        RECT 56.100 604.050 57.900 605.850 ;
        RECT 62.700 604.050 63.900 611.400 ;
        RECT 67.950 606.450 70.050 607.050 ;
        RECT 67.950 605.550 75.450 606.450 ;
        RECT 67.950 604.950 70.050 605.550 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 19.950 601.950 22.050 604.050 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 8.550 599.550 13.050 601.050 ;
        RECT 14.100 600.150 15.900 601.950 ;
        RECT 9.000 598.950 13.050 599.550 ;
        RECT 17.700 596.700 18.900 601.950 ;
        RECT 19.950 600.150 21.750 601.950 ;
        RECT 32.100 600.150 33.900 601.950 ;
        RECT 35.100 597.600 36.300 601.950 ;
        RECT 38.100 600.150 39.900 601.950 ;
        RECT 59.100 600.150 60.900 601.950 ;
        RECT 14.700 595.800 18.900 596.700 ;
        RECT 32.700 596.700 36.300 597.600 ;
        RECT 62.700 597.600 63.900 601.950 ;
        RECT 65.100 600.150 66.900 601.950 ;
        RECT 74.550 601.050 75.450 605.550 ;
        RECT 80.700 604.050 81.900 617.400 ;
        RECT 95.100 612.300 96.900 623.400 ;
        RECT 98.100 613.200 99.900 624.000 ;
        RECT 101.100 612.300 102.900 623.400 ;
        RECT 95.100 611.400 102.900 612.300 ;
        RECT 104.100 611.400 105.900 623.400 ;
        RECT 116.100 617.400 117.900 624.000 ;
        RECT 119.100 617.400 120.900 623.400 ;
        RECT 134.700 617.400 136.500 624.000 ;
        RECT 88.950 607.950 91.050 610.050 ;
        RECT 83.100 604.050 84.900 605.850 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 74.550 599.550 79.050 601.050 ;
        RECT 75.000 598.950 79.050 599.550 ;
        RECT 62.700 596.700 66.300 597.600 ;
        RECT 14.700 588.600 16.500 595.800 ;
        RECT 32.700 594.600 33.900 596.700 ;
        RECT 19.800 588.000 21.600 594.600 ;
        RECT 32.100 588.600 33.900 594.600 ;
        RECT 35.100 593.700 42.900 595.050 ;
        RECT 35.100 588.600 36.900 593.700 ;
        RECT 38.100 588.000 39.900 592.800 ;
        RECT 41.100 588.600 42.900 593.700 ;
        RECT 56.100 593.700 63.900 595.050 ;
        RECT 56.100 588.600 57.900 593.700 ;
        RECT 59.100 588.000 60.900 592.800 ;
        RECT 62.100 588.600 63.900 593.700 ;
        RECT 65.100 594.600 66.300 596.700 ;
        RECT 65.100 588.600 66.900 594.600 ;
        RECT 80.700 591.600 81.900 601.950 ;
        RECT 89.550 601.050 90.450 607.950 ;
        RECT 98.250 604.050 100.050 605.850 ;
        RECT 104.700 604.050 105.600 611.400 ;
        RECT 106.950 606.450 111.000 607.050 ;
        RECT 106.950 604.950 111.450 606.450 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 85.950 599.550 90.450 601.050 ;
        RECT 95.100 600.150 96.900 601.950 ;
        RECT 101.250 600.150 103.050 601.950 ;
        RECT 85.950 598.950 90.000 599.550 ;
        RECT 104.700 594.600 105.600 601.950 ;
        RECT 110.550 601.050 111.450 604.950 ;
        RECT 116.100 604.050 117.900 605.850 ;
        RECT 119.100 604.050 120.300 617.400 ;
        RECT 135.000 614.100 136.800 615.900 ;
        RECT 137.700 612.900 139.500 623.400 ;
        RECT 137.100 611.400 139.500 612.900 ;
        RECT 142.800 611.400 144.600 624.000 ;
        RECT 155.100 617.400 156.900 624.000 ;
        RECT 158.100 617.400 159.900 623.400 ;
        RECT 161.100 617.400 162.900 624.000 ;
        RECT 173.700 617.400 175.500 624.000 ;
        RECT 137.100 604.050 138.300 611.400 ;
        RECT 143.100 604.050 144.900 605.850 ;
        RECT 158.100 604.050 159.300 617.400 ;
        RECT 174.000 614.100 175.800 615.900 ;
        RECT 176.700 612.900 178.500 623.400 ;
        RECT 176.100 611.400 178.500 612.900 ;
        RECT 181.800 611.400 183.600 624.000 ;
        RECT 197.400 611.400 199.200 624.000 ;
        RECT 202.500 612.900 204.300 623.400 ;
        RECT 205.500 617.400 207.300 624.000 ;
        RECT 221.700 617.400 223.500 624.000 ;
        RECT 205.200 614.100 207.000 615.900 ;
        RECT 222.000 614.100 223.800 615.900 ;
        RECT 202.500 611.400 204.900 612.900 ;
        RECT 168.000 606.450 172.050 607.050 ;
        RECT 167.550 604.950 172.050 606.450 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 154.950 601.950 157.050 604.050 ;
        RECT 157.950 601.950 160.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 109.950 598.950 112.050 601.050 ;
        RECT 80.100 588.600 81.900 591.600 ;
        RECT 83.100 588.000 84.900 591.600 ;
        RECT 96.000 588.000 97.800 594.600 ;
        RECT 100.500 593.400 105.600 594.600 ;
        RECT 100.500 588.600 102.300 593.400 ;
        RECT 119.100 591.600 120.300 601.950 ;
        RECT 134.100 600.150 135.900 601.950 ;
        RECT 137.100 597.600 138.300 601.950 ;
        RECT 140.100 600.150 141.900 601.950 ;
        RECT 155.250 600.150 157.050 601.950 ;
        RECT 134.700 596.700 138.300 597.600 ;
        RECT 158.100 596.700 159.300 601.950 ;
        RECT 161.100 600.150 162.900 601.950 ;
        RECT 167.550 601.050 168.450 604.950 ;
        RECT 176.100 604.050 177.300 611.400 ;
        RECT 184.950 606.450 189.000 607.050 ;
        RECT 182.100 604.050 183.900 605.850 ;
        RECT 184.950 604.950 189.450 606.450 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 175.950 601.950 178.050 604.050 ;
        RECT 178.950 601.950 181.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 163.950 599.550 168.450 601.050 ;
        RECT 173.100 600.150 174.900 601.950 ;
        RECT 163.950 598.950 168.000 599.550 ;
        RECT 176.100 597.600 177.300 601.950 ;
        RECT 179.100 600.150 180.900 601.950 ;
        RECT 188.550 601.050 189.450 604.950 ;
        RECT 197.100 604.050 198.900 605.850 ;
        RECT 203.700 604.050 204.900 611.400 ;
        RECT 205.950 612.450 208.050 613.050 ;
        RECT 217.950 612.450 220.050 613.050 ;
        RECT 224.700 612.900 226.500 623.400 ;
        RECT 205.950 611.550 220.050 612.450 ;
        RECT 205.950 610.950 208.050 611.550 ;
        RECT 217.950 610.950 220.050 611.550 ;
        RECT 224.100 611.400 226.500 612.900 ;
        RECT 229.800 611.400 231.600 624.000 ;
        RECT 242.100 612.600 243.900 623.400 ;
        RECT 245.100 613.500 246.900 624.000 ;
        RECT 248.100 622.500 255.900 623.400 ;
        RECT 248.100 612.600 249.900 622.500 ;
        RECT 242.100 611.700 249.900 612.600 ;
        RECT 208.950 606.450 211.050 607.050 ;
        RECT 208.950 605.550 216.450 606.450 ;
        RECT 208.950 604.950 211.050 605.550 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 184.950 599.550 189.450 601.050 ;
        RECT 200.100 600.150 201.900 601.950 ;
        RECT 184.950 598.950 189.000 599.550 ;
        RECT 173.700 596.700 177.300 597.600 ;
        RECT 203.700 597.600 204.900 601.950 ;
        RECT 206.100 600.150 207.900 601.950 ;
        RECT 215.550 601.050 216.450 605.550 ;
        RECT 224.100 604.050 225.300 611.400 ;
        RECT 251.100 610.500 252.900 621.600 ;
        RECT 254.100 611.400 255.900 622.500 ;
        RECT 269.100 617.400 270.900 623.400 ;
        RECT 272.100 617.400 273.900 624.000 ;
        RECT 287.100 617.400 288.900 624.000 ;
        RECT 290.100 617.400 291.900 623.400 ;
        RECT 302.100 617.400 303.900 624.000 ;
        RECT 305.100 617.400 306.900 623.400 ;
        RECT 308.100 617.400 309.900 624.000 ;
        RECT 323.100 617.400 324.900 624.000 ;
        RECT 326.100 617.400 327.900 623.400 ;
        RECT 329.100 617.400 330.900 624.000 ;
        RECT 341.700 617.400 343.500 624.000 ;
        RECT 248.100 609.600 252.900 610.500 ;
        RECT 232.950 606.450 237.000 607.050 ;
        RECT 230.100 604.050 231.900 605.850 ;
        RECT 232.950 604.950 237.450 606.450 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 226.950 601.950 229.050 604.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 215.550 599.550 220.050 601.050 ;
        RECT 221.100 600.150 222.900 601.950 ;
        RECT 216.000 598.950 220.050 599.550 ;
        RECT 224.100 597.600 225.300 601.950 ;
        RECT 227.100 600.150 228.900 601.950 ;
        RECT 236.550 601.050 237.450 604.950 ;
        RECT 245.250 604.050 247.050 605.850 ;
        RECT 248.100 604.050 249.000 609.600 ;
        RECT 251.100 604.050 252.900 605.850 ;
        RECT 269.700 604.050 270.900 617.400 ;
        RECT 282.000 606.450 286.050 607.050 ;
        RECT 272.100 604.050 273.900 605.850 ;
        RECT 281.550 604.950 286.050 606.450 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 232.950 599.550 237.450 601.050 ;
        RECT 242.250 600.150 244.050 601.950 ;
        RECT 232.950 598.950 237.000 599.550 ;
        RECT 203.700 596.700 207.300 597.600 ;
        RECT 134.700 594.600 135.900 596.700 ;
        RECT 158.100 595.800 162.300 596.700 ;
        RECT 103.500 588.000 105.300 591.600 ;
        RECT 116.100 588.000 117.900 591.600 ;
        RECT 119.100 588.600 120.900 591.600 ;
        RECT 134.100 588.600 135.900 594.600 ;
        RECT 137.100 593.700 144.900 595.050 ;
        RECT 137.100 588.600 138.900 593.700 ;
        RECT 140.100 588.000 141.900 592.800 ;
        RECT 143.100 588.600 144.900 593.700 ;
        RECT 155.400 588.000 157.200 594.600 ;
        RECT 160.500 588.600 162.300 595.800 ;
        RECT 173.700 594.600 174.900 596.700 ;
        RECT 173.100 588.600 174.900 594.600 ;
        RECT 176.100 593.700 183.900 595.050 ;
        RECT 176.100 588.600 177.900 593.700 ;
        RECT 179.100 588.000 180.900 592.800 ;
        RECT 182.100 588.600 183.900 593.700 ;
        RECT 197.100 593.700 204.900 595.050 ;
        RECT 197.100 588.600 198.900 593.700 ;
        RECT 200.100 588.000 201.900 592.800 ;
        RECT 203.100 588.600 204.900 593.700 ;
        RECT 206.100 594.600 207.300 596.700 ;
        RECT 221.700 596.700 225.300 597.600 ;
        RECT 221.700 594.600 222.900 596.700 ;
        RECT 206.100 588.600 207.900 594.600 ;
        RECT 221.100 588.600 222.900 594.600 ;
        RECT 224.100 593.700 231.900 595.050 ;
        RECT 248.100 594.600 249.300 601.950 ;
        RECT 254.100 600.150 255.900 601.950 ;
        RECT 250.950 597.450 253.050 598.050 ;
        RECT 265.950 597.450 268.050 598.050 ;
        RECT 250.950 596.550 268.050 597.450 ;
        RECT 250.950 595.950 253.050 596.550 ;
        RECT 265.950 595.950 268.050 596.550 ;
        RECT 224.100 588.600 225.900 593.700 ;
        RECT 227.100 588.000 228.900 592.800 ;
        RECT 230.100 588.600 231.900 593.700 ;
        RECT 242.700 588.000 244.500 594.600 ;
        RECT 247.200 588.600 249.000 594.600 ;
        RECT 251.700 588.000 253.500 594.600 ;
        RECT 269.700 591.600 270.900 601.950 ;
        RECT 274.950 600.450 277.050 601.050 ;
        RECT 281.550 600.450 282.450 604.950 ;
        RECT 287.100 604.050 288.900 605.850 ;
        RECT 290.100 604.050 291.300 617.400 ;
        RECT 292.950 606.450 297.000 607.050 ;
        RECT 292.950 604.950 297.450 606.450 ;
        RECT 286.950 601.950 289.050 604.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 274.950 599.550 282.450 600.450 ;
        RECT 274.950 598.950 277.050 599.550 ;
        RECT 290.100 591.600 291.300 601.950 ;
        RECT 296.550 601.050 297.450 604.950 ;
        RECT 305.100 604.050 306.300 617.400 ;
        RECT 326.700 604.050 327.900 617.400 ;
        RECT 342.000 614.100 343.800 615.900 ;
        RECT 344.700 612.900 346.500 623.400 ;
        RECT 344.100 611.400 346.500 612.900 ;
        RECT 349.800 611.400 351.600 624.000 ;
        RECT 362.100 617.400 363.900 624.000 ;
        RECT 365.100 617.400 366.900 623.400 ;
        RECT 368.100 617.400 369.900 624.000 ;
        RECT 336.000 606.450 340.050 607.050 ;
        RECT 335.550 604.950 340.050 606.450 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 307.950 601.950 310.050 604.050 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 296.550 599.550 301.050 601.050 ;
        RECT 302.250 600.150 304.050 601.950 ;
        RECT 297.000 598.950 301.050 599.550 ;
        RECT 305.100 596.700 306.300 601.950 ;
        RECT 308.100 600.150 309.900 601.950 ;
        RECT 323.100 600.150 324.900 601.950 ;
        RECT 326.700 596.700 327.900 601.950 ;
        RECT 328.950 600.150 330.750 601.950 ;
        RECT 335.550 600.450 336.450 604.950 ;
        RECT 344.100 604.050 345.300 611.400 ;
        RECT 350.100 604.050 351.900 605.850 ;
        RECT 365.700 604.050 366.900 617.400 ;
        RECT 383.100 612.300 384.900 623.400 ;
        RECT 386.100 613.200 387.900 624.000 ;
        RECT 389.100 612.300 390.900 623.400 ;
        RECT 383.100 611.400 390.900 612.300 ;
        RECT 392.100 611.400 393.900 623.400 ;
        RECT 407.100 611.400 408.900 624.000 ;
        RECT 410.100 611.400 411.900 623.400 ;
        RECT 413.100 611.400 414.900 624.000 ;
        RECT 428.400 611.400 430.200 624.000 ;
        RECT 433.500 612.900 435.300 623.400 ;
        RECT 436.500 617.400 438.300 624.000 ;
        RECT 440.700 617.400 442.500 624.000 ;
        RECT 443.700 617.400 445.500 623.400 ;
        RECT 447.000 617.400 448.800 624.000 ;
        RECT 450.000 617.400 451.800 623.400 ;
        RECT 453.000 617.400 454.800 624.000 ;
        RECT 456.000 617.400 457.800 623.400 ;
        RECT 459.000 617.400 460.800 624.000 ;
        RECT 462.000 620.400 463.800 623.400 ;
        RECT 465.000 620.400 466.800 623.400 ;
        RECT 468.000 620.400 469.800 623.400 ;
        RECT 461.700 618.300 463.800 620.400 ;
        RECT 464.700 618.300 466.800 620.400 ;
        RECT 467.700 618.300 469.800 620.400 ;
        RECT 471.000 617.400 472.800 623.400 ;
        RECT 474.000 617.400 475.800 624.000 ;
        RECT 436.200 614.100 438.000 615.900 ;
        RECT 433.500 611.400 435.900 612.900 ;
        RECT 386.250 604.050 388.050 605.850 ;
        RECT 392.700 604.050 393.600 611.400 ;
        RECT 410.550 604.050 411.600 611.400 ;
        RECT 412.950 609.450 415.050 610.050 ;
        RECT 430.950 609.450 433.050 610.200 ;
        RECT 412.950 608.550 433.050 609.450 ;
        RECT 412.950 607.950 415.050 608.550 ;
        RECT 430.950 608.100 433.050 608.550 ;
        RECT 428.100 604.050 429.900 605.850 ;
        RECT 434.700 604.050 435.900 611.400 ;
        RECT 444.000 607.050 445.500 617.400 ;
        RECT 450.000 616.500 451.200 617.400 ;
        RECT 443.100 604.950 445.500 607.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 407.400 601.950 411.600 604.050 ;
        RECT 412.500 601.950 414.600 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 332.550 599.550 336.450 600.450 ;
        RECT 341.100 600.150 342.900 601.950 ;
        RECT 332.550 598.050 333.450 599.550 ;
        RECT 305.100 595.800 309.300 596.700 ;
        RECT 269.100 588.600 270.900 591.600 ;
        RECT 272.100 588.000 273.900 591.600 ;
        RECT 287.100 588.000 288.900 591.600 ;
        RECT 290.100 588.600 291.900 591.600 ;
        RECT 302.400 588.000 304.200 594.600 ;
        RECT 307.500 588.600 309.300 595.800 ;
        RECT 323.700 595.800 327.900 596.700 ;
        RECT 328.950 596.550 333.450 598.050 ;
        RECT 344.100 597.600 345.300 601.950 ;
        RECT 347.100 600.150 348.900 601.950 ;
        RECT 362.100 600.150 363.900 601.950 ;
        RECT 341.700 596.700 345.300 597.600 ;
        RECT 365.700 596.700 366.900 601.950 ;
        RECT 367.950 600.150 369.750 601.950 ;
        RECT 383.100 600.150 384.900 601.950 ;
        RECT 389.250 600.150 391.050 601.950 ;
        RECT 328.950 595.950 333.000 596.550 ;
        RECT 323.700 588.600 325.500 595.800 ;
        RECT 341.700 594.600 342.900 596.700 ;
        RECT 362.700 595.800 366.900 596.700 ;
        RECT 328.800 588.000 330.600 594.600 ;
        RECT 341.100 588.600 342.900 594.600 ;
        RECT 344.100 593.700 351.900 595.050 ;
        RECT 344.100 588.600 345.900 593.700 ;
        RECT 347.100 588.000 348.900 592.800 ;
        RECT 350.100 588.600 351.900 593.700 ;
        RECT 362.700 588.600 364.500 595.800 ;
        RECT 392.700 594.600 393.600 601.950 ;
        RECT 410.550 594.600 411.600 601.950 ;
        RECT 412.800 600.150 414.600 601.950 ;
        RECT 415.950 600.450 418.050 601.050 ;
        RECT 424.950 600.450 427.050 601.050 ;
        RECT 415.950 599.550 427.050 600.450 ;
        RECT 431.100 600.150 432.900 601.950 ;
        RECT 415.950 598.950 418.050 599.550 ;
        RECT 424.950 598.950 427.050 599.550 ;
        RECT 434.700 597.600 435.900 601.950 ;
        RECT 437.100 600.150 438.900 601.950 ;
        RECT 434.700 596.700 438.300 597.600 ;
        RECT 367.800 588.000 369.600 594.600 ;
        RECT 384.000 588.000 385.800 594.600 ;
        RECT 388.500 593.400 393.600 594.600 ;
        RECT 388.500 588.600 390.300 593.400 ;
        RECT 391.500 588.000 393.300 591.600 ;
        RECT 407.100 588.000 408.900 594.600 ;
        RECT 410.100 588.600 411.900 594.600 ;
        RECT 413.100 588.000 414.900 594.600 ;
        RECT 428.100 593.700 435.900 595.050 ;
        RECT 428.100 588.600 429.900 593.700 ;
        RECT 431.100 588.000 432.900 592.800 ;
        RECT 434.100 588.600 435.900 593.700 ;
        RECT 437.100 594.600 438.300 596.700 ;
        RECT 437.100 588.600 438.900 594.600 ;
        RECT 444.000 591.600 445.500 604.950 ;
        RECT 440.700 588.000 442.500 591.600 ;
        RECT 443.700 588.600 445.500 591.600 ;
        RECT 447.300 615.600 451.200 616.500 ;
        RECT 447.300 612.300 448.200 615.600 ;
        RECT 452.100 614.400 453.900 615.000 ;
        RECT 456.600 614.400 457.800 617.400 ;
        RECT 464.700 616.500 466.800 617.400 ;
        RECT 458.700 615.300 466.800 616.500 ;
        RECT 458.700 614.700 460.500 615.300 ;
        RECT 452.100 613.200 457.800 614.400 ;
        RECT 470.100 613.500 472.800 617.400 ;
        RECT 477.000 615.900 478.800 623.400 ;
        RECT 480.900 617.400 482.700 624.000 ;
        RECT 483.900 617.400 485.700 623.400 ;
        RECT 486.900 620.400 488.700 623.400 ;
        RECT 489.900 620.400 491.700 623.400 ;
        RECT 486.600 618.300 488.700 620.400 ;
        RECT 489.600 618.300 491.700 620.400 ;
        RECT 493.500 617.400 495.300 624.000 ;
        RECT 475.500 613.800 478.800 615.900 ;
        RECT 484.200 615.300 486.300 617.400 ;
        RECT 496.500 614.400 498.300 623.400 ;
        RECT 499.500 617.400 501.300 624.000 ;
        RECT 502.500 618.300 504.300 623.400 ;
        RECT 502.500 617.400 504.600 618.300 ;
        RECT 505.500 617.400 507.300 624.000 ;
        RECT 509.700 617.400 511.500 624.000 ;
        RECT 512.700 617.400 514.500 623.400 ;
        RECT 516.000 617.400 517.800 624.000 ;
        RECT 519.000 617.400 520.800 623.400 ;
        RECT 522.000 617.400 523.800 624.000 ;
        RECT 525.000 617.400 526.800 623.400 ;
        RECT 528.000 617.400 529.800 624.000 ;
        RECT 531.000 620.400 532.800 623.400 ;
        RECT 534.000 620.400 535.800 623.400 ;
        RECT 537.000 620.400 538.800 623.400 ;
        RECT 530.700 618.300 532.800 620.400 ;
        RECT 533.700 618.300 535.800 620.400 ;
        RECT 536.700 618.300 538.800 620.400 ;
        RECT 540.000 617.400 541.800 623.400 ;
        RECT 543.000 617.400 544.800 624.000 ;
        RECT 503.700 616.500 504.600 617.400 ;
        RECT 503.700 615.600 507.300 616.500 ;
        RECT 501.000 614.400 502.800 614.700 ;
        RECT 461.700 612.300 463.800 613.500 ;
        RECT 447.300 611.400 463.800 612.300 ;
        RECT 467.100 612.600 469.200 613.500 ;
        RECT 483.600 613.200 502.800 614.400 ;
        RECT 483.600 612.600 484.800 613.200 ;
        RECT 501.000 612.900 502.800 613.200 ;
        RECT 467.100 611.400 484.800 612.600 ;
        RECT 487.500 611.700 489.600 612.300 ;
        RECT 497.700 611.700 499.500 612.300 ;
        RECT 447.300 594.600 448.200 611.400 ;
        RECT 487.500 610.500 499.500 611.700 ;
        RECT 449.100 609.300 484.800 610.500 ;
        RECT 487.500 610.200 489.600 610.500 ;
        RECT 449.100 608.700 450.900 609.300 ;
        RECT 483.600 608.700 484.800 609.300 ;
        RECT 452.100 604.950 454.200 607.050 ;
        RECT 452.700 602.100 454.200 604.950 ;
        RECT 456.300 604.800 461.400 606.600 ;
        RECT 460.500 603.300 461.400 604.800 ;
        RECT 464.100 606.300 465.900 608.100 ;
        RECT 470.100 607.800 472.200 608.100 ;
        RECT 483.600 607.800 497.100 608.700 ;
        RECT 464.100 605.100 465.000 606.300 ;
        RECT 470.100 606.000 474.000 607.800 ;
        RECT 475.500 606.300 477.600 607.200 ;
        RECT 495.300 607.050 497.100 607.800 ;
        RECT 475.500 605.100 486.600 606.300 ;
        RECT 495.300 605.250 499.200 607.050 ;
        RECT 464.100 604.200 477.600 605.100 ;
        RECT 484.800 604.500 486.600 605.100 ;
        RECT 497.100 604.950 499.200 605.250 ;
        RECT 503.100 604.950 505.200 607.050 ;
        RECT 503.100 603.300 504.900 604.950 ;
        RECT 460.500 602.100 504.900 603.300 ;
        RECT 452.700 600.600 459.300 602.100 ;
        RECT 449.100 597.900 456.900 599.700 ;
        RECT 457.800 599.100 474.900 600.600 ;
        RECT 472.800 598.500 474.900 599.100 ;
        RECT 479.100 600.000 481.200 601.050 ;
        RECT 479.100 599.100 484.200 600.000 ;
        RECT 487.800 599.400 489.600 601.200 ;
        RECT 506.100 599.400 507.300 615.600 ;
        RECT 513.000 607.050 514.500 617.400 ;
        RECT 519.000 616.500 520.200 617.400 ;
        RECT 512.100 604.950 514.500 607.050 ;
        RECT 479.100 598.950 481.200 599.100 ;
        RECT 455.400 594.600 456.900 597.900 ;
        RECT 473.100 596.700 474.900 598.500 ;
        RECT 482.400 598.200 484.200 599.100 ;
        RECT 488.700 596.400 489.600 599.400 ;
        RECT 490.500 598.200 507.300 599.400 ;
        RECT 490.500 597.300 492.600 598.200 ;
        RECT 501.300 596.700 503.100 597.300 ;
        RECT 461.100 594.600 467.700 596.400 ;
        RECT 482.400 595.200 489.600 596.400 ;
        RECT 494.700 595.500 503.100 596.700 ;
        RECT 482.400 594.600 483.300 595.200 ;
        RECT 485.400 594.600 487.200 595.200 ;
        RECT 494.700 594.600 496.200 595.500 ;
        RECT 506.100 594.600 507.300 598.200 ;
        RECT 447.300 588.600 449.100 594.600 ;
        RECT 452.700 588.000 454.500 594.600 ;
        RECT 455.400 593.400 459.600 594.600 ;
        RECT 457.800 588.600 459.600 593.400 ;
        RECT 461.700 591.600 463.800 593.700 ;
        RECT 464.700 591.600 466.800 593.700 ;
        RECT 467.700 591.600 469.800 593.700 ;
        RECT 470.700 591.600 472.800 593.700 ;
        RECT 476.100 592.500 478.800 594.600 ;
        RECT 480.600 593.400 483.300 594.600 ;
        RECT 480.600 592.500 482.400 593.400 ;
        RECT 462.000 588.600 463.800 591.600 ;
        RECT 465.000 588.600 466.800 591.600 ;
        RECT 468.000 588.600 469.800 591.600 ;
        RECT 471.000 588.600 472.800 591.600 ;
        RECT 474.000 588.000 475.800 591.600 ;
        RECT 477.000 588.600 478.800 592.500 ;
        RECT 484.200 591.600 486.300 593.700 ;
        RECT 487.200 591.600 489.300 593.700 ;
        RECT 490.200 591.600 492.300 593.700 ;
        RECT 481.500 588.000 483.300 591.600 ;
        RECT 484.500 588.600 486.300 591.600 ;
        RECT 487.500 588.600 489.300 591.600 ;
        RECT 490.500 588.600 492.300 591.600 ;
        RECT 494.700 588.600 496.500 594.600 ;
        RECT 500.100 588.000 501.900 594.600 ;
        RECT 505.500 588.600 507.300 594.600 ;
        RECT 513.000 591.600 514.500 604.950 ;
        RECT 509.700 588.000 511.500 591.600 ;
        RECT 512.700 588.600 514.500 591.600 ;
        RECT 516.300 615.600 520.200 616.500 ;
        RECT 516.300 612.300 517.200 615.600 ;
        RECT 521.100 614.400 522.900 615.000 ;
        RECT 525.600 614.400 526.800 617.400 ;
        RECT 533.700 616.500 535.800 617.400 ;
        RECT 527.700 615.300 535.800 616.500 ;
        RECT 527.700 614.700 529.500 615.300 ;
        RECT 521.100 613.200 526.800 614.400 ;
        RECT 539.100 613.500 541.800 617.400 ;
        RECT 546.000 615.900 547.800 623.400 ;
        RECT 549.900 617.400 551.700 624.000 ;
        RECT 552.900 617.400 554.700 623.400 ;
        RECT 555.900 620.400 557.700 623.400 ;
        RECT 558.900 620.400 560.700 623.400 ;
        RECT 555.600 618.300 557.700 620.400 ;
        RECT 558.600 618.300 560.700 620.400 ;
        RECT 562.500 617.400 564.300 624.000 ;
        RECT 544.500 613.800 547.800 615.900 ;
        RECT 553.200 615.300 555.300 617.400 ;
        RECT 565.500 614.400 567.300 623.400 ;
        RECT 568.500 617.400 570.300 624.000 ;
        RECT 571.500 618.300 573.300 623.400 ;
        RECT 571.500 617.400 573.600 618.300 ;
        RECT 574.500 617.400 576.300 624.000 ;
        RECT 577.950 621.450 580.050 622.050 ;
        RECT 586.950 621.450 589.050 622.050 ;
        RECT 577.950 620.550 589.050 621.450 ;
        RECT 577.950 619.950 580.050 620.550 ;
        RECT 586.950 619.950 589.050 620.550 ;
        RECT 572.700 616.500 573.600 617.400 ;
        RECT 572.700 615.600 576.300 616.500 ;
        RECT 570.000 614.400 571.800 614.700 ;
        RECT 530.700 612.300 532.800 613.500 ;
        RECT 516.300 611.400 532.800 612.300 ;
        RECT 536.100 612.600 538.200 613.500 ;
        RECT 552.600 613.200 571.800 614.400 ;
        RECT 552.600 612.600 553.800 613.200 ;
        RECT 570.000 612.900 571.800 613.200 ;
        RECT 536.100 611.400 553.800 612.600 ;
        RECT 556.500 611.700 558.600 612.300 ;
        RECT 566.700 611.700 568.500 612.300 ;
        RECT 516.300 594.600 517.200 611.400 ;
        RECT 556.500 610.500 568.500 611.700 ;
        RECT 518.100 609.300 553.800 610.500 ;
        RECT 556.500 610.200 558.600 610.500 ;
        RECT 518.100 608.700 519.900 609.300 ;
        RECT 552.600 608.700 553.800 609.300 ;
        RECT 521.100 604.950 523.200 607.050 ;
        RECT 521.700 602.100 523.200 604.950 ;
        RECT 525.300 604.800 530.400 606.600 ;
        RECT 529.500 603.300 530.400 604.800 ;
        RECT 533.100 606.300 534.900 608.100 ;
        RECT 539.100 607.800 541.200 608.100 ;
        RECT 552.600 607.800 566.100 608.700 ;
        RECT 533.100 605.100 534.000 606.300 ;
        RECT 539.100 606.000 543.000 607.800 ;
        RECT 544.500 606.300 546.600 607.200 ;
        RECT 564.300 607.050 566.100 607.800 ;
        RECT 544.500 605.100 555.600 606.300 ;
        RECT 564.300 605.250 568.200 607.050 ;
        RECT 533.100 604.200 546.600 605.100 ;
        RECT 553.800 604.500 555.600 605.100 ;
        RECT 566.100 604.950 568.200 605.250 ;
        RECT 572.100 604.950 574.200 607.050 ;
        RECT 572.100 603.300 573.900 604.950 ;
        RECT 529.500 602.100 573.900 603.300 ;
        RECT 521.700 600.600 528.300 602.100 ;
        RECT 518.100 597.900 525.900 599.700 ;
        RECT 526.800 599.100 543.900 600.600 ;
        RECT 541.800 598.500 543.900 599.100 ;
        RECT 548.100 600.000 550.200 601.050 ;
        RECT 548.100 599.100 553.200 600.000 ;
        RECT 556.800 599.400 558.600 601.200 ;
        RECT 575.100 599.400 576.300 615.600 ;
        RECT 590.400 611.400 592.200 624.000 ;
        RECT 595.500 612.900 597.300 623.400 ;
        RECT 598.500 617.400 600.300 624.000 ;
        RECT 598.200 614.100 600.000 615.900 ;
        RECT 595.500 611.400 597.900 612.900 ;
        RECT 614.100 611.400 615.900 624.000 ;
        RECT 619.200 612.600 621.000 623.400 ;
        RECT 617.400 611.400 621.000 612.600 ;
        RECT 633.600 611.400 635.400 624.000 ;
        RECT 638.100 611.400 641.400 623.400 ;
        RECT 644.100 611.400 645.900 624.000 ;
        RECT 659.100 617.400 660.900 624.000 ;
        RECT 662.100 617.400 663.900 623.400 ;
        RECT 665.100 617.400 666.900 624.000 ;
        RECT 590.100 604.050 591.900 605.850 ;
        RECT 596.700 604.050 597.900 611.400 ;
        RECT 609.000 606.450 613.050 607.050 ;
        RECT 608.550 604.950 613.050 606.450 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 593.100 600.150 594.900 601.950 ;
        RECT 548.100 598.950 550.200 599.100 ;
        RECT 524.400 594.600 525.900 597.900 ;
        RECT 542.100 596.700 543.900 598.500 ;
        RECT 551.400 598.200 553.200 599.100 ;
        RECT 557.700 596.400 558.600 599.400 ;
        RECT 559.500 598.200 576.300 599.400 ;
        RECT 559.500 597.300 561.600 598.200 ;
        RECT 570.300 596.700 572.100 597.300 ;
        RECT 530.100 594.600 536.700 596.400 ;
        RECT 551.400 595.200 558.600 596.400 ;
        RECT 563.700 595.500 572.100 596.700 ;
        RECT 551.400 594.600 552.300 595.200 ;
        RECT 554.400 594.600 556.200 595.200 ;
        RECT 563.700 594.600 565.200 595.500 ;
        RECT 575.100 594.600 576.300 598.200 ;
        RECT 596.700 597.600 597.900 601.950 ;
        RECT 599.100 600.150 600.900 601.950 ;
        RECT 608.550 601.050 609.450 604.950 ;
        RECT 614.250 604.050 616.050 605.850 ;
        RECT 617.400 604.050 618.300 611.400 ;
        RECT 625.950 609.450 628.050 610.050 ;
        RECT 634.950 609.450 637.050 610.050 ;
        RECT 625.950 608.550 637.050 609.450 ;
        RECT 625.950 607.950 628.050 608.550 ;
        RECT 634.950 607.950 637.050 608.550 ;
        RECT 620.100 604.050 621.900 605.850 ;
        RECT 632.250 604.050 634.050 605.850 ;
        RECT 639.000 604.050 640.050 611.400 ;
        RECT 654.000 606.450 658.050 607.050 ;
        RECT 644.100 604.050 645.900 605.850 ;
        RECT 653.550 604.950 658.050 606.450 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 608.550 599.550 613.050 601.050 ;
        RECT 609.000 598.950 613.050 599.550 ;
        RECT 596.700 596.700 600.300 597.600 ;
        RECT 516.300 588.600 518.100 594.600 ;
        RECT 521.700 588.000 523.500 594.600 ;
        RECT 524.400 593.400 528.600 594.600 ;
        RECT 526.800 588.600 528.600 593.400 ;
        RECT 530.700 591.600 532.800 593.700 ;
        RECT 533.700 591.600 535.800 593.700 ;
        RECT 536.700 591.600 538.800 593.700 ;
        RECT 539.700 591.600 541.800 593.700 ;
        RECT 545.100 592.500 547.800 594.600 ;
        RECT 549.600 593.400 552.300 594.600 ;
        RECT 549.600 592.500 551.400 593.400 ;
        RECT 531.000 588.600 532.800 591.600 ;
        RECT 534.000 588.600 535.800 591.600 ;
        RECT 537.000 588.600 538.800 591.600 ;
        RECT 540.000 588.600 541.800 591.600 ;
        RECT 543.000 588.000 544.800 591.600 ;
        RECT 546.000 588.600 547.800 592.500 ;
        RECT 553.200 591.600 555.300 593.700 ;
        RECT 556.200 591.600 558.300 593.700 ;
        RECT 559.200 591.600 561.300 593.700 ;
        RECT 550.500 588.000 552.300 591.600 ;
        RECT 553.500 588.600 555.300 591.600 ;
        RECT 556.500 588.600 558.300 591.600 ;
        RECT 559.500 588.600 561.300 591.600 ;
        RECT 563.700 588.600 565.500 594.600 ;
        RECT 569.100 588.000 570.900 594.600 ;
        RECT 574.500 588.600 576.300 594.600 ;
        RECT 590.100 593.700 597.900 595.050 ;
        RECT 590.100 588.600 591.900 593.700 ;
        RECT 593.100 588.000 594.900 592.800 ;
        RECT 596.100 588.600 597.900 593.700 ;
        RECT 599.100 594.600 600.300 596.700 ;
        RECT 599.100 588.600 600.900 594.600 ;
        RECT 617.400 591.600 618.300 601.950 ;
        RECT 635.250 600.150 637.050 601.950 ;
        RECT 639.000 597.300 640.050 601.950 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 640.950 600.150 642.750 601.950 ;
        RECT 653.550 601.050 654.450 604.950 ;
        RECT 662.100 604.050 663.300 617.400 ;
        RECT 680.400 611.400 682.200 624.000 ;
        RECT 685.500 612.900 687.300 623.400 ;
        RECT 688.500 617.400 690.300 624.000 ;
        RECT 701.100 617.400 702.900 624.000 ;
        RECT 704.100 617.400 705.900 623.400 ;
        RECT 707.100 617.400 708.900 624.000 ;
        RECT 722.100 617.400 723.900 624.000 ;
        RECT 725.100 617.400 726.900 623.400 ;
        RECT 737.100 617.400 738.900 624.000 ;
        RECT 740.100 617.400 741.900 623.400 ;
        RECT 755.100 617.400 756.900 624.000 ;
        RECT 758.100 617.400 759.900 623.400 ;
        RECT 770.700 617.400 772.500 624.000 ;
        RECT 688.200 614.100 690.000 615.900 ;
        RECT 685.500 611.400 687.900 612.900 ;
        RECT 670.950 609.450 673.050 610.050 ;
        RECT 682.950 609.450 685.050 610.200 ;
        RECT 670.950 608.550 685.050 609.450 ;
        RECT 670.950 607.950 673.050 608.550 ;
        RECT 682.950 608.100 685.050 608.550 ;
        RECT 680.100 604.050 681.900 605.850 ;
        RECT 686.700 604.050 687.900 611.400 ;
        RECT 704.100 604.050 705.300 617.400 ;
        RECT 722.100 604.050 723.900 605.850 ;
        RECT 725.100 604.050 726.300 617.400 ;
        RECT 737.100 604.050 738.900 605.850 ;
        RECT 740.100 604.050 741.300 617.400 ;
        RECT 755.100 604.050 756.900 605.850 ;
        RECT 758.100 604.050 759.300 617.400 ;
        RECT 771.000 614.100 772.800 615.900 ;
        RECT 773.700 612.900 775.500 623.400 ;
        RECT 773.100 611.400 775.500 612.900 ;
        RECT 778.800 611.400 780.600 624.000 ;
        RECT 794.100 612.300 795.900 623.400 ;
        RECT 797.100 613.200 798.900 624.000 ;
        RECT 800.100 612.300 801.900 623.400 ;
        RECT 794.100 611.400 801.900 612.300 ;
        RECT 803.100 611.400 804.900 623.400 ;
        RECT 818.100 617.400 819.900 624.000 ;
        RECT 821.100 617.400 822.900 623.400 ;
        RECT 824.100 617.400 825.900 624.000 ;
        RECT 839.100 617.400 840.900 624.000 ;
        RECT 842.100 617.400 843.900 623.400 ;
        RECT 845.100 618.000 846.900 624.000 ;
        RECT 773.100 604.050 774.300 611.400 ;
        RECT 784.950 609.450 787.050 610.050 ;
        RECT 799.950 609.450 802.050 610.050 ;
        RECT 784.950 608.550 802.050 609.450 ;
        RECT 784.950 607.950 787.050 608.550 ;
        RECT 799.950 607.950 802.050 608.550 ;
        RECT 779.100 604.050 780.900 605.850 ;
        RECT 797.250 604.050 799.050 605.850 ;
        RECT 803.700 604.050 804.600 611.400 ;
        RECT 821.700 604.050 822.900 617.400 ;
        RECT 842.400 617.100 843.900 617.400 ;
        RECT 848.100 617.400 849.900 623.400 ;
        RECT 863.100 617.400 864.900 623.400 ;
        RECT 866.100 617.400 867.900 624.000 ;
        RECT 848.100 617.100 849.000 617.400 ;
        RECT 842.400 616.200 849.000 617.100 ;
        RECT 842.100 604.050 843.900 605.850 ;
        RECT 848.100 604.050 849.000 616.200 ;
        RECT 858.000 606.450 862.050 607.050 ;
        RECT 857.550 604.950 862.050 606.450 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 721.950 601.950 724.050 604.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 653.550 599.550 658.050 601.050 ;
        RECT 659.250 600.150 661.050 601.950 ;
        RECT 654.000 598.950 658.050 599.550 ;
        RECT 635.700 596.100 640.050 597.300 ;
        RECT 662.100 596.700 663.300 601.950 ;
        RECT 665.100 600.150 666.900 601.950 ;
        RECT 683.100 600.150 684.900 601.950 ;
        RECT 686.700 597.600 687.900 601.950 ;
        RECT 689.100 600.150 690.900 601.950 ;
        RECT 701.250 600.150 703.050 601.950 ;
        RECT 686.700 596.700 690.300 597.600 ;
        RECT 635.700 594.600 636.600 596.100 ;
        RECT 662.100 595.800 666.300 596.700 ;
        RECT 614.100 588.000 615.900 591.600 ;
        RECT 617.100 588.600 618.900 591.600 ;
        RECT 620.100 588.000 621.900 591.600 ;
        RECT 632.100 589.500 633.900 594.600 ;
        RECT 635.100 590.400 636.900 594.600 ;
        RECT 638.100 594.000 645.900 594.900 ;
        RECT 638.100 589.500 639.900 594.000 ;
        RECT 632.100 588.600 639.900 589.500 ;
        RECT 641.100 588.000 642.900 593.100 ;
        RECT 644.100 588.600 645.900 594.000 ;
        RECT 659.400 588.000 661.200 594.600 ;
        RECT 664.500 588.600 666.300 595.800 ;
        RECT 680.100 593.700 687.900 595.050 ;
        RECT 680.100 588.600 681.900 593.700 ;
        RECT 683.100 588.000 684.900 592.800 ;
        RECT 686.100 588.600 687.900 593.700 ;
        RECT 689.100 594.600 690.300 596.700 ;
        RECT 704.100 596.700 705.300 601.950 ;
        RECT 707.100 600.150 708.900 601.950 ;
        RECT 704.100 595.800 708.300 596.700 ;
        RECT 689.100 588.600 690.900 594.600 ;
        RECT 701.400 588.000 703.200 594.600 ;
        RECT 706.500 588.600 708.300 595.800 ;
        RECT 725.100 591.600 726.300 601.950 ;
        RECT 740.100 591.600 741.300 601.950 ;
        RECT 758.100 591.600 759.300 601.950 ;
        RECT 770.100 600.150 771.900 601.950 ;
        RECT 773.100 597.600 774.300 601.950 ;
        RECT 776.100 600.150 777.900 601.950 ;
        RECT 794.100 600.150 795.900 601.950 ;
        RECT 800.250 600.150 802.050 601.950 ;
        RECT 770.700 596.700 774.300 597.600 ;
        RECT 770.700 594.600 771.900 596.700 ;
        RECT 722.100 588.000 723.900 591.600 ;
        RECT 725.100 588.600 726.900 591.600 ;
        RECT 737.100 588.000 738.900 591.600 ;
        RECT 740.100 588.600 741.900 591.600 ;
        RECT 755.100 588.000 756.900 591.600 ;
        RECT 758.100 588.600 759.900 591.600 ;
        RECT 770.100 588.600 771.900 594.600 ;
        RECT 773.100 593.700 780.900 595.050 ;
        RECT 803.700 594.600 804.600 601.950 ;
        RECT 818.100 600.150 819.900 601.950 ;
        RECT 821.700 596.700 822.900 601.950 ;
        RECT 823.950 600.150 825.750 601.950 ;
        RECT 839.100 600.150 840.900 601.950 ;
        RECT 845.100 600.150 846.900 601.950 ;
        RECT 848.100 598.200 849.000 601.950 ;
        RECT 857.550 601.050 858.450 604.950 ;
        RECT 863.700 604.050 864.900 617.400 ;
        RECT 878.400 611.400 880.200 624.000 ;
        RECT 883.500 612.900 885.300 623.400 ;
        RECT 886.500 617.400 888.300 624.000 ;
        RECT 902.100 622.500 909.900 623.400 ;
        RECT 886.200 614.100 888.000 615.900 ;
        RECT 902.100 613.200 903.900 622.500 ;
        RECT 905.100 613.800 906.900 621.600 ;
        RECT 883.500 611.400 885.900 612.900 ;
        RECT 868.950 606.450 873.000 607.050 ;
        RECT 866.100 604.050 867.900 605.850 ;
        RECT 868.950 604.950 873.450 606.450 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 857.550 599.550 862.050 601.050 ;
        RECT 858.000 598.950 862.050 599.550 ;
        RECT 773.100 588.600 774.900 593.700 ;
        RECT 776.100 588.000 777.900 592.800 ;
        RECT 779.100 588.600 780.900 593.700 ;
        RECT 795.000 588.000 796.800 594.600 ;
        RECT 799.500 593.400 804.600 594.600 ;
        RECT 818.700 595.800 822.900 596.700 ;
        RECT 799.500 588.600 801.300 593.400 ;
        RECT 802.500 588.000 804.300 591.600 ;
        RECT 818.700 588.600 820.500 595.800 ;
        RECT 823.800 588.000 825.600 594.600 ;
        RECT 839.100 588.000 840.900 597.600 ;
        RECT 845.700 597.000 849.000 598.200 ;
        RECT 845.700 588.600 847.500 597.000 ;
        RECT 850.950 591.450 853.050 592.050 ;
        RECT 859.950 591.450 862.050 592.050 ;
        RECT 863.700 591.600 864.900 601.950 ;
        RECT 872.550 601.050 873.450 604.950 ;
        RECT 878.100 604.050 879.900 605.850 ;
        RECT 884.700 604.050 885.900 611.400 ;
        RECT 905.700 604.050 906.900 613.800 ;
        RECT 908.100 613.800 909.900 622.500 ;
        RECT 911.100 622.500 918.900 623.400 ;
        RECT 911.100 614.700 912.900 622.500 ;
        RECT 914.100 613.800 915.900 621.600 ;
        RECT 908.100 612.900 915.900 613.800 ;
        RECT 917.100 613.500 918.900 622.500 ;
        RECT 920.100 614.400 921.900 624.000 ;
        RECT 923.100 613.500 924.900 623.400 ;
        RECT 917.100 612.600 924.900 613.500 ;
        RECT 910.950 604.050 912.750 605.850 ;
        RECT 920.100 604.050 921.900 605.850 ;
        RECT 877.950 601.950 880.050 604.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 905.400 601.950 907.500 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 920.100 601.950 922.200 604.050 ;
        RECT 868.950 599.550 873.450 601.050 ;
        RECT 881.100 600.150 882.900 601.950 ;
        RECT 868.950 598.950 873.000 599.550 ;
        RECT 884.700 597.600 885.900 601.950 ;
        RECT 887.100 600.150 888.900 601.950 ;
        RECT 884.700 596.700 888.300 597.600 ;
        RECT 865.950 594.450 868.050 594.900 ;
        RECT 874.950 594.450 877.050 595.050 ;
        RECT 865.950 593.550 877.050 594.450 ;
        RECT 865.950 592.800 868.050 593.550 ;
        RECT 874.950 592.950 877.050 593.550 ;
        RECT 878.100 593.700 885.900 595.050 ;
        RECT 850.950 590.550 862.050 591.450 ;
        RECT 850.950 589.950 853.050 590.550 ;
        RECT 859.950 589.950 862.050 590.550 ;
        RECT 863.100 588.600 864.900 591.600 ;
        RECT 866.100 588.000 867.900 591.600 ;
        RECT 878.100 588.600 879.900 593.700 ;
        RECT 881.100 588.000 882.900 592.800 ;
        RECT 884.100 588.600 885.900 593.700 ;
        RECT 887.100 594.600 888.300 596.700 ;
        RECT 887.100 588.600 888.900 594.600 ;
        RECT 905.700 593.400 906.900 601.950 ;
        RECT 914.250 600.150 916.050 601.950 ;
        RECT 910.950 597.450 913.050 597.750 ;
        RECT 934.950 597.450 937.050 598.050 ;
        RECT 910.950 596.550 937.050 597.450 ;
        RECT 910.950 595.650 913.050 596.550 ;
        RECT 934.950 595.950 937.050 596.550 ;
        RECT 905.700 592.500 918.300 593.400 ;
        RECT 910.200 591.600 911.100 592.500 ;
        RECT 917.400 591.600 918.300 592.500 ;
        RECT 910.200 588.600 912.900 591.600 ;
        RECT 914.100 588.000 915.900 591.600 ;
        RECT 917.100 588.600 918.900 591.600 ;
        RECT 920.100 588.000 922.200 591.600 ;
        RECT 14.100 581.400 15.900 584.400 ;
        RECT 17.100 581.400 18.900 585.000 ;
        RECT 14.700 571.050 15.900 581.400 ;
        RECT 29.400 578.400 31.200 585.000 ;
        RECT 34.500 577.200 36.300 584.400 ;
        RECT 52.500 578.400 54.300 585.000 ;
        RECT 57.000 578.400 58.800 584.400 ;
        RECT 61.500 578.400 63.300 585.000 ;
        RECT 74.400 578.400 76.200 585.000 ;
        RECT 32.100 576.300 36.300 577.200 ;
        RECT 43.950 576.450 46.050 577.050 ;
        RECT 49.950 576.450 52.050 577.050 ;
        RECT 29.250 571.050 31.050 572.850 ;
        RECT 32.100 571.050 33.300 576.300 ;
        RECT 43.950 575.550 52.050 576.450 ;
        RECT 43.950 574.950 46.050 575.550 ;
        RECT 49.950 574.950 52.050 575.550 ;
        RECT 35.100 571.050 36.900 572.850 ;
        RECT 50.100 571.050 51.900 572.850 ;
        RECT 56.700 571.050 57.900 578.400 ;
        RECT 79.500 577.200 81.300 584.400 ;
        RECT 95.100 579.300 96.900 584.400 ;
        RECT 98.100 580.200 99.900 585.000 ;
        RECT 101.100 579.300 102.900 584.400 ;
        RECT 95.100 577.950 102.900 579.300 ;
        RECT 104.100 578.400 105.900 584.400 ;
        RECT 116.100 581.400 117.900 585.000 ;
        RECT 119.100 581.400 120.900 584.400 ;
        RECT 134.100 581.400 135.900 585.000 ;
        RECT 137.100 581.400 138.900 584.400 ;
        RECT 140.100 581.400 141.900 585.000 ;
        RECT 67.950 574.950 70.050 577.050 ;
        RECT 77.100 576.300 81.300 577.200 ;
        RECT 104.100 576.300 105.300 578.400 ;
        RECT 61.950 571.050 63.750 572.850 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 14.700 555.600 15.900 568.950 ;
        RECT 17.100 567.150 18.900 568.950 ;
        RECT 32.100 555.600 33.300 568.950 ;
        RECT 53.100 567.150 54.900 568.950 ;
        RECT 37.950 564.450 40.050 565.050 ;
        RECT 49.950 564.450 52.050 565.050 ;
        RECT 37.950 563.550 52.050 564.450 ;
        RECT 37.950 562.950 40.050 563.550 ;
        RECT 49.950 562.950 52.050 563.550 ;
        RECT 57.000 563.400 57.900 568.950 ;
        RECT 58.950 567.150 60.750 568.950 ;
        RECT 68.550 568.050 69.450 574.950 ;
        RECT 74.250 571.050 76.050 572.850 ;
        RECT 77.100 571.050 78.300 576.300 ;
        RECT 101.700 575.400 105.300 576.300 ;
        RECT 82.950 573.450 85.050 574.050 ;
        RECT 80.100 571.050 81.900 572.850 ;
        RECT 82.950 572.550 90.450 573.450 ;
        RECT 82.950 571.950 85.050 572.550 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 64.950 566.550 69.450 568.050 ;
        RECT 64.950 565.950 69.000 566.550 ;
        RECT 53.100 562.500 57.900 563.400 ;
        RECT 14.100 549.600 15.900 555.600 ;
        RECT 17.100 549.000 18.900 555.600 ;
        RECT 29.100 549.000 30.900 555.600 ;
        RECT 32.100 549.600 33.900 555.600 ;
        RECT 35.100 549.000 36.900 555.600 ;
        RECT 50.100 550.500 51.900 561.600 ;
        RECT 53.100 551.400 54.900 562.500 ;
        RECT 56.100 560.400 63.900 561.300 ;
        RECT 56.100 550.500 57.900 560.400 ;
        RECT 50.100 549.600 57.900 550.500 ;
        RECT 59.100 549.000 60.900 559.500 ;
        RECT 62.100 549.600 63.900 560.400 ;
        RECT 77.100 555.600 78.300 568.950 ;
        RECT 89.550 568.050 90.450 572.550 ;
        RECT 98.100 571.050 99.900 572.850 ;
        RECT 101.700 571.050 102.900 575.400 ;
        RECT 104.100 571.050 105.900 572.850 ;
        RECT 119.100 571.050 120.300 581.400 ;
        RECT 137.700 571.050 138.600 581.400 ;
        RECT 155.100 578.400 156.900 584.400 ;
        RECT 155.700 576.300 156.900 578.400 ;
        RECT 158.100 579.300 159.900 584.400 ;
        RECT 161.100 580.200 162.900 585.000 ;
        RECT 164.100 579.300 165.900 584.400 ;
        RECT 158.100 577.950 165.900 579.300 ;
        RECT 179.700 578.400 181.500 585.000 ;
        RECT 184.200 578.400 186.000 584.400 ;
        RECT 188.700 578.400 190.500 585.000 ;
        RECT 155.700 575.400 159.300 576.300 ;
        RECT 155.100 571.050 156.900 572.850 ;
        RECT 158.100 571.050 159.300 575.400 ;
        RECT 161.100 571.050 162.900 572.850 ;
        RECT 179.250 571.050 181.050 572.850 ;
        RECT 185.100 571.050 186.300 578.400 ;
        RECT 196.950 576.450 201.000 577.050 ;
        RECT 196.950 574.950 201.450 576.450 ;
        RECT 208.500 576.000 210.300 584.400 ;
        RECT 193.950 573.450 198.000 574.050 ;
        RECT 191.100 571.050 192.900 572.850 ;
        RECT 193.950 571.950 198.450 573.450 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 89.550 566.550 94.050 568.050 ;
        RECT 95.100 567.150 96.900 568.950 ;
        RECT 90.000 565.950 94.050 566.550 ;
        RECT 101.700 561.600 102.900 568.950 ;
        RECT 116.100 567.150 117.900 568.950 ;
        RECT 74.100 549.000 75.900 555.600 ;
        RECT 77.100 549.600 78.900 555.600 ;
        RECT 80.100 549.000 81.900 555.600 ;
        RECT 95.400 549.000 97.200 561.600 ;
        RECT 100.500 560.100 102.900 561.600 ;
        RECT 100.500 549.600 102.300 560.100 ;
        RECT 103.200 557.100 105.000 558.900 ;
        RECT 119.100 555.600 120.300 568.950 ;
        RECT 121.950 567.450 124.050 568.050 ;
        RECT 127.950 567.450 130.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 178.950 568.950 181.050 571.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 184.950 568.950 187.050 571.050 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 121.950 567.000 130.050 567.450 ;
        RECT 134.100 567.150 135.900 568.950 ;
        RECT 121.950 566.550 129.450 567.000 ;
        RECT 121.950 565.950 124.050 566.550 ;
        RECT 137.700 561.600 138.600 568.950 ;
        RECT 139.950 567.150 141.750 568.950 ;
        RECT 145.950 567.450 148.050 568.050 ;
        RECT 151.950 567.450 154.050 568.050 ;
        RECT 145.950 566.550 154.050 567.450 ;
        RECT 145.950 565.950 148.050 566.550 ;
        RECT 151.950 565.950 154.050 566.550 ;
        RECT 158.100 561.600 159.300 568.950 ;
        RECT 164.100 567.150 165.900 568.950 ;
        RECT 182.250 567.150 184.050 568.950 ;
        RECT 185.100 563.400 186.000 568.950 ;
        RECT 188.100 567.150 189.900 568.950 ;
        RECT 190.950 564.450 193.050 564.750 ;
        RECT 197.550 564.450 198.450 571.950 ;
        RECT 200.550 568.050 201.450 574.950 ;
        RECT 207.000 574.800 210.300 576.000 ;
        RECT 215.100 575.400 216.900 585.000 ;
        RECT 230.100 578.400 231.900 584.400 ;
        RECT 233.100 579.300 234.900 585.000 ;
        RECT 237.600 578.400 239.400 584.400 ;
        RECT 242.100 579.300 243.900 585.000 ;
        RECT 245.100 578.400 246.900 584.400 ;
        RECT 230.700 576.600 231.900 578.400 ;
        RECT 237.900 576.900 239.100 578.400 ;
        RECT 242.100 577.500 246.900 578.400 ;
        RECT 230.700 575.700 237.000 576.600 ;
        RECT 207.000 571.050 207.900 574.800 ;
        RECT 234.900 573.600 237.000 575.700 ;
        RECT 209.100 571.050 210.900 572.850 ;
        RECT 215.100 571.050 216.900 572.850 ;
        RECT 230.400 571.050 232.200 572.850 ;
        RECT 235.200 571.800 237.000 573.600 ;
        RECT 237.900 574.800 240.900 576.900 ;
        RECT 242.100 576.300 244.200 577.500 ;
        RECT 262.500 576.000 264.300 584.400 ;
        RECT 261.000 574.800 264.300 576.000 ;
        RECT 269.100 575.400 270.900 585.000 ;
        RECT 284.400 578.400 286.200 585.000 ;
        RECT 289.500 577.200 291.300 584.400 ;
        RECT 305.100 581.400 306.900 585.000 ;
        RECT 308.100 581.400 309.900 584.400 ;
        RECT 287.100 576.300 291.300 577.200 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 230.100 570.300 232.200 571.050 ;
        RECT 230.100 568.950 237.000 570.300 ;
        RECT 200.550 566.550 205.050 568.050 ;
        RECT 201.000 565.950 205.050 566.550 ;
        RECT 190.950 563.550 198.450 564.450 ;
        RECT 185.100 562.500 189.900 563.400 ;
        RECT 190.950 562.650 193.050 563.550 ;
        RECT 135.000 560.400 138.600 561.600 ;
        RECT 103.500 549.000 105.300 555.600 ;
        RECT 116.100 549.000 117.900 555.600 ;
        RECT 119.100 549.600 120.900 555.600 ;
        RECT 135.000 549.600 136.800 560.400 ;
        RECT 140.100 549.000 141.900 561.600 ;
        RECT 158.100 560.100 160.500 561.600 ;
        RECT 156.000 557.100 157.800 558.900 ;
        RECT 155.700 549.000 157.500 555.600 ;
        RECT 158.700 549.600 160.500 560.100 ;
        RECT 163.800 549.000 165.600 561.600 ;
        RECT 179.100 560.400 186.900 561.300 ;
        RECT 179.100 549.600 180.900 560.400 ;
        RECT 182.100 549.000 183.900 559.500 ;
        RECT 185.100 550.500 186.900 560.400 ;
        RECT 188.100 551.400 189.900 562.500 ;
        RECT 191.100 550.500 192.900 561.600 ;
        RECT 207.000 556.800 207.900 568.950 ;
        RECT 212.100 567.150 213.900 568.950 ;
        RECT 235.200 568.500 237.000 568.950 ;
        RECT 237.900 569.100 239.100 574.800 ;
        RECT 240.000 571.800 242.100 573.900 ;
        RECT 240.300 570.000 242.100 571.800 ;
        RECT 261.000 571.050 261.900 574.800 ;
        RECT 263.100 571.050 264.900 572.850 ;
        RECT 269.100 571.050 270.900 572.850 ;
        RECT 284.250 571.050 286.050 572.850 ;
        RECT 287.100 571.050 288.300 576.300 ;
        RECT 290.100 571.050 291.900 572.850 ;
        RECT 308.100 571.050 309.300 581.400 ;
        RECT 323.100 578.400 324.900 584.400 ;
        RECT 326.100 578.400 327.900 585.000 ;
        RECT 329.100 581.400 330.900 584.400 ;
        RECT 332.700 581.400 334.500 585.000 ;
        RECT 335.700 581.400 337.500 584.400 ;
        RECT 319.950 571.950 322.050 574.050 ;
        RECT 237.900 568.200 240.300 569.100 ;
        RECT 238.800 568.050 240.300 568.200 ;
        RECT 244.800 568.950 246.900 571.050 ;
        RECT 259.950 568.950 262.050 571.050 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 226.950 565.950 229.050 568.050 ;
        RECT 227.550 559.050 228.450 565.950 ;
        RECT 234.000 565.500 237.900 567.300 ;
        RECT 235.800 565.200 237.900 565.500 ;
        RECT 238.800 565.950 240.900 568.050 ;
        RECT 244.800 567.150 246.600 568.950 ;
        RECT 238.800 564.000 239.700 565.950 ;
        RECT 232.500 561.600 234.600 563.700 ;
        RECT 238.200 562.950 239.700 564.000 ;
        RECT 238.200 561.600 239.400 562.950 ;
        RECT 230.100 560.700 234.600 561.600 ;
        RECT 226.950 556.950 229.050 559.050 ;
        RECT 207.000 555.900 213.600 556.800 ;
        RECT 207.000 555.600 207.900 555.900 ;
        RECT 185.100 549.600 192.900 550.500 ;
        RECT 206.100 549.600 207.900 555.600 ;
        RECT 212.100 555.600 213.600 555.900 ;
        RECT 209.100 549.000 210.900 555.000 ;
        RECT 212.100 549.600 213.900 555.600 ;
        RECT 215.100 549.000 216.900 555.600 ;
        RECT 230.100 549.600 231.900 560.700 ;
        RECT 233.100 549.000 234.900 559.500 ;
        RECT 237.600 549.600 239.400 561.600 ;
        RECT 242.100 561.600 244.200 562.500 ;
        RECT 242.100 560.400 246.900 561.600 ;
        RECT 242.100 549.000 243.900 559.500 ;
        RECT 245.100 549.600 246.900 560.400 ;
        RECT 261.000 556.800 261.900 568.950 ;
        RECT 266.100 567.150 267.900 568.950 ;
        RECT 274.950 567.450 277.050 571.050 ;
        RECT 283.950 568.950 286.050 571.050 ;
        RECT 286.950 568.950 289.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 304.950 568.950 307.050 571.050 ;
        RECT 307.950 568.950 310.050 571.050 ;
        RECT 280.950 567.450 283.050 568.050 ;
        RECT 274.950 567.000 283.050 567.450 ;
        RECT 275.550 566.550 283.050 567.000 ;
        RECT 280.950 565.950 283.050 566.550 ;
        RECT 261.000 555.900 267.600 556.800 ;
        RECT 261.000 555.600 261.900 555.900 ;
        RECT 260.100 549.600 261.900 555.600 ;
        RECT 266.100 555.600 267.600 555.900 ;
        RECT 287.100 555.600 288.300 568.950 ;
        RECT 305.100 567.150 306.900 568.950 ;
        RECT 308.100 555.600 309.300 568.950 ;
        RECT 320.550 568.050 321.450 571.950 ;
        RECT 316.950 566.550 321.450 568.050 ;
        RECT 323.100 571.050 324.300 578.400 ;
        RECT 329.700 577.500 330.900 581.400 ;
        RECT 325.200 576.600 330.900 577.500 ;
        RECT 325.200 575.700 327.000 576.600 ;
        RECT 323.100 568.950 325.200 571.050 ;
        RECT 316.950 565.950 321.000 566.550 ;
        RECT 323.100 561.600 324.300 568.950 ;
        RECT 326.100 564.300 327.000 575.700 ;
        RECT 328.500 568.950 330.600 571.050 ;
        RECT 328.800 567.150 330.600 568.950 ;
        RECT 336.000 568.050 337.500 581.400 ;
        RECT 335.100 565.950 337.500 568.050 ;
        RECT 325.200 563.400 327.000 564.300 ;
        RECT 325.200 562.500 330.900 563.400 ;
        RECT 263.100 549.000 264.900 555.000 ;
        RECT 266.100 549.600 267.900 555.600 ;
        RECT 269.100 549.000 270.900 555.600 ;
        RECT 284.100 549.000 285.900 555.600 ;
        RECT 287.100 549.600 288.900 555.600 ;
        RECT 290.100 549.000 291.900 555.600 ;
        RECT 305.100 549.000 306.900 555.600 ;
        RECT 308.100 549.600 309.900 555.600 ;
        RECT 323.100 549.600 324.900 561.600 ;
        RECT 326.100 549.000 327.900 559.800 ;
        RECT 329.700 555.600 330.900 562.500 ;
        RECT 336.000 555.600 337.500 565.950 ;
        RECT 339.300 578.400 341.100 584.400 ;
        RECT 344.700 578.400 346.500 585.000 ;
        RECT 349.800 579.600 351.600 584.400 ;
        RECT 354.000 581.400 355.800 584.400 ;
        RECT 357.000 581.400 358.800 584.400 ;
        RECT 360.000 581.400 361.800 584.400 ;
        RECT 363.000 581.400 364.800 584.400 ;
        RECT 366.000 581.400 367.800 585.000 ;
        RECT 347.400 578.400 351.600 579.600 ;
        RECT 353.700 579.300 355.800 581.400 ;
        RECT 356.700 579.300 358.800 581.400 ;
        RECT 359.700 579.300 361.800 581.400 ;
        RECT 362.700 579.300 364.800 581.400 ;
        RECT 369.000 580.500 370.800 584.400 ;
        RECT 373.500 581.400 375.300 585.000 ;
        RECT 376.500 581.400 378.300 584.400 ;
        RECT 379.500 581.400 381.300 584.400 ;
        RECT 382.500 581.400 384.300 584.400 ;
        RECT 368.100 578.400 370.800 580.500 ;
        RECT 372.600 579.600 374.400 580.500 ;
        RECT 372.600 578.400 375.300 579.600 ;
        RECT 376.200 579.300 378.300 581.400 ;
        RECT 379.200 579.300 381.300 581.400 ;
        RECT 382.200 579.300 384.300 581.400 ;
        RECT 386.700 578.400 388.500 584.400 ;
        RECT 392.100 578.400 393.900 585.000 ;
        RECT 397.500 578.400 399.300 584.400 ;
        RECT 413.100 578.400 414.900 584.400 ;
        RECT 339.300 561.600 340.200 578.400 ;
        RECT 347.400 575.100 348.900 578.400 ;
        RECT 353.100 576.600 359.700 578.400 ;
        RECT 374.400 577.800 375.300 578.400 ;
        RECT 377.400 577.800 379.200 578.400 ;
        RECT 374.400 576.600 381.600 577.800 ;
        RECT 341.100 573.300 348.900 575.100 ;
        RECT 365.100 574.500 366.900 576.300 ;
        RECT 364.800 573.900 366.900 574.500 ;
        RECT 349.800 572.400 366.900 573.900 ;
        RECT 371.100 573.900 373.200 574.050 ;
        RECT 374.400 573.900 376.200 574.800 ;
        RECT 371.100 573.000 376.200 573.900 ;
        RECT 380.700 573.600 381.600 576.600 ;
        RECT 386.700 577.500 388.200 578.400 ;
        RECT 386.700 576.300 395.100 577.500 ;
        RECT 393.300 575.700 395.100 576.300 ;
        RECT 382.500 574.800 384.600 575.700 ;
        RECT 398.100 574.800 399.300 578.400 ;
        RECT 413.700 576.300 414.900 578.400 ;
        RECT 416.100 579.300 417.900 584.400 ;
        RECT 419.100 580.200 420.900 585.000 ;
        RECT 422.100 579.300 423.900 584.400 ;
        RECT 416.100 577.950 423.900 579.300 ;
        RECT 434.100 579.300 435.900 584.400 ;
        RECT 437.100 580.200 438.900 585.000 ;
        RECT 440.100 579.300 441.900 584.400 ;
        RECT 434.100 577.950 441.900 579.300 ;
        RECT 443.100 578.400 444.900 584.400 ;
        RECT 458.100 578.400 459.900 584.400 ;
        RECT 461.100 578.400 462.900 585.000 ;
        RECT 464.100 581.400 465.900 584.400 ;
        RECT 443.100 576.300 444.300 578.400 ;
        RECT 413.700 575.400 417.300 576.300 ;
        RECT 382.500 573.600 399.300 574.800 ;
        RECT 344.700 570.900 351.300 572.400 ;
        RECT 371.100 571.950 373.200 573.000 ;
        RECT 379.800 571.800 381.600 573.600 ;
        RECT 344.700 568.050 346.200 570.900 ;
        RECT 352.500 569.700 396.900 570.900 ;
        RECT 352.500 568.200 353.400 569.700 ;
        RECT 344.100 565.950 346.200 568.050 ;
        RECT 348.300 566.400 353.400 568.200 ;
        RECT 356.100 567.900 369.600 568.800 ;
        RECT 376.800 567.900 378.600 568.500 ;
        RECT 395.100 568.050 396.900 569.700 ;
        RECT 356.100 566.700 357.000 567.900 ;
        RECT 356.100 564.900 357.900 566.700 ;
        RECT 362.100 565.200 366.000 567.000 ;
        RECT 367.500 566.700 378.600 567.900 ;
        RECT 389.100 567.750 391.200 568.050 ;
        RECT 367.500 565.800 369.600 566.700 ;
        RECT 387.300 565.950 391.200 567.750 ;
        RECT 395.100 565.950 397.200 568.050 ;
        RECT 387.300 565.200 389.100 565.950 ;
        RECT 362.100 564.900 364.200 565.200 ;
        RECT 375.600 564.300 389.100 565.200 ;
        RECT 341.100 563.700 342.900 564.300 ;
        RECT 375.600 563.700 376.800 564.300 ;
        RECT 341.100 562.500 376.800 563.700 ;
        RECT 379.500 562.500 381.600 562.800 ;
        RECT 339.300 560.700 355.800 561.600 ;
        RECT 339.300 557.400 340.200 560.700 ;
        RECT 344.100 558.600 349.800 559.800 ;
        RECT 353.700 559.500 355.800 560.700 ;
        RECT 359.100 560.400 376.800 561.600 ;
        RECT 379.500 561.300 391.500 562.500 ;
        RECT 379.500 560.700 381.600 561.300 ;
        RECT 389.700 560.700 391.500 561.300 ;
        RECT 359.100 559.500 361.200 560.400 ;
        RECT 375.600 559.800 376.800 560.400 ;
        RECT 393.000 559.800 394.800 560.100 ;
        RECT 344.100 558.000 345.900 558.600 ;
        RECT 339.300 556.500 343.200 557.400 ;
        RECT 342.000 555.600 343.200 556.500 ;
        RECT 348.600 555.600 349.800 558.600 ;
        RECT 350.700 557.700 352.500 558.300 ;
        RECT 350.700 556.500 358.800 557.700 ;
        RECT 356.700 555.600 358.800 556.500 ;
        RECT 362.100 555.600 364.800 559.500 ;
        RECT 367.500 557.100 370.800 559.200 ;
        RECT 375.600 558.600 394.800 559.800 ;
        RECT 329.100 549.600 330.900 555.600 ;
        RECT 332.700 549.000 334.500 555.600 ;
        RECT 335.700 549.600 337.500 555.600 ;
        RECT 339.000 549.000 340.800 555.600 ;
        RECT 342.000 549.600 343.800 555.600 ;
        RECT 345.000 549.000 346.800 555.600 ;
        RECT 348.000 549.600 349.800 555.600 ;
        RECT 351.000 549.000 352.800 555.600 ;
        RECT 353.700 552.600 355.800 554.700 ;
        RECT 356.700 552.600 358.800 554.700 ;
        RECT 359.700 552.600 361.800 554.700 ;
        RECT 354.000 549.600 355.800 552.600 ;
        RECT 357.000 549.600 358.800 552.600 ;
        RECT 360.000 549.600 361.800 552.600 ;
        RECT 363.000 549.600 364.800 555.600 ;
        RECT 366.000 549.000 367.800 555.600 ;
        RECT 369.000 549.600 370.800 557.100 ;
        RECT 376.200 555.600 378.300 557.700 ;
        RECT 372.900 549.000 374.700 555.600 ;
        RECT 375.900 549.600 377.700 555.600 ;
        RECT 378.600 552.600 380.700 554.700 ;
        RECT 381.600 552.600 383.700 554.700 ;
        RECT 378.900 549.600 380.700 552.600 ;
        RECT 381.900 549.600 383.700 552.600 ;
        RECT 385.500 549.000 387.300 555.600 ;
        RECT 388.500 549.600 390.300 558.600 ;
        RECT 393.000 558.300 394.800 558.600 ;
        RECT 398.100 557.400 399.300 573.600 ;
        RECT 413.100 571.050 414.900 572.850 ;
        RECT 416.100 571.050 417.300 575.400 ;
        RECT 440.700 575.400 444.300 576.300 ;
        RECT 419.100 571.050 420.900 572.850 ;
        RECT 437.100 571.050 438.900 572.850 ;
        RECT 440.700 571.050 441.900 575.400 ;
        RECT 445.950 573.450 448.050 574.050 ;
        RECT 445.950 573.000 453.450 573.450 ;
        RECT 443.100 571.050 444.900 572.850 ;
        RECT 445.950 572.550 454.050 573.000 ;
        RECT 445.950 571.950 448.050 572.550 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 418.950 568.950 421.050 571.050 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 451.950 568.950 454.050 572.550 ;
        RECT 458.100 571.050 459.300 578.400 ;
        RECT 464.700 577.500 465.900 581.400 ;
        RECT 460.200 576.600 465.900 577.500 ;
        RECT 467.700 578.400 469.500 584.400 ;
        RECT 473.100 578.400 474.900 585.000 ;
        RECT 478.500 578.400 480.300 584.400 ;
        RECT 482.700 581.400 484.500 584.400 ;
        RECT 485.700 581.400 487.500 584.400 ;
        RECT 488.700 581.400 490.500 584.400 ;
        RECT 491.700 581.400 493.500 585.000 ;
        RECT 482.700 579.300 484.800 581.400 ;
        RECT 485.700 579.300 487.800 581.400 ;
        RECT 488.700 579.300 490.800 581.400 ;
        RECT 496.200 580.500 498.000 584.400 ;
        RECT 499.200 581.400 501.000 585.000 ;
        RECT 502.200 581.400 504.000 584.400 ;
        RECT 505.200 581.400 507.000 584.400 ;
        RECT 508.200 581.400 510.000 584.400 ;
        RECT 511.200 581.400 513.000 584.400 ;
        RECT 492.600 579.600 494.400 580.500 ;
        RECT 491.700 578.400 494.400 579.600 ;
        RECT 496.200 578.400 498.900 580.500 ;
        RECT 502.200 579.300 504.300 581.400 ;
        RECT 505.200 579.300 507.300 581.400 ;
        RECT 508.200 579.300 510.300 581.400 ;
        RECT 511.200 579.300 513.300 581.400 ;
        RECT 515.400 579.600 517.200 584.400 ;
        RECT 515.400 578.400 519.600 579.600 ;
        RECT 520.500 578.400 522.300 585.000 ;
        RECT 525.900 578.400 527.700 584.400 ;
        RECT 460.200 575.700 462.000 576.600 ;
        RECT 458.100 568.950 460.200 571.050 ;
        RECT 406.950 567.450 409.050 568.050 ;
        RECT 401.550 567.000 409.050 567.450 ;
        RECT 400.950 566.550 409.050 567.000 ;
        RECT 400.950 562.800 403.050 566.550 ;
        RECT 406.950 565.950 409.050 566.550 ;
        RECT 416.100 561.600 417.300 568.950 ;
        RECT 422.100 567.150 423.900 568.950 ;
        RECT 434.100 567.150 435.900 568.950 ;
        RECT 440.700 561.600 441.900 568.950 ;
        RECT 416.100 560.100 418.500 561.600 ;
        RECT 395.700 556.500 399.300 557.400 ;
        RECT 414.000 557.100 415.800 558.900 ;
        RECT 395.700 555.600 396.600 556.500 ;
        RECT 391.500 549.000 393.300 555.600 ;
        RECT 394.500 554.700 396.600 555.600 ;
        RECT 394.500 549.600 396.300 554.700 ;
        RECT 397.500 549.000 399.300 555.600 ;
        RECT 413.700 549.000 415.500 555.600 ;
        RECT 416.700 549.600 418.500 560.100 ;
        RECT 421.800 549.000 423.600 561.600 ;
        RECT 434.400 549.000 436.200 561.600 ;
        RECT 439.500 560.100 441.900 561.600 ;
        RECT 458.100 561.600 459.300 568.950 ;
        RECT 461.100 564.300 462.000 575.700 ;
        RECT 467.700 574.800 468.900 578.400 ;
        RECT 478.800 577.500 480.300 578.400 ;
        RECT 487.800 577.800 489.600 578.400 ;
        RECT 491.700 577.800 492.600 578.400 ;
        RECT 471.900 576.300 480.300 577.500 ;
        RECT 485.400 576.600 492.600 577.800 ;
        RECT 507.300 576.600 513.900 578.400 ;
        RECT 471.900 575.700 473.700 576.300 ;
        RECT 482.400 574.800 484.500 575.700 ;
        RECT 467.700 573.600 484.500 574.800 ;
        RECT 485.400 573.600 486.300 576.600 ;
        RECT 490.800 573.900 492.600 574.800 ;
        RECT 500.100 574.500 501.900 576.300 ;
        RECT 518.100 575.100 519.600 578.400 ;
        RECT 493.800 573.900 495.900 574.050 ;
        RECT 463.500 568.950 465.600 571.050 ;
        RECT 463.800 567.150 465.600 568.950 ;
        RECT 460.200 563.400 462.000 564.300 ;
        RECT 460.200 562.500 465.900 563.400 ;
        RECT 439.500 549.600 441.300 560.100 ;
        RECT 442.200 557.100 444.000 558.900 ;
        RECT 442.500 549.000 444.300 555.600 ;
        RECT 458.100 549.600 459.900 561.600 ;
        RECT 461.100 549.000 462.900 559.800 ;
        RECT 464.700 555.600 465.900 562.500 ;
        RECT 467.700 557.400 468.900 573.600 ;
        RECT 485.400 571.800 487.200 573.600 ;
        RECT 490.800 573.000 495.900 573.900 ;
        RECT 493.800 571.950 495.900 573.000 ;
        RECT 500.100 573.900 502.200 574.500 ;
        RECT 500.100 572.400 517.200 573.900 ;
        RECT 518.100 573.300 525.900 575.100 ;
        RECT 515.700 570.900 522.300 572.400 ;
        RECT 470.100 569.700 514.500 570.900 ;
        RECT 470.100 568.050 471.900 569.700 ;
        RECT 469.800 565.950 471.900 568.050 ;
        RECT 475.800 567.750 477.900 568.050 ;
        RECT 488.400 567.900 490.200 568.500 ;
        RECT 497.400 567.900 510.900 568.800 ;
        RECT 475.800 565.950 479.700 567.750 ;
        RECT 488.400 566.700 499.500 567.900 ;
        RECT 477.900 565.200 479.700 565.950 ;
        RECT 497.400 565.800 499.500 566.700 ;
        RECT 501.000 565.200 504.900 567.000 ;
        RECT 510.000 566.700 510.900 567.900 ;
        RECT 477.900 564.300 491.400 565.200 ;
        RECT 502.800 564.900 504.900 565.200 ;
        RECT 509.100 564.900 510.900 566.700 ;
        RECT 513.600 568.200 514.500 569.700 ;
        RECT 513.600 566.400 518.700 568.200 ;
        RECT 520.800 568.050 522.300 570.900 ;
        RECT 520.800 565.950 522.900 568.050 ;
        RECT 490.200 563.700 491.400 564.300 ;
        RECT 524.100 563.700 525.900 564.300 ;
        RECT 485.400 562.500 487.500 562.800 ;
        RECT 490.200 562.500 525.900 563.700 ;
        RECT 475.500 561.300 487.500 562.500 ;
        RECT 526.800 561.600 527.700 578.400 ;
        RECT 475.500 560.700 477.300 561.300 ;
        RECT 485.400 560.700 487.500 561.300 ;
        RECT 490.200 560.400 507.900 561.600 ;
        RECT 472.200 559.800 474.000 560.100 ;
        RECT 490.200 559.800 491.400 560.400 ;
        RECT 472.200 558.600 491.400 559.800 ;
        RECT 505.800 559.500 507.900 560.400 ;
        RECT 511.200 560.700 527.700 561.600 ;
        RECT 511.200 559.500 513.300 560.700 ;
        RECT 472.200 558.300 474.000 558.600 ;
        RECT 467.700 556.500 471.300 557.400 ;
        RECT 470.400 555.600 471.300 556.500 ;
        RECT 464.100 549.600 465.900 555.600 ;
        RECT 467.700 549.000 469.500 555.600 ;
        RECT 470.400 554.700 472.500 555.600 ;
        RECT 470.700 549.600 472.500 554.700 ;
        RECT 473.700 549.000 475.500 555.600 ;
        RECT 476.700 549.600 478.500 558.600 ;
        RECT 488.700 555.600 490.800 557.700 ;
        RECT 496.200 557.100 499.500 559.200 ;
        RECT 479.700 549.000 481.500 555.600 ;
        RECT 483.300 552.600 485.400 554.700 ;
        RECT 486.300 552.600 488.400 554.700 ;
        RECT 483.300 549.600 485.100 552.600 ;
        RECT 486.300 549.600 488.100 552.600 ;
        RECT 489.300 549.600 491.100 555.600 ;
        RECT 492.300 549.000 494.100 555.600 ;
        RECT 496.200 549.600 498.000 557.100 ;
        RECT 502.200 555.600 504.900 559.500 ;
        RECT 517.200 558.600 522.900 559.800 ;
        RECT 514.500 557.700 516.300 558.300 ;
        RECT 508.200 556.500 516.300 557.700 ;
        RECT 508.200 555.600 510.300 556.500 ;
        RECT 517.200 555.600 518.400 558.600 ;
        RECT 521.100 558.000 522.900 558.600 ;
        RECT 526.800 557.400 527.700 560.700 ;
        RECT 523.800 556.500 527.700 557.400 ;
        RECT 529.500 581.400 531.300 584.400 ;
        RECT 532.500 581.400 534.300 585.000 ;
        RECT 529.500 568.050 531.000 581.400 ;
        RECT 545.100 579.300 546.900 584.400 ;
        RECT 548.100 580.200 549.900 585.000 ;
        RECT 551.100 579.300 552.900 584.400 ;
        RECT 545.100 577.950 552.900 579.300 ;
        RECT 554.100 578.400 555.900 584.400 ;
        RECT 569.400 578.400 571.200 585.000 ;
        RECT 554.100 576.300 555.300 578.400 ;
        RECT 574.500 577.200 576.300 584.400 ;
        RECT 590.100 581.400 591.900 585.000 ;
        RECT 593.100 581.400 594.900 584.400 ;
        RECT 608.100 581.400 609.900 584.400 ;
        RECT 577.950 579.450 580.050 580.050 ;
        RECT 589.950 579.450 592.050 580.050 ;
        RECT 577.950 578.550 592.050 579.450 ;
        RECT 577.950 577.950 580.050 578.550 ;
        RECT 589.950 577.950 592.050 578.550 ;
        RECT 551.700 575.400 555.300 576.300 ;
        RECT 559.950 576.450 562.050 576.900 ;
        RECT 568.950 576.450 571.050 577.050 ;
        RECT 559.950 575.550 571.050 576.450 ;
        RECT 548.100 571.050 549.900 572.850 ;
        RECT 551.700 571.050 552.900 575.400 ;
        RECT 559.950 574.800 562.050 575.550 ;
        RECT 568.950 574.950 571.050 575.550 ;
        RECT 572.100 576.300 576.300 577.200 ;
        RECT 554.100 571.050 555.900 572.850 ;
        RECT 569.250 571.050 571.050 572.850 ;
        RECT 572.100 571.050 573.300 576.300 ;
        RECT 575.100 571.050 576.900 572.850 ;
        RECT 593.100 571.050 594.300 581.400 ;
        RECT 608.100 577.500 609.300 581.400 ;
        RECT 611.100 578.400 612.900 585.000 ;
        RECT 614.100 578.400 615.900 584.400 ;
        RECT 629.100 581.400 630.900 584.400 ;
        RECT 632.100 581.400 633.900 585.000 ;
        RECT 644.100 581.400 645.900 585.000 ;
        RECT 647.100 581.400 648.900 584.400 ;
        RECT 608.100 576.600 613.800 577.500 ;
        RECT 612.000 575.700 613.800 576.600 ;
        RECT 544.950 568.950 547.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 608.400 568.950 610.500 571.050 ;
        RECT 529.500 565.950 531.900 568.050 ;
        RECT 545.100 567.150 546.900 568.950 ;
        RECT 523.800 555.600 525.000 556.500 ;
        RECT 529.500 555.600 531.000 565.950 ;
        RECT 551.700 561.600 552.900 568.950 ;
        RECT 499.200 549.000 501.000 555.600 ;
        RECT 502.200 549.600 504.000 555.600 ;
        RECT 505.200 552.600 507.300 554.700 ;
        RECT 508.200 552.600 510.300 554.700 ;
        RECT 511.200 552.600 513.300 554.700 ;
        RECT 505.200 549.600 507.000 552.600 ;
        RECT 508.200 549.600 510.000 552.600 ;
        RECT 511.200 549.600 513.000 552.600 ;
        RECT 514.200 549.000 516.000 555.600 ;
        RECT 517.200 549.600 519.000 555.600 ;
        RECT 520.200 549.000 522.000 555.600 ;
        RECT 523.200 549.600 525.000 555.600 ;
        RECT 526.200 549.000 528.000 555.600 ;
        RECT 529.500 549.600 531.300 555.600 ;
        RECT 532.500 549.000 534.300 555.600 ;
        RECT 545.400 549.000 547.200 561.600 ;
        RECT 550.500 560.100 552.900 561.600 ;
        RECT 550.500 549.600 552.300 560.100 ;
        RECT 553.200 557.100 555.000 558.900 ;
        RECT 572.100 555.600 573.300 568.950 ;
        RECT 590.100 567.150 591.900 568.950 ;
        RECT 580.950 564.450 583.050 565.050 ;
        RECT 589.950 564.450 592.050 565.050 ;
        RECT 580.950 563.550 592.050 564.450 ;
        RECT 580.950 562.950 583.050 563.550 ;
        RECT 589.950 562.950 592.050 563.550 ;
        RECT 593.100 555.600 594.300 568.950 ;
        RECT 608.400 567.150 610.200 568.950 ;
        RECT 612.000 564.300 612.900 575.700 ;
        RECT 614.700 571.050 615.900 578.400 ;
        RECT 629.700 571.050 630.900 581.400 ;
        RECT 647.100 571.050 648.300 581.400 ;
        RECT 662.100 579.300 663.900 584.400 ;
        RECT 665.100 580.200 666.900 585.000 ;
        RECT 668.100 579.300 669.900 584.400 ;
        RECT 662.100 577.950 669.900 579.300 ;
        RECT 671.100 578.400 672.900 584.400 ;
        RECT 683.400 578.400 685.200 585.000 ;
        RECT 671.100 576.300 672.300 578.400 ;
        RECT 688.500 577.200 690.300 584.400 ;
        RECT 701.100 578.400 702.900 584.400 ;
        RECT 704.400 579.300 706.200 585.000 ;
        RECT 708.900 579.000 710.700 584.400 ;
        RECT 713.100 579.300 714.900 585.000 ;
        RECT 701.100 577.500 705.600 578.400 ;
        RECT 668.700 575.400 672.300 576.300 ;
        RECT 686.100 576.300 690.300 577.200 ;
        RECT 665.100 571.050 666.900 572.850 ;
        RECT 668.700 571.050 669.900 575.400 ;
        RECT 671.100 571.050 672.900 572.850 ;
        RECT 683.250 571.050 685.050 572.850 ;
        RECT 686.100 571.050 687.300 576.300 ;
        RECT 703.500 575.100 705.600 577.500 ;
        RECT 708.900 576.900 709.800 579.000 ;
        RECT 716.100 578.400 717.900 584.400 ;
        RECT 731.400 578.400 733.200 585.000 ;
        RECT 716.400 577.500 717.900 578.400 ;
        RECT 706.800 574.800 709.800 576.900 ;
        RECT 713.400 576.000 717.900 577.500 ;
        RECT 736.500 577.200 738.300 584.400 ;
        RECT 734.100 576.300 738.300 577.200 ;
        RECT 752.700 577.200 754.500 584.400 ;
        RECT 757.800 578.400 759.600 585.000 ;
        RECT 770.100 581.400 771.900 585.000 ;
        RECT 773.100 581.400 774.900 584.400 ;
        RECT 776.100 581.400 777.900 585.000 ;
        RECT 791.100 584.400 792.300 585.000 ;
        RECT 791.100 581.400 792.900 584.400 ;
        RECT 794.100 581.400 795.900 584.400 ;
        RECT 752.700 576.300 756.900 577.200 ;
        RECT 689.100 571.050 690.900 572.850 ;
        RECT 613.800 568.950 615.900 571.050 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 661.950 568.950 664.050 571.050 ;
        RECT 664.950 568.950 667.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 685.950 568.950 688.050 571.050 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 701.100 568.950 703.200 571.050 ;
        RECT 705.900 570.900 708.000 573.000 ;
        RECT 706.200 569.100 708.000 570.900 ;
        RECT 612.000 563.400 613.800 564.300 ;
        RECT 608.100 562.500 613.800 563.400 ;
        RECT 608.100 555.600 609.300 562.500 ;
        RECT 614.700 561.600 615.900 568.950 ;
        RECT 553.500 549.000 555.300 555.600 ;
        RECT 569.100 549.000 570.900 555.600 ;
        RECT 572.100 549.600 573.900 555.600 ;
        RECT 575.100 549.000 576.900 555.600 ;
        RECT 590.100 549.000 591.900 555.600 ;
        RECT 593.100 549.600 594.900 555.600 ;
        RECT 608.100 549.600 609.900 555.600 ;
        RECT 611.100 549.000 612.900 559.800 ;
        RECT 614.100 549.600 615.900 561.600 ;
        RECT 629.700 555.600 630.900 568.950 ;
        RECT 632.100 567.150 633.900 568.950 ;
        RECT 644.100 567.150 645.900 568.950 ;
        RECT 647.100 555.600 648.300 568.950 ;
        RECT 662.100 567.150 663.900 568.950 ;
        RECT 652.950 564.450 655.050 565.050 ;
        RECT 661.950 564.450 664.050 565.050 ;
        RECT 652.950 563.550 664.050 564.450 ;
        RECT 652.950 562.950 655.050 563.550 ;
        RECT 661.950 562.950 664.050 563.550 ;
        RECT 668.700 561.600 669.900 568.950 ;
        RECT 629.100 549.600 630.900 555.600 ;
        RECT 632.100 549.000 633.900 555.600 ;
        RECT 644.100 549.000 645.900 555.600 ;
        RECT 647.100 549.600 648.900 555.600 ;
        RECT 662.400 549.000 664.200 561.600 ;
        RECT 667.500 560.100 669.900 561.600 ;
        RECT 667.500 549.600 669.300 560.100 ;
        RECT 670.200 557.100 672.000 558.900 ;
        RECT 686.100 555.600 687.300 568.950 ;
        RECT 701.400 567.150 703.200 568.950 ;
        RECT 708.900 568.050 709.800 574.800 ;
        RECT 710.700 573.900 712.500 575.700 ;
        RECT 713.400 575.400 715.500 576.000 ;
        RECT 711.000 573.000 713.100 573.900 ;
        RECT 711.000 571.800 717.600 573.000 ;
        RECT 715.800 571.200 717.600 571.800 ;
        RECT 711.000 568.800 713.100 570.900 ;
        RECT 715.800 568.950 717.900 571.200 ;
        RECT 731.250 571.050 733.050 572.850 ;
        RECT 734.100 571.050 735.300 576.300 ;
        RECT 737.100 571.050 738.900 572.850 ;
        RECT 752.100 571.050 753.900 572.850 ;
        RECT 755.700 571.050 756.900 576.300 ;
        RECT 760.950 576.450 763.050 577.050 ;
        RECT 769.950 576.450 772.050 577.050 ;
        RECT 760.950 575.550 772.050 576.450 ;
        RECT 760.950 574.950 763.050 575.550 ;
        RECT 769.950 574.950 772.050 575.550 ;
        RECT 757.950 571.050 759.750 572.850 ;
        RECT 773.700 571.050 774.600 581.400 ;
        RECT 794.400 577.200 795.300 581.400 ;
        RECT 797.100 579.000 798.900 585.000 ;
        RECT 800.100 578.400 801.900 584.400 ;
        RECT 794.400 576.300 799.800 577.200 ;
        RECT 797.700 575.400 799.800 576.300 ;
        RECT 791.400 571.050 793.200 572.850 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 733.950 568.950 736.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 791.100 568.950 793.200 571.050 ;
        RECT 794.400 568.950 796.500 571.050 ;
        RECT 706.800 566.700 709.800 568.050 ;
        RECT 711.300 567.000 713.100 568.800 ;
        RECT 706.800 565.950 708.900 566.700 ;
        RECT 704.100 561.600 706.200 562.500 ;
        RECT 701.100 560.400 706.200 561.600 ;
        RECT 707.100 561.600 708.300 565.950 ;
        RECT 709.800 563.700 711.600 565.500 ;
        RECT 709.800 562.800 715.200 563.700 ;
        RECT 713.100 561.900 715.200 562.800 ;
        RECT 707.100 560.700 710.400 561.600 ;
        RECT 713.100 560.700 717.900 561.900 ;
        RECT 670.500 549.000 672.300 555.600 ;
        RECT 683.100 549.000 684.900 555.600 ;
        RECT 686.100 549.600 687.900 555.600 ;
        RECT 689.100 549.000 690.900 555.600 ;
        RECT 701.100 549.600 702.900 560.400 ;
        RECT 704.100 549.000 706.200 559.500 ;
        RECT 708.600 549.600 710.400 560.700 ;
        RECT 713.100 549.000 714.900 559.500 ;
        RECT 716.100 549.600 717.900 560.700 ;
        RECT 734.100 555.600 735.300 568.950 ;
        RECT 755.700 555.600 756.900 568.950 ;
        RECT 770.100 567.150 771.900 568.950 ;
        RECT 773.700 561.600 774.600 568.950 ;
        RECT 775.950 567.150 777.750 568.950 ;
        RECT 795.000 567.150 796.800 568.950 ;
        RECT 797.700 564.900 798.600 575.400 ;
        RECT 801.000 571.050 801.900 578.400 ;
        RECT 812.100 575.400 813.900 585.000 ;
        RECT 818.700 576.000 820.500 584.400 ;
        RECT 833.700 577.200 835.500 584.400 ;
        RECT 838.800 578.400 840.600 585.000 ;
        RECT 833.700 576.300 837.900 577.200 ;
        RECT 818.700 574.800 822.000 576.000 ;
        RECT 812.100 571.050 813.900 572.850 ;
        RECT 818.100 571.050 819.900 572.850 ;
        RECT 821.100 571.050 822.000 574.800 ;
        RECT 828.000 573.450 832.050 574.050 ;
        RECT 827.550 571.950 832.050 573.450 ;
        RECT 799.800 568.950 801.900 571.050 ;
        RECT 811.950 568.950 814.050 571.050 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 797.100 564.300 798.900 564.900 ;
        RECT 791.100 563.100 798.900 564.300 ;
        RECT 791.100 561.600 792.300 563.100 ;
        RECT 799.800 561.600 801.000 568.950 ;
        RECT 815.100 567.150 816.900 568.950 ;
        RECT 802.950 564.450 805.050 565.050 ;
        RECT 817.950 564.450 820.050 565.050 ;
        RECT 802.950 563.550 820.050 564.450 ;
        RECT 802.950 562.950 805.050 563.550 ;
        RECT 817.950 562.950 820.050 563.550 ;
        RECT 771.000 560.400 774.600 561.600 ;
        RECT 731.100 549.000 732.900 555.600 ;
        RECT 734.100 549.600 735.900 555.600 ;
        RECT 737.100 549.000 738.900 555.600 ;
        RECT 752.100 549.000 753.900 555.600 ;
        RECT 755.100 549.600 756.900 555.600 ;
        RECT 758.100 549.000 759.900 555.600 ;
        RECT 771.000 549.600 772.800 560.400 ;
        RECT 776.100 549.000 777.900 561.600 ;
        RECT 791.100 549.600 792.900 561.600 ;
        RECT 795.600 549.000 797.400 561.600 ;
        RECT 798.600 560.100 801.000 561.600 ;
        RECT 798.600 549.600 800.400 560.100 ;
        RECT 821.100 556.800 822.000 568.950 ;
        RECT 827.550 564.450 828.450 571.950 ;
        RECT 833.100 571.050 834.900 572.850 ;
        RECT 836.700 571.050 837.900 576.300 ;
        RECT 854.100 575.400 855.900 585.000 ;
        RECT 860.700 576.000 862.500 584.400 ;
        RECT 875.100 578.400 876.900 584.400 ;
        RECT 875.700 576.300 876.900 578.400 ;
        RECT 878.100 579.300 879.900 584.400 ;
        RECT 881.100 580.200 882.900 585.000 ;
        RECT 884.100 579.300 885.900 584.400 ;
        RECT 899.100 581.400 900.900 585.000 ;
        RECT 902.100 581.400 903.900 584.400 ;
        RECT 905.100 581.400 906.900 585.000 ;
        RECT 917.700 581.400 919.500 585.000 ;
        RECT 878.100 577.950 885.900 579.300 ;
        RECT 860.700 574.800 864.000 576.000 ;
        RECT 875.700 575.400 879.300 576.300 ;
        RECT 838.950 571.050 840.750 572.850 ;
        RECT 854.100 571.050 855.900 572.850 ;
        RECT 860.100 571.050 861.900 572.850 ;
        RECT 863.100 571.050 864.000 574.800 ;
        RECT 875.100 571.050 876.900 572.850 ;
        RECT 878.100 571.050 879.300 575.400 ;
        RECT 881.100 571.050 882.900 572.850 ;
        RECT 902.700 571.050 903.600 581.400 ;
        RECT 920.700 579.600 922.500 584.400 ;
        RECT 917.400 578.400 922.500 579.600 ;
        RECT 925.200 578.400 927.000 585.000 ;
        RECT 941.100 581.400 942.900 584.400 ;
        RECT 944.100 581.400 945.900 585.000 ;
        RECT 917.400 571.050 918.300 578.400 ;
        RECT 919.950 571.050 921.750 572.850 ;
        RECT 926.100 571.050 927.900 572.850 ;
        RECT 941.700 571.050 942.900 581.400 ;
        RECT 832.950 568.950 835.050 571.050 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 874.950 568.950 877.050 571.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 898.950 568.950 901.050 571.050 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 916.950 568.950 919.050 571.050 ;
        RECT 919.950 568.950 922.050 571.050 ;
        RECT 922.950 568.950 925.050 571.050 ;
        RECT 925.950 568.950 928.050 571.050 ;
        RECT 940.950 568.950 943.050 571.050 ;
        RECT 943.950 568.950 946.050 571.050 ;
        RECT 832.950 564.450 835.050 565.050 ;
        RECT 827.550 563.550 835.050 564.450 ;
        RECT 832.950 562.950 835.050 563.550 ;
        RECT 815.400 555.900 822.000 556.800 ;
        RECT 815.400 555.600 816.900 555.900 ;
        RECT 812.100 549.000 813.900 555.600 ;
        RECT 815.100 549.600 816.900 555.600 ;
        RECT 821.100 555.600 822.000 555.900 ;
        RECT 836.700 555.600 837.900 568.950 ;
        RECT 857.100 567.150 858.900 568.950 ;
        RECT 844.950 564.450 847.050 565.050 ;
        RECT 859.950 564.450 862.050 565.050 ;
        RECT 844.950 563.550 862.050 564.450 ;
        RECT 844.950 562.950 847.050 563.550 ;
        RECT 859.950 562.950 862.050 563.550 ;
        RECT 863.100 556.800 864.000 568.950 ;
        RECT 878.100 561.600 879.300 568.950 ;
        RECT 884.100 567.150 885.900 568.950 ;
        RECT 899.100 567.150 900.900 568.950 ;
        RECT 902.700 561.600 903.600 568.950 ;
        RECT 904.950 567.150 906.750 568.950 ;
        RECT 917.400 561.600 918.300 568.950 ;
        RECT 922.950 567.150 924.750 568.950 ;
        RECT 878.100 560.100 880.500 561.600 ;
        RECT 876.000 557.100 877.800 558.900 ;
        RECT 857.400 555.900 864.000 556.800 ;
        RECT 857.400 555.600 858.900 555.900 ;
        RECT 818.100 549.000 819.900 555.000 ;
        RECT 821.100 549.600 822.900 555.600 ;
        RECT 833.100 549.000 834.900 555.600 ;
        RECT 836.100 549.600 837.900 555.600 ;
        RECT 839.100 549.000 840.900 555.600 ;
        RECT 854.100 549.000 855.900 555.600 ;
        RECT 857.100 549.600 858.900 555.600 ;
        RECT 863.100 555.600 864.000 555.900 ;
        RECT 860.100 549.000 861.900 555.000 ;
        RECT 863.100 549.600 864.900 555.600 ;
        RECT 875.700 549.000 877.500 555.600 ;
        RECT 878.700 549.600 880.500 560.100 ;
        RECT 883.800 549.000 885.600 561.600 ;
        RECT 900.000 560.400 903.600 561.600 ;
        RECT 900.000 549.600 901.800 560.400 ;
        RECT 905.100 549.000 906.900 561.600 ;
        RECT 917.100 549.600 918.900 561.600 ;
        RECT 920.100 560.700 927.900 561.600 ;
        RECT 920.100 549.600 921.900 560.700 ;
        RECT 923.100 549.000 924.900 559.800 ;
        RECT 926.100 549.600 927.900 560.700 ;
        RECT 941.700 555.600 942.900 568.950 ;
        RECT 944.100 567.150 945.900 568.950 ;
        RECT 941.100 549.600 942.900 555.600 ;
        RECT 944.100 549.000 945.900 555.600 ;
        RECT 14.700 539.400 16.500 546.000 ;
        RECT 15.000 536.100 16.800 537.900 ;
        RECT 17.700 534.900 19.500 545.400 ;
        RECT 17.100 533.400 19.500 534.900 ;
        RECT 22.800 533.400 24.600 546.000 ;
        RECT 38.100 539.400 39.900 545.400 ;
        RECT 41.100 539.400 42.900 546.000 ;
        RECT 56.100 539.400 57.900 545.400 ;
        RECT 59.100 539.400 60.900 546.000 ;
        RECT 74.700 539.400 76.500 546.000 ;
        RECT 17.100 526.050 18.300 533.400 ;
        RECT 23.100 526.050 24.900 527.850 ;
        RECT 38.700 526.050 39.900 539.400 ;
        RECT 41.100 526.050 42.900 527.850 ;
        RECT 56.700 526.050 57.900 539.400 ;
        RECT 75.000 536.100 76.800 537.900 ;
        RECT 77.700 534.900 79.500 545.400 ;
        RECT 77.100 533.400 79.500 534.900 ;
        RECT 82.800 533.400 84.600 546.000 ;
        RECT 95.100 534.300 96.900 545.400 ;
        RECT 98.100 535.200 99.900 546.000 ;
        RECT 101.100 534.300 102.900 545.400 ;
        RECT 95.100 533.400 102.900 534.300 ;
        RECT 104.100 533.400 105.900 545.400 ;
        RECT 116.100 539.400 117.900 546.000 ;
        RECT 119.100 539.400 120.900 545.400 ;
        RECT 59.100 526.050 60.900 527.850 ;
        RECT 77.100 526.050 78.300 533.400 ;
        RECT 79.950 531.450 82.050 532.050 ;
        RECT 79.950 530.550 90.450 531.450 ;
        RECT 79.950 529.950 82.050 530.550 ;
        RECT 83.100 526.050 84.900 527.850 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 19.950 523.950 22.050 526.050 ;
        RECT 22.950 523.950 25.050 526.050 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 14.100 522.150 15.900 523.950 ;
        RECT 17.100 519.600 18.300 523.950 ;
        RECT 20.100 522.150 21.900 523.950 ;
        RECT 14.700 518.700 18.300 519.600 ;
        RECT 14.700 516.600 15.900 518.700 ;
        RECT 14.100 510.600 15.900 516.600 ;
        RECT 17.100 515.700 24.900 517.050 ;
        RECT 17.100 510.600 18.900 515.700 ;
        RECT 20.100 510.000 21.900 514.800 ;
        RECT 23.100 510.600 24.900 515.700 ;
        RECT 38.700 513.600 39.900 523.950 ;
        RECT 56.700 513.600 57.900 523.950 ;
        RECT 74.100 522.150 75.900 523.950 ;
        RECT 67.950 519.450 70.050 520.050 ;
        RECT 77.100 519.600 78.300 523.950 ;
        RECT 80.100 522.150 81.900 523.950 ;
        RECT 89.550 522.450 90.450 530.550 ;
        RECT 98.250 526.050 100.050 527.850 ;
        RECT 104.700 526.050 105.600 533.400 ;
        RECT 106.950 528.450 111.000 529.050 ;
        RECT 106.950 526.950 111.450 528.450 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 89.550 521.550 93.450 522.450 ;
        RECT 95.100 522.150 96.900 523.950 ;
        RECT 101.250 522.150 103.050 523.950 ;
        RECT 59.550 519.000 70.050 519.450 ;
        RECT 58.950 518.550 70.050 519.000 ;
        RECT 58.950 514.950 61.050 518.550 ;
        RECT 67.950 517.950 70.050 518.550 ;
        RECT 74.700 518.700 78.300 519.600 ;
        RECT 92.550 519.450 93.450 521.550 ;
        RECT 97.950 519.450 100.050 520.050 ;
        RECT 74.700 516.600 75.900 518.700 ;
        RECT 92.550 518.550 100.050 519.450 ;
        RECT 97.950 517.950 100.050 518.550 ;
        RECT 38.100 510.600 39.900 513.600 ;
        RECT 41.100 510.000 42.900 513.600 ;
        RECT 56.100 510.600 57.900 513.600 ;
        RECT 59.100 510.000 60.900 513.600 ;
        RECT 74.100 510.600 75.900 516.600 ;
        RECT 77.100 515.700 84.900 517.050 ;
        RECT 104.700 516.600 105.600 523.950 ;
        RECT 110.550 523.050 111.450 526.950 ;
        RECT 116.100 526.050 117.900 527.850 ;
        RECT 119.100 526.050 120.300 539.400 ;
        RECT 134.400 533.400 136.200 546.000 ;
        RECT 139.500 534.900 141.300 545.400 ;
        RECT 142.500 539.400 144.300 546.000 ;
        RECT 142.200 536.100 144.000 537.900 ;
        RECT 139.500 533.400 141.900 534.900 ;
        RECT 159.000 534.600 160.800 545.400 ;
        RECT 159.000 533.400 162.600 534.600 ;
        RECT 164.100 533.400 165.900 546.000 ;
        RECT 176.400 533.400 178.200 546.000 ;
        RECT 181.500 534.900 183.300 545.400 ;
        RECT 184.500 539.400 186.300 546.000 ;
        RECT 197.700 539.400 199.500 546.000 ;
        RECT 184.200 536.100 186.000 537.900 ;
        RECT 198.000 536.100 199.800 537.900 ;
        RECT 200.700 534.900 202.500 545.400 ;
        RECT 181.500 533.400 183.900 534.900 ;
        RECT 129.000 528.450 133.050 529.050 ;
        RECT 128.550 526.950 133.050 528.450 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 110.550 521.550 115.050 523.050 ;
        RECT 111.000 520.950 115.050 521.550 ;
        RECT 77.100 510.600 78.900 515.700 ;
        RECT 80.100 510.000 81.900 514.800 ;
        RECT 83.100 510.600 84.900 515.700 ;
        RECT 96.000 510.000 97.800 516.600 ;
        RECT 100.500 515.400 105.600 516.600 ;
        RECT 100.500 510.600 102.300 515.400 ;
        RECT 119.100 513.600 120.300 523.950 ;
        RECT 128.550 523.050 129.450 526.950 ;
        RECT 134.100 526.050 135.900 527.850 ;
        RECT 140.700 526.050 141.900 533.400 ;
        RECT 145.950 528.450 150.000 529.050 ;
        RECT 153.000 528.450 157.050 529.050 ;
        RECT 145.950 526.950 150.450 528.450 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 128.550 521.550 133.050 523.050 ;
        RECT 137.100 522.150 138.900 523.950 ;
        RECT 129.000 520.950 133.050 521.550 ;
        RECT 140.700 519.600 141.900 523.950 ;
        RECT 143.100 522.150 144.900 523.950 ;
        RECT 140.700 518.700 144.300 519.600 ;
        RECT 134.100 515.700 141.900 517.050 ;
        RECT 103.500 510.000 105.300 513.600 ;
        RECT 116.100 510.000 117.900 513.600 ;
        RECT 119.100 510.600 120.900 513.600 ;
        RECT 134.100 510.600 135.900 515.700 ;
        RECT 137.100 510.000 138.900 514.800 ;
        RECT 140.100 510.600 141.900 515.700 ;
        RECT 143.100 516.600 144.300 518.700 ;
        RECT 149.550 519.450 150.450 526.950 ;
        RECT 152.550 526.950 157.050 528.450 ;
        RECT 152.550 523.050 153.450 526.950 ;
        RECT 158.100 526.050 159.900 527.850 ;
        RECT 161.700 526.050 162.600 533.400 ;
        RECT 163.950 526.050 165.750 527.850 ;
        RECT 176.100 526.050 177.900 527.850 ;
        RECT 182.700 526.050 183.900 533.400 ;
        RECT 200.100 533.400 202.500 534.900 ;
        RECT 205.800 533.400 207.600 546.000 ;
        RECT 218.100 539.400 219.900 546.000 ;
        RECT 221.100 539.400 222.900 545.400 ;
        RECT 224.100 539.400 225.900 546.000 ;
        RECT 187.950 528.450 192.000 529.050 ;
        RECT 187.950 526.950 192.450 528.450 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 152.550 521.550 157.050 523.050 ;
        RECT 153.000 520.950 157.050 521.550 ;
        RECT 157.950 519.450 160.050 519.750 ;
        RECT 149.550 518.550 160.050 519.450 ;
        RECT 157.950 517.650 160.050 518.550 ;
        RECT 143.100 510.600 144.900 516.600 ;
        RECT 161.700 513.600 162.600 523.950 ;
        RECT 179.100 522.150 180.900 523.950 ;
        RECT 182.700 519.600 183.900 523.950 ;
        RECT 185.100 522.150 186.900 523.950 ;
        RECT 191.550 523.050 192.450 526.950 ;
        RECT 200.100 526.050 201.300 533.400 ;
        RECT 211.950 531.450 214.050 532.050 ;
        RECT 217.950 531.450 220.050 532.050 ;
        RECT 211.950 530.550 220.050 531.450 ;
        RECT 211.950 529.950 214.050 530.550 ;
        RECT 217.950 529.950 220.050 530.550 ;
        RECT 206.100 526.050 207.900 527.850 ;
        RECT 221.700 526.050 222.900 539.400 ;
        RECT 239.400 533.400 241.200 546.000 ;
        RECT 244.500 534.900 246.300 545.400 ;
        RECT 247.500 539.400 249.300 546.000 ;
        RECT 247.200 536.100 249.000 537.900 ;
        RECT 244.500 533.400 246.900 534.900 ;
        RECT 261.000 534.600 262.800 545.400 ;
        RECT 261.000 533.400 264.600 534.600 ;
        RECT 266.100 533.400 267.900 546.000 ;
        RECT 281.400 533.400 283.200 546.000 ;
        RECT 286.500 534.900 288.300 545.400 ;
        RECT 289.500 539.400 291.300 546.000 ;
        RECT 302.100 539.400 303.900 546.000 ;
        RECT 305.100 539.400 306.900 545.400 ;
        RECT 308.100 539.400 309.900 546.000 ;
        RECT 289.200 536.100 291.000 537.900 ;
        RECT 286.500 533.400 288.900 534.900 ;
        RECT 239.100 526.050 240.900 527.850 ;
        RECT 245.700 526.050 246.900 533.400 ;
        RECT 250.950 528.450 255.000 529.050 ;
        RECT 250.950 526.950 255.450 528.450 ;
        RECT 196.950 523.950 199.050 526.050 ;
        RECT 199.950 523.950 202.050 526.050 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 217.950 523.950 220.050 526.050 ;
        RECT 220.950 523.950 223.050 526.050 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 244.950 523.950 247.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 187.950 521.550 192.450 523.050 ;
        RECT 197.100 522.150 198.900 523.950 ;
        RECT 187.950 520.950 192.000 521.550 ;
        RECT 200.100 519.600 201.300 523.950 ;
        RECT 203.100 522.150 204.900 523.950 ;
        RECT 218.100 522.150 219.900 523.950 ;
        RECT 182.700 518.700 186.300 519.600 ;
        RECT 176.100 515.700 183.900 517.050 ;
        RECT 158.100 510.000 159.900 513.600 ;
        RECT 161.100 510.600 162.900 513.600 ;
        RECT 164.100 510.000 165.900 513.600 ;
        RECT 176.100 510.600 177.900 515.700 ;
        RECT 179.100 510.000 180.900 514.800 ;
        RECT 182.100 510.600 183.900 515.700 ;
        RECT 185.100 516.600 186.300 518.700 ;
        RECT 197.700 518.700 201.300 519.600 ;
        RECT 221.700 518.700 222.900 523.950 ;
        RECT 223.950 522.150 225.750 523.950 ;
        RECT 232.950 522.450 235.050 523.050 ;
        RECT 197.700 516.600 198.900 518.700 ;
        RECT 218.700 517.800 222.900 518.700 ;
        RECT 227.550 521.550 235.050 522.450 ;
        RECT 242.100 522.150 243.900 523.950 ;
        RECT 185.100 510.600 186.900 516.600 ;
        RECT 197.100 510.600 198.900 516.600 ;
        RECT 200.100 515.700 207.900 517.050 ;
        RECT 200.100 510.600 201.900 515.700 ;
        RECT 203.100 510.000 204.900 514.800 ;
        RECT 206.100 510.600 207.900 515.700 ;
        RECT 218.700 510.600 220.500 517.800 ;
        RECT 223.800 510.000 225.600 516.600 ;
        RECT 227.550 516.450 228.450 521.550 ;
        RECT 232.950 520.950 235.050 521.550 ;
        RECT 245.700 519.600 246.900 523.950 ;
        RECT 248.100 522.150 249.900 523.950 ;
        RECT 254.550 523.050 255.450 526.950 ;
        RECT 260.100 526.050 261.900 527.850 ;
        RECT 263.700 526.050 264.600 533.400 ;
        RECT 283.950 531.450 286.050 532.050 ;
        RECT 278.550 530.550 286.050 531.450 ;
        RECT 268.950 528.450 273.000 529.050 ;
        RECT 278.550 528.450 279.450 530.550 ;
        RECT 283.950 529.950 286.050 530.550 ;
        RECT 265.950 526.050 267.750 527.850 ;
        RECT 268.950 526.950 273.450 528.450 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 254.550 521.550 259.050 523.050 ;
        RECT 255.000 520.950 259.050 521.550 ;
        RECT 245.700 518.700 249.300 519.600 ;
        RECT 232.950 516.450 235.050 517.050 ;
        RECT 227.550 515.550 235.050 516.450 ;
        RECT 232.950 514.950 235.050 515.550 ;
        RECT 239.100 515.700 246.900 517.050 ;
        RECT 239.100 510.600 240.900 515.700 ;
        RECT 242.100 510.000 243.900 514.800 ;
        RECT 245.100 510.600 246.900 515.700 ;
        RECT 248.100 516.600 249.300 518.700 ;
        RECT 248.100 510.600 249.900 516.600 ;
        RECT 263.700 513.600 264.600 523.950 ;
        RECT 272.550 523.050 273.450 526.950 ;
        RECT 268.950 521.550 273.450 523.050 ;
        RECT 275.550 527.550 279.450 528.450 ;
        RECT 275.550 523.050 276.450 527.550 ;
        RECT 281.100 526.050 282.900 527.850 ;
        RECT 287.700 526.050 288.900 533.400 ;
        RECT 305.100 526.050 306.300 539.400 ;
        RECT 323.100 533.400 324.900 545.400 ;
        RECT 326.100 535.200 327.900 546.000 ;
        RECT 329.100 539.400 330.900 545.400 ;
        RECT 332.700 539.400 334.500 546.000 ;
        RECT 335.700 539.400 337.500 545.400 ;
        RECT 339.000 539.400 340.800 546.000 ;
        RECT 342.000 539.400 343.800 545.400 ;
        RECT 345.000 539.400 346.800 546.000 ;
        RECT 348.000 539.400 349.800 545.400 ;
        RECT 351.000 539.400 352.800 546.000 ;
        RECT 354.000 542.400 355.800 545.400 ;
        RECT 357.000 542.400 358.800 545.400 ;
        RECT 360.000 542.400 361.800 545.400 ;
        RECT 353.700 540.300 355.800 542.400 ;
        RECT 356.700 540.300 358.800 542.400 ;
        RECT 359.700 540.300 361.800 542.400 ;
        RECT 363.000 539.400 364.800 545.400 ;
        RECT 366.000 539.400 367.800 546.000 ;
        RECT 310.950 528.450 315.000 529.050 ;
        RECT 310.950 526.950 315.450 528.450 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 304.950 523.950 307.050 526.050 ;
        RECT 307.950 523.950 310.050 526.050 ;
        RECT 275.550 521.550 280.050 523.050 ;
        RECT 284.100 522.150 285.900 523.950 ;
        RECT 268.950 520.950 273.000 521.550 ;
        RECT 276.000 520.950 280.050 521.550 ;
        RECT 287.700 519.600 288.900 523.950 ;
        RECT 290.100 522.150 291.900 523.950 ;
        RECT 302.250 522.150 304.050 523.950 ;
        RECT 287.700 518.700 291.300 519.600 ;
        RECT 281.100 515.700 288.900 517.050 ;
        RECT 260.100 510.000 261.900 513.600 ;
        RECT 263.100 510.600 264.900 513.600 ;
        RECT 266.100 510.000 267.900 513.600 ;
        RECT 281.100 510.600 282.900 515.700 ;
        RECT 284.100 510.000 285.900 514.800 ;
        RECT 287.100 510.600 288.900 515.700 ;
        RECT 290.100 516.600 291.300 518.700 ;
        RECT 305.100 518.700 306.300 523.950 ;
        RECT 308.100 522.150 309.900 523.950 ;
        RECT 314.550 523.050 315.450 526.950 ;
        RECT 310.950 521.550 315.450 523.050 ;
        RECT 323.100 526.050 324.300 533.400 ;
        RECT 329.700 532.500 330.900 539.400 ;
        RECT 325.200 531.600 330.900 532.500 ;
        RECT 325.200 530.700 327.000 531.600 ;
        RECT 323.100 523.950 325.200 526.050 ;
        RECT 310.950 520.950 315.000 521.550 ;
        RECT 305.100 517.800 309.300 518.700 ;
        RECT 290.100 510.600 291.900 516.600 ;
        RECT 302.400 510.000 304.200 516.600 ;
        RECT 307.500 510.600 309.300 517.800 ;
        RECT 323.100 516.600 324.300 523.950 ;
        RECT 326.100 519.300 327.000 530.700 ;
        RECT 336.000 529.050 337.500 539.400 ;
        RECT 342.000 538.500 343.200 539.400 ;
        RECT 328.800 526.050 330.600 527.850 ;
        RECT 335.100 526.950 337.500 529.050 ;
        RECT 328.500 523.950 330.600 526.050 ;
        RECT 325.200 518.400 327.000 519.300 ;
        RECT 325.200 517.500 330.900 518.400 ;
        RECT 323.100 510.600 324.900 516.600 ;
        RECT 326.100 510.000 327.900 516.600 ;
        RECT 329.700 513.600 330.900 517.500 ;
        RECT 336.000 513.600 337.500 526.950 ;
        RECT 329.100 510.600 330.900 513.600 ;
        RECT 332.700 510.000 334.500 513.600 ;
        RECT 335.700 510.600 337.500 513.600 ;
        RECT 339.300 537.600 343.200 538.500 ;
        RECT 339.300 534.300 340.200 537.600 ;
        RECT 344.100 536.400 345.900 537.000 ;
        RECT 348.600 536.400 349.800 539.400 ;
        RECT 356.700 538.500 358.800 539.400 ;
        RECT 350.700 537.300 358.800 538.500 ;
        RECT 350.700 536.700 352.500 537.300 ;
        RECT 344.100 535.200 349.800 536.400 ;
        RECT 362.100 535.500 364.800 539.400 ;
        RECT 369.000 537.900 370.800 545.400 ;
        RECT 372.900 539.400 374.700 546.000 ;
        RECT 375.900 539.400 377.700 545.400 ;
        RECT 378.900 542.400 380.700 545.400 ;
        RECT 381.900 542.400 383.700 545.400 ;
        RECT 378.600 540.300 380.700 542.400 ;
        RECT 381.600 540.300 383.700 542.400 ;
        RECT 385.500 539.400 387.300 546.000 ;
        RECT 367.500 535.800 370.800 537.900 ;
        RECT 376.200 537.300 378.300 539.400 ;
        RECT 388.500 536.400 390.300 545.400 ;
        RECT 391.500 539.400 393.300 546.000 ;
        RECT 394.500 540.300 396.300 545.400 ;
        RECT 394.500 539.400 396.600 540.300 ;
        RECT 397.500 539.400 399.300 546.000 ;
        RECT 400.950 543.450 403.050 544.050 ;
        RECT 409.950 543.450 412.050 544.050 ;
        RECT 400.950 542.550 412.050 543.450 ;
        RECT 400.950 541.950 403.050 542.550 ;
        RECT 409.950 541.950 412.050 542.550 ;
        RECT 413.100 539.400 414.900 546.000 ;
        RECT 416.100 539.400 417.900 545.400 ;
        RECT 419.100 539.400 420.900 546.000 ;
        RECT 422.700 539.400 424.500 546.000 ;
        RECT 425.700 540.300 427.500 545.400 ;
        RECT 425.400 539.400 427.500 540.300 ;
        RECT 428.700 539.400 430.500 546.000 ;
        RECT 395.700 538.500 396.600 539.400 ;
        RECT 395.700 537.600 399.300 538.500 ;
        RECT 393.000 536.400 394.800 536.700 ;
        RECT 353.700 534.300 355.800 535.500 ;
        RECT 339.300 533.400 355.800 534.300 ;
        RECT 359.100 534.600 361.200 535.500 ;
        RECT 375.600 535.200 394.800 536.400 ;
        RECT 375.600 534.600 376.800 535.200 ;
        RECT 393.000 534.900 394.800 535.200 ;
        RECT 359.100 533.400 376.800 534.600 ;
        RECT 379.500 533.700 381.600 534.300 ;
        RECT 389.700 533.700 391.500 534.300 ;
        RECT 339.300 516.600 340.200 533.400 ;
        RECT 379.500 532.500 391.500 533.700 ;
        RECT 341.100 531.300 376.800 532.500 ;
        RECT 379.500 532.200 381.600 532.500 ;
        RECT 341.100 530.700 342.900 531.300 ;
        RECT 375.600 530.700 376.800 531.300 ;
        RECT 344.100 526.950 346.200 529.050 ;
        RECT 344.700 524.100 346.200 526.950 ;
        RECT 348.300 526.800 353.400 528.600 ;
        RECT 352.500 525.300 353.400 526.800 ;
        RECT 356.100 528.300 357.900 530.100 ;
        RECT 362.100 529.800 364.200 530.100 ;
        RECT 375.600 529.800 389.100 530.700 ;
        RECT 356.100 527.100 357.000 528.300 ;
        RECT 362.100 528.000 366.000 529.800 ;
        RECT 367.500 528.300 369.600 529.200 ;
        RECT 387.300 529.050 389.100 529.800 ;
        RECT 367.500 527.100 378.600 528.300 ;
        RECT 387.300 527.250 391.200 529.050 ;
        RECT 356.100 526.200 369.600 527.100 ;
        RECT 376.800 526.500 378.600 527.100 ;
        RECT 389.100 526.950 391.200 527.250 ;
        RECT 395.100 526.950 397.200 529.050 ;
        RECT 395.100 525.300 396.900 526.950 ;
        RECT 352.500 524.100 396.900 525.300 ;
        RECT 344.700 522.600 351.300 524.100 ;
        RECT 341.100 519.900 348.900 521.700 ;
        RECT 349.800 521.100 366.900 522.600 ;
        RECT 364.800 520.500 366.900 521.100 ;
        RECT 371.100 522.000 373.200 523.050 ;
        RECT 371.100 521.100 376.200 522.000 ;
        RECT 379.800 521.400 381.600 523.200 ;
        RECT 398.100 521.400 399.300 537.600 ;
        RECT 400.950 534.450 403.050 535.050 ;
        RECT 400.950 534.000 414.450 534.450 ;
        RECT 400.950 533.550 415.050 534.000 ;
        RECT 400.950 532.950 403.050 533.550 ;
        RECT 412.950 530.100 415.050 533.550 ;
        RECT 408.000 528.450 412.050 529.050 ;
        RECT 407.550 526.950 412.050 528.450 ;
        RECT 371.100 520.950 373.200 521.100 ;
        RECT 347.400 516.600 348.900 519.900 ;
        RECT 365.100 518.700 366.900 520.500 ;
        RECT 374.400 520.200 376.200 521.100 ;
        RECT 380.700 518.400 381.600 521.400 ;
        RECT 382.500 520.200 399.300 521.400 ;
        RECT 400.950 522.450 403.050 522.900 ;
        RECT 407.550 522.450 408.450 526.950 ;
        RECT 416.700 526.050 417.900 539.400 ;
        RECT 425.400 538.500 426.300 539.400 ;
        RECT 422.700 537.600 426.300 538.500 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 400.950 521.550 408.450 522.450 ;
        RECT 413.100 522.150 414.900 523.950 ;
        RECT 400.950 520.800 403.050 521.550 ;
        RECT 382.500 519.300 384.600 520.200 ;
        RECT 393.300 518.700 395.100 519.300 ;
        RECT 353.100 516.600 359.700 518.400 ;
        RECT 374.400 517.200 381.600 518.400 ;
        RECT 386.700 517.500 395.100 518.700 ;
        RECT 374.400 516.600 375.300 517.200 ;
        RECT 377.400 516.600 379.200 517.200 ;
        RECT 386.700 516.600 388.200 517.500 ;
        RECT 398.100 516.600 399.300 520.200 ;
        RECT 416.700 518.700 417.900 523.950 ;
        RECT 418.950 522.150 420.750 523.950 ;
        RECT 339.300 510.600 341.100 516.600 ;
        RECT 344.700 510.000 346.500 516.600 ;
        RECT 347.400 515.400 351.600 516.600 ;
        RECT 349.800 510.600 351.600 515.400 ;
        RECT 353.700 513.600 355.800 515.700 ;
        RECT 356.700 513.600 358.800 515.700 ;
        RECT 359.700 513.600 361.800 515.700 ;
        RECT 362.700 513.600 364.800 515.700 ;
        RECT 368.100 514.500 370.800 516.600 ;
        RECT 372.600 515.400 375.300 516.600 ;
        RECT 372.600 514.500 374.400 515.400 ;
        RECT 354.000 510.600 355.800 513.600 ;
        RECT 357.000 510.600 358.800 513.600 ;
        RECT 360.000 510.600 361.800 513.600 ;
        RECT 363.000 510.600 364.800 513.600 ;
        RECT 366.000 510.000 367.800 513.600 ;
        RECT 369.000 510.600 370.800 514.500 ;
        RECT 376.200 513.600 378.300 515.700 ;
        RECT 379.200 513.600 381.300 515.700 ;
        RECT 382.200 513.600 384.300 515.700 ;
        RECT 373.500 510.000 375.300 513.600 ;
        RECT 376.500 510.600 378.300 513.600 ;
        RECT 379.500 510.600 381.300 513.600 ;
        RECT 382.500 510.600 384.300 513.600 ;
        RECT 386.700 510.600 388.500 516.600 ;
        RECT 392.100 510.000 393.900 516.600 ;
        RECT 397.500 510.600 399.300 516.600 ;
        RECT 413.700 517.800 417.900 518.700 ;
        RECT 422.700 521.400 423.900 537.600 ;
        RECT 427.200 536.400 429.000 536.700 ;
        RECT 431.700 536.400 433.500 545.400 ;
        RECT 434.700 539.400 436.500 546.000 ;
        RECT 438.300 542.400 440.100 545.400 ;
        RECT 441.300 542.400 443.100 545.400 ;
        RECT 438.300 540.300 440.400 542.400 ;
        RECT 441.300 540.300 443.400 542.400 ;
        RECT 444.300 539.400 446.100 545.400 ;
        RECT 447.300 539.400 449.100 546.000 ;
        RECT 443.700 537.300 445.800 539.400 ;
        RECT 451.200 537.900 453.000 545.400 ;
        RECT 454.200 539.400 456.000 546.000 ;
        RECT 457.200 539.400 459.000 545.400 ;
        RECT 460.200 542.400 462.000 545.400 ;
        RECT 463.200 542.400 465.000 545.400 ;
        RECT 466.200 542.400 468.000 545.400 ;
        RECT 460.200 540.300 462.300 542.400 ;
        RECT 463.200 540.300 465.300 542.400 ;
        RECT 466.200 540.300 468.300 542.400 ;
        RECT 469.200 539.400 471.000 546.000 ;
        RECT 472.200 539.400 474.000 545.400 ;
        RECT 475.200 539.400 477.000 546.000 ;
        RECT 478.200 539.400 480.000 545.400 ;
        RECT 481.200 539.400 483.000 546.000 ;
        RECT 484.500 539.400 486.300 545.400 ;
        RECT 487.500 539.400 489.300 546.000 ;
        RECT 491.700 539.400 493.500 546.000 ;
        RECT 494.700 540.300 496.500 545.400 ;
        RECT 494.400 539.400 496.500 540.300 ;
        RECT 497.700 539.400 499.500 546.000 ;
        RECT 427.200 535.200 446.400 536.400 ;
        RECT 451.200 535.800 454.500 537.900 ;
        RECT 457.200 535.500 459.900 539.400 ;
        RECT 463.200 538.500 465.300 539.400 ;
        RECT 463.200 537.300 471.300 538.500 ;
        RECT 469.500 536.700 471.300 537.300 ;
        RECT 472.200 536.400 473.400 539.400 ;
        RECT 478.800 538.500 480.000 539.400 ;
        RECT 478.800 537.600 482.700 538.500 ;
        RECT 476.100 536.400 477.900 537.000 ;
        RECT 427.200 534.900 429.000 535.200 ;
        RECT 445.200 534.600 446.400 535.200 ;
        RECT 460.800 534.600 462.900 535.500 ;
        RECT 430.500 533.700 432.300 534.300 ;
        RECT 440.400 533.700 442.500 534.300 ;
        RECT 430.500 532.500 442.500 533.700 ;
        RECT 445.200 533.400 462.900 534.600 ;
        RECT 466.200 534.300 468.300 535.500 ;
        RECT 472.200 535.200 477.900 536.400 ;
        RECT 481.800 534.300 482.700 537.600 ;
        RECT 466.200 533.400 482.700 534.300 ;
        RECT 440.400 532.200 442.500 532.500 ;
        RECT 445.200 531.300 480.900 532.500 ;
        RECT 445.200 530.700 446.400 531.300 ;
        RECT 479.100 530.700 480.900 531.300 ;
        RECT 432.900 529.800 446.400 530.700 ;
        RECT 457.800 529.800 459.900 530.100 ;
        RECT 432.900 529.050 434.700 529.800 ;
        RECT 424.800 526.950 426.900 529.050 ;
        RECT 430.800 527.250 434.700 529.050 ;
        RECT 452.400 528.300 454.500 529.200 ;
        RECT 430.800 526.950 432.900 527.250 ;
        RECT 443.400 527.100 454.500 528.300 ;
        RECT 456.000 528.000 459.900 529.800 ;
        RECT 464.100 528.300 465.900 530.100 ;
        RECT 465.000 527.100 465.900 528.300 ;
        RECT 425.100 525.300 426.900 526.950 ;
        RECT 443.400 526.500 445.200 527.100 ;
        RECT 452.400 526.200 465.900 527.100 ;
        RECT 468.600 526.800 473.700 528.600 ;
        RECT 475.800 526.950 477.900 529.050 ;
        RECT 468.600 525.300 469.500 526.800 ;
        RECT 425.100 524.100 469.500 525.300 ;
        RECT 475.800 524.100 477.300 526.950 ;
        RECT 440.400 521.400 442.200 523.200 ;
        RECT 448.800 522.000 450.900 523.050 ;
        RECT 470.700 522.600 477.300 524.100 ;
        RECT 422.700 520.200 439.500 521.400 ;
        RECT 413.700 510.600 415.500 517.800 ;
        RECT 422.700 516.600 423.900 520.200 ;
        RECT 437.400 519.300 439.500 520.200 ;
        RECT 426.900 518.700 428.700 519.300 ;
        RECT 426.900 517.500 435.300 518.700 ;
        RECT 433.800 516.600 435.300 517.500 ;
        RECT 440.400 518.400 441.300 521.400 ;
        RECT 445.800 521.100 450.900 522.000 ;
        RECT 445.800 520.200 447.600 521.100 ;
        RECT 448.800 520.950 450.900 521.100 ;
        RECT 455.100 521.100 472.200 522.600 ;
        RECT 455.100 520.500 457.200 521.100 ;
        RECT 455.100 518.700 456.900 520.500 ;
        RECT 473.100 519.900 480.900 521.700 ;
        RECT 440.400 517.200 447.600 518.400 ;
        RECT 442.800 516.600 444.600 517.200 ;
        RECT 446.700 516.600 447.600 517.200 ;
        RECT 462.300 516.600 468.900 518.400 ;
        RECT 473.100 516.600 474.600 519.900 ;
        RECT 481.800 516.600 482.700 533.400 ;
        RECT 418.800 510.000 420.600 516.600 ;
        RECT 422.700 510.600 424.500 516.600 ;
        RECT 428.100 510.000 429.900 516.600 ;
        RECT 433.500 510.600 435.300 516.600 ;
        RECT 437.700 513.600 439.800 515.700 ;
        RECT 440.700 513.600 442.800 515.700 ;
        RECT 443.700 513.600 445.800 515.700 ;
        RECT 446.700 515.400 449.400 516.600 ;
        RECT 447.600 514.500 449.400 515.400 ;
        RECT 451.200 514.500 453.900 516.600 ;
        RECT 437.700 510.600 439.500 513.600 ;
        RECT 440.700 510.600 442.500 513.600 ;
        RECT 443.700 510.600 445.500 513.600 ;
        RECT 446.700 510.000 448.500 513.600 ;
        RECT 451.200 510.600 453.000 514.500 ;
        RECT 457.200 513.600 459.300 515.700 ;
        RECT 460.200 513.600 462.300 515.700 ;
        RECT 463.200 513.600 465.300 515.700 ;
        RECT 466.200 513.600 468.300 515.700 ;
        RECT 470.400 515.400 474.600 516.600 ;
        RECT 454.200 510.000 456.000 513.600 ;
        RECT 457.200 510.600 459.000 513.600 ;
        RECT 460.200 510.600 462.000 513.600 ;
        RECT 463.200 510.600 465.000 513.600 ;
        RECT 466.200 510.600 468.000 513.600 ;
        RECT 470.400 510.600 472.200 515.400 ;
        RECT 475.500 510.000 477.300 516.600 ;
        RECT 480.900 510.600 482.700 516.600 ;
        RECT 484.500 529.050 486.000 539.400 ;
        RECT 494.400 538.500 495.300 539.400 ;
        RECT 491.700 537.600 495.300 538.500 ;
        RECT 484.500 526.950 486.900 529.050 ;
        RECT 484.500 513.600 486.000 526.950 ;
        RECT 491.700 521.400 492.900 537.600 ;
        RECT 496.200 536.400 498.000 536.700 ;
        RECT 500.700 536.400 502.500 545.400 ;
        RECT 503.700 539.400 505.500 546.000 ;
        RECT 507.300 542.400 509.100 545.400 ;
        RECT 510.300 542.400 512.100 545.400 ;
        RECT 507.300 540.300 509.400 542.400 ;
        RECT 510.300 540.300 512.400 542.400 ;
        RECT 513.300 539.400 515.100 545.400 ;
        RECT 516.300 539.400 518.100 546.000 ;
        RECT 512.700 537.300 514.800 539.400 ;
        RECT 520.200 537.900 522.000 545.400 ;
        RECT 523.200 539.400 525.000 546.000 ;
        RECT 526.200 539.400 528.000 545.400 ;
        RECT 529.200 542.400 531.000 545.400 ;
        RECT 532.200 542.400 534.000 545.400 ;
        RECT 535.200 542.400 537.000 545.400 ;
        RECT 529.200 540.300 531.300 542.400 ;
        RECT 532.200 540.300 534.300 542.400 ;
        RECT 535.200 540.300 537.300 542.400 ;
        RECT 538.200 539.400 540.000 546.000 ;
        RECT 541.200 539.400 543.000 545.400 ;
        RECT 544.200 539.400 546.000 546.000 ;
        RECT 547.200 539.400 549.000 545.400 ;
        RECT 550.200 539.400 552.000 546.000 ;
        RECT 553.500 539.400 555.300 545.400 ;
        RECT 556.500 539.400 558.300 546.000 ;
        RECT 569.100 539.400 570.900 546.000 ;
        RECT 572.100 539.400 573.900 545.400 ;
        RECT 575.100 539.400 576.900 546.000 ;
        RECT 590.100 539.400 591.900 546.000 ;
        RECT 593.100 539.400 594.900 545.400 ;
        RECT 596.100 539.400 597.900 546.000 ;
        RECT 496.200 535.200 515.400 536.400 ;
        RECT 520.200 535.800 523.500 537.900 ;
        RECT 526.200 535.500 528.900 539.400 ;
        RECT 532.200 538.500 534.300 539.400 ;
        RECT 532.200 537.300 540.300 538.500 ;
        RECT 538.500 536.700 540.300 537.300 ;
        RECT 541.200 536.400 542.400 539.400 ;
        RECT 547.800 538.500 549.000 539.400 ;
        RECT 547.800 537.600 551.700 538.500 ;
        RECT 545.100 536.400 546.900 537.000 ;
        RECT 496.200 534.900 498.000 535.200 ;
        RECT 514.200 534.600 515.400 535.200 ;
        RECT 529.800 534.600 531.900 535.500 ;
        RECT 499.500 533.700 501.300 534.300 ;
        RECT 509.400 533.700 511.500 534.300 ;
        RECT 499.500 532.500 511.500 533.700 ;
        RECT 514.200 533.400 531.900 534.600 ;
        RECT 535.200 534.300 537.300 535.500 ;
        RECT 541.200 535.200 546.900 536.400 ;
        RECT 550.800 534.300 551.700 537.600 ;
        RECT 535.200 533.400 551.700 534.300 ;
        RECT 509.400 532.200 511.500 532.500 ;
        RECT 514.200 531.300 549.900 532.500 ;
        RECT 514.200 530.700 515.400 531.300 ;
        RECT 548.100 530.700 549.900 531.300 ;
        RECT 501.900 529.800 515.400 530.700 ;
        RECT 526.800 529.800 528.900 530.100 ;
        RECT 501.900 529.050 503.700 529.800 ;
        RECT 493.800 526.950 495.900 529.050 ;
        RECT 499.800 527.250 503.700 529.050 ;
        RECT 521.400 528.300 523.500 529.200 ;
        RECT 499.800 526.950 501.900 527.250 ;
        RECT 512.400 527.100 523.500 528.300 ;
        RECT 525.000 528.000 528.900 529.800 ;
        RECT 533.100 528.300 534.900 530.100 ;
        RECT 534.000 527.100 534.900 528.300 ;
        RECT 494.100 525.300 495.900 526.950 ;
        RECT 512.400 526.500 514.200 527.100 ;
        RECT 521.400 526.200 534.900 527.100 ;
        RECT 537.600 526.800 542.700 528.600 ;
        RECT 544.800 526.950 546.900 529.050 ;
        RECT 537.600 525.300 538.500 526.800 ;
        RECT 494.100 524.100 538.500 525.300 ;
        RECT 544.800 524.100 546.300 526.950 ;
        RECT 509.400 521.400 511.200 523.200 ;
        RECT 517.800 522.000 519.900 523.050 ;
        RECT 539.700 522.600 546.300 524.100 ;
        RECT 491.700 520.200 508.500 521.400 ;
        RECT 491.700 516.600 492.900 520.200 ;
        RECT 506.400 519.300 508.500 520.200 ;
        RECT 495.900 518.700 497.700 519.300 ;
        RECT 495.900 517.500 504.300 518.700 ;
        RECT 502.800 516.600 504.300 517.500 ;
        RECT 509.400 518.400 510.300 521.400 ;
        RECT 514.800 521.100 519.900 522.000 ;
        RECT 514.800 520.200 516.600 521.100 ;
        RECT 517.800 520.950 519.900 521.100 ;
        RECT 524.100 521.100 541.200 522.600 ;
        RECT 524.100 520.500 526.200 521.100 ;
        RECT 524.100 518.700 525.900 520.500 ;
        RECT 542.100 519.900 549.900 521.700 ;
        RECT 509.400 517.200 516.600 518.400 ;
        RECT 511.800 516.600 513.600 517.200 ;
        RECT 515.700 516.600 516.600 517.200 ;
        RECT 531.300 516.600 537.900 518.400 ;
        RECT 542.100 516.600 543.600 519.900 ;
        RECT 550.800 516.600 551.700 533.400 ;
        RECT 484.500 510.600 486.300 513.600 ;
        RECT 487.500 510.000 489.300 513.600 ;
        RECT 491.700 510.600 493.500 516.600 ;
        RECT 497.100 510.000 498.900 516.600 ;
        RECT 502.500 510.600 504.300 516.600 ;
        RECT 506.700 513.600 508.800 515.700 ;
        RECT 509.700 513.600 511.800 515.700 ;
        RECT 512.700 513.600 514.800 515.700 ;
        RECT 515.700 515.400 518.400 516.600 ;
        RECT 516.600 514.500 518.400 515.400 ;
        RECT 520.200 514.500 522.900 516.600 ;
        RECT 506.700 510.600 508.500 513.600 ;
        RECT 509.700 510.600 511.500 513.600 ;
        RECT 512.700 510.600 514.500 513.600 ;
        RECT 515.700 510.000 517.500 513.600 ;
        RECT 520.200 510.600 522.000 514.500 ;
        RECT 526.200 513.600 528.300 515.700 ;
        RECT 529.200 513.600 531.300 515.700 ;
        RECT 532.200 513.600 534.300 515.700 ;
        RECT 535.200 513.600 537.300 515.700 ;
        RECT 539.400 515.400 543.600 516.600 ;
        RECT 523.200 510.000 525.000 513.600 ;
        RECT 526.200 510.600 528.000 513.600 ;
        RECT 529.200 510.600 531.000 513.600 ;
        RECT 532.200 510.600 534.000 513.600 ;
        RECT 535.200 510.600 537.000 513.600 ;
        RECT 539.400 510.600 541.200 515.400 ;
        RECT 544.500 510.000 546.300 516.600 ;
        RECT 549.900 510.600 551.700 516.600 ;
        RECT 553.500 529.050 555.000 539.400 ;
        RECT 553.500 526.950 555.900 529.050 ;
        RECT 553.500 513.600 555.000 526.950 ;
        RECT 572.100 526.050 573.300 539.400 ;
        RECT 593.100 526.050 594.300 539.400 ;
        RECT 608.100 533.400 609.900 546.000 ;
        RECT 611.100 533.400 612.900 545.400 ;
        RECT 626.400 533.400 628.200 546.000 ;
        RECT 631.500 534.900 633.300 545.400 ;
        RECT 634.500 539.400 636.300 546.000 ;
        RECT 634.200 536.100 636.000 537.900 ;
        RECT 631.500 533.400 633.900 534.900 ;
        RECT 650.400 533.400 652.200 546.000 ;
        RECT 655.500 534.900 657.300 545.400 ;
        RECT 658.500 539.400 660.300 546.000 ;
        RECT 671.100 539.400 672.900 546.000 ;
        RECT 674.100 539.400 675.900 545.400 ;
        RECT 689.100 539.400 690.900 546.000 ;
        RECT 692.100 539.400 693.900 545.400 ;
        RECT 695.100 540.000 696.900 546.000 ;
        RECT 658.200 536.100 660.000 537.900 ;
        RECT 655.500 533.400 657.900 534.900 ;
        RECT 611.100 526.050 612.300 533.400 ;
        RECT 626.100 526.050 627.900 527.850 ;
        RECT 632.700 526.050 633.900 533.400 ;
        RECT 650.100 526.050 651.900 527.850 ;
        RECT 656.700 526.050 657.900 533.400 ;
        RECT 661.950 528.450 666.000 529.050 ;
        RECT 661.950 526.950 666.450 528.450 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 607.950 523.950 610.050 526.050 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 631.950 523.950 634.050 526.050 ;
        RECT 634.950 523.950 637.050 526.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 569.250 522.150 571.050 523.950 ;
        RECT 572.100 518.700 573.300 523.950 ;
        RECT 575.100 522.150 576.900 523.950 ;
        RECT 590.250 522.150 592.050 523.950 ;
        RECT 593.100 518.700 594.300 523.950 ;
        RECT 596.100 522.150 597.900 523.950 ;
        RECT 608.100 522.150 609.900 523.950 ;
        RECT 572.100 517.800 576.300 518.700 ;
        RECT 593.100 517.800 597.300 518.700 ;
        RECT 553.500 510.600 555.300 513.600 ;
        RECT 556.500 510.000 558.300 513.600 ;
        RECT 569.400 510.000 571.200 516.600 ;
        RECT 574.500 510.600 576.300 517.800 ;
        RECT 590.400 510.000 592.200 516.600 ;
        RECT 595.500 510.600 597.300 517.800 ;
        RECT 611.100 516.600 612.300 523.950 ;
        RECT 629.100 522.150 630.900 523.950 ;
        RECT 632.700 519.600 633.900 523.950 ;
        RECT 635.100 522.150 636.900 523.950 ;
        RECT 653.100 522.150 654.900 523.950 ;
        RECT 656.700 519.600 657.900 523.950 ;
        RECT 659.100 522.150 660.900 523.950 ;
        RECT 665.550 523.050 666.450 526.950 ;
        RECT 671.100 526.050 672.900 527.850 ;
        RECT 674.100 526.050 675.300 539.400 ;
        RECT 692.400 539.100 693.900 539.400 ;
        RECT 698.100 539.400 699.900 545.400 ;
        RECT 698.100 539.100 699.000 539.400 ;
        RECT 692.400 538.200 699.000 539.100 ;
        RECT 676.950 531.450 679.050 532.050 ;
        RECT 688.950 531.450 691.050 532.050 ;
        RECT 676.950 530.550 691.050 531.450 ;
        RECT 676.950 529.950 679.050 530.550 ;
        RECT 688.950 529.950 691.050 530.550 ;
        RECT 692.100 526.050 693.900 527.850 ;
        RECT 698.100 526.050 699.000 538.200 ;
        RECT 713.400 533.400 715.200 546.000 ;
        RECT 718.500 534.900 720.300 545.400 ;
        RECT 721.500 539.400 723.300 546.000 ;
        RECT 737.700 539.400 739.500 546.000 ;
        RECT 721.200 536.100 723.000 537.900 ;
        RECT 738.000 536.100 739.800 537.900 ;
        RECT 740.700 534.900 742.500 545.400 ;
        RECT 718.500 533.400 720.900 534.900 ;
        RECT 713.100 526.050 714.900 527.850 ;
        RECT 719.700 526.050 720.900 533.400 ;
        RECT 740.100 533.400 742.500 534.900 ;
        RECT 745.800 533.400 747.600 546.000 ;
        RECT 758.100 539.400 759.900 545.400 ;
        RECT 761.100 539.400 762.900 546.000 ;
        RECT 724.950 528.450 729.000 529.050 ;
        RECT 724.950 526.950 729.450 528.450 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 694.950 523.950 697.050 526.050 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 665.550 521.550 670.050 523.050 ;
        RECT 666.000 520.950 670.050 521.550 ;
        RECT 632.700 518.700 636.300 519.600 ;
        RECT 656.700 518.700 660.300 519.600 ;
        RECT 608.100 510.000 609.900 516.600 ;
        RECT 611.100 510.600 612.900 516.600 ;
        RECT 626.100 515.700 633.900 517.050 ;
        RECT 626.100 510.600 627.900 515.700 ;
        RECT 629.100 510.000 630.900 514.800 ;
        RECT 632.100 510.600 633.900 515.700 ;
        RECT 635.100 516.600 636.300 518.700 ;
        RECT 635.100 510.600 636.900 516.600 ;
        RECT 650.100 515.700 657.900 517.050 ;
        RECT 650.100 510.600 651.900 515.700 ;
        RECT 653.100 510.000 654.900 514.800 ;
        RECT 656.100 510.600 657.900 515.700 ;
        RECT 659.100 516.600 660.300 518.700 ;
        RECT 659.100 510.600 660.900 516.600 ;
        RECT 674.100 513.600 675.300 523.950 ;
        RECT 689.100 522.150 690.900 523.950 ;
        RECT 695.100 522.150 696.900 523.950 ;
        RECT 698.100 520.200 699.000 523.950 ;
        RECT 716.100 522.150 717.900 523.950 ;
        RECT 671.100 510.000 672.900 513.600 ;
        RECT 674.100 510.600 675.900 513.600 ;
        RECT 689.100 510.000 690.900 519.600 ;
        RECT 695.700 519.000 699.000 520.200 ;
        RECT 719.700 519.600 720.900 523.950 ;
        RECT 722.100 522.150 723.900 523.950 ;
        RECT 728.550 522.450 729.450 526.950 ;
        RECT 740.100 526.050 741.300 533.400 ;
        RECT 748.950 528.450 753.000 529.050 ;
        RECT 746.100 526.050 747.900 527.850 ;
        RECT 748.950 526.950 753.450 528.450 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 725.550 522.000 729.450 522.450 ;
        RECT 737.100 522.150 738.900 523.950 ;
        RECT 724.950 521.550 729.450 522.000 ;
        RECT 695.700 510.600 697.500 519.000 ;
        RECT 719.700 518.700 723.300 519.600 ;
        RECT 713.100 515.700 720.900 517.050 ;
        RECT 713.100 510.600 714.900 515.700 ;
        RECT 716.100 510.000 717.900 514.800 ;
        RECT 719.100 510.600 720.900 515.700 ;
        RECT 722.100 516.600 723.300 518.700 ;
        RECT 724.950 517.950 727.050 521.550 ;
        RECT 740.100 519.600 741.300 523.950 ;
        RECT 743.100 522.150 744.900 523.950 ;
        RECT 752.550 523.050 753.450 526.950 ;
        RECT 758.700 526.050 759.900 539.400 ;
        RECT 773.100 534.300 774.900 545.400 ;
        RECT 776.100 535.500 777.900 546.000 ;
        RECT 773.100 533.400 777.600 534.300 ;
        RECT 780.600 533.400 782.400 545.400 ;
        RECT 785.100 535.500 786.900 546.000 ;
        RECT 788.100 534.600 789.900 545.400 ;
        RECT 800.700 539.400 802.500 546.000 ;
        RECT 801.000 536.100 802.800 537.900 ;
        RECT 803.700 534.900 805.500 545.400 ;
        RECT 775.500 531.300 777.600 533.400 ;
        RECT 781.200 532.050 782.400 533.400 ;
        RECT 785.100 533.400 789.900 534.600 ;
        RECT 803.100 533.400 805.500 534.900 ;
        RECT 808.800 533.400 810.600 546.000 ;
        RECT 824.100 539.400 825.900 546.000 ;
        RECT 827.100 539.400 828.900 545.400 ;
        RECT 785.100 532.500 787.200 533.400 ;
        RECT 781.200 531.000 782.700 532.050 ;
        RECT 778.800 529.500 780.900 529.800 ;
        RECT 761.100 526.050 762.900 527.850 ;
        RECT 777.000 527.700 780.900 529.500 ;
        RECT 781.800 529.050 782.700 531.000 ;
        RECT 781.800 526.950 783.900 529.050 ;
        RECT 781.800 526.800 783.300 526.950 ;
        RECT 778.200 526.050 780.000 526.500 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 773.100 524.700 780.000 526.050 ;
        RECT 780.900 525.900 783.300 526.800 ;
        RECT 787.800 526.050 789.600 527.850 ;
        RECT 803.100 526.050 804.300 533.400 ;
        RECT 809.100 526.050 810.900 527.850 ;
        RECT 773.100 523.950 775.200 524.700 ;
        RECT 752.550 521.550 757.050 523.050 ;
        RECT 753.000 520.950 757.050 521.550 ;
        RECT 737.700 518.700 741.300 519.600 ;
        RECT 737.700 516.600 738.900 518.700 ;
        RECT 722.100 510.600 723.900 516.600 ;
        RECT 737.100 510.600 738.900 516.600 ;
        RECT 740.100 515.700 747.900 517.050 ;
        RECT 740.100 510.600 741.900 515.700 ;
        RECT 743.100 510.000 744.900 514.800 ;
        RECT 746.100 510.600 747.900 515.700 ;
        RECT 758.700 513.600 759.900 523.950 ;
        RECT 773.400 522.150 775.200 523.950 ;
        RECT 778.200 521.400 780.000 523.200 ;
        RECT 763.950 519.450 766.050 519.900 ;
        RECT 769.950 519.450 772.050 520.050 ;
        RECT 763.950 518.550 772.050 519.450 ;
        RECT 777.900 519.300 780.000 521.400 ;
        RECT 763.950 517.800 766.050 518.550 ;
        RECT 769.950 517.950 772.050 518.550 ;
        RECT 773.700 518.400 780.000 519.300 ;
        RECT 780.900 520.200 782.100 525.900 ;
        RECT 783.300 523.200 785.100 525.000 ;
        RECT 787.800 523.950 789.900 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 808.950 523.950 811.050 526.050 ;
        RECT 824.100 523.950 826.200 526.050 ;
        RECT 783.000 521.100 785.100 523.200 ;
        RECT 800.100 522.150 801.900 523.950 ;
        RECT 773.700 516.600 774.900 518.400 ;
        RECT 780.900 518.100 783.900 520.200 ;
        RECT 803.100 519.600 804.300 523.950 ;
        RECT 806.100 522.150 807.900 523.950 ;
        RECT 824.250 522.150 826.050 523.950 ;
        RECT 800.700 518.700 804.300 519.600 ;
        RECT 827.100 519.300 828.000 539.400 ;
        RECT 830.100 534.000 831.900 546.000 ;
        RECT 833.100 533.400 834.900 545.400 ;
        RECT 845.100 539.400 846.900 546.000 ;
        RECT 848.100 539.400 849.900 545.400 ;
        RECT 851.100 540.000 852.900 546.000 ;
        RECT 848.400 539.100 849.900 539.400 ;
        RECT 854.100 539.400 855.900 545.400 ;
        RECT 854.100 539.100 855.000 539.400 ;
        RECT 848.400 538.200 855.000 539.100 ;
        RECT 829.200 526.050 831.000 527.850 ;
        RECT 833.400 526.050 834.300 533.400 ;
        RECT 848.100 526.050 849.900 527.850 ;
        RECT 854.100 526.050 855.000 538.200 ;
        RECT 869.100 534.600 870.900 545.400 ;
        RECT 872.100 535.500 873.900 546.000 ;
        RECT 875.100 544.500 882.900 545.400 ;
        RECT 875.100 534.600 876.900 544.500 ;
        RECT 869.100 533.700 876.900 534.600 ;
        RECT 878.100 532.500 879.900 543.600 ;
        RECT 881.100 533.400 882.900 544.500 ;
        RECT 896.100 533.400 897.900 546.000 ;
        RECT 901.200 534.600 903.000 545.400 ;
        RECT 917.100 539.400 918.900 545.400 ;
        RECT 920.100 539.400 921.900 546.000 ;
        RECT 935.100 539.400 936.900 546.000 ;
        RECT 938.100 539.400 939.900 545.400 ;
        RECT 941.100 539.400 942.900 546.000 ;
        RECT 899.400 533.400 903.000 534.600 ;
        RECT 875.100 531.600 879.900 532.500 ;
        RECT 872.250 526.050 874.050 527.850 ;
        RECT 875.100 526.050 876.000 531.600 ;
        RECT 880.950 531.450 883.050 532.050 ;
        RECT 886.950 531.450 889.050 532.050 ;
        RECT 895.950 531.450 898.050 532.050 ;
        RECT 880.950 530.550 898.050 531.450 ;
        RECT 880.950 529.950 883.050 530.550 ;
        RECT 886.950 529.950 889.050 530.550 ;
        RECT 895.950 529.950 898.050 530.550 ;
        RECT 878.100 526.050 879.900 527.850 ;
        RECT 896.250 526.050 898.050 527.850 ;
        RECT 899.400 526.050 900.300 533.400 ;
        RECT 902.100 526.050 903.900 527.850 ;
        RECT 917.700 526.050 918.900 539.400 ;
        RECT 920.100 526.050 921.900 527.850 ;
        RECT 938.100 526.050 939.300 539.400 ;
        RECT 829.500 523.950 831.600 526.050 ;
        RECT 832.800 523.950 834.900 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 850.950 523.950 853.050 526.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 880.950 523.950 883.050 526.050 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 916.950 523.950 919.050 526.050 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 934.950 523.950 937.050 526.050 ;
        RECT 937.950 523.950 940.050 526.050 ;
        RECT 940.950 523.950 943.050 526.050 ;
        RECT 780.900 516.600 782.100 518.100 ;
        RECT 785.100 517.500 787.200 518.700 ;
        RECT 785.100 516.600 789.900 517.500 ;
        RECT 800.700 516.600 801.900 518.700 ;
        RECT 824.100 518.400 832.500 519.300 ;
        RECT 758.100 510.600 759.900 513.600 ;
        RECT 761.100 510.000 762.900 513.600 ;
        RECT 773.100 510.600 774.900 516.600 ;
        RECT 776.100 510.000 777.900 515.700 ;
        RECT 780.600 510.600 782.400 516.600 ;
        RECT 785.100 510.000 786.900 515.700 ;
        RECT 788.100 510.600 789.900 516.600 ;
        RECT 800.100 510.600 801.900 516.600 ;
        RECT 803.100 515.700 810.900 517.050 ;
        RECT 803.100 510.600 804.900 515.700 ;
        RECT 806.100 510.000 807.900 514.800 ;
        RECT 809.100 510.600 810.900 515.700 ;
        RECT 824.100 510.600 825.900 518.400 ;
        RECT 830.700 517.500 832.500 518.400 ;
        RECT 833.400 516.600 834.300 523.950 ;
        RECT 845.100 522.150 846.900 523.950 ;
        RECT 851.100 522.150 852.900 523.950 ;
        RECT 854.100 520.200 855.000 523.950 ;
        RECT 869.250 522.150 871.050 523.950 ;
        RECT 828.600 510.000 830.400 516.600 ;
        RECT 831.600 514.800 834.300 516.600 ;
        RECT 831.600 510.600 833.400 514.800 ;
        RECT 845.100 510.000 846.900 519.600 ;
        RECT 851.700 519.000 855.000 520.200 ;
        RECT 851.700 510.600 853.500 519.000 ;
        RECT 875.100 516.600 876.300 523.950 ;
        RECT 881.100 522.150 882.900 523.950 ;
        RECT 869.700 510.000 871.500 516.600 ;
        RECT 874.200 510.600 876.000 516.600 ;
        RECT 878.700 510.000 880.500 516.600 ;
        RECT 899.400 513.600 900.300 523.950 ;
        RECT 917.700 513.600 918.900 523.950 ;
        RECT 935.250 522.150 937.050 523.950 ;
        RECT 919.950 519.450 922.050 520.050 ;
        RECT 925.950 519.450 928.050 519.900 ;
        RECT 919.950 518.550 928.050 519.450 ;
        RECT 919.950 517.950 922.050 518.550 ;
        RECT 925.950 517.800 928.050 518.550 ;
        RECT 938.100 518.700 939.300 523.950 ;
        RECT 941.100 522.150 942.900 523.950 ;
        RECT 938.100 517.800 942.300 518.700 ;
        RECT 896.100 510.000 897.900 513.600 ;
        RECT 899.100 510.600 900.900 513.600 ;
        RECT 902.100 510.000 903.900 513.600 ;
        RECT 917.100 510.600 918.900 513.600 ;
        RECT 920.100 510.000 921.900 513.600 ;
        RECT 935.400 510.000 937.200 516.600 ;
        RECT 940.500 510.600 942.300 517.800 ;
        RECT 14.100 503.400 15.900 507.000 ;
        RECT 17.100 503.400 18.900 506.400 ;
        RECT 20.100 503.400 21.900 507.000 ;
        RECT 17.700 493.050 18.600 503.400 ;
        RECT 32.100 501.300 33.900 506.400 ;
        RECT 35.100 502.200 36.900 507.000 ;
        RECT 38.100 501.300 39.900 506.400 ;
        RECT 32.100 499.950 39.900 501.300 ;
        RECT 41.100 500.400 42.900 506.400 ;
        RECT 41.100 498.300 42.300 500.400 ;
        RECT 56.700 499.200 58.500 506.400 ;
        RECT 61.800 500.400 63.600 507.000 ;
        RECT 56.700 498.300 60.900 499.200 ;
        RECT 38.700 497.400 42.300 498.300 ;
        RECT 35.100 493.050 36.900 494.850 ;
        RECT 38.700 493.050 39.900 497.400 ;
        RECT 52.950 495.450 55.050 496.050 ;
        RECT 41.100 493.050 42.900 494.850 ;
        RECT 47.550 494.550 55.050 495.450 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 31.950 490.950 34.050 493.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 14.100 489.150 15.900 490.950 ;
        RECT 17.700 483.600 18.600 490.950 ;
        RECT 19.950 489.150 21.750 490.950 ;
        RECT 32.100 489.150 33.900 490.950 ;
        RECT 38.700 483.600 39.900 490.950 ;
        RECT 47.550 490.050 48.450 494.550 ;
        RECT 52.950 493.950 55.050 494.550 ;
        RECT 56.100 493.050 57.900 494.850 ;
        RECT 59.700 493.050 60.900 498.300 ;
        RECT 77.100 497.400 78.900 507.000 ;
        RECT 83.700 498.000 85.500 506.400 ;
        RECT 100.500 500.400 102.300 507.000 ;
        RECT 105.000 500.400 106.800 506.400 ;
        RECT 109.500 500.400 111.300 507.000 ;
        RECT 125.100 500.400 126.900 506.400 ;
        RECT 83.700 496.800 87.000 498.000 ;
        RECT 64.950 495.450 67.050 496.050 ;
        RECT 70.950 495.450 73.050 496.050 ;
        RECT 61.950 493.050 63.750 494.850 ;
        RECT 64.950 494.550 73.050 495.450 ;
        RECT 64.950 493.950 67.050 494.550 ;
        RECT 70.950 493.950 73.050 494.550 ;
        RECT 77.100 493.050 78.900 494.850 ;
        RECT 83.100 493.050 84.900 494.850 ;
        RECT 86.100 493.050 87.000 496.800 ;
        RECT 98.100 493.050 99.900 494.850 ;
        RECT 104.700 493.050 105.900 500.400 ;
        RECT 125.700 498.300 126.900 500.400 ;
        RECT 128.100 501.300 129.900 506.400 ;
        RECT 131.100 502.200 132.900 507.000 ;
        RECT 134.100 501.300 135.900 506.400 ;
        RECT 128.100 499.950 135.900 501.300 ;
        RECT 149.100 500.400 150.900 506.400 ;
        RECT 152.100 500.400 153.900 507.000 ;
        RECT 164.100 501.300 165.900 506.400 ;
        RECT 167.100 502.200 168.900 507.000 ;
        RECT 170.100 501.300 171.900 506.400 ;
        RECT 136.950 498.450 139.050 499.050 ;
        RECT 142.950 498.450 145.050 499.050 ;
        RECT 125.700 497.400 129.300 498.300 ;
        RECT 109.950 493.050 111.750 494.850 ;
        RECT 125.100 493.050 126.900 494.850 ;
        RECT 128.100 493.050 129.300 497.400 ;
        RECT 136.950 497.550 145.050 498.450 ;
        RECT 136.950 496.950 139.050 497.550 ;
        RECT 142.950 496.950 145.050 497.550 ;
        RECT 131.100 493.050 132.900 494.850 ;
        RECT 149.700 493.050 150.900 500.400 ;
        RECT 164.100 499.950 171.900 501.300 ;
        RECT 173.100 500.400 174.900 506.400 ;
        RECT 189.000 500.400 190.800 507.000 ;
        RECT 193.500 501.600 195.300 506.400 ;
        RECT 196.500 503.400 198.300 507.000 ;
        RECT 193.500 500.400 198.600 501.600 ;
        RECT 173.100 498.300 174.300 500.400 ;
        RECT 170.700 497.400 174.300 498.300 ;
        RECT 152.100 493.050 153.900 494.850 ;
        RECT 167.100 493.050 168.900 494.850 ;
        RECT 170.700 493.050 171.900 497.400 ;
        RECT 175.950 495.450 178.050 499.050 ;
        RECT 175.950 495.000 183.450 495.450 ;
        RECT 173.100 493.050 174.900 494.850 ;
        RECT 176.550 494.550 183.450 495.000 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 133.950 490.950 136.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 163.950 490.950 166.050 493.050 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 43.950 488.550 48.450 490.050 ;
        RECT 43.950 487.950 48.000 488.550 ;
        RECT 15.000 482.400 18.600 483.600 ;
        RECT 15.000 471.600 16.800 482.400 ;
        RECT 20.100 471.000 21.900 483.600 ;
        RECT 32.400 471.000 34.200 483.600 ;
        RECT 37.500 482.100 39.900 483.600 ;
        RECT 37.500 471.600 39.300 482.100 ;
        RECT 40.200 479.100 42.000 480.900 ;
        RECT 59.700 477.600 60.900 490.950 ;
        RECT 80.100 489.150 81.900 490.950 ;
        RECT 61.950 486.450 64.050 487.050 ;
        RECT 82.950 486.450 85.050 487.050 ;
        RECT 61.950 485.550 85.050 486.450 ;
        RECT 61.950 484.950 64.050 485.550 ;
        RECT 82.950 484.950 85.050 485.550 ;
        RECT 86.100 478.800 87.000 490.950 ;
        RECT 101.100 489.150 102.900 490.950 ;
        RECT 105.000 485.400 105.900 490.950 ;
        RECT 106.950 489.150 108.750 490.950 ;
        RECT 101.100 484.500 105.900 485.400 ;
        RECT 80.400 477.900 87.000 478.800 ;
        RECT 80.400 477.600 81.900 477.900 ;
        RECT 40.500 471.000 42.300 477.600 ;
        RECT 56.100 471.000 57.900 477.600 ;
        RECT 59.100 471.600 60.900 477.600 ;
        RECT 62.100 471.000 63.900 477.600 ;
        RECT 77.100 471.000 78.900 477.600 ;
        RECT 80.100 471.600 81.900 477.600 ;
        RECT 86.100 477.600 87.000 477.900 ;
        RECT 83.100 471.000 84.900 477.000 ;
        RECT 86.100 471.600 87.900 477.600 ;
        RECT 98.100 472.500 99.900 483.600 ;
        RECT 101.100 473.400 102.900 484.500 ;
        RECT 112.950 483.450 115.050 484.050 ;
        RECT 121.950 483.450 124.050 484.050 ;
        RECT 104.100 482.400 111.900 483.300 ;
        RECT 104.100 472.500 105.900 482.400 ;
        RECT 98.100 471.600 105.900 472.500 ;
        RECT 107.100 471.000 108.900 481.500 ;
        RECT 110.100 471.600 111.900 482.400 ;
        RECT 112.950 482.550 124.050 483.450 ;
        RECT 112.950 481.950 115.050 482.550 ;
        RECT 121.950 481.950 124.050 482.550 ;
        RECT 128.100 483.600 129.300 490.950 ;
        RECT 134.100 489.150 135.900 490.950 ;
        RECT 130.950 486.450 133.050 487.050 ;
        RECT 145.950 486.450 148.050 487.050 ;
        RECT 130.950 485.550 148.050 486.450 ;
        RECT 130.950 484.950 133.050 485.550 ;
        RECT 145.950 484.950 148.050 485.550 ;
        RECT 149.700 483.600 150.900 490.950 ;
        RECT 164.100 489.150 165.900 490.950 ;
        RECT 170.700 483.600 171.900 490.950 ;
        RECT 182.550 489.450 183.450 494.550 ;
        RECT 188.100 493.050 189.900 494.850 ;
        RECT 194.250 493.050 196.050 494.850 ;
        RECT 197.700 493.050 198.600 500.400 ;
        RECT 212.100 501.300 213.900 506.400 ;
        RECT 215.100 502.200 216.900 507.000 ;
        RECT 218.100 501.300 219.900 506.400 ;
        RECT 212.100 499.950 219.900 501.300 ;
        RECT 221.100 500.400 222.900 506.400 ;
        RECT 236.700 505.200 237.900 507.000 ;
        RECT 221.100 498.300 222.300 500.400 ;
        RECT 236.100 499.200 237.900 505.200 ;
        RECT 240.600 500.700 242.400 505.200 ;
        RECT 245.700 504.600 246.900 507.000 ;
        RECT 240.300 499.800 242.400 500.700 ;
        RECT 245.100 499.800 246.900 504.600 ;
        RECT 248.100 502.200 249.900 505.200 ;
        RECT 260.100 503.400 261.900 506.400 ;
        RECT 263.100 503.400 264.900 507.000 ;
        RECT 218.700 497.400 222.300 498.300 ;
        RECT 215.100 493.050 216.900 494.850 ;
        RECT 218.700 493.050 219.900 497.400 ;
        RECT 221.100 493.050 222.900 494.850 ;
        RECT 240.300 493.050 241.200 499.800 ;
        RECT 249.000 498.900 249.900 502.200 ;
        RECT 187.950 490.950 190.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 211.950 490.950 214.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 236.100 490.950 238.200 493.050 ;
        RECT 239.100 490.950 241.200 493.050 ;
        RECT 242.700 498.000 249.900 498.900 ;
        RECT 242.700 490.950 243.900 498.000 ;
        RECT 255.000 495.450 259.050 496.050 ;
        RECT 248.100 493.050 249.900 494.850 ;
        RECT 244.800 490.950 246.900 493.050 ;
        RECT 247.800 490.950 249.900 493.050 ;
        RECT 254.550 493.950 259.050 495.450 ;
        RECT 182.550 488.550 186.450 489.450 ;
        RECT 191.250 489.150 193.050 490.950 ;
        RECT 185.550 486.450 186.450 488.550 ;
        RECT 193.950 486.450 196.050 487.050 ;
        RECT 185.550 485.550 196.050 486.450 ;
        RECT 193.950 484.950 196.050 485.550 ;
        RECT 197.700 483.600 198.600 490.950 ;
        RECT 212.100 489.150 213.900 490.950 ;
        RECT 218.700 483.600 219.900 490.950 ;
        RECT 236.400 489.150 238.200 490.950 ;
        RECT 128.100 482.100 130.500 483.600 ;
        RECT 126.000 479.100 127.800 480.900 ;
        RECT 125.700 471.000 127.500 477.600 ;
        RECT 128.700 471.600 130.500 482.100 ;
        RECT 133.800 471.000 135.600 483.600 ;
        RECT 149.100 471.600 150.900 483.600 ;
        RECT 152.100 471.000 153.900 483.600 ;
        RECT 164.400 471.000 166.200 483.600 ;
        RECT 169.500 482.100 171.900 483.600 ;
        RECT 188.100 482.700 195.900 483.600 ;
        RECT 169.500 471.600 171.300 482.100 ;
        RECT 172.200 479.100 174.000 480.900 ;
        RECT 172.500 471.000 174.300 477.600 ;
        RECT 188.100 471.600 189.900 482.700 ;
        RECT 191.100 471.000 192.900 481.800 ;
        RECT 194.100 471.600 195.900 482.700 ;
        RECT 197.100 471.600 198.900 483.600 ;
        RECT 212.400 471.000 214.200 483.600 ;
        RECT 217.500 482.100 219.900 483.600 ;
        RECT 217.500 471.600 219.300 482.100 ;
        RECT 220.200 479.100 222.000 480.900 ;
        RECT 220.500 471.000 222.300 477.600 ;
        RECT 236.100 471.000 237.900 483.600 ;
        RECT 240.300 483.000 241.200 490.950 ;
        RECT 242.100 489.150 243.900 490.950 ;
        RECT 245.100 489.150 246.900 490.950 ;
        RECT 254.550 490.050 255.450 493.950 ;
        RECT 260.700 493.050 261.900 503.400 ;
        RECT 278.100 501.300 279.900 506.400 ;
        RECT 281.100 502.200 282.900 507.000 ;
        RECT 284.100 501.300 285.900 506.400 ;
        RECT 278.100 499.950 285.900 501.300 ;
        RECT 287.100 500.400 288.900 506.400 ;
        RECT 292.950 501.450 295.050 502.050 ;
        RECT 298.950 501.450 301.050 502.050 ;
        RECT 292.950 500.550 301.050 501.450 ;
        RECT 287.100 498.300 288.300 500.400 ;
        RECT 292.950 499.950 295.050 500.550 ;
        RECT 298.950 499.950 301.050 500.550 ;
        RECT 302.100 500.400 303.900 506.400 ;
        RECT 284.700 497.400 288.300 498.300 ;
        RECT 302.700 498.300 303.900 500.400 ;
        RECT 305.100 501.300 306.900 506.400 ;
        RECT 308.100 502.200 309.900 507.000 ;
        RECT 311.100 501.300 312.900 506.400 ;
        RECT 305.100 499.950 312.900 501.300 ;
        RECT 323.700 499.200 325.500 506.400 ;
        RECT 328.800 500.400 330.600 507.000 ;
        RECT 344.100 500.400 345.900 506.400 ;
        RECT 323.700 498.300 327.900 499.200 ;
        RECT 302.700 497.400 306.300 498.300 ;
        RECT 281.100 493.050 282.900 494.850 ;
        RECT 284.700 493.050 285.900 497.400 ;
        RECT 287.100 493.050 288.900 494.850 ;
        RECT 302.100 493.050 303.900 494.850 ;
        RECT 305.100 493.050 306.300 497.400 ;
        RECT 308.100 493.050 309.900 494.850 ;
        RECT 323.100 493.050 324.900 494.850 ;
        RECT 326.700 493.050 327.900 498.300 ;
        RECT 328.950 498.450 331.050 499.050 ;
        RECT 337.950 498.450 340.050 499.050 ;
        RECT 328.950 497.550 340.050 498.450 ;
        RECT 328.950 496.950 331.050 497.550 ;
        RECT 337.950 496.950 340.050 497.550 ;
        RECT 344.700 498.300 345.900 500.400 ;
        RECT 347.100 501.300 348.900 506.400 ;
        RECT 350.100 502.200 351.900 507.000 ;
        RECT 353.100 501.300 354.900 506.400 ;
        RECT 347.100 499.950 354.900 501.300 ;
        RECT 368.100 501.300 369.900 506.400 ;
        RECT 371.100 502.200 372.900 507.000 ;
        RECT 374.100 501.300 375.900 506.400 ;
        RECT 368.100 499.950 375.900 501.300 ;
        RECT 377.100 500.400 378.900 506.400 ;
        RECT 392.400 500.400 394.200 507.000 ;
        RECT 377.100 498.300 378.300 500.400 ;
        RECT 397.500 499.200 399.300 506.400 ;
        RECT 344.700 497.400 348.300 498.300 ;
        RECT 328.950 493.050 330.750 494.850 ;
        RECT 344.100 493.050 345.900 494.850 ;
        RECT 347.100 493.050 348.300 497.400 ;
        RECT 374.700 497.400 378.300 498.300 ;
        RECT 395.100 498.300 399.300 499.200 ;
        RECT 413.100 503.400 414.900 506.400 ;
        RECT 413.100 499.500 414.300 503.400 ;
        RECT 416.100 500.400 417.900 507.000 ;
        RECT 419.100 500.400 420.900 506.400 ;
        RECT 413.100 498.600 418.800 499.500 ;
        RECT 350.100 493.050 351.900 494.850 ;
        RECT 371.100 493.050 372.900 494.850 ;
        RECT 374.700 493.050 375.900 497.400 ;
        RECT 377.100 493.050 378.900 494.850 ;
        RECT 392.250 493.050 394.050 494.850 ;
        RECT 395.100 493.050 396.300 498.300 ;
        RECT 417.000 497.700 418.800 498.600 ;
        RECT 398.100 493.050 399.900 494.850 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 304.950 490.950 307.050 493.050 ;
        RECT 307.950 490.950 310.050 493.050 ;
        RECT 310.950 490.950 313.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 349.950 490.950 352.050 493.050 ;
        RECT 352.950 490.950 355.050 493.050 ;
        RECT 367.950 490.950 370.050 493.050 ;
        RECT 370.950 490.950 373.050 493.050 ;
        RECT 373.950 490.950 376.050 493.050 ;
        RECT 376.950 490.950 379.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 413.400 490.950 415.500 493.050 ;
        RECT 242.100 484.800 243.300 489.150 ;
        RECT 254.550 488.550 259.050 490.050 ;
        RECT 255.000 487.950 259.050 488.550 ;
        RECT 242.100 483.900 249.900 484.800 ;
        RECT 240.300 482.100 242.400 483.000 ;
        RECT 240.600 471.600 242.400 482.100 ;
        RECT 245.100 471.000 246.900 483.000 ;
        RECT 249.000 478.800 249.900 483.900 ;
        RECT 248.100 472.800 249.900 478.800 ;
        RECT 260.700 477.600 261.900 490.950 ;
        RECT 263.100 489.150 264.900 490.950 ;
        RECT 278.100 489.150 279.900 490.950 ;
        RECT 284.700 483.600 285.900 490.950 ;
        RECT 260.100 471.600 261.900 477.600 ;
        RECT 263.100 471.000 264.900 477.600 ;
        RECT 278.400 471.000 280.200 483.600 ;
        RECT 283.500 482.100 285.900 483.600 ;
        RECT 305.100 483.600 306.300 490.950 ;
        RECT 311.100 489.150 312.900 490.950 ;
        RECT 305.100 482.100 307.500 483.600 ;
        RECT 283.500 471.600 285.300 482.100 ;
        RECT 286.200 479.100 288.000 480.900 ;
        RECT 303.000 479.100 304.800 480.900 ;
        RECT 286.500 471.000 288.300 477.600 ;
        RECT 302.700 471.000 304.500 477.600 ;
        RECT 305.700 471.600 307.500 482.100 ;
        RECT 310.800 471.000 312.600 483.600 ;
        RECT 326.700 477.600 327.900 490.950 ;
        RECT 328.950 483.450 331.050 484.050 ;
        RECT 343.950 483.450 346.050 484.050 ;
        RECT 328.950 482.550 346.050 483.450 ;
        RECT 328.950 481.950 331.050 482.550 ;
        RECT 343.950 481.950 346.050 482.550 ;
        RECT 347.100 483.600 348.300 490.950 ;
        RECT 353.100 489.150 354.900 490.950 ;
        RECT 368.100 489.150 369.900 490.950 ;
        RECT 374.700 483.600 375.900 490.950 ;
        RECT 376.950 486.450 379.050 486.750 ;
        RECT 391.950 486.450 394.050 487.050 ;
        RECT 376.950 485.550 394.050 486.450 ;
        RECT 376.950 484.650 379.050 485.550 ;
        RECT 391.950 484.950 394.050 485.550 ;
        RECT 347.100 482.100 349.500 483.600 ;
        RECT 345.000 479.100 346.800 480.900 ;
        RECT 323.100 471.000 324.900 477.600 ;
        RECT 326.100 471.600 327.900 477.600 ;
        RECT 329.100 471.000 330.900 477.600 ;
        RECT 344.700 471.000 346.500 477.600 ;
        RECT 347.700 471.600 349.500 482.100 ;
        RECT 352.800 471.000 354.600 483.600 ;
        RECT 368.400 471.000 370.200 483.600 ;
        RECT 373.500 482.100 375.900 483.600 ;
        RECT 373.500 471.600 375.300 482.100 ;
        RECT 376.200 479.100 378.000 480.900 ;
        RECT 395.100 477.600 396.300 490.950 ;
        RECT 413.400 489.150 415.200 490.950 ;
        RECT 417.000 486.300 417.900 497.700 ;
        RECT 419.700 493.050 420.900 500.400 ;
        RECT 418.800 490.950 420.900 493.050 ;
        RECT 417.000 485.400 418.800 486.300 ;
        RECT 413.100 484.500 418.800 485.400 ;
        RECT 413.100 477.600 414.300 484.500 ;
        RECT 419.700 483.600 420.900 490.950 ;
        RECT 376.500 471.000 378.300 477.600 ;
        RECT 392.100 471.000 393.900 477.600 ;
        RECT 395.100 471.600 396.900 477.600 ;
        RECT 398.100 471.000 399.900 477.600 ;
        RECT 413.100 471.600 414.900 477.600 ;
        RECT 416.100 471.000 417.900 481.800 ;
        RECT 419.100 471.600 420.900 483.600 ;
        RECT 434.100 500.400 435.900 506.400 ;
        RECT 437.100 500.400 438.900 507.000 ;
        RECT 440.100 503.400 441.900 506.400 ;
        RECT 434.100 493.050 435.300 500.400 ;
        RECT 440.700 499.500 441.900 503.400 ;
        RECT 436.200 498.600 441.900 499.500 ;
        RECT 455.100 503.400 456.900 506.400 ;
        RECT 455.100 499.500 456.300 503.400 ;
        RECT 458.100 500.400 459.900 507.000 ;
        RECT 461.100 500.400 462.900 506.400 ;
        RECT 455.100 498.600 460.800 499.500 ;
        RECT 436.200 497.700 438.000 498.600 ;
        RECT 434.100 490.950 436.200 493.050 ;
        RECT 434.100 483.600 435.300 490.950 ;
        RECT 437.100 486.300 438.000 497.700 ;
        RECT 459.000 497.700 460.800 498.600 ;
        RECT 439.500 490.950 441.600 493.050 ;
        RECT 439.800 489.150 441.600 490.950 ;
        RECT 455.400 490.950 457.500 493.050 ;
        RECT 455.400 489.150 457.200 490.950 ;
        RECT 436.200 485.400 438.000 486.300 ;
        RECT 459.000 486.300 459.900 497.700 ;
        RECT 461.700 493.050 462.900 500.400 ;
        RECT 473.100 503.400 474.900 506.400 ;
        RECT 473.100 499.500 474.300 503.400 ;
        RECT 476.100 500.400 477.900 507.000 ;
        RECT 479.100 500.400 480.900 506.400 ;
        RECT 494.100 500.400 495.900 507.000 ;
        RECT 497.100 500.400 498.900 506.400 ;
        RECT 473.100 498.600 478.800 499.500 ;
        RECT 477.000 497.700 478.800 498.600 ;
        RECT 460.800 490.950 462.900 493.050 ;
        RECT 459.000 485.400 460.800 486.300 ;
        RECT 436.200 484.500 441.900 485.400 ;
        RECT 434.100 471.600 435.900 483.600 ;
        RECT 437.100 471.000 438.900 481.800 ;
        RECT 440.700 477.600 441.900 484.500 ;
        RECT 440.100 471.600 441.900 477.600 ;
        RECT 455.100 484.500 460.800 485.400 ;
        RECT 455.100 477.600 456.300 484.500 ;
        RECT 461.700 483.600 462.900 490.950 ;
        RECT 473.400 490.950 475.500 493.050 ;
        RECT 473.400 489.150 475.200 490.950 ;
        RECT 477.000 486.300 477.900 497.700 ;
        RECT 479.700 493.050 480.900 500.400 ;
        RECT 481.950 498.450 484.050 499.050 ;
        RECT 493.950 498.450 496.050 499.050 ;
        RECT 481.950 497.550 496.050 498.450 ;
        RECT 481.950 496.950 484.050 497.550 ;
        RECT 493.950 496.950 496.050 497.550 ;
        RECT 494.100 493.050 495.900 494.850 ;
        RECT 497.100 493.050 498.300 500.400 ;
        RECT 512.700 499.200 514.500 506.400 ;
        RECT 517.800 500.400 519.600 507.000 ;
        RECT 533.700 499.200 535.500 506.400 ;
        RECT 538.800 500.400 540.600 507.000 ;
        RECT 551.700 499.200 553.500 506.400 ;
        RECT 556.800 500.400 558.600 507.000 ;
        RECT 572.100 506.400 573.300 507.000 ;
        RECT 572.100 503.400 573.900 506.400 ;
        RECT 575.100 503.400 576.900 506.400 ;
        RECT 575.400 499.200 576.300 503.400 ;
        RECT 578.100 501.000 579.900 507.000 ;
        RECT 581.100 500.400 582.900 506.400 ;
        RECT 512.700 498.300 516.900 499.200 ;
        RECT 533.700 498.300 537.900 499.200 ;
        RECT 551.700 498.300 555.900 499.200 ;
        RECT 575.400 498.300 580.800 499.200 ;
        RECT 512.100 493.050 513.900 494.850 ;
        RECT 515.700 493.050 516.900 498.300 ;
        RECT 517.950 493.050 519.750 494.850 ;
        RECT 533.100 493.050 534.900 494.850 ;
        RECT 536.700 493.050 537.900 498.300 ;
        RECT 538.950 493.050 540.750 494.850 ;
        RECT 551.100 493.050 552.900 494.850 ;
        RECT 554.700 493.050 555.900 498.300 ;
        RECT 578.700 497.400 580.800 498.300 ;
        RECT 556.950 493.050 558.750 494.850 ;
        RECT 572.400 493.050 574.200 494.850 ;
        RECT 478.800 490.950 480.900 493.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 572.100 490.950 574.200 493.050 ;
        RECT 575.400 490.950 577.500 493.050 ;
        RECT 477.000 485.400 478.800 486.300 ;
        RECT 455.100 471.600 456.900 477.600 ;
        RECT 458.100 471.000 459.900 481.800 ;
        RECT 461.100 471.600 462.900 483.600 ;
        RECT 473.100 484.500 478.800 485.400 ;
        RECT 473.100 477.600 474.300 484.500 ;
        RECT 479.700 483.600 480.900 490.950 ;
        RECT 497.100 483.600 498.300 490.950 ;
        RECT 473.100 471.600 474.900 477.600 ;
        RECT 476.100 471.000 477.900 481.800 ;
        RECT 479.100 471.600 480.900 483.600 ;
        RECT 494.100 471.000 495.900 483.600 ;
        RECT 497.100 471.600 498.900 483.600 ;
        RECT 515.700 477.600 516.900 490.950 ;
        RECT 536.700 477.600 537.900 490.950 ;
        RECT 554.700 477.600 555.900 490.950 ;
        RECT 576.000 489.150 577.800 490.950 ;
        RECT 578.700 486.900 579.600 497.400 ;
        RECT 582.000 493.050 582.900 500.400 ;
        RECT 593.100 501.300 594.900 506.400 ;
        RECT 596.100 502.200 597.900 507.000 ;
        RECT 599.100 501.300 600.900 506.400 ;
        RECT 593.100 499.950 600.900 501.300 ;
        RECT 602.100 500.400 603.900 506.400 ;
        RECT 617.100 500.400 618.900 506.400 ;
        RECT 602.100 498.300 603.300 500.400 ;
        RECT 599.700 497.400 603.300 498.300 ;
        RECT 617.700 498.300 618.900 500.400 ;
        RECT 620.100 501.300 621.900 506.400 ;
        RECT 623.100 502.200 624.900 507.000 ;
        RECT 638.100 506.400 639.300 507.000 ;
        RECT 626.100 501.300 627.900 506.400 ;
        RECT 638.100 503.400 639.900 506.400 ;
        RECT 641.100 503.400 642.900 506.400 ;
        RECT 620.100 499.950 627.900 501.300 ;
        RECT 641.400 499.200 642.300 503.400 ;
        RECT 644.100 501.000 645.900 507.000 ;
        RECT 647.100 500.400 648.900 506.400 ;
        RECT 636.000 498.450 640.050 499.050 ;
        RECT 617.700 497.400 621.300 498.300 ;
        RECT 596.100 493.050 597.900 494.850 ;
        RECT 599.700 493.050 600.900 497.400 ;
        RECT 604.950 495.450 607.050 496.050 ;
        RECT 602.100 493.050 603.900 494.850 ;
        RECT 604.950 494.550 612.450 495.450 ;
        RECT 604.950 493.950 607.050 494.550 ;
        RECT 580.800 490.950 582.900 493.050 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 578.100 486.300 579.900 486.900 ;
        RECT 572.100 485.100 579.900 486.300 ;
        RECT 572.100 483.600 573.300 485.100 ;
        RECT 580.800 483.600 582.000 490.950 ;
        RECT 593.100 489.150 594.900 490.950 ;
        RECT 599.700 483.600 600.900 490.950 ;
        RECT 611.550 490.050 612.450 494.550 ;
        RECT 617.100 493.050 618.900 494.850 ;
        RECT 620.100 493.050 621.300 497.400 ;
        RECT 635.550 496.950 640.050 498.450 ;
        RECT 641.400 498.300 646.800 499.200 ;
        RECT 644.700 497.400 646.800 498.300 ;
        RECT 623.100 493.050 624.900 494.850 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 625.950 490.950 628.050 493.050 ;
        RECT 611.550 488.550 616.050 490.050 ;
        RECT 612.000 487.950 616.050 488.550 ;
        RECT 512.100 471.000 513.900 477.600 ;
        RECT 515.100 471.600 516.900 477.600 ;
        RECT 518.100 471.000 519.900 477.600 ;
        RECT 533.100 471.000 534.900 477.600 ;
        RECT 536.100 471.600 537.900 477.600 ;
        RECT 539.100 471.000 540.900 477.600 ;
        RECT 551.100 471.000 552.900 477.600 ;
        RECT 554.100 471.600 555.900 477.600 ;
        RECT 557.100 471.000 558.900 477.600 ;
        RECT 572.100 471.600 573.900 483.600 ;
        RECT 576.600 471.000 578.400 483.600 ;
        RECT 579.600 482.100 582.000 483.600 ;
        RECT 579.600 471.600 581.400 482.100 ;
        RECT 593.400 471.000 595.200 483.600 ;
        RECT 598.500 482.100 600.900 483.600 ;
        RECT 620.100 483.600 621.300 490.950 ;
        RECT 626.100 489.150 627.900 490.950 ;
        RECT 628.950 489.450 631.050 490.050 ;
        RECT 635.550 489.450 636.450 496.950 ;
        RECT 638.400 493.050 640.200 494.850 ;
        RECT 638.100 490.950 640.200 493.050 ;
        RECT 641.400 490.950 643.500 493.050 ;
        RECT 628.950 488.550 636.450 489.450 ;
        RECT 642.000 489.150 643.800 490.950 ;
        RECT 628.950 487.950 631.050 488.550 ;
        RECT 644.700 486.900 645.600 497.400 ;
        RECT 648.000 493.050 648.900 500.400 ;
        RECT 659.100 498.600 660.900 506.400 ;
        RECT 663.600 500.400 665.400 507.000 ;
        RECT 666.600 502.200 668.400 506.400 ;
        RECT 666.600 500.400 669.300 502.200 ;
        RECT 665.700 498.600 667.500 499.500 ;
        RECT 659.100 497.700 667.500 498.600 ;
        RECT 659.250 493.050 661.050 494.850 ;
        RECT 646.800 490.950 648.900 493.050 ;
        RECT 659.100 490.950 661.200 493.050 ;
        RECT 644.100 486.300 645.900 486.900 ;
        RECT 638.100 485.100 645.900 486.300 ;
        RECT 638.100 483.600 639.300 485.100 ;
        RECT 646.800 483.600 648.000 490.950 ;
        RECT 620.100 482.100 622.500 483.600 ;
        RECT 598.500 471.600 600.300 482.100 ;
        RECT 601.200 479.100 603.000 480.900 ;
        RECT 618.000 479.100 619.800 480.900 ;
        RECT 601.500 471.000 603.300 477.600 ;
        RECT 617.700 471.000 619.500 477.600 ;
        RECT 620.700 471.600 622.500 482.100 ;
        RECT 625.800 471.000 627.600 483.600 ;
        RECT 638.100 471.600 639.900 483.600 ;
        RECT 642.600 471.000 644.400 483.600 ;
        RECT 645.600 482.100 648.000 483.600 ;
        RECT 645.600 471.600 647.400 482.100 ;
        RECT 662.100 477.600 663.000 497.700 ;
        RECT 668.400 493.050 669.300 500.400 ;
        RECT 680.100 501.300 681.900 506.400 ;
        RECT 683.100 502.200 684.900 507.000 ;
        RECT 686.100 501.300 687.900 506.400 ;
        RECT 680.100 499.950 687.900 501.300 ;
        RECT 689.100 500.400 690.900 506.400 ;
        RECT 704.100 503.400 705.900 507.000 ;
        RECT 707.100 503.400 708.900 506.400 ;
        RECT 722.700 503.400 724.500 507.000 ;
        RECT 689.100 498.300 690.300 500.400 ;
        RECT 686.700 497.400 690.300 498.300 ;
        RECT 683.100 493.050 684.900 494.850 ;
        RECT 686.700 493.050 687.900 497.400 ;
        RECT 689.100 493.050 690.900 494.850 ;
        RECT 707.100 493.050 708.300 503.400 ;
        RECT 725.700 501.600 727.500 506.400 ;
        RECT 722.400 500.400 727.500 501.600 ;
        RECT 730.200 500.400 732.000 507.000 ;
        RECT 722.400 493.050 723.300 500.400 ;
        RECT 724.950 498.450 727.050 499.050 ;
        RECT 739.950 498.450 742.050 499.050 ;
        RECT 724.950 497.550 742.050 498.450 ;
        RECT 724.950 496.950 727.050 497.550 ;
        RECT 739.950 496.950 742.050 497.550 ;
        RECT 743.100 497.400 744.900 507.000 ;
        RECT 749.700 498.000 751.500 506.400 ;
        RECT 749.700 496.800 753.000 498.000 ;
        RECT 767.100 497.400 768.900 507.000 ;
        RECT 773.700 498.000 775.500 506.400 ;
        RECT 773.700 496.800 777.000 498.000 ;
        RECT 788.100 497.400 789.900 507.000 ;
        RECT 794.700 498.000 796.500 506.400 ;
        RECT 812.700 499.200 814.500 506.400 ;
        RECT 817.800 500.400 819.600 507.000 ;
        RECT 812.700 498.300 816.900 499.200 ;
        RECT 794.700 496.800 798.000 498.000 ;
        RECT 724.950 493.050 726.750 494.850 ;
        RECT 731.100 493.050 732.900 494.850 ;
        RECT 743.100 493.050 744.900 494.850 ;
        RECT 749.100 493.050 750.900 494.850 ;
        RECT 752.100 493.050 753.000 496.800 ;
        RECT 767.100 493.050 768.900 494.850 ;
        RECT 773.100 493.050 774.900 494.850 ;
        RECT 776.100 493.050 777.000 496.800 ;
        RECT 788.100 493.050 789.900 494.850 ;
        RECT 794.100 493.050 795.900 494.850 ;
        RECT 797.100 493.050 798.000 496.800 ;
        RECT 812.100 493.050 813.900 494.850 ;
        RECT 815.700 493.050 816.900 498.300 ;
        RECT 830.100 497.400 831.900 507.000 ;
        RECT 836.700 498.000 838.500 506.400 ;
        RECT 851.100 503.400 852.900 507.000 ;
        RECT 854.100 503.400 855.900 506.400 ;
        RECT 857.100 503.400 858.900 507.000 ;
        RECT 836.700 496.800 840.000 498.000 ;
        RECT 817.950 493.050 819.750 494.850 ;
        RECT 830.100 493.050 831.900 494.850 ;
        RECT 836.100 493.050 837.900 494.850 ;
        RECT 839.100 493.050 840.000 496.800 ;
        RECT 854.400 493.050 855.300 503.400 ;
        RECT 870.000 500.400 871.800 507.000 ;
        RECT 874.500 501.600 876.300 506.400 ;
        RECT 877.500 503.400 879.300 507.000 ;
        RECT 874.500 500.400 879.600 501.600 ;
        RECT 893.100 500.400 894.900 506.400 ;
        RECT 856.950 498.450 861.000 499.050 ;
        RECT 856.950 496.950 861.450 498.450 ;
        RECT 860.550 495.450 861.450 496.950 ;
        RECT 860.550 494.550 864.450 495.450 ;
        RECT 664.500 490.950 666.600 493.050 ;
        RECT 667.800 490.950 669.900 493.050 ;
        RECT 679.950 490.950 682.050 493.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 745.950 490.950 748.050 493.050 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 829.950 490.950 832.050 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 664.200 489.150 666.000 490.950 ;
        RECT 668.400 483.600 669.300 490.950 ;
        RECT 680.100 489.150 681.900 490.950 ;
        RECT 686.700 483.600 687.900 490.950 ;
        RECT 704.100 489.150 705.900 490.950 ;
        RECT 659.100 471.000 660.900 477.600 ;
        RECT 662.100 471.600 663.900 477.600 ;
        RECT 665.100 471.000 666.900 483.000 ;
        RECT 668.100 471.600 669.900 483.600 ;
        RECT 680.400 471.000 682.200 483.600 ;
        RECT 685.500 482.100 687.900 483.600 ;
        RECT 685.500 471.600 687.300 482.100 ;
        RECT 688.200 479.100 690.000 480.900 ;
        RECT 707.100 477.600 708.300 490.950 ;
        RECT 722.400 483.600 723.300 490.950 ;
        RECT 727.950 489.150 729.750 490.950 ;
        RECT 746.100 489.150 747.900 490.950 ;
        RECT 724.950 486.450 727.050 487.050 ;
        RECT 742.950 486.450 745.050 487.050 ;
        RECT 724.950 485.550 745.050 486.450 ;
        RECT 724.950 484.950 727.050 485.550 ;
        RECT 742.950 484.950 745.050 485.550 ;
        RECT 688.500 471.000 690.300 477.600 ;
        RECT 704.100 471.000 705.900 477.600 ;
        RECT 707.100 471.600 708.900 477.600 ;
        RECT 722.100 471.600 723.900 483.600 ;
        RECT 725.100 482.700 732.900 483.600 ;
        RECT 725.100 471.600 726.900 482.700 ;
        RECT 728.100 471.000 729.900 481.800 ;
        RECT 731.100 471.600 732.900 482.700 ;
        RECT 752.100 478.800 753.000 490.950 ;
        RECT 770.100 489.150 771.900 490.950 ;
        RECT 776.100 478.800 777.000 490.950 ;
        RECT 791.100 489.150 792.900 490.950 ;
        RECT 797.100 478.800 798.000 490.950 ;
        RECT 746.400 477.900 753.000 478.800 ;
        RECT 746.400 477.600 747.900 477.900 ;
        RECT 743.100 471.000 744.900 477.600 ;
        RECT 746.100 471.600 747.900 477.600 ;
        RECT 752.100 477.600 753.000 477.900 ;
        RECT 770.400 477.900 777.000 478.800 ;
        RECT 770.400 477.600 771.900 477.900 ;
        RECT 749.100 471.000 750.900 477.000 ;
        RECT 752.100 471.600 753.900 477.600 ;
        RECT 767.100 471.000 768.900 477.600 ;
        RECT 770.100 471.600 771.900 477.600 ;
        RECT 776.100 477.600 777.000 477.900 ;
        RECT 791.400 477.900 798.000 478.800 ;
        RECT 791.400 477.600 792.900 477.900 ;
        RECT 773.100 471.000 774.900 477.000 ;
        RECT 776.100 471.600 777.900 477.600 ;
        RECT 788.100 471.000 789.900 477.600 ;
        RECT 791.100 471.600 792.900 477.600 ;
        RECT 797.100 477.600 798.000 477.900 ;
        RECT 815.700 477.600 816.900 490.950 ;
        RECT 833.100 489.150 834.900 490.950 ;
        RECT 820.950 486.450 823.050 487.050 ;
        RECT 829.950 486.450 832.050 487.050 ;
        RECT 820.950 485.550 832.050 486.450 ;
        RECT 820.950 484.950 823.050 485.550 ;
        RECT 829.950 484.950 832.050 485.550 ;
        RECT 839.100 478.800 840.000 490.950 ;
        RECT 851.250 489.150 853.050 490.950 ;
        RECT 854.400 483.600 855.300 490.950 ;
        RECT 857.100 489.150 858.900 490.950 ;
        RECT 863.550 490.050 864.450 494.550 ;
        RECT 869.100 493.050 870.900 494.850 ;
        RECT 875.250 493.050 877.050 494.850 ;
        RECT 878.700 493.050 879.600 500.400 ;
        RECT 893.700 498.300 894.900 500.400 ;
        RECT 896.100 501.300 897.900 506.400 ;
        RECT 899.100 502.200 900.900 507.000 ;
        RECT 902.100 501.300 903.900 506.400 ;
        RECT 896.100 499.950 903.900 501.300 ;
        RECT 917.700 499.200 919.500 506.400 ;
        RECT 922.800 500.400 924.600 507.000 ;
        RECT 938.700 499.200 940.500 506.400 ;
        RECT 943.800 500.400 945.600 507.000 ;
        RECT 917.700 498.300 921.900 499.200 ;
        RECT 938.700 498.300 942.900 499.200 ;
        RECT 893.700 497.400 897.300 498.300 ;
        RECT 893.100 493.050 894.900 494.850 ;
        RECT 896.100 493.050 897.300 497.400 ;
        RECT 904.950 495.450 909.000 496.050 ;
        RECT 899.100 493.050 900.900 494.850 ;
        RECT 904.950 493.950 909.450 495.450 ;
        RECT 868.950 490.950 871.050 493.050 ;
        RECT 871.950 490.950 874.050 493.050 ;
        RECT 874.950 490.950 877.050 493.050 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 895.950 490.950 898.050 493.050 ;
        RECT 898.950 490.950 901.050 493.050 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 859.950 488.550 864.450 490.050 ;
        RECT 872.250 489.150 874.050 490.950 ;
        RECT 859.950 487.950 864.000 488.550 ;
        RECT 865.950 486.450 868.050 487.050 ;
        RECT 874.950 486.450 877.050 487.050 ;
        RECT 865.950 485.550 877.050 486.450 ;
        RECT 865.950 484.950 868.050 485.550 ;
        RECT 874.950 484.950 877.050 485.550 ;
        RECT 878.700 483.600 879.600 490.950 ;
        RECT 883.950 489.450 886.050 490.050 ;
        RECT 889.950 489.450 892.050 490.050 ;
        RECT 883.950 488.550 892.050 489.450 ;
        RECT 883.950 487.950 886.050 488.550 ;
        RECT 889.950 487.950 892.050 488.550 ;
        RECT 896.100 483.600 897.300 490.950 ;
        RECT 902.100 489.150 903.900 490.950 ;
        RECT 901.950 486.450 904.050 487.050 ;
        RECT 908.550 486.450 909.450 493.950 ;
        RECT 917.100 493.050 918.900 494.850 ;
        RECT 920.700 493.050 921.900 498.300 ;
        RECT 922.950 493.050 924.750 494.850 ;
        RECT 938.100 493.050 939.900 494.850 ;
        RECT 941.700 493.050 942.900 498.300 ;
        RECT 943.950 493.050 945.750 494.850 ;
        RECT 916.950 490.950 919.050 493.050 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 922.950 490.950 925.050 493.050 ;
        RECT 937.950 490.950 940.050 493.050 ;
        RECT 940.950 490.950 943.050 493.050 ;
        RECT 943.950 490.950 946.050 493.050 ;
        RECT 901.950 485.550 909.450 486.450 ;
        RECT 901.950 484.950 904.050 485.550 ;
        RECT 833.400 477.900 840.000 478.800 ;
        RECT 833.400 477.600 834.900 477.900 ;
        RECT 794.100 471.000 795.900 477.000 ;
        RECT 797.100 471.600 798.900 477.600 ;
        RECT 812.100 471.000 813.900 477.600 ;
        RECT 815.100 471.600 816.900 477.600 ;
        RECT 818.100 471.000 819.900 477.600 ;
        RECT 830.100 471.000 831.900 477.600 ;
        RECT 833.100 471.600 834.900 477.600 ;
        RECT 839.100 477.600 840.000 477.900 ;
        RECT 836.100 471.000 837.900 477.000 ;
        RECT 839.100 471.600 840.900 477.600 ;
        RECT 851.100 471.000 852.900 483.600 ;
        RECT 854.400 482.400 858.000 483.600 ;
        RECT 856.200 471.600 858.000 482.400 ;
        RECT 869.100 482.700 876.900 483.600 ;
        RECT 869.100 471.600 870.900 482.700 ;
        RECT 872.100 471.000 873.900 481.800 ;
        RECT 875.100 471.600 876.900 482.700 ;
        RECT 878.100 471.600 879.900 483.600 ;
        RECT 896.100 482.100 898.500 483.600 ;
        RECT 894.000 479.100 895.800 480.900 ;
        RECT 893.700 471.000 895.500 477.600 ;
        RECT 896.700 471.600 898.500 482.100 ;
        RECT 901.800 471.000 903.600 483.600 ;
        RECT 920.700 477.600 921.900 490.950 ;
        RECT 925.950 489.450 928.050 490.050 ;
        RECT 931.950 489.450 934.050 490.050 ;
        RECT 925.950 488.550 934.050 489.450 ;
        RECT 925.950 487.950 928.050 488.550 ;
        RECT 931.950 487.950 934.050 488.550 ;
        RECT 931.950 486.450 934.050 486.900 ;
        RECT 937.950 486.450 940.050 487.050 ;
        RECT 931.950 485.550 940.050 486.450 ;
        RECT 931.950 484.800 934.050 485.550 ;
        RECT 937.950 484.950 940.050 485.550 ;
        RECT 941.700 477.600 942.900 490.950 ;
        RECT 917.100 471.000 918.900 477.600 ;
        RECT 920.100 471.600 921.900 477.600 ;
        RECT 923.100 471.000 924.900 477.600 ;
        RECT 938.100 471.000 939.900 477.600 ;
        RECT 941.100 471.600 942.900 477.600 ;
        RECT 944.100 471.000 945.900 477.600 ;
        RECT 11.400 455.400 13.200 468.000 ;
        RECT 16.500 456.900 18.300 467.400 ;
        RECT 19.500 461.400 21.300 468.000 ;
        RECT 35.100 461.400 36.900 468.000 ;
        RECT 38.100 461.400 39.900 467.400 ;
        RECT 41.100 461.400 42.900 468.000 ;
        RECT 53.100 461.400 54.900 468.000 ;
        RECT 56.100 461.400 57.900 467.400 ;
        RECT 59.100 461.400 60.900 468.000 ;
        RECT 19.200 458.100 21.000 459.900 ;
        RECT 16.500 455.400 18.900 456.900 ;
        RECT 11.100 448.050 12.900 449.850 ;
        RECT 17.700 448.050 18.900 455.400 ;
        RECT 38.700 448.050 39.900 461.400 ;
        RECT 48.000 450.900 51.000 451.050 ;
        RECT 48.000 450.450 52.050 450.900 ;
        RECT 47.550 448.950 52.050 450.450 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 34.950 445.950 37.050 448.050 ;
        RECT 37.950 445.950 40.050 448.050 ;
        RECT 40.950 445.950 43.050 448.050 ;
        RECT 14.100 444.150 15.900 445.950 ;
        RECT 17.700 441.600 18.900 445.950 ;
        RECT 20.100 444.150 21.900 445.950 ;
        RECT 25.950 444.450 28.050 445.050 ;
        RECT 31.950 444.450 34.050 445.050 ;
        RECT 25.950 443.550 34.050 444.450 ;
        RECT 35.100 444.150 36.900 445.950 ;
        RECT 25.950 442.950 28.050 443.550 ;
        RECT 31.950 442.950 34.050 443.550 ;
        RECT 17.700 440.700 21.300 441.600 ;
        RECT 38.700 440.700 39.900 445.950 ;
        RECT 40.950 444.150 42.750 445.950 ;
        RECT 47.550 445.050 48.450 448.950 ;
        RECT 49.950 448.800 52.050 448.950 ;
        RECT 56.700 448.050 57.900 461.400 ;
        RECT 74.100 455.400 75.900 467.400 ;
        RECT 77.100 456.300 78.900 467.400 ;
        RECT 80.100 457.200 81.900 468.000 ;
        RECT 83.100 456.300 84.900 467.400 ;
        RECT 95.700 461.400 97.500 468.000 ;
        RECT 96.000 458.100 97.800 459.900 ;
        RECT 98.700 456.900 100.500 467.400 ;
        RECT 77.100 455.400 84.900 456.300 ;
        RECT 98.100 455.400 100.500 456.900 ;
        RECT 103.800 455.400 105.600 468.000 ;
        RECT 119.100 456.600 120.900 467.400 ;
        RECT 122.100 457.500 123.900 468.000 ;
        RECT 125.100 466.500 132.900 467.400 ;
        RECT 125.100 456.600 126.900 466.500 ;
        RECT 119.100 455.700 126.900 456.600 ;
        RECT 74.400 448.050 75.300 455.400 ;
        RECT 82.950 453.450 85.050 454.050 ;
        RECT 88.950 453.450 91.050 454.050 ;
        RECT 82.950 452.550 91.050 453.450 ;
        RECT 82.950 451.950 85.050 452.550 ;
        RECT 88.950 451.950 91.050 452.550 ;
        RECT 79.950 448.050 81.750 449.850 ;
        RECT 98.100 448.050 99.300 455.400 ;
        RECT 128.100 454.500 129.900 465.600 ;
        RECT 131.100 455.400 132.900 466.500 ;
        RECT 146.100 461.400 147.900 468.000 ;
        RECT 149.100 461.400 150.900 467.400 ;
        RECT 152.100 461.400 153.900 468.000 ;
        RECT 125.100 453.600 129.900 454.500 ;
        RECT 104.100 448.050 105.900 449.850 ;
        RECT 122.250 448.050 124.050 449.850 ;
        RECT 125.100 448.050 126.000 453.600 ;
        RECT 141.000 450.450 145.050 451.050 ;
        RECT 128.100 448.050 129.900 449.850 ;
        RECT 140.550 448.950 145.050 450.450 ;
        RECT 52.950 445.950 55.050 448.050 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 73.950 445.950 76.050 448.050 ;
        RECT 76.950 445.950 79.050 448.050 ;
        RECT 79.950 445.950 82.050 448.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 94.950 445.950 97.050 448.050 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 118.950 445.950 121.050 448.050 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 127.950 445.950 130.050 448.050 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 47.550 443.550 52.050 445.050 ;
        RECT 53.100 444.150 54.900 445.950 ;
        RECT 48.000 442.950 52.050 443.550 ;
        RECT 56.700 440.700 57.900 445.950 ;
        RECT 58.950 444.150 60.750 445.950 ;
        RECT 11.100 437.700 18.900 439.050 ;
        RECT 11.100 432.600 12.900 437.700 ;
        RECT 14.100 432.000 15.900 436.800 ;
        RECT 17.100 432.600 18.900 437.700 ;
        RECT 20.100 438.600 21.300 440.700 ;
        RECT 35.700 439.800 39.900 440.700 ;
        RECT 53.700 439.800 57.900 440.700 ;
        RECT 20.100 432.600 21.900 438.600 ;
        RECT 35.700 432.600 37.500 439.800 ;
        RECT 40.800 432.000 42.600 438.600 ;
        RECT 53.700 432.600 55.500 439.800 ;
        RECT 74.400 438.600 75.300 445.950 ;
        RECT 76.950 444.150 78.750 445.950 ;
        RECT 83.100 444.150 84.900 445.950 ;
        RECT 95.100 444.150 96.900 445.950 ;
        RECT 98.100 441.600 99.300 445.950 ;
        RECT 101.100 444.150 102.900 445.950 ;
        RECT 119.250 444.150 121.050 445.950 ;
        RECT 95.700 440.700 99.300 441.600 ;
        RECT 95.700 438.600 96.900 440.700 ;
        RECT 58.800 432.000 60.600 438.600 ;
        RECT 74.400 437.400 79.500 438.600 ;
        RECT 74.700 432.000 76.500 435.600 ;
        RECT 77.700 432.600 79.500 437.400 ;
        RECT 82.200 432.000 84.000 438.600 ;
        RECT 95.100 432.600 96.900 438.600 ;
        RECT 98.100 437.700 105.900 439.050 ;
        RECT 125.100 438.600 126.300 445.950 ;
        RECT 131.100 444.150 132.900 445.950 ;
        RECT 133.950 444.450 136.050 445.050 ;
        RECT 140.550 444.450 141.450 448.950 ;
        RECT 149.100 448.050 150.300 461.400 ;
        RECT 167.100 455.400 168.900 468.000 ;
        RECT 170.100 455.400 171.900 467.400 ;
        RECT 185.100 461.400 186.900 468.000 ;
        RECT 188.100 461.400 189.900 467.400 ;
        RECT 170.100 448.050 171.300 455.400 ;
        RECT 185.100 448.050 186.900 449.850 ;
        RECT 188.100 448.050 189.300 461.400 ;
        RECT 203.100 456.600 204.900 467.400 ;
        RECT 206.100 457.500 207.900 468.000 ;
        RECT 209.100 466.500 216.900 467.400 ;
        RECT 209.100 456.600 210.900 466.500 ;
        RECT 203.100 455.700 210.900 456.600 ;
        RECT 212.100 454.500 213.900 465.600 ;
        RECT 215.100 455.400 216.900 466.500 ;
        RECT 227.100 461.400 228.900 467.400 ;
        RECT 230.100 462.000 231.900 468.000 ;
        RECT 228.000 461.100 228.900 461.400 ;
        RECT 233.100 461.400 234.900 467.400 ;
        RECT 236.100 461.400 237.900 468.000 ;
        RECT 233.100 461.100 234.600 461.400 ;
        RECT 228.000 460.200 234.600 461.100 ;
        RECT 209.100 453.600 213.900 454.500 ;
        RECT 206.250 448.050 208.050 449.850 ;
        RECT 209.100 448.050 210.000 453.600 ;
        RECT 212.100 448.050 213.900 449.850 ;
        RECT 228.000 448.050 228.900 460.200 ;
        RECT 251.400 455.400 253.200 468.000 ;
        RECT 256.500 456.900 258.300 467.400 ;
        RECT 259.500 461.400 261.300 468.000 ;
        RECT 275.100 461.400 276.900 468.000 ;
        RECT 278.100 461.400 279.900 467.400 ;
        RECT 281.100 461.400 282.900 468.000 ;
        RECT 296.100 461.400 297.900 468.000 ;
        RECT 299.100 461.400 300.900 467.400 ;
        RECT 259.200 458.100 261.000 459.900 ;
        RECT 256.500 455.400 258.900 456.900 ;
        RECT 253.950 453.450 256.050 454.050 ;
        RECT 248.550 452.550 256.050 453.450 ;
        RECT 238.950 450.450 243.000 451.050 ;
        RECT 248.550 450.450 249.450 452.550 ;
        RECT 253.950 451.950 256.050 452.550 ;
        RECT 233.100 448.050 234.900 449.850 ;
        RECT 238.950 448.950 243.450 450.450 ;
        RECT 145.950 445.950 148.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 205.950 445.950 208.050 448.050 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 211.950 445.950 214.050 448.050 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 226.950 445.950 229.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 232.950 445.950 235.050 448.050 ;
        RECT 235.950 445.950 238.050 448.050 ;
        RECT 133.950 443.550 141.450 444.450 ;
        RECT 146.250 444.150 148.050 445.950 ;
        RECT 133.950 442.950 136.050 443.550 ;
        RECT 149.100 440.700 150.300 445.950 ;
        RECT 152.100 444.150 153.900 445.950 ;
        RECT 167.100 444.150 168.900 445.950 ;
        RECT 149.100 439.800 153.300 440.700 ;
        RECT 98.100 432.600 99.900 437.700 ;
        RECT 101.100 432.000 102.900 436.800 ;
        RECT 104.100 432.600 105.900 437.700 ;
        RECT 119.700 432.000 121.500 438.600 ;
        RECT 124.200 432.600 126.000 438.600 ;
        RECT 128.700 432.000 130.500 438.600 ;
        RECT 146.400 432.000 148.200 438.600 ;
        RECT 151.500 432.600 153.300 439.800 ;
        RECT 170.100 438.600 171.300 445.950 ;
        RECT 167.100 432.000 168.900 438.600 ;
        RECT 170.100 432.600 171.900 438.600 ;
        RECT 188.100 435.600 189.300 445.950 ;
        RECT 203.250 444.150 205.050 445.950 ;
        RECT 209.100 438.600 210.300 445.950 ;
        RECT 215.100 444.150 216.900 445.950 ;
        RECT 228.000 442.200 228.900 445.950 ;
        RECT 230.100 444.150 231.900 445.950 ;
        RECT 236.100 444.150 237.900 445.950 ;
        RECT 242.550 444.450 243.450 448.950 ;
        RECT 239.550 444.000 243.450 444.450 ;
        RECT 238.950 443.550 243.450 444.000 ;
        RECT 245.550 449.550 249.450 450.450 ;
        RECT 245.550 445.050 246.450 449.550 ;
        RECT 251.100 448.050 252.900 449.850 ;
        RECT 257.700 448.050 258.900 455.400 ;
        RECT 278.100 448.050 279.300 461.400 ;
        RECT 280.950 453.450 283.050 454.050 ;
        RECT 289.950 453.450 292.050 454.050 ;
        RECT 280.950 452.550 292.050 453.450 ;
        RECT 280.950 451.950 283.050 452.550 ;
        RECT 289.950 451.950 292.050 452.550 ;
        RECT 250.950 445.950 253.050 448.050 ;
        RECT 253.950 445.950 256.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 296.100 445.950 298.200 448.050 ;
        RECT 245.550 443.550 250.050 445.050 ;
        RECT 254.100 444.150 255.900 445.950 ;
        RECT 228.000 441.000 231.300 442.200 ;
        RECT 185.100 432.000 186.900 435.600 ;
        RECT 188.100 432.600 189.900 435.600 ;
        RECT 203.700 432.000 205.500 438.600 ;
        RECT 208.200 432.600 210.000 438.600 ;
        RECT 212.700 432.000 214.500 438.600 ;
        RECT 229.500 432.600 231.300 441.000 ;
        RECT 236.100 432.000 237.900 441.600 ;
        RECT 238.950 439.950 241.050 443.550 ;
        RECT 246.000 442.950 250.050 443.550 ;
        RECT 257.700 441.600 258.900 445.950 ;
        RECT 260.100 444.150 261.900 445.950 ;
        RECT 275.250 444.150 277.050 445.950 ;
        RECT 257.700 440.700 261.300 441.600 ;
        RECT 251.100 437.700 258.900 439.050 ;
        RECT 251.100 432.600 252.900 437.700 ;
        RECT 254.100 432.000 255.900 436.800 ;
        RECT 257.100 432.600 258.900 437.700 ;
        RECT 260.100 438.600 261.300 440.700 ;
        RECT 278.100 440.700 279.300 445.950 ;
        RECT 281.100 444.150 282.900 445.950 ;
        RECT 296.250 444.150 298.050 445.950 ;
        RECT 299.100 441.300 300.000 461.400 ;
        RECT 302.100 456.000 303.900 468.000 ;
        RECT 305.100 455.400 306.900 467.400 ;
        RECT 320.400 455.400 322.200 468.000 ;
        RECT 325.500 456.900 327.300 467.400 ;
        RECT 328.500 461.400 330.300 468.000 ;
        RECT 328.200 458.100 330.000 459.900 ;
        RECT 325.500 455.400 327.900 456.900 ;
        RECT 301.200 448.050 303.000 449.850 ;
        RECT 305.400 448.050 306.300 455.400 ;
        RECT 320.100 448.050 321.900 449.850 ;
        RECT 326.700 448.050 327.900 455.400 ;
        RECT 344.100 455.400 345.900 467.400 ;
        RECT 347.100 457.200 348.900 468.000 ;
        RECT 350.100 461.400 351.900 467.400 ;
        RECT 344.100 448.050 345.300 455.400 ;
        RECT 350.700 454.500 351.900 461.400 ;
        RECT 346.200 453.600 351.900 454.500 ;
        RECT 362.100 461.400 363.900 467.400 ;
        RECT 362.100 454.500 363.300 461.400 ;
        RECT 365.100 457.200 366.900 468.000 ;
        RECT 368.100 455.400 369.900 467.400 ;
        RECT 383.100 455.400 384.900 467.400 ;
        RECT 386.100 455.400 387.900 468.000 ;
        RECT 398.100 461.400 399.900 468.000 ;
        RECT 401.100 461.400 402.900 467.400 ;
        RECT 404.100 461.400 405.900 468.000 ;
        RECT 362.100 453.600 367.800 454.500 ;
        RECT 346.200 452.700 348.000 453.600 ;
        RECT 301.500 445.950 303.600 448.050 ;
        RECT 304.800 445.950 306.900 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 344.100 445.950 346.200 448.050 ;
        RECT 278.100 439.800 282.300 440.700 ;
        RECT 260.100 432.600 261.900 438.600 ;
        RECT 275.400 432.000 277.200 438.600 ;
        RECT 280.500 432.600 282.300 439.800 ;
        RECT 296.100 440.400 304.500 441.300 ;
        RECT 296.100 432.600 297.900 440.400 ;
        RECT 302.700 439.500 304.500 440.400 ;
        RECT 305.400 438.600 306.300 445.950 ;
        RECT 323.100 444.150 324.900 445.950 ;
        RECT 326.700 441.600 327.900 445.950 ;
        RECT 329.100 444.150 330.900 445.950 ;
        RECT 326.700 440.700 330.300 441.600 ;
        RECT 300.600 432.000 302.400 438.600 ;
        RECT 303.600 436.800 306.300 438.600 ;
        RECT 320.100 437.700 327.900 439.050 ;
        RECT 303.600 432.600 305.400 436.800 ;
        RECT 320.100 432.600 321.900 437.700 ;
        RECT 323.100 432.000 324.900 436.800 ;
        RECT 326.100 432.600 327.900 437.700 ;
        RECT 329.100 438.600 330.300 440.700 ;
        RECT 344.100 438.600 345.300 445.950 ;
        RECT 347.100 441.300 348.000 452.700 ;
        RECT 366.000 452.700 367.800 453.600 ;
        RECT 349.800 448.050 351.600 449.850 ;
        RECT 349.500 445.950 351.600 448.050 ;
        RECT 362.400 448.050 364.200 449.850 ;
        RECT 362.400 445.950 364.500 448.050 ;
        RECT 346.200 440.400 348.000 441.300 ;
        RECT 366.000 441.300 366.900 452.700 ;
        RECT 368.700 448.050 369.900 455.400 ;
        RECT 383.700 448.050 384.900 455.400 ;
        RECT 401.700 448.050 402.900 461.400 ;
        RECT 416.100 456.600 417.900 467.400 ;
        RECT 419.100 457.500 420.900 468.000 ;
        RECT 422.100 466.500 429.900 467.400 ;
        RECT 422.100 456.600 423.900 466.500 ;
        RECT 416.100 455.700 423.900 456.600 ;
        RECT 425.100 454.500 426.900 465.600 ;
        RECT 428.100 455.400 429.900 466.500 ;
        RECT 443.100 461.400 444.900 468.000 ;
        RECT 446.100 461.400 447.900 467.400 ;
        RECT 409.950 453.450 412.050 454.050 ;
        RECT 415.950 453.450 418.050 454.050 ;
        RECT 409.950 452.550 418.050 453.450 ;
        RECT 409.950 451.950 412.050 452.550 ;
        RECT 415.950 451.950 418.050 452.550 ;
        RECT 422.100 453.600 426.900 454.500 ;
        RECT 419.250 448.050 421.050 449.850 ;
        RECT 422.100 448.050 423.000 453.600 ;
        RECT 439.950 450.450 442.050 454.050 ;
        RECT 437.550 450.000 442.050 450.450 ;
        RECT 425.100 448.050 426.900 449.850 ;
        RECT 437.550 449.550 441.450 450.000 ;
        RECT 367.800 445.950 369.900 448.050 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 400.950 445.950 403.050 448.050 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 424.950 445.950 427.050 448.050 ;
        RECT 427.950 445.950 430.050 448.050 ;
        RECT 366.000 440.400 367.800 441.300 ;
        RECT 346.200 439.500 351.900 440.400 ;
        RECT 329.100 432.600 330.900 438.600 ;
        RECT 344.100 432.600 345.900 438.600 ;
        RECT 347.100 432.000 348.900 438.600 ;
        RECT 350.700 435.600 351.900 439.500 ;
        RECT 350.100 432.600 351.900 435.600 ;
        RECT 362.100 439.500 367.800 440.400 ;
        RECT 362.100 435.600 363.300 439.500 ;
        RECT 368.700 438.600 369.900 445.950 ;
        RECT 383.700 438.600 384.900 445.950 ;
        RECT 386.100 444.150 387.900 445.950 ;
        RECT 398.100 444.150 399.900 445.950 ;
        RECT 401.700 440.700 402.900 445.950 ;
        RECT 403.950 444.150 405.750 445.950 ;
        RECT 416.250 444.150 418.050 445.950 ;
        RECT 398.700 439.800 402.900 440.700 ;
        RECT 362.100 432.600 363.900 435.600 ;
        RECT 365.100 432.000 366.900 438.600 ;
        RECT 368.100 432.600 369.900 438.600 ;
        RECT 383.100 432.600 384.900 438.600 ;
        RECT 386.100 432.000 387.900 438.600 ;
        RECT 398.700 432.600 400.500 439.800 ;
        RECT 422.100 438.600 423.300 445.950 ;
        RECT 428.100 444.150 429.900 445.950 ;
        RECT 437.550 445.050 438.450 449.550 ;
        RECT 443.100 448.050 444.900 449.850 ;
        RECT 446.100 448.050 447.300 461.400 ;
        RECT 461.100 455.400 462.900 467.400 ;
        RECT 464.100 456.000 465.900 468.000 ;
        RECT 467.100 461.400 468.900 467.400 ;
        RECT 470.100 461.400 471.900 468.000 ;
        RECT 485.100 461.400 486.900 468.000 ;
        RECT 488.100 461.400 489.900 467.400 ;
        RECT 491.100 461.400 492.900 468.000 ;
        RECT 461.700 448.050 462.600 455.400 ;
        RECT 465.000 448.050 466.800 449.850 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 461.100 445.950 463.200 448.050 ;
        RECT 464.400 445.950 466.500 448.050 ;
        RECT 437.550 443.550 442.050 445.050 ;
        RECT 438.000 442.950 442.050 443.550 ;
        RECT 403.800 432.000 405.600 438.600 ;
        RECT 416.700 432.000 418.500 438.600 ;
        RECT 421.200 432.600 423.000 438.600 ;
        RECT 425.700 432.000 427.500 438.600 ;
        RECT 446.100 435.600 447.300 445.950 ;
        RECT 461.700 438.600 462.600 445.950 ;
        RECT 468.000 441.300 468.900 461.400 ;
        RECT 480.000 450.450 484.050 451.050 ;
        RECT 479.550 448.950 484.050 450.450 ;
        RECT 469.800 445.950 471.900 448.050 ;
        RECT 469.950 444.150 471.750 445.950 ;
        RECT 472.950 444.450 475.050 444.900 ;
        RECT 479.550 444.450 480.450 448.950 ;
        RECT 488.100 448.050 489.300 461.400 ;
        RECT 503.100 455.400 504.900 467.400 ;
        RECT 506.100 456.300 507.900 467.400 ;
        RECT 509.100 457.200 510.900 468.000 ;
        RECT 512.100 456.300 513.900 467.400 ;
        RECT 524.100 461.400 525.900 468.000 ;
        RECT 527.100 461.400 528.900 467.400 ;
        RECT 530.100 462.000 531.900 468.000 ;
        RECT 527.400 461.100 528.900 461.400 ;
        RECT 533.100 461.400 534.900 467.400 ;
        RECT 548.700 461.400 550.500 468.000 ;
        RECT 533.100 461.100 534.000 461.400 ;
        RECT 527.400 460.200 534.000 461.100 ;
        RECT 506.100 455.400 513.900 456.300 ;
        RECT 503.400 448.050 504.300 455.400 ;
        RECT 508.950 448.050 510.750 449.850 ;
        RECT 527.100 448.050 528.900 449.850 ;
        RECT 533.100 448.050 534.000 460.200 ;
        RECT 549.000 458.100 550.800 459.900 ;
        RECT 551.700 456.900 553.500 467.400 ;
        RECT 551.100 455.400 553.500 456.900 ;
        RECT 556.800 455.400 558.600 468.000 ;
        RECT 572.100 466.500 579.900 467.400 ;
        RECT 572.100 455.400 573.900 466.500 ;
        RECT 551.100 448.050 552.300 455.400 ;
        RECT 575.100 454.500 576.900 465.600 ;
        RECT 578.100 456.600 579.900 466.500 ;
        RECT 581.100 457.500 582.900 468.000 ;
        RECT 584.100 456.600 585.900 467.400 ;
        RECT 596.100 461.400 597.900 468.000 ;
        RECT 599.100 461.400 600.900 467.400 ;
        RECT 602.100 461.400 603.900 468.000 ;
        RECT 578.100 455.700 585.900 456.600 ;
        RECT 575.100 453.600 579.900 454.500 ;
        RECT 557.100 448.050 558.900 449.850 ;
        RECT 575.100 448.050 576.900 449.850 ;
        RECT 579.000 448.050 579.900 453.600 ;
        RECT 586.950 450.450 591.000 451.050 ;
        RECT 580.950 448.050 582.750 449.850 ;
        RECT 586.950 448.950 591.450 450.450 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 556.950 445.950 559.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 577.950 445.950 580.050 448.050 ;
        RECT 580.950 445.950 583.050 448.050 ;
        RECT 583.950 445.950 586.050 448.050 ;
        RECT 472.950 443.550 480.450 444.450 ;
        RECT 485.250 444.150 487.050 445.950 ;
        RECT 472.950 442.800 475.050 443.550 ;
        RECT 463.500 440.400 471.900 441.300 ;
        RECT 463.500 439.500 465.300 440.400 ;
        RECT 461.700 436.800 464.400 438.600 ;
        RECT 443.100 432.000 444.900 435.600 ;
        RECT 446.100 432.600 447.900 435.600 ;
        RECT 462.600 432.600 464.400 436.800 ;
        RECT 465.600 432.000 467.400 438.600 ;
        RECT 470.100 432.600 471.900 440.400 ;
        RECT 488.100 440.700 489.300 445.950 ;
        RECT 491.100 444.150 492.900 445.950 ;
        RECT 488.100 439.800 492.300 440.700 ;
        RECT 485.400 432.000 487.200 438.600 ;
        RECT 490.500 432.600 492.300 439.800 ;
        RECT 503.400 438.600 504.300 445.950 ;
        RECT 505.950 444.150 507.750 445.950 ;
        RECT 512.100 444.150 513.900 445.950 ;
        RECT 524.100 444.150 525.900 445.950 ;
        RECT 530.100 444.150 531.900 445.950 ;
        RECT 533.100 442.200 534.000 445.950 ;
        RECT 548.100 444.150 549.900 445.950 ;
        RECT 503.400 437.400 508.500 438.600 ;
        RECT 503.700 432.000 505.500 435.600 ;
        RECT 506.700 432.600 508.500 437.400 ;
        RECT 511.200 432.000 513.000 438.600 ;
        RECT 524.100 432.000 525.900 441.600 ;
        RECT 530.700 441.000 534.000 442.200 ;
        RECT 551.100 441.600 552.300 445.950 ;
        RECT 554.100 444.150 555.900 445.950 ;
        RECT 572.100 444.150 573.900 445.950 ;
        RECT 530.700 432.600 532.500 441.000 ;
        RECT 548.700 440.700 552.300 441.600 ;
        RECT 548.700 438.600 549.900 440.700 ;
        RECT 548.100 432.600 549.900 438.600 ;
        RECT 551.100 437.700 558.900 439.050 ;
        RECT 578.700 438.600 579.900 445.950 ;
        RECT 583.950 444.150 585.750 445.950 ;
        RECT 590.550 445.050 591.450 448.950 ;
        RECT 599.100 448.050 600.300 461.400 ;
        RECT 617.100 455.400 618.900 468.000 ;
        RECT 621.600 455.400 624.900 467.400 ;
        RECT 627.600 455.400 629.400 468.000 ;
        RECT 644.400 455.400 646.200 468.000 ;
        RECT 649.500 456.900 651.300 467.400 ;
        RECT 652.500 461.400 654.300 468.000 ;
        RECT 665.100 461.400 666.900 468.000 ;
        RECT 668.100 461.400 669.900 467.400 ;
        RECT 652.200 458.100 654.000 459.900 ;
        RECT 649.500 455.400 651.900 456.900 ;
        RECT 617.100 448.050 618.900 449.850 ;
        RECT 622.950 448.050 624.000 455.400 ;
        RECT 628.950 448.050 630.750 449.850 ;
        RECT 644.100 448.050 645.900 449.850 ;
        RECT 650.700 448.050 651.900 455.400 ;
        RECT 665.100 448.050 666.900 449.850 ;
        RECT 668.100 448.050 669.300 461.400 ;
        RECT 680.100 455.400 681.900 468.000 ;
        RECT 685.200 456.600 687.000 467.400 ;
        RECT 683.400 455.400 687.000 456.600 ;
        RECT 698.100 455.400 699.900 468.000 ;
        RECT 703.200 456.600 705.000 467.400 ;
        RECT 719.100 461.400 720.900 468.000 ;
        RECT 722.100 461.400 723.900 467.400 ;
        RECT 725.100 461.400 726.900 468.000 ;
        RECT 740.100 461.400 741.900 468.000 ;
        RECT 743.100 461.400 744.900 467.400 ;
        RECT 746.100 462.000 747.900 468.000 ;
        RECT 701.400 455.400 705.000 456.600 ;
        RECT 680.250 448.050 682.050 449.850 ;
        RECT 683.400 448.050 684.300 455.400 ;
        RECT 686.100 448.050 687.900 449.850 ;
        RECT 698.250 448.050 700.050 449.850 ;
        RECT 701.400 448.050 702.300 455.400 ;
        RECT 704.100 448.050 705.900 449.850 ;
        RECT 722.100 448.050 723.300 461.400 ;
        RECT 743.400 461.100 744.900 461.400 ;
        RECT 749.100 461.400 750.900 467.400 ;
        RECT 764.100 461.400 765.900 468.000 ;
        RECT 767.100 461.400 768.900 467.400 ;
        RECT 749.100 461.100 750.000 461.400 ;
        RECT 743.400 460.200 750.000 461.100 ;
        RECT 727.950 450.450 732.000 451.050 ;
        RECT 727.950 448.950 732.450 450.450 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 598.950 445.950 601.050 448.050 ;
        RECT 601.950 445.950 604.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 586.950 443.550 591.450 445.050 ;
        RECT 596.250 444.150 598.050 445.950 ;
        RECT 586.950 442.950 591.000 443.550 ;
        RECT 599.100 440.700 600.300 445.950 ;
        RECT 602.100 444.150 603.900 445.950 ;
        RECT 620.250 444.150 622.050 445.950 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 697.950 445.950 700.050 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 622.950 441.300 624.000 445.950 ;
        RECT 625.950 444.150 627.750 445.950 ;
        RECT 647.100 444.150 648.900 445.950 ;
        RECT 628.950 441.450 631.050 441.750 ;
        RECT 637.950 441.450 640.050 442.050 ;
        RECT 599.100 439.800 603.300 440.700 ;
        RECT 622.950 440.100 627.300 441.300 ;
        RECT 551.100 432.600 552.900 437.700 ;
        RECT 554.100 432.000 555.900 436.800 ;
        RECT 557.100 432.600 558.900 437.700 ;
        RECT 574.500 432.000 576.300 438.600 ;
        RECT 579.000 432.600 580.800 438.600 ;
        RECT 583.500 432.000 585.300 438.600 ;
        RECT 596.400 432.000 598.200 438.600 ;
        RECT 601.500 432.600 603.300 439.800 ;
        RECT 617.100 438.000 624.900 438.900 ;
        RECT 626.400 438.600 627.300 440.100 ;
        RECT 628.950 440.550 640.050 441.450 ;
        RECT 650.700 441.600 651.900 445.950 ;
        RECT 653.100 444.150 654.900 445.950 ;
        RECT 650.700 440.700 654.300 441.600 ;
        RECT 628.950 439.650 631.050 440.550 ;
        RECT 637.950 439.950 640.050 440.550 ;
        RECT 617.100 432.600 618.900 438.000 ;
        RECT 620.100 432.000 621.900 437.100 ;
        RECT 623.100 433.500 624.900 438.000 ;
        RECT 626.100 434.400 627.900 438.600 ;
        RECT 629.100 433.500 630.900 438.600 ;
        RECT 623.100 432.600 630.900 433.500 ;
        RECT 644.100 437.700 651.900 439.050 ;
        RECT 644.100 432.600 645.900 437.700 ;
        RECT 647.100 432.000 648.900 436.800 ;
        RECT 650.100 432.600 651.900 437.700 ;
        RECT 653.100 438.600 654.300 440.700 ;
        RECT 653.100 432.600 654.900 438.600 ;
        RECT 668.100 435.600 669.300 445.950 ;
        RECT 683.400 435.600 684.300 445.950 ;
        RECT 701.400 435.600 702.300 445.950 ;
        RECT 719.250 444.150 721.050 445.950 ;
        RECT 722.100 440.700 723.300 445.950 ;
        RECT 725.100 444.150 726.900 445.950 ;
        RECT 731.550 445.050 732.450 448.950 ;
        RECT 743.100 448.050 744.900 449.850 ;
        RECT 749.100 448.050 750.000 460.200 ;
        RECT 759.000 450.450 763.050 451.050 ;
        RECT 758.550 448.950 763.050 450.450 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 727.950 443.550 732.450 445.050 ;
        RECT 740.100 444.150 741.900 445.950 ;
        RECT 746.100 444.150 747.900 445.950 ;
        RECT 727.950 442.950 732.000 443.550 ;
        RECT 749.100 442.200 750.000 445.950 ;
        RECT 758.550 445.050 759.450 448.950 ;
        RECT 764.100 448.050 765.900 449.850 ;
        RECT 767.100 448.050 768.300 461.400 ;
        RECT 782.400 455.400 784.200 468.000 ;
        RECT 787.500 456.900 789.300 467.400 ;
        RECT 790.500 461.400 792.300 468.000 ;
        RECT 806.100 461.400 807.900 468.000 ;
        RECT 809.100 461.400 810.900 467.400 ;
        RECT 812.100 462.000 813.900 468.000 ;
        RECT 809.400 461.100 810.900 461.400 ;
        RECT 815.100 461.400 816.900 467.400 ;
        RECT 827.100 461.400 828.900 468.000 ;
        RECT 830.100 461.400 831.900 467.400 ;
        RECT 833.100 462.000 834.900 468.000 ;
        RECT 815.100 461.100 816.000 461.400 ;
        RECT 809.400 460.200 816.000 461.100 ;
        RECT 830.400 461.100 831.900 461.400 ;
        RECT 836.100 461.400 837.900 467.400 ;
        RECT 836.100 461.100 837.000 461.400 ;
        RECT 830.400 460.200 837.000 461.100 ;
        RECT 790.200 458.100 792.000 459.900 ;
        RECT 787.500 455.400 789.900 456.900 ;
        RECT 777.000 450.450 781.050 451.050 ;
        RECT 776.550 448.950 781.050 450.450 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 766.950 445.950 769.050 448.050 ;
        RECT 758.550 443.550 763.050 445.050 ;
        RECT 759.000 442.950 763.050 443.550 ;
        RECT 722.100 439.800 726.300 440.700 ;
        RECT 665.100 432.000 666.900 435.600 ;
        RECT 668.100 432.600 669.900 435.600 ;
        RECT 680.100 432.000 681.900 435.600 ;
        RECT 683.100 432.600 684.900 435.600 ;
        RECT 686.100 432.000 687.900 435.600 ;
        RECT 698.100 432.000 699.900 435.600 ;
        RECT 701.100 432.600 702.900 435.600 ;
        RECT 704.100 432.000 705.900 435.600 ;
        RECT 719.400 432.000 721.200 438.600 ;
        RECT 724.500 432.600 726.300 439.800 ;
        RECT 740.100 432.000 741.900 441.600 ;
        RECT 746.700 441.000 750.000 442.200 ;
        RECT 746.700 432.600 748.500 441.000 ;
        RECT 767.100 435.600 768.300 445.950 ;
        RECT 776.550 445.050 777.450 448.950 ;
        RECT 782.100 448.050 783.900 449.850 ;
        RECT 788.700 448.050 789.900 455.400 ;
        RECT 793.950 456.450 796.050 457.050 ;
        RECT 805.950 456.450 808.050 456.900 ;
        RECT 793.950 455.550 808.050 456.450 ;
        RECT 793.950 454.950 796.050 455.550 ;
        RECT 805.950 454.800 808.050 455.550 ;
        RECT 799.950 453.450 802.050 454.050 ;
        RECT 811.950 453.450 814.050 454.050 ;
        RECT 799.950 452.550 814.050 453.450 ;
        RECT 799.950 451.950 802.050 452.550 ;
        RECT 811.950 451.950 814.050 452.550 ;
        RECT 809.100 448.050 810.900 449.850 ;
        RECT 815.100 448.050 816.000 460.200 ;
        RECT 832.950 453.450 835.050 454.050 ;
        RECT 824.550 452.550 835.050 453.450 ;
        RECT 824.550 450.450 825.450 452.550 ;
        RECT 832.950 451.950 835.050 452.550 ;
        RECT 821.550 449.550 825.450 450.450 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 787.950 445.950 790.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 805.950 445.950 808.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 776.550 443.550 781.050 445.050 ;
        RECT 785.100 444.150 786.900 445.950 ;
        RECT 777.000 442.950 781.050 443.550 ;
        RECT 788.700 441.600 789.900 445.950 ;
        RECT 791.100 444.150 792.900 445.950 ;
        RECT 806.100 444.150 807.900 445.950 ;
        RECT 812.100 444.150 813.900 445.950 ;
        RECT 815.100 442.200 816.000 445.950 ;
        RECT 821.550 445.050 822.450 449.550 ;
        RECT 830.100 448.050 831.900 449.850 ;
        RECT 836.100 448.050 837.000 460.200 ;
        RECT 851.400 455.400 853.200 468.000 ;
        RECT 856.500 456.900 858.300 467.400 ;
        RECT 859.500 461.400 861.300 468.000 ;
        RECT 875.100 461.400 876.900 468.000 ;
        RECT 878.100 461.400 879.900 467.400 ;
        RECT 881.100 462.000 882.900 468.000 ;
        RECT 878.400 461.100 879.900 461.400 ;
        RECT 884.100 461.400 885.900 467.400 ;
        RECT 884.100 461.100 885.000 461.400 ;
        RECT 878.400 460.200 885.000 461.100 ;
        RECT 859.200 458.100 861.000 459.900 ;
        RECT 856.500 455.400 858.900 456.900 ;
        RECT 838.950 450.450 843.000 451.050 ;
        RECT 846.000 450.450 850.050 451.050 ;
        RECT 838.950 448.950 843.450 450.450 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 817.950 443.550 822.450 445.050 ;
        RECT 827.100 444.150 828.900 445.950 ;
        RECT 833.100 444.150 834.900 445.950 ;
        RECT 817.950 442.950 822.000 443.550 ;
        RECT 836.100 442.200 837.000 445.950 ;
        RECT 788.700 440.700 792.300 441.600 ;
        RECT 782.100 437.700 789.900 439.050 ;
        RECT 764.100 432.000 765.900 435.600 ;
        RECT 767.100 432.600 768.900 435.600 ;
        RECT 782.100 432.600 783.900 437.700 ;
        RECT 785.100 432.000 786.900 436.800 ;
        RECT 788.100 432.600 789.900 437.700 ;
        RECT 791.100 438.600 792.300 440.700 ;
        RECT 791.100 432.600 792.900 438.600 ;
        RECT 806.100 432.000 807.900 441.600 ;
        RECT 812.700 441.000 816.000 442.200 ;
        RECT 812.700 432.600 814.500 441.000 ;
        RECT 827.100 432.000 828.900 441.600 ;
        RECT 833.700 441.000 837.000 442.200 ;
        RECT 842.550 442.050 843.450 448.950 ;
        RECT 845.550 448.950 850.050 450.450 ;
        RECT 845.550 445.050 846.450 448.950 ;
        RECT 851.100 448.050 852.900 449.850 ;
        RECT 857.700 448.050 858.900 455.400 ;
        RECT 868.950 453.450 871.050 454.050 ;
        RECT 874.950 453.450 877.050 454.050 ;
        RECT 868.950 452.550 877.050 453.450 ;
        RECT 868.950 451.950 871.050 452.550 ;
        RECT 874.950 451.950 877.050 452.550 ;
        RECT 862.950 450.450 867.000 451.050 ;
        RECT 862.950 448.950 867.450 450.450 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 845.550 443.550 850.050 445.050 ;
        RECT 854.100 444.150 855.900 445.950 ;
        RECT 846.000 442.950 850.050 443.550 ;
        RECT 833.700 432.600 835.500 441.000 ;
        RECT 841.950 439.950 844.050 442.050 ;
        RECT 857.700 441.600 858.900 445.950 ;
        RECT 860.100 444.150 861.900 445.950 ;
        RECT 866.550 444.450 867.450 448.950 ;
        RECT 878.100 448.050 879.900 449.850 ;
        RECT 884.100 448.050 885.000 460.200 ;
        RECT 896.400 455.400 898.200 468.000 ;
        RECT 901.500 456.900 903.300 467.400 ;
        RECT 904.500 461.400 906.300 468.000 ;
        RECT 904.200 458.100 906.000 459.900 ;
        RECT 901.500 455.400 903.900 456.900 ;
        RECT 917.100 455.400 918.900 467.400 ;
        RECT 920.100 456.300 921.900 467.400 ;
        RECT 923.100 457.200 924.900 468.000 ;
        RECT 926.100 456.300 927.900 467.400 ;
        RECT 938.100 461.400 939.900 467.400 ;
        RECT 941.100 461.400 942.900 468.000 ;
        RECT 920.100 455.400 927.900 456.300 ;
        RECT 898.950 453.450 901.050 454.050 ;
        RECT 893.550 452.550 901.050 453.450 ;
        RECT 893.550 450.450 894.450 452.550 ;
        RECT 898.950 451.950 901.050 452.550 ;
        RECT 890.550 449.550 894.450 450.450 ;
        RECT 874.950 445.950 877.050 448.050 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 871.950 444.450 874.050 445.050 ;
        RECT 866.550 443.550 874.050 444.450 ;
        RECT 875.100 444.150 876.900 445.950 ;
        RECT 881.100 444.150 882.900 445.950 ;
        RECT 871.950 442.950 874.050 443.550 ;
        RECT 884.100 442.200 885.000 445.950 ;
        RECT 890.550 445.050 891.450 449.550 ;
        RECT 896.100 448.050 897.900 449.850 ;
        RECT 902.700 448.050 903.900 455.400 ;
        RECT 917.400 448.050 918.300 455.400 ;
        RECT 919.950 453.450 922.050 454.050 ;
        RECT 934.950 453.450 937.050 454.050 ;
        RECT 919.950 452.550 937.050 453.450 ;
        RECT 919.950 451.950 922.050 452.550 ;
        RECT 934.950 451.950 937.050 452.550 ;
        RECT 928.950 450.450 933.000 451.050 ;
        RECT 922.950 448.050 924.750 449.850 ;
        RECT 928.950 448.950 933.450 450.450 ;
        RECT 895.950 445.950 898.050 448.050 ;
        RECT 898.950 445.950 901.050 448.050 ;
        RECT 901.950 445.950 904.050 448.050 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 916.950 445.950 919.050 448.050 ;
        RECT 919.950 445.950 922.050 448.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 925.950 445.950 928.050 448.050 ;
        RECT 890.550 443.550 895.050 445.050 ;
        RECT 899.100 444.150 900.900 445.950 ;
        RECT 891.000 442.950 895.050 443.550 ;
        RECT 857.700 440.700 861.300 441.600 ;
        RECT 851.100 437.700 858.900 439.050 ;
        RECT 851.100 432.600 852.900 437.700 ;
        RECT 854.100 432.000 855.900 436.800 ;
        RECT 857.100 432.600 858.900 437.700 ;
        RECT 860.100 438.600 861.300 440.700 ;
        RECT 860.100 432.600 861.900 438.600 ;
        RECT 875.100 432.000 876.900 441.600 ;
        RECT 881.700 441.000 885.000 442.200 ;
        RECT 902.700 441.600 903.900 445.950 ;
        RECT 905.100 444.150 906.900 445.950 ;
        RECT 881.700 432.600 883.500 441.000 ;
        RECT 902.700 440.700 906.300 441.600 ;
        RECT 896.100 437.700 903.900 439.050 ;
        RECT 896.100 432.600 897.900 437.700 ;
        RECT 899.100 432.000 900.900 436.800 ;
        RECT 902.100 432.600 903.900 437.700 ;
        RECT 905.100 438.600 906.300 440.700 ;
        RECT 917.400 438.600 918.300 445.950 ;
        RECT 919.950 444.150 921.750 445.950 ;
        RECT 926.100 444.150 927.900 445.950 ;
        RECT 932.550 442.050 933.450 448.950 ;
        RECT 938.700 448.050 939.900 461.400 ;
        RECT 941.100 448.050 942.900 449.850 ;
        RECT 937.950 445.950 940.050 448.050 ;
        RECT 940.950 445.950 943.050 448.050 ;
        RECT 931.950 439.950 934.050 442.050 ;
        RECT 905.100 432.600 906.900 438.600 ;
        RECT 917.400 437.400 922.500 438.600 ;
        RECT 917.700 432.000 919.500 435.600 ;
        RECT 920.700 432.600 922.500 437.400 ;
        RECT 925.200 432.000 927.000 438.600 ;
        RECT 938.700 435.600 939.900 445.950 ;
        RECT 938.100 432.600 939.900 435.600 ;
        RECT 941.100 432.000 942.900 435.600 ;
        RECT 14.100 424.200 15.900 427.200 ;
        RECT 17.100 426.600 18.300 429.000 ;
        RECT 26.100 427.200 27.300 429.000 ;
        RECT 14.100 420.900 15.000 424.200 ;
        RECT 17.100 421.800 18.900 426.600 ;
        RECT 21.600 422.700 23.400 427.200 ;
        RECT 21.600 421.800 23.700 422.700 ;
        RECT 14.100 420.000 21.300 420.900 ;
        RECT 14.100 415.050 15.900 416.850 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 17.100 412.950 19.200 415.050 ;
        RECT 20.100 412.950 21.300 420.000 ;
        RECT 22.800 415.050 23.700 421.800 ;
        RECT 26.100 421.200 27.900 427.200 ;
        RECT 38.100 425.400 39.900 428.400 ;
        RECT 41.100 425.400 42.900 429.000 ;
        RECT 38.700 415.050 39.900 425.400 ;
        RECT 56.700 421.200 58.500 428.400 ;
        RECT 61.800 422.400 63.600 429.000 ;
        RECT 74.400 422.400 76.200 429.000 ;
        RECT 79.500 421.200 81.300 428.400 ;
        RECT 56.700 420.300 60.900 421.200 ;
        RECT 56.100 415.050 57.900 416.850 ;
        RECT 59.700 415.050 60.900 420.300 ;
        RECT 77.100 420.300 81.300 421.200 ;
        RECT 92.700 421.200 94.500 428.400 ;
        RECT 97.800 422.400 99.600 429.000 ;
        RECT 114.000 422.400 115.800 429.000 ;
        RECT 118.500 423.600 120.300 428.400 ;
        RECT 121.500 425.400 123.300 429.000 ;
        RECT 118.500 422.400 123.600 423.600 ;
        RECT 92.700 420.300 96.900 421.200 ;
        RECT 61.950 415.050 63.750 416.850 ;
        RECT 74.250 415.050 76.050 416.850 ;
        RECT 77.100 415.050 78.300 420.300 ;
        RECT 80.100 415.050 81.900 416.850 ;
        RECT 92.100 415.050 93.900 416.850 ;
        RECT 95.700 415.050 96.900 420.300 ;
        RECT 97.950 415.050 99.750 416.850 ;
        RECT 113.100 415.050 114.900 416.850 ;
        RECT 119.250 415.050 121.050 416.850 ;
        RECT 122.700 415.050 123.600 422.400 ;
        RECT 137.100 422.400 138.900 428.400 ;
        RECT 140.100 422.400 141.900 429.000 ;
        RECT 143.100 425.400 144.900 428.400 ;
        RECT 137.100 415.050 138.300 422.400 ;
        RECT 143.700 421.500 144.900 425.400 ;
        RECT 139.200 420.600 144.900 421.500 ;
        RECT 155.100 425.400 156.900 428.400 ;
        RECT 155.100 421.500 156.300 425.400 ;
        RECT 158.100 422.400 159.900 429.000 ;
        RECT 161.100 422.400 162.900 428.400 ;
        RECT 155.100 420.600 160.800 421.500 ;
        RECT 139.200 419.700 141.000 420.600 ;
        RECT 22.800 412.950 24.900 415.050 ;
        RECT 25.800 412.950 27.900 415.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 55.950 412.950 58.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 97.950 412.950 100.050 415.050 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 118.950 412.950 121.050 415.050 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 137.100 412.950 139.200 415.050 ;
        RECT 17.100 411.150 18.900 412.950 ;
        RECT 20.100 411.150 21.900 412.950 ;
        RECT 20.700 406.800 21.900 411.150 ;
        RECT 14.100 405.900 21.900 406.800 ;
        RECT 14.100 400.800 15.000 405.900 ;
        RECT 22.800 405.000 23.700 412.950 ;
        RECT 25.800 411.150 27.600 412.950 ;
        RECT 14.100 394.800 15.900 400.800 ;
        RECT 17.100 393.000 18.900 405.000 ;
        RECT 21.600 404.100 23.700 405.000 ;
        RECT 21.600 393.600 23.400 404.100 ;
        RECT 26.100 393.000 27.900 405.600 ;
        RECT 38.700 399.600 39.900 412.950 ;
        RECT 41.100 411.150 42.900 412.950 ;
        RECT 59.700 399.600 60.900 412.950 ;
        RECT 77.100 399.600 78.300 412.950 ;
        RECT 95.700 399.600 96.900 412.950 ;
        RECT 116.250 411.150 118.050 412.950 ;
        RECT 122.700 405.600 123.600 412.950 ;
        RECT 137.100 405.600 138.300 412.950 ;
        RECT 140.100 408.300 141.000 419.700 ;
        RECT 159.000 419.700 160.800 420.600 ;
        RECT 142.500 412.950 144.600 415.050 ;
        RECT 142.800 411.150 144.600 412.950 ;
        RECT 155.400 412.950 157.500 415.050 ;
        RECT 155.400 411.150 157.200 412.950 ;
        RECT 139.200 407.400 141.000 408.300 ;
        RECT 159.000 408.300 159.900 419.700 ;
        RECT 161.700 415.050 162.900 422.400 ;
        RECT 176.100 423.300 177.900 428.400 ;
        RECT 179.100 424.200 180.900 429.000 ;
        RECT 182.100 423.300 183.900 428.400 ;
        RECT 176.100 421.950 183.900 423.300 ;
        RECT 185.100 422.400 186.900 428.400 ;
        RECT 200.100 425.400 201.900 429.000 ;
        RECT 203.100 425.400 204.900 428.400 ;
        RECT 206.100 425.400 207.900 429.000 ;
        RECT 185.100 420.300 186.300 422.400 ;
        RECT 182.700 419.400 186.300 420.300 ;
        RECT 179.100 415.050 180.900 416.850 ;
        RECT 182.700 415.050 183.900 419.400 ;
        RECT 185.100 415.050 186.900 416.850 ;
        RECT 203.400 415.050 204.300 425.400 ;
        RECT 221.100 423.300 222.900 428.400 ;
        RECT 224.100 424.200 225.900 429.000 ;
        RECT 227.100 423.300 228.900 428.400 ;
        RECT 221.100 421.950 228.900 423.300 ;
        RECT 230.100 422.400 231.900 428.400 ;
        RECT 242.100 425.400 243.900 429.000 ;
        RECT 245.100 425.400 246.900 428.400 ;
        RECT 248.100 425.400 249.900 429.000 ;
        RECT 263.100 425.400 264.900 428.400 ;
        RECT 266.100 425.400 267.900 429.000 ;
        RECT 205.950 420.450 208.050 421.050 ;
        RECT 217.950 420.450 220.050 421.050 ;
        RECT 205.950 419.550 220.050 420.450 ;
        RECT 230.100 420.300 231.300 422.400 ;
        RECT 205.950 418.950 208.050 419.550 ;
        RECT 217.950 418.950 220.050 419.550 ;
        RECT 227.700 419.400 231.300 420.300 ;
        RECT 224.100 415.050 225.900 416.850 ;
        RECT 227.700 415.050 228.900 419.400 ;
        RECT 230.100 415.050 231.900 416.850 ;
        RECT 245.400 415.050 246.300 425.400 ;
        RECT 247.950 420.450 250.050 421.050 ;
        RECT 253.950 420.450 256.050 421.050 ;
        RECT 247.950 419.550 256.050 420.450 ;
        RECT 247.950 418.950 250.050 419.550 ;
        RECT 253.950 418.950 256.050 419.550 ;
        RECT 263.700 415.050 264.900 425.400 ;
        RECT 281.700 421.200 283.500 428.400 ;
        RECT 286.800 422.400 288.600 429.000 ;
        RECT 299.700 421.200 301.500 428.400 ;
        RECT 304.800 422.400 306.600 429.000 ;
        RECT 317.100 425.400 318.900 429.000 ;
        RECT 320.100 425.400 321.900 428.400 ;
        RECT 281.700 420.300 285.900 421.200 ;
        RECT 299.700 420.300 303.900 421.200 ;
        RECT 281.100 415.050 282.900 416.850 ;
        RECT 284.700 415.050 285.900 420.300 ;
        RECT 286.950 415.050 288.750 416.850 ;
        RECT 299.100 415.050 300.900 416.850 ;
        RECT 302.700 415.050 303.900 420.300 ;
        RECT 304.950 415.050 306.750 416.850 ;
        RECT 320.100 415.050 321.300 425.400 ;
        RECT 335.100 423.300 336.900 428.400 ;
        RECT 338.100 424.200 339.900 429.000 ;
        RECT 341.100 423.300 342.900 428.400 ;
        RECT 335.100 421.950 342.900 423.300 ;
        RECT 344.100 422.400 345.900 428.400 ;
        RECT 356.100 423.300 357.900 428.400 ;
        RECT 359.100 424.200 360.900 429.000 ;
        RECT 362.100 423.300 363.900 428.400 ;
        RECT 344.100 420.300 345.300 422.400 ;
        RECT 356.100 421.950 363.900 423.300 ;
        RECT 365.100 422.400 366.900 428.400 ;
        RECT 380.100 425.400 381.900 428.400 ;
        RECT 365.100 420.300 366.300 422.400 ;
        RECT 380.100 421.500 381.300 425.400 ;
        RECT 383.100 422.400 384.900 429.000 ;
        RECT 386.100 422.400 387.900 428.400 ;
        RECT 401.100 425.400 402.900 429.000 ;
        RECT 404.100 425.400 405.900 428.400 ;
        RECT 419.700 425.400 421.500 429.000 ;
        RECT 380.100 420.600 385.800 421.500 ;
        RECT 341.700 419.400 345.300 420.300 ;
        RECT 362.700 419.400 366.300 420.300 ;
        RECT 384.000 419.700 385.800 420.600 ;
        RECT 338.100 415.050 339.900 416.850 ;
        RECT 341.700 415.050 342.900 419.400 ;
        RECT 344.100 415.050 345.900 416.850 ;
        RECT 359.100 415.050 360.900 416.850 ;
        RECT 362.700 415.050 363.900 419.400 ;
        RECT 367.950 417.450 372.000 418.050 ;
        RECT 365.100 415.050 366.900 416.850 ;
        RECT 367.950 415.950 372.450 417.450 ;
        RECT 160.800 412.950 162.900 415.050 ;
        RECT 175.950 412.950 178.050 415.050 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 244.950 412.950 247.050 415.050 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 358.950 412.950 361.050 415.050 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 159.000 407.400 160.800 408.300 ;
        RECT 139.200 406.500 144.900 407.400 ;
        RECT 113.100 404.700 120.900 405.600 ;
        RECT 38.100 393.600 39.900 399.600 ;
        RECT 41.100 393.000 42.900 399.600 ;
        RECT 56.100 393.000 57.900 399.600 ;
        RECT 59.100 393.600 60.900 399.600 ;
        RECT 62.100 393.000 63.900 399.600 ;
        RECT 74.100 393.000 75.900 399.600 ;
        RECT 77.100 393.600 78.900 399.600 ;
        RECT 80.100 393.000 81.900 399.600 ;
        RECT 92.100 393.000 93.900 399.600 ;
        RECT 95.100 393.600 96.900 399.600 ;
        RECT 98.100 393.000 99.900 399.600 ;
        RECT 113.100 393.600 114.900 404.700 ;
        RECT 116.100 393.000 117.900 403.800 ;
        RECT 119.100 393.600 120.900 404.700 ;
        RECT 122.100 393.600 123.900 405.600 ;
        RECT 137.100 393.600 138.900 405.600 ;
        RECT 140.100 393.000 141.900 403.800 ;
        RECT 143.700 399.600 144.900 406.500 ;
        RECT 143.100 393.600 144.900 399.600 ;
        RECT 155.100 406.500 160.800 407.400 ;
        RECT 155.100 399.600 156.300 406.500 ;
        RECT 161.700 405.600 162.900 412.950 ;
        RECT 176.100 411.150 177.900 412.950 ;
        RECT 182.700 405.600 183.900 412.950 ;
        RECT 200.250 411.150 202.050 412.950 ;
        RECT 203.400 405.600 204.300 412.950 ;
        RECT 206.100 411.150 207.900 412.950 ;
        RECT 221.100 411.150 222.900 412.950 ;
        RECT 227.700 405.600 228.900 412.950 ;
        RECT 242.250 411.150 244.050 412.950 ;
        RECT 245.400 405.600 246.300 412.950 ;
        RECT 248.100 411.150 249.900 412.950 ;
        RECT 155.100 393.600 156.900 399.600 ;
        RECT 158.100 393.000 159.900 403.800 ;
        RECT 161.100 393.600 162.900 405.600 ;
        RECT 176.400 393.000 178.200 405.600 ;
        RECT 181.500 404.100 183.900 405.600 ;
        RECT 181.500 393.600 183.300 404.100 ;
        RECT 184.200 401.100 186.000 402.900 ;
        RECT 184.500 393.000 186.300 399.600 ;
        RECT 200.100 393.000 201.900 405.600 ;
        RECT 203.400 404.400 207.000 405.600 ;
        RECT 205.200 393.600 207.000 404.400 ;
        RECT 221.400 393.000 223.200 405.600 ;
        RECT 226.500 404.100 228.900 405.600 ;
        RECT 226.500 393.600 228.300 404.100 ;
        RECT 229.200 401.100 231.000 402.900 ;
        RECT 229.500 393.000 231.300 399.600 ;
        RECT 242.100 393.000 243.900 405.600 ;
        RECT 245.400 404.400 249.000 405.600 ;
        RECT 247.200 393.600 249.000 404.400 ;
        RECT 263.700 399.600 264.900 412.950 ;
        RECT 266.100 411.150 267.900 412.950 ;
        RECT 284.700 399.600 285.900 412.950 ;
        RECT 302.700 399.600 303.900 412.950 ;
        RECT 317.100 411.150 318.900 412.950 ;
        RECT 320.100 399.600 321.300 412.950 ;
        RECT 335.100 411.150 336.900 412.950 ;
        RECT 341.700 405.600 342.900 412.950 ;
        RECT 356.100 411.150 357.900 412.950 ;
        RECT 362.700 405.600 363.900 412.950 ;
        RECT 371.550 412.050 372.450 415.950 ;
        RECT 367.950 410.550 372.450 412.050 ;
        RECT 380.400 412.950 382.500 415.050 ;
        RECT 380.400 411.150 382.200 412.950 ;
        RECT 367.950 409.950 372.000 410.550 ;
        RECT 384.000 408.300 384.900 419.700 ;
        RECT 386.700 415.050 387.900 422.400 ;
        RECT 404.100 415.050 405.300 425.400 ;
        RECT 422.700 423.600 424.500 428.400 ;
        RECT 419.400 422.400 424.500 423.600 ;
        RECT 427.200 422.400 429.000 429.000 ;
        RECT 419.400 415.050 420.300 422.400 ;
        RECT 443.100 419.400 444.900 429.000 ;
        RECT 449.700 420.000 451.500 428.400 ;
        RECT 467.100 422.400 468.900 428.400 ;
        RECT 467.700 420.300 468.900 422.400 ;
        RECT 470.100 423.300 471.900 428.400 ;
        RECT 473.100 424.200 474.900 429.000 ;
        RECT 476.100 423.300 477.900 428.400 ;
        RECT 470.100 421.950 477.900 423.300 ;
        RECT 491.100 427.500 498.900 428.400 ;
        RECT 491.100 422.400 492.900 427.500 ;
        RECT 494.100 422.400 495.900 426.600 ;
        RECT 497.100 423.000 498.900 427.500 ;
        RECT 500.100 423.900 501.900 429.000 ;
        RECT 503.100 423.000 504.900 428.400 ;
        RECT 518.100 425.400 519.900 429.000 ;
        RECT 521.100 425.400 522.900 428.400 ;
        RECT 524.100 425.400 525.900 429.000 ;
        RECT 494.700 420.900 495.600 422.400 ;
        RECT 497.100 422.100 504.900 423.000 ;
        RECT 449.700 418.800 453.000 420.000 ;
        RECT 467.700 419.400 471.300 420.300 ;
        RECT 494.700 419.700 499.050 420.900 ;
        RECT 421.950 415.050 423.750 416.850 ;
        RECT 428.100 415.050 429.900 416.850 ;
        RECT 443.100 415.050 444.900 416.850 ;
        RECT 449.100 415.050 450.900 416.850 ;
        RECT 452.100 415.050 453.000 418.800 ;
        RECT 467.100 415.050 468.900 416.850 ;
        RECT 470.100 415.050 471.300 419.400 ;
        RECT 478.950 417.450 483.000 418.050 ;
        RECT 486.000 417.450 490.050 418.050 ;
        RECT 473.100 415.050 474.900 416.850 ;
        RECT 478.950 415.950 483.450 417.450 ;
        RECT 485.550 417.000 490.050 417.450 ;
        RECT 385.800 412.950 387.900 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 472.950 412.950 475.050 415.050 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 384.000 407.400 385.800 408.300 ;
        RECT 263.100 393.600 264.900 399.600 ;
        RECT 266.100 393.000 267.900 399.600 ;
        RECT 281.100 393.000 282.900 399.600 ;
        RECT 284.100 393.600 285.900 399.600 ;
        RECT 287.100 393.000 288.900 399.600 ;
        RECT 299.100 393.000 300.900 399.600 ;
        RECT 302.100 393.600 303.900 399.600 ;
        RECT 305.100 393.000 306.900 399.600 ;
        RECT 317.100 393.000 318.900 399.600 ;
        RECT 320.100 393.600 321.900 399.600 ;
        RECT 335.400 393.000 337.200 405.600 ;
        RECT 340.500 404.100 342.900 405.600 ;
        RECT 340.500 393.600 342.300 404.100 ;
        RECT 343.200 401.100 345.000 402.900 ;
        RECT 343.500 393.000 345.300 399.600 ;
        RECT 356.400 393.000 358.200 405.600 ;
        RECT 361.500 404.100 363.900 405.600 ;
        RECT 380.100 406.500 385.800 407.400 ;
        RECT 361.500 393.600 363.300 404.100 ;
        RECT 364.200 401.100 366.000 402.900 ;
        RECT 380.100 399.600 381.300 406.500 ;
        RECT 386.700 405.600 387.900 412.950 ;
        RECT 401.100 411.150 402.900 412.950 ;
        RECT 364.500 393.000 366.300 399.600 ;
        RECT 380.100 393.600 381.900 399.600 ;
        RECT 383.100 393.000 384.900 403.800 ;
        RECT 386.100 393.600 387.900 405.600 ;
        RECT 404.100 399.600 405.300 412.950 ;
        RECT 419.400 405.600 420.300 412.950 ;
        RECT 424.950 411.150 426.750 412.950 ;
        RECT 446.100 411.150 447.900 412.950 ;
        RECT 421.950 408.450 424.050 409.050 ;
        RECT 442.950 408.450 445.050 409.050 ;
        RECT 421.950 407.550 445.050 408.450 ;
        RECT 421.950 406.950 424.050 407.550 ;
        RECT 442.950 406.950 445.050 407.550 ;
        RECT 401.100 393.000 402.900 399.600 ;
        RECT 404.100 393.600 405.900 399.600 ;
        RECT 419.100 393.600 420.900 405.600 ;
        RECT 422.100 404.700 429.900 405.600 ;
        RECT 422.100 393.600 423.900 404.700 ;
        RECT 425.100 393.000 426.900 403.800 ;
        RECT 428.100 393.600 429.900 404.700 ;
        RECT 452.100 400.800 453.000 412.950 ;
        RECT 470.100 405.600 471.300 412.950 ;
        RECT 476.100 411.150 477.900 412.950 ;
        RECT 482.550 411.450 483.450 415.950 ;
        RECT 484.950 415.950 490.050 417.000 ;
        RECT 484.950 412.800 487.050 415.950 ;
        RECT 494.250 415.050 496.050 416.850 ;
        RECT 498.000 415.050 499.050 419.700 ;
        RECT 505.950 417.450 510.000 418.050 ;
        RECT 513.000 417.450 517.050 418.050 ;
        RECT 490.950 412.950 493.050 415.050 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 499.950 415.050 501.750 416.850 ;
        RECT 505.950 415.950 510.450 417.450 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 479.550 410.550 483.450 411.450 ;
        RECT 491.250 411.150 493.050 412.950 ;
        RECT 472.950 408.450 475.050 409.050 ;
        RECT 479.550 408.450 480.450 410.550 ;
        RECT 472.950 407.550 480.450 408.450 ;
        RECT 472.950 406.950 475.050 407.550 ;
        RECT 498.000 405.600 499.050 412.950 ;
        RECT 503.100 411.150 504.900 412.950 ;
        RECT 509.550 412.050 510.450 415.950 ;
        RECT 505.950 410.550 510.450 412.050 ;
        RECT 512.550 415.950 517.050 417.450 ;
        RECT 512.550 412.050 513.450 415.950 ;
        RECT 521.400 415.050 522.300 425.400 ;
        RECT 536.100 419.400 537.900 429.000 ;
        RECT 542.700 420.000 544.500 428.400 ;
        RECT 560.400 422.400 562.200 429.000 ;
        RECT 565.500 421.200 567.300 428.400 ;
        RECT 578.400 422.400 580.200 429.000 ;
        RECT 583.500 421.200 585.300 428.400 ;
        RECT 563.100 420.300 567.300 421.200 ;
        RECT 581.100 420.300 585.300 421.200 ;
        RECT 599.700 421.200 601.500 428.400 ;
        RECT 604.800 422.400 606.600 429.000 ;
        RECT 617.100 428.400 618.300 429.000 ;
        RECT 617.100 425.400 618.900 428.400 ;
        RECT 620.100 425.400 621.900 428.400 ;
        RECT 620.400 421.200 621.300 425.400 ;
        RECT 623.100 423.000 624.900 429.000 ;
        RECT 626.100 422.400 627.900 428.400 ;
        RECT 599.700 420.300 603.900 421.200 ;
        RECT 620.400 420.300 625.800 421.200 ;
        RECT 542.700 418.800 546.000 420.000 ;
        RECT 531.000 417.450 535.050 418.050 ;
        RECT 530.550 415.950 535.050 417.450 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 512.550 410.550 517.050 412.050 ;
        RECT 518.250 411.150 520.050 412.950 ;
        RECT 505.950 409.950 510.000 410.550 ;
        RECT 513.000 409.950 517.050 410.550 ;
        RECT 521.400 405.600 522.300 412.950 ;
        RECT 524.100 411.150 525.900 412.950 ;
        RECT 530.550 412.050 531.450 415.950 ;
        RECT 536.100 415.050 537.900 416.850 ;
        RECT 542.100 415.050 543.900 416.850 ;
        RECT 545.100 415.050 546.000 418.800 ;
        RECT 547.950 417.450 550.050 418.050 ;
        RECT 547.950 416.550 555.450 417.450 ;
        RECT 547.950 415.950 550.050 416.550 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 530.550 410.550 535.050 412.050 ;
        RECT 539.100 411.150 540.900 412.950 ;
        RECT 531.000 409.950 535.050 410.550 ;
        RECT 523.950 408.450 526.050 409.050 ;
        RECT 535.950 408.450 538.050 409.050 ;
        RECT 523.950 407.550 538.050 408.450 ;
        RECT 523.950 406.950 526.050 407.550 ;
        RECT 535.950 406.950 538.050 407.550 ;
        RECT 470.100 404.100 472.500 405.600 ;
        RECT 468.000 401.100 469.800 402.900 ;
        RECT 446.400 399.900 453.000 400.800 ;
        RECT 446.400 399.600 447.900 399.900 ;
        RECT 443.100 393.000 444.900 399.600 ;
        RECT 446.100 393.600 447.900 399.600 ;
        RECT 452.100 399.600 453.000 399.900 ;
        RECT 449.100 393.000 450.900 399.000 ;
        RECT 452.100 393.600 453.900 399.600 ;
        RECT 467.700 393.000 469.500 399.600 ;
        RECT 470.700 393.600 472.500 404.100 ;
        RECT 475.800 393.000 477.600 405.600 ;
        RECT 492.600 393.000 494.400 405.600 ;
        RECT 497.100 393.600 500.400 405.600 ;
        RECT 503.100 393.000 504.900 405.600 ;
        RECT 518.100 393.000 519.900 405.600 ;
        RECT 521.400 404.400 525.000 405.600 ;
        RECT 523.200 393.600 525.000 404.400 ;
        RECT 545.100 400.800 546.000 412.950 ;
        RECT 554.550 412.050 555.450 416.550 ;
        RECT 560.250 415.050 562.050 416.850 ;
        RECT 563.100 415.050 564.300 420.300 ;
        RECT 566.100 415.050 567.900 416.850 ;
        RECT 578.250 415.050 580.050 416.850 ;
        RECT 581.100 415.050 582.300 420.300 ;
        RECT 584.100 415.050 585.900 416.850 ;
        RECT 599.100 415.050 600.900 416.850 ;
        RECT 602.700 415.050 603.900 420.300 ;
        RECT 623.700 419.400 625.800 420.300 ;
        RECT 604.950 415.050 606.750 416.850 ;
        RECT 617.400 415.050 619.200 416.850 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 580.950 412.950 583.050 415.050 ;
        RECT 583.950 412.950 586.050 415.050 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 617.100 412.950 619.200 415.050 ;
        RECT 620.400 412.950 622.500 415.050 ;
        RECT 554.550 410.550 559.050 412.050 ;
        RECT 555.000 409.950 559.050 410.550 ;
        RECT 539.400 399.900 546.000 400.800 ;
        RECT 539.400 399.600 540.900 399.900 ;
        RECT 536.100 393.000 537.900 399.600 ;
        RECT 539.100 393.600 540.900 399.600 ;
        RECT 545.100 399.600 546.000 399.900 ;
        RECT 563.100 399.600 564.300 412.950 ;
        RECT 581.100 399.600 582.300 412.950 ;
        RECT 583.950 408.450 586.050 408.750 ;
        RECT 592.950 408.450 595.050 409.050 ;
        RECT 583.950 407.550 595.050 408.450 ;
        RECT 583.950 406.650 586.050 407.550 ;
        RECT 592.950 406.950 595.050 407.550 ;
        RECT 583.950 402.450 586.050 403.050 ;
        RECT 595.950 402.450 598.050 403.050 ;
        RECT 583.950 401.550 598.050 402.450 ;
        RECT 583.950 400.950 586.050 401.550 ;
        RECT 595.950 400.950 598.050 401.550 ;
        RECT 602.700 399.600 603.900 412.950 ;
        RECT 621.000 411.150 622.800 412.950 ;
        RECT 623.700 408.900 624.600 419.400 ;
        RECT 627.000 415.050 627.900 422.400 ;
        RECT 638.100 422.400 639.900 428.400 ;
        RECT 641.400 423.300 643.200 429.000 ;
        RECT 645.900 423.000 647.700 428.400 ;
        RECT 650.100 423.300 651.900 429.000 ;
        RECT 638.100 421.500 642.600 422.400 ;
        RECT 640.500 419.100 642.600 421.500 ;
        RECT 645.900 420.900 646.800 423.000 ;
        RECT 653.100 422.400 654.900 428.400 ;
        RECT 653.400 421.500 654.900 422.400 ;
        RECT 665.100 423.300 666.900 428.400 ;
        RECT 668.100 424.200 669.900 429.000 ;
        RECT 671.100 423.300 672.900 428.400 ;
        RECT 665.100 421.950 672.900 423.300 ;
        RECT 674.100 422.400 675.900 428.400 ;
        RECT 689.100 425.400 690.900 429.000 ;
        RECT 692.100 425.400 693.900 428.400 ;
        RECT 643.800 418.800 646.800 420.900 ;
        RECT 650.400 420.000 654.900 421.500 ;
        RECT 674.100 420.300 675.300 422.400 ;
        RECT 625.800 412.950 627.900 415.050 ;
        RECT 638.100 412.950 640.200 415.050 ;
        RECT 642.900 414.900 645.000 417.000 ;
        RECT 643.200 413.100 645.000 414.900 ;
        RECT 623.100 408.300 624.900 408.900 ;
        RECT 617.100 407.100 624.900 408.300 ;
        RECT 617.100 405.600 618.300 407.100 ;
        RECT 625.800 405.600 627.000 412.950 ;
        RECT 638.400 411.150 640.200 412.950 ;
        RECT 645.900 412.050 646.800 418.800 ;
        RECT 647.700 417.900 649.500 419.700 ;
        RECT 650.400 419.400 652.500 420.000 ;
        RECT 671.700 419.400 675.300 420.300 ;
        RECT 648.000 417.000 650.100 417.900 ;
        RECT 648.000 415.800 654.600 417.000 ;
        RECT 652.800 415.200 654.600 415.800 ;
        RECT 648.000 412.800 650.100 414.900 ;
        RECT 652.800 412.950 654.900 415.200 ;
        RECT 668.100 415.050 669.900 416.850 ;
        RECT 671.700 415.050 672.900 419.400 ;
        RECT 674.100 415.050 675.900 416.850 ;
        RECT 692.100 415.050 693.300 425.400 ;
        RECT 707.100 419.400 708.900 429.000 ;
        RECT 713.700 420.000 715.500 428.400 ;
        RECT 728.400 422.400 730.200 429.000 ;
        RECT 733.500 421.200 735.300 428.400 ;
        RECT 749.100 425.400 750.900 429.000 ;
        RECT 752.100 425.400 753.900 428.400 ;
        RECT 764.100 425.400 765.900 429.000 ;
        RECT 767.100 425.400 768.900 428.400 ;
        RECT 731.100 420.300 735.300 421.200 ;
        RECT 713.700 418.800 717.000 420.000 ;
        RECT 707.100 415.050 708.900 416.850 ;
        RECT 713.100 415.050 714.900 416.850 ;
        RECT 716.100 415.050 717.000 418.800 ;
        RECT 728.250 415.050 730.050 416.850 ;
        RECT 731.100 415.050 732.300 420.300 ;
        RECT 734.100 415.050 735.900 416.850 ;
        RECT 752.100 415.050 753.300 425.400 ;
        RECT 767.100 415.050 768.300 425.400 ;
        RECT 782.100 423.300 783.900 428.400 ;
        RECT 785.100 424.200 786.900 429.000 ;
        RECT 788.100 423.300 789.900 428.400 ;
        RECT 782.100 421.950 789.900 423.300 ;
        RECT 791.100 422.400 792.900 428.400 ;
        RECT 806.100 425.400 807.900 429.000 ;
        RECT 809.100 425.400 810.900 428.400 ;
        RECT 791.100 420.300 792.300 422.400 ;
        RECT 788.700 419.400 792.300 420.300 ;
        RECT 785.100 415.050 786.900 416.850 ;
        RECT 788.700 415.050 789.900 419.400 ;
        RECT 791.100 415.050 792.900 416.850 ;
        RECT 809.100 415.050 810.300 425.400 ;
        RECT 824.100 423.300 825.900 428.400 ;
        RECT 827.100 424.200 828.900 429.000 ;
        RECT 830.100 423.300 831.900 428.400 ;
        RECT 824.100 421.950 831.900 423.300 ;
        RECT 833.100 422.400 834.900 428.400 ;
        RECT 833.100 420.300 834.300 422.400 ;
        RECT 845.700 421.200 847.500 428.400 ;
        RECT 850.800 422.400 852.600 429.000 ;
        RECT 845.700 420.300 849.900 421.200 ;
        RECT 830.700 419.400 834.300 420.300 ;
        RECT 827.100 415.050 828.900 416.850 ;
        RECT 830.700 415.050 831.900 419.400 ;
        RECT 833.100 415.050 834.900 416.850 ;
        RECT 845.100 415.050 846.900 416.850 ;
        RECT 848.700 415.050 849.900 420.300 ;
        RECT 866.100 420.600 867.900 428.400 ;
        RECT 870.600 422.400 872.400 429.000 ;
        RECT 873.600 424.200 875.400 428.400 ;
        RECT 873.600 422.400 876.300 424.200 ;
        RECT 890.400 422.400 892.200 429.000 ;
        RECT 872.700 420.600 874.500 421.500 ;
        RECT 866.100 419.700 874.500 420.600 ;
        RECT 850.950 415.050 852.750 416.850 ;
        RECT 866.250 415.050 868.050 416.850 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 763.950 412.950 766.050 415.050 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 787.950 412.950 790.050 415.050 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 866.100 412.950 868.200 415.050 ;
        RECT 643.800 410.700 646.800 412.050 ;
        RECT 648.300 411.000 650.100 412.800 ;
        RECT 665.100 411.150 666.900 412.950 ;
        RECT 643.800 409.950 645.900 410.700 ;
        RECT 641.100 405.600 643.200 406.500 ;
        RECT 542.100 393.000 543.900 399.000 ;
        RECT 545.100 393.600 546.900 399.600 ;
        RECT 560.100 393.000 561.900 399.600 ;
        RECT 563.100 393.600 564.900 399.600 ;
        RECT 566.100 393.000 567.900 399.600 ;
        RECT 578.100 393.000 579.900 399.600 ;
        RECT 581.100 393.600 582.900 399.600 ;
        RECT 584.100 393.000 585.900 399.600 ;
        RECT 599.100 393.000 600.900 399.600 ;
        RECT 602.100 393.600 603.900 399.600 ;
        RECT 605.100 393.000 606.900 399.600 ;
        RECT 617.100 393.600 618.900 405.600 ;
        RECT 621.600 393.000 623.400 405.600 ;
        RECT 624.600 404.100 627.000 405.600 ;
        RECT 638.100 404.400 643.200 405.600 ;
        RECT 644.100 405.600 645.300 409.950 ;
        RECT 646.800 407.700 648.600 409.500 ;
        RECT 646.800 406.800 652.200 407.700 ;
        RECT 650.100 405.900 652.200 406.800 ;
        RECT 644.100 404.700 647.400 405.600 ;
        RECT 650.100 404.700 654.900 405.900 ;
        RECT 671.700 405.600 672.900 412.950 ;
        RECT 689.100 411.150 690.900 412.950 ;
        RECT 624.600 393.600 626.400 404.100 ;
        RECT 638.100 393.600 639.900 404.400 ;
        RECT 641.100 393.000 643.200 403.500 ;
        RECT 645.600 393.600 647.400 404.700 ;
        RECT 650.100 393.000 651.900 403.500 ;
        RECT 653.100 393.600 654.900 404.700 ;
        RECT 665.400 393.000 667.200 405.600 ;
        RECT 670.500 404.100 672.900 405.600 ;
        RECT 670.500 393.600 672.300 404.100 ;
        RECT 673.200 401.100 675.000 402.900 ;
        RECT 692.100 399.600 693.300 412.950 ;
        RECT 710.100 411.150 711.900 412.950 ;
        RECT 694.950 408.450 697.050 409.050 ;
        RECT 706.950 408.450 709.050 409.050 ;
        RECT 694.950 407.550 709.050 408.450 ;
        RECT 694.950 406.950 697.050 407.550 ;
        RECT 706.950 406.950 709.050 407.550 ;
        RECT 716.100 400.800 717.000 412.950 ;
        RECT 710.400 399.900 717.000 400.800 ;
        RECT 710.400 399.600 711.900 399.900 ;
        RECT 673.500 393.000 675.300 399.600 ;
        RECT 689.100 393.000 690.900 399.600 ;
        RECT 692.100 393.600 693.900 399.600 ;
        RECT 707.100 393.000 708.900 399.600 ;
        RECT 710.100 393.600 711.900 399.600 ;
        RECT 716.100 399.600 717.000 399.900 ;
        RECT 731.100 399.600 732.300 412.950 ;
        RECT 749.100 411.150 750.900 412.950 ;
        RECT 752.100 399.600 753.300 412.950 ;
        RECT 764.100 411.150 765.900 412.950 ;
        RECT 767.100 399.600 768.300 412.950 ;
        RECT 782.100 411.150 783.900 412.950 ;
        RECT 769.950 408.450 772.050 409.050 ;
        RECT 784.950 408.450 787.050 409.050 ;
        RECT 769.950 407.550 787.050 408.450 ;
        RECT 769.950 406.950 772.050 407.550 ;
        RECT 784.950 406.950 787.050 407.550 ;
        RECT 788.700 405.600 789.900 412.950 ;
        RECT 806.100 411.150 807.900 412.950 ;
        RECT 713.100 393.000 714.900 399.000 ;
        RECT 716.100 393.600 717.900 399.600 ;
        RECT 728.100 393.000 729.900 399.600 ;
        RECT 731.100 393.600 732.900 399.600 ;
        RECT 734.100 393.000 735.900 399.600 ;
        RECT 749.100 393.000 750.900 399.600 ;
        RECT 752.100 393.600 753.900 399.600 ;
        RECT 764.100 393.000 765.900 399.600 ;
        RECT 767.100 393.600 768.900 399.600 ;
        RECT 782.400 393.000 784.200 405.600 ;
        RECT 787.500 404.100 789.900 405.600 ;
        RECT 787.500 393.600 789.300 404.100 ;
        RECT 790.200 401.100 792.000 402.900 ;
        RECT 809.100 399.600 810.300 412.950 ;
        RECT 824.100 411.150 825.900 412.950 ;
        RECT 830.700 405.600 831.900 412.950 ;
        RECT 790.500 393.000 792.300 399.600 ;
        RECT 806.100 393.000 807.900 399.600 ;
        RECT 809.100 393.600 810.900 399.600 ;
        RECT 824.400 393.000 826.200 405.600 ;
        RECT 829.500 404.100 831.900 405.600 ;
        RECT 832.950 405.450 835.050 406.050 ;
        RECT 844.950 405.450 847.050 406.050 ;
        RECT 832.950 404.550 847.050 405.450 ;
        RECT 829.500 393.600 831.300 404.100 ;
        RECT 832.950 403.950 835.050 404.550 ;
        RECT 844.950 403.950 847.050 404.550 ;
        RECT 832.200 401.100 834.000 402.900 ;
        RECT 848.700 399.600 849.900 412.950 ;
        RECT 869.100 399.600 870.000 419.700 ;
        RECT 875.400 415.050 876.300 422.400 ;
        RECT 895.500 421.200 897.300 428.400 ;
        RECT 893.100 420.300 897.300 421.200 ;
        RECT 890.250 415.050 892.050 416.850 ;
        RECT 893.100 415.050 894.300 420.300 ;
        RECT 911.100 419.400 912.900 429.000 ;
        RECT 917.700 420.000 919.500 428.400 ;
        RECT 935.700 421.200 937.500 428.400 ;
        RECT 940.800 422.400 942.600 429.000 ;
        RECT 935.700 420.300 939.900 421.200 ;
        RECT 917.700 418.800 921.000 420.000 ;
        RECT 896.100 415.050 897.900 416.850 ;
        RECT 911.100 415.050 912.900 416.850 ;
        RECT 917.100 415.050 918.900 416.850 ;
        RECT 920.100 415.050 921.000 418.800 ;
        RECT 931.950 417.450 934.050 418.050 ;
        RECT 926.550 416.550 934.050 417.450 ;
        RECT 871.500 412.950 873.600 415.050 ;
        RECT 874.800 412.950 876.900 415.050 ;
        RECT 889.950 412.950 892.050 415.050 ;
        RECT 892.950 412.950 895.050 415.050 ;
        RECT 895.950 412.950 898.050 415.050 ;
        RECT 910.950 412.950 913.050 415.050 ;
        RECT 913.950 412.950 916.050 415.050 ;
        RECT 916.950 412.950 919.050 415.050 ;
        RECT 919.950 412.950 922.050 415.050 ;
        RECT 871.200 411.150 873.000 412.950 ;
        RECT 875.400 405.600 876.300 412.950 ;
        RECT 832.500 393.000 834.300 399.600 ;
        RECT 845.100 393.000 846.900 399.600 ;
        RECT 848.100 393.600 849.900 399.600 ;
        RECT 851.100 393.000 852.900 399.600 ;
        RECT 866.100 393.000 867.900 399.600 ;
        RECT 869.100 393.600 870.900 399.600 ;
        RECT 872.100 393.000 873.900 405.000 ;
        RECT 875.100 393.600 876.900 405.600 ;
        RECT 893.100 399.600 894.300 412.950 ;
        RECT 914.100 411.150 915.900 412.950 ;
        RECT 895.950 408.450 898.050 409.050 ;
        RECT 904.950 408.450 907.050 409.050 ;
        RECT 895.950 407.550 907.050 408.450 ;
        RECT 895.950 406.950 898.050 407.550 ;
        RECT 904.950 406.950 907.050 407.550 ;
        RECT 920.100 400.800 921.000 412.950 ;
        RECT 926.550 412.050 927.450 416.550 ;
        RECT 931.950 415.950 934.050 416.550 ;
        RECT 935.100 415.050 936.900 416.850 ;
        RECT 938.700 415.050 939.900 420.300 ;
        RECT 940.950 415.050 942.750 416.850 ;
        RECT 934.950 412.950 937.050 415.050 ;
        RECT 937.950 412.950 940.050 415.050 ;
        RECT 940.950 412.950 943.050 415.050 ;
        RECT 922.950 410.550 927.450 412.050 ;
        RECT 922.950 409.950 927.000 410.550 ;
        RECT 914.400 399.900 921.000 400.800 ;
        RECT 914.400 399.600 915.900 399.900 ;
        RECT 890.100 393.000 891.900 399.600 ;
        RECT 893.100 393.600 894.900 399.600 ;
        RECT 896.100 393.000 897.900 399.600 ;
        RECT 911.100 393.000 912.900 399.600 ;
        RECT 914.100 393.600 915.900 399.600 ;
        RECT 920.100 399.600 921.000 399.900 ;
        RECT 938.700 399.600 939.900 412.950 ;
        RECT 917.100 393.000 918.900 399.000 ;
        RECT 920.100 393.600 921.900 399.600 ;
        RECT 935.100 393.000 936.900 399.600 ;
        RECT 938.100 393.600 939.900 399.600 ;
        RECT 941.100 393.000 942.900 399.600 ;
        RECT 14.100 377.400 15.900 389.400 ;
        RECT 18.600 377.400 20.400 390.000 ;
        RECT 21.600 378.900 23.400 389.400 ;
        RECT 38.100 383.400 39.900 390.000 ;
        RECT 41.100 383.400 42.900 389.400 ;
        RECT 44.100 383.400 45.900 390.000 ;
        RECT 21.600 377.400 24.000 378.900 ;
        RECT 14.100 375.900 15.300 377.400 ;
        RECT 14.100 374.700 21.900 375.900 ;
        RECT 20.100 374.100 21.900 374.700 ;
        RECT 18.000 370.050 19.800 371.850 ;
        RECT 14.100 367.950 16.200 370.050 ;
        RECT 17.400 367.950 19.500 370.050 ;
        RECT 14.400 366.150 16.200 367.950 ;
        RECT 20.700 363.600 21.600 374.100 ;
        RECT 22.800 370.050 24.000 377.400 ;
        RECT 41.100 370.050 42.300 383.400 ;
        RECT 59.400 377.400 61.200 390.000 ;
        RECT 64.500 378.900 66.300 389.400 ;
        RECT 67.500 383.400 69.300 390.000 ;
        RECT 67.200 380.100 69.000 381.900 ;
        RECT 64.500 377.400 66.900 378.900 ;
        RECT 59.100 370.050 60.900 371.850 ;
        RECT 65.700 370.050 66.900 377.400 ;
        RECT 80.100 377.400 81.900 389.400 ;
        RECT 84.600 377.400 86.400 390.000 ;
        RECT 87.600 378.900 89.400 389.400 ;
        RECT 104.100 383.400 105.900 389.400 ;
        RECT 107.100 384.000 108.900 390.000 ;
        RECT 105.000 383.100 105.900 383.400 ;
        RECT 110.100 383.400 111.900 389.400 ;
        RECT 113.100 383.400 114.900 390.000 ;
        RECT 125.100 383.400 126.900 390.000 ;
        RECT 128.100 383.400 129.900 389.400 ;
        RECT 140.100 383.400 141.900 390.000 ;
        RECT 143.100 383.400 144.900 389.400 ;
        RECT 146.100 383.400 147.900 390.000 ;
        RECT 161.100 383.400 162.900 390.000 ;
        RECT 164.100 383.400 165.900 389.400 ;
        RECT 167.100 383.400 168.900 390.000 ;
        RECT 110.100 383.100 111.600 383.400 ;
        RECT 105.000 382.200 111.600 383.100 ;
        RECT 87.600 377.400 90.000 378.900 ;
        RECT 80.100 375.900 81.300 377.400 ;
        RECT 80.100 374.700 87.900 375.900 ;
        RECT 86.100 374.100 87.900 374.700 ;
        RECT 84.000 370.050 85.800 371.850 ;
        RECT 22.800 367.950 24.900 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 67.950 367.950 70.050 370.050 ;
        RECT 80.100 367.950 82.200 370.050 ;
        RECT 83.400 367.950 85.500 370.050 ;
        RECT 20.700 362.700 22.800 363.600 ;
        RECT 17.400 361.800 22.800 362.700 ;
        RECT 17.400 357.600 18.300 361.800 ;
        RECT 24.000 360.600 24.900 367.950 ;
        RECT 38.250 366.150 40.050 367.950 ;
        RECT 41.100 362.700 42.300 367.950 ;
        RECT 44.100 366.150 45.900 367.950 ;
        RECT 62.100 366.150 63.900 367.950 ;
        RECT 65.700 363.600 66.900 367.950 ;
        RECT 68.100 366.150 69.900 367.950 ;
        RECT 80.400 366.150 82.200 367.950 ;
        RECT 86.700 363.600 87.600 374.100 ;
        RECT 88.800 370.050 90.000 377.400 ;
        RECT 105.000 370.050 105.900 382.200 ;
        RECT 110.100 370.050 111.900 371.850 ;
        RECT 125.100 370.050 126.900 371.850 ;
        RECT 128.100 370.050 129.300 383.400 ;
        RECT 143.100 370.050 144.300 383.400 ;
        RECT 145.950 375.450 148.050 376.050 ;
        RECT 151.950 375.450 154.050 376.050 ;
        RECT 145.950 374.550 154.050 375.450 ;
        RECT 145.950 373.950 148.050 374.550 ;
        RECT 151.950 373.950 154.050 374.550 ;
        RECT 164.700 370.050 165.900 383.400 ;
        RECT 182.100 377.400 183.900 389.400 ;
        RECT 185.100 379.200 186.900 390.000 ;
        RECT 188.100 383.400 189.900 389.400 ;
        RECT 203.100 383.400 204.900 390.000 ;
        RECT 206.100 383.400 207.900 389.400 ;
        RECT 209.100 383.400 210.900 390.000 ;
        RECT 224.100 388.500 231.900 389.400 ;
        RECT 182.100 370.050 183.300 377.400 ;
        RECT 188.700 376.500 189.900 383.400 ;
        RECT 184.200 375.600 189.900 376.500 ;
        RECT 184.200 374.700 186.000 375.600 ;
        RECT 88.800 367.950 90.900 370.050 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 106.950 367.950 109.050 370.050 ;
        RECT 109.950 367.950 112.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 182.100 367.950 184.200 370.050 ;
        RECT 65.700 362.700 69.300 363.600 ;
        RECT 86.700 362.700 88.800 363.600 ;
        RECT 41.100 361.800 45.300 362.700 ;
        RECT 14.100 354.600 15.900 357.600 ;
        RECT 17.100 354.600 18.900 357.600 ;
        RECT 14.100 354.000 15.300 354.600 ;
        RECT 20.100 354.000 21.900 360.000 ;
        RECT 23.100 354.600 24.900 360.600 ;
        RECT 38.400 354.000 40.200 360.600 ;
        RECT 43.500 354.600 45.300 361.800 ;
        RECT 59.100 359.700 66.900 361.050 ;
        RECT 59.100 354.600 60.900 359.700 ;
        RECT 62.100 354.000 63.900 358.800 ;
        RECT 65.100 354.600 66.900 359.700 ;
        RECT 68.100 360.600 69.300 362.700 ;
        RECT 83.400 361.800 88.800 362.700 ;
        RECT 68.100 354.600 69.900 360.600 ;
        RECT 83.400 357.600 84.300 361.800 ;
        RECT 90.000 360.600 90.900 367.950 ;
        RECT 105.000 364.200 105.900 367.950 ;
        RECT 107.100 366.150 108.900 367.950 ;
        RECT 113.100 366.150 114.900 367.950 ;
        RECT 105.000 363.000 108.300 364.200 ;
        RECT 80.100 354.600 81.900 357.600 ;
        RECT 83.100 354.600 84.900 357.600 ;
        RECT 80.100 354.000 81.300 354.600 ;
        RECT 86.100 354.000 87.900 360.000 ;
        RECT 89.100 354.600 90.900 360.600 ;
        RECT 106.500 354.600 108.300 363.000 ;
        RECT 113.100 354.000 114.900 363.600 ;
        RECT 128.100 357.600 129.300 367.950 ;
        RECT 140.250 366.150 142.050 367.950 ;
        RECT 143.100 362.700 144.300 367.950 ;
        RECT 146.100 366.150 147.900 367.950 ;
        RECT 161.100 366.150 162.900 367.950 ;
        RECT 164.700 362.700 165.900 367.950 ;
        RECT 166.950 366.150 168.750 367.950 ;
        RECT 143.100 361.800 147.300 362.700 ;
        RECT 125.100 354.000 126.900 357.600 ;
        RECT 128.100 354.600 129.900 357.600 ;
        RECT 140.400 354.000 142.200 360.600 ;
        RECT 145.500 354.600 147.300 361.800 ;
        RECT 161.700 361.800 165.900 362.700 ;
        RECT 161.700 354.600 163.500 361.800 ;
        RECT 182.100 360.600 183.300 367.950 ;
        RECT 185.100 363.300 186.000 374.700 ;
        RECT 187.800 370.050 189.600 371.850 ;
        RECT 206.100 370.050 207.300 383.400 ;
        RECT 224.100 377.400 225.900 388.500 ;
        RECT 227.100 376.500 228.900 387.600 ;
        RECT 230.100 378.600 231.900 388.500 ;
        RECT 233.100 379.500 234.900 390.000 ;
        RECT 236.100 378.600 237.900 389.400 ;
        RECT 230.100 377.700 237.900 378.600 ;
        RECT 251.100 377.400 252.900 389.400 ;
        RECT 254.100 378.000 255.900 390.000 ;
        RECT 257.100 383.400 258.900 389.400 ;
        RECT 260.100 383.400 261.900 390.000 ;
        RECT 227.100 375.600 231.900 376.500 ;
        RECT 227.100 370.050 228.900 371.850 ;
        RECT 231.000 370.050 231.900 375.600 ;
        RECT 235.950 375.450 238.050 376.050 ;
        RECT 247.950 375.450 250.050 376.050 ;
        RECT 235.950 374.550 250.050 375.450 ;
        RECT 235.950 373.950 238.050 374.550 ;
        RECT 247.950 373.950 250.050 374.550 ;
        RECT 232.950 370.050 234.750 371.850 ;
        RECT 251.700 370.050 252.600 377.400 ;
        RECT 255.000 370.050 256.800 371.850 ;
        RECT 187.500 367.950 189.600 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 205.950 367.950 208.050 370.050 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 226.950 367.950 229.050 370.050 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 251.100 367.950 253.200 370.050 ;
        RECT 254.400 367.950 256.500 370.050 ;
        RECT 203.250 366.150 205.050 367.950 ;
        RECT 184.200 362.400 186.000 363.300 ;
        RECT 206.100 362.700 207.300 367.950 ;
        RECT 209.100 366.150 210.900 367.950 ;
        RECT 224.100 366.150 225.900 367.950 ;
        RECT 217.950 363.450 220.050 364.050 ;
        RECT 223.950 363.450 226.050 364.050 ;
        RECT 184.200 361.500 189.900 362.400 ;
        RECT 206.100 361.800 210.300 362.700 ;
        RECT 217.950 362.550 226.050 363.450 ;
        RECT 217.950 361.950 220.050 362.550 ;
        RECT 223.950 361.950 226.050 362.550 ;
        RECT 166.800 354.000 168.600 360.600 ;
        RECT 182.100 354.600 183.900 360.600 ;
        RECT 185.100 354.000 186.900 360.600 ;
        RECT 188.700 357.600 189.900 361.500 ;
        RECT 188.100 354.600 189.900 357.600 ;
        RECT 203.400 354.000 205.200 360.600 ;
        RECT 208.500 354.600 210.300 361.800 ;
        RECT 230.700 360.600 231.900 367.950 ;
        RECT 235.950 366.150 237.750 367.950 ;
        RECT 251.700 360.600 252.600 367.950 ;
        RECT 258.000 363.300 258.900 383.400 ;
        RECT 272.100 377.400 273.900 389.400 ;
        RECT 275.100 379.200 276.900 390.000 ;
        RECT 278.100 383.400 279.900 389.400 ;
        RECT 272.100 370.050 273.300 377.400 ;
        RECT 278.700 376.500 279.900 383.400 ;
        RECT 274.200 375.600 279.900 376.500 ;
        RECT 293.100 383.400 294.900 389.400 ;
        RECT 293.100 376.500 294.300 383.400 ;
        RECT 296.100 379.200 297.900 390.000 ;
        RECT 299.100 377.400 300.900 389.400 ;
        RECT 314.100 377.400 315.900 390.000 ;
        RECT 319.200 378.600 321.000 389.400 ;
        RECT 317.400 377.400 321.000 378.600 ;
        RECT 332.100 377.400 333.900 389.400 ;
        RECT 335.100 378.300 336.900 389.400 ;
        RECT 338.100 379.200 339.900 390.000 ;
        RECT 341.100 378.300 342.900 389.400 ;
        RECT 335.100 377.400 342.900 378.300 ;
        RECT 356.100 377.400 357.900 389.400 ;
        RECT 359.100 378.000 360.900 390.000 ;
        RECT 362.100 383.400 363.900 389.400 ;
        RECT 365.100 383.400 366.900 390.000 ;
        RECT 380.100 383.400 381.900 390.000 ;
        RECT 383.100 383.400 384.900 389.400 ;
        RECT 293.100 375.600 298.800 376.500 ;
        RECT 274.200 374.700 276.000 375.600 ;
        RECT 259.800 367.950 261.900 370.050 ;
        RECT 272.100 367.950 274.200 370.050 ;
        RECT 259.950 366.150 261.750 367.950 ;
        RECT 253.500 362.400 261.900 363.300 ;
        RECT 253.500 361.500 255.300 362.400 ;
        RECT 226.500 354.000 228.300 360.600 ;
        RECT 231.000 354.600 232.800 360.600 ;
        RECT 235.500 354.000 237.300 360.600 ;
        RECT 251.700 358.800 254.400 360.600 ;
        RECT 252.600 354.600 254.400 358.800 ;
        RECT 255.600 354.000 257.400 360.600 ;
        RECT 260.100 354.600 261.900 362.400 ;
        RECT 272.100 360.600 273.300 367.950 ;
        RECT 275.100 363.300 276.000 374.700 ;
        RECT 297.000 374.700 298.800 375.600 ;
        RECT 277.800 370.050 279.600 371.850 ;
        RECT 277.500 367.950 279.600 370.050 ;
        RECT 293.400 370.050 295.200 371.850 ;
        RECT 293.400 367.950 295.500 370.050 ;
        RECT 274.200 362.400 276.000 363.300 ;
        RECT 297.000 363.300 297.900 374.700 ;
        RECT 299.700 370.050 300.900 377.400 ;
        RECT 314.250 370.050 316.050 371.850 ;
        RECT 317.400 370.050 318.300 377.400 ;
        RECT 327.000 372.450 331.050 373.050 ;
        RECT 320.100 370.050 321.900 371.850 ;
        RECT 326.550 370.950 331.050 372.450 ;
        RECT 298.800 367.950 300.900 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 297.000 362.400 298.800 363.300 ;
        RECT 274.200 361.500 279.900 362.400 ;
        RECT 272.100 354.600 273.900 360.600 ;
        RECT 275.100 354.000 276.900 360.600 ;
        RECT 278.700 357.600 279.900 361.500 ;
        RECT 278.100 354.600 279.900 357.600 ;
        RECT 293.100 361.500 298.800 362.400 ;
        RECT 293.100 357.600 294.300 361.500 ;
        RECT 299.700 360.600 300.900 367.950 ;
        RECT 293.100 354.600 294.900 357.600 ;
        RECT 296.100 354.000 297.900 360.600 ;
        RECT 299.100 354.600 300.900 360.600 ;
        RECT 317.400 357.600 318.300 367.950 ;
        RECT 326.550 367.050 327.450 370.950 ;
        RECT 332.400 370.050 333.300 377.400 ;
        RECT 343.950 372.450 348.000 373.050 ;
        RECT 337.950 370.050 339.750 371.850 ;
        RECT 343.950 370.950 348.450 372.450 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 326.550 365.550 331.050 367.050 ;
        RECT 327.000 364.950 331.050 365.550 ;
        RECT 332.400 360.600 333.300 367.950 ;
        RECT 334.950 366.150 336.750 367.950 ;
        RECT 341.100 366.150 342.900 367.950 ;
        RECT 334.950 363.450 337.050 364.050 ;
        RECT 347.550 363.450 348.450 370.950 ;
        RECT 356.700 370.050 357.600 377.400 ;
        RECT 360.000 370.050 361.800 371.850 ;
        RECT 356.100 367.950 358.200 370.050 ;
        RECT 359.400 367.950 361.500 370.050 ;
        RECT 334.950 362.550 348.450 363.450 ;
        RECT 334.950 361.950 337.050 362.550 ;
        RECT 356.700 360.600 357.600 367.950 ;
        RECT 363.000 363.300 363.900 383.400 ;
        RECT 364.800 367.950 366.900 370.050 ;
        RECT 380.100 367.950 382.200 370.050 ;
        RECT 364.950 366.150 366.750 367.950 ;
        RECT 380.250 366.150 382.050 367.950 ;
        RECT 383.100 363.300 384.000 383.400 ;
        RECT 386.100 378.000 387.900 390.000 ;
        RECT 389.100 377.400 390.900 389.400 ;
        RECT 401.100 383.400 402.900 390.000 ;
        RECT 404.100 383.400 405.900 389.400 ;
        RECT 385.200 370.050 387.000 371.850 ;
        RECT 389.400 370.050 390.300 377.400 ;
        RECT 385.500 367.950 387.600 370.050 ;
        RECT 388.800 367.950 390.900 370.050 ;
        RECT 401.100 367.950 403.200 370.050 ;
        RECT 358.500 362.400 366.900 363.300 ;
        RECT 358.500 361.500 360.300 362.400 ;
        RECT 332.400 359.400 337.500 360.600 ;
        RECT 314.100 354.000 315.900 357.600 ;
        RECT 317.100 354.600 318.900 357.600 ;
        RECT 320.100 354.000 321.900 357.600 ;
        RECT 332.700 354.000 334.500 357.600 ;
        RECT 335.700 354.600 337.500 359.400 ;
        RECT 340.200 354.000 342.000 360.600 ;
        RECT 356.700 358.800 359.400 360.600 ;
        RECT 357.600 354.600 359.400 358.800 ;
        RECT 360.600 354.000 362.400 360.600 ;
        RECT 365.100 354.600 366.900 362.400 ;
        RECT 380.100 362.400 388.500 363.300 ;
        RECT 380.100 354.600 381.900 362.400 ;
        RECT 386.700 361.500 388.500 362.400 ;
        RECT 389.400 360.600 390.300 367.950 ;
        RECT 401.250 366.150 403.050 367.950 ;
        RECT 404.100 363.300 405.000 383.400 ;
        RECT 407.100 378.000 408.900 390.000 ;
        RECT 410.100 377.400 411.900 389.400 ;
        RECT 425.100 383.400 426.900 390.000 ;
        RECT 428.100 383.400 429.900 389.400 ;
        RECT 431.100 383.400 432.900 390.000 ;
        RECT 446.700 383.400 448.500 390.000 ;
        RECT 406.200 370.050 408.000 371.850 ;
        RECT 410.400 370.050 411.300 377.400 ;
        RECT 428.700 370.050 429.900 383.400 ;
        RECT 430.950 381.450 433.050 382.050 ;
        RECT 442.950 381.450 445.050 382.050 ;
        RECT 430.950 380.550 445.050 381.450 ;
        RECT 430.950 379.950 433.050 380.550 ;
        RECT 442.950 379.950 445.050 380.550 ;
        RECT 447.000 380.100 448.800 381.900 ;
        RECT 430.950 378.450 433.050 378.900 ;
        RECT 436.950 378.450 439.050 379.050 ;
        RECT 449.700 378.900 451.500 389.400 ;
        RECT 430.950 377.550 439.050 378.450 ;
        RECT 430.950 376.800 433.050 377.550 ;
        RECT 436.950 376.950 439.050 377.550 ;
        RECT 449.100 377.400 451.500 378.900 ;
        RECT 454.800 377.400 456.600 390.000 ;
        RECT 470.100 388.500 477.900 389.400 ;
        RECT 470.100 377.400 471.900 388.500 ;
        RECT 449.100 370.050 450.300 377.400 ;
        RECT 473.100 376.500 474.900 387.600 ;
        RECT 476.100 378.600 477.900 388.500 ;
        RECT 479.100 379.500 480.900 390.000 ;
        RECT 482.100 378.600 483.900 389.400 ;
        RECT 497.100 383.400 498.900 390.000 ;
        RECT 500.100 383.400 501.900 389.400 ;
        RECT 503.100 383.400 504.900 390.000 ;
        RECT 515.100 383.400 516.900 390.000 ;
        RECT 518.100 383.400 519.900 389.400 ;
        RECT 521.100 383.400 522.900 390.000 ;
        RECT 476.100 377.700 483.900 378.600 ;
        RECT 473.100 375.600 477.900 376.500 ;
        RECT 455.100 370.050 456.900 371.850 ;
        RECT 473.100 370.050 474.900 371.850 ;
        RECT 477.000 370.050 477.900 375.600 ;
        RECT 478.950 370.050 480.750 371.850 ;
        RECT 500.700 370.050 501.900 383.400 ;
        RECT 502.950 375.450 505.050 376.050 ;
        RECT 514.950 375.450 517.050 376.050 ;
        RECT 502.950 374.550 517.050 375.450 ;
        RECT 502.950 373.950 505.050 374.550 ;
        RECT 514.950 373.950 517.050 374.550 ;
        RECT 505.950 372.450 510.000 373.050 ;
        RECT 505.950 370.950 510.450 372.450 ;
        RECT 406.500 367.950 408.600 370.050 ;
        RECT 409.800 367.950 411.900 370.050 ;
        RECT 424.950 367.950 427.050 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 469.950 367.950 472.050 370.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 384.600 354.000 386.400 360.600 ;
        RECT 387.600 358.800 390.300 360.600 ;
        RECT 401.100 362.400 409.500 363.300 ;
        RECT 387.600 354.600 389.400 358.800 ;
        RECT 401.100 354.600 402.900 362.400 ;
        RECT 407.700 361.500 409.500 362.400 ;
        RECT 410.400 360.600 411.300 367.950 ;
        RECT 425.100 366.150 426.900 367.950 ;
        RECT 428.700 362.700 429.900 367.950 ;
        RECT 430.950 366.150 432.750 367.950 ;
        RECT 446.100 366.150 447.900 367.950 ;
        RECT 449.100 363.600 450.300 367.950 ;
        RECT 452.100 366.150 453.900 367.950 ;
        RECT 470.100 366.150 471.900 367.950 ;
        RECT 405.600 354.000 407.400 360.600 ;
        RECT 408.600 358.800 411.300 360.600 ;
        RECT 425.700 361.800 429.900 362.700 ;
        RECT 446.700 362.700 450.300 363.600 ;
        RECT 408.600 354.600 410.400 358.800 ;
        RECT 425.700 354.600 427.500 361.800 ;
        RECT 446.700 360.600 447.900 362.700 ;
        RECT 430.800 354.000 432.600 360.600 ;
        RECT 446.100 354.600 447.900 360.600 ;
        RECT 449.100 359.700 456.900 361.050 ;
        RECT 476.700 360.600 477.900 367.950 ;
        RECT 481.950 366.150 483.750 367.950 ;
        RECT 486.000 366.450 490.050 367.050 ;
        RECT 485.550 364.950 490.050 366.450 ;
        RECT 497.100 366.150 498.900 367.950 ;
        RECT 485.550 364.050 486.450 364.950 ;
        RECT 481.950 362.550 486.450 364.050 ;
        RECT 500.700 362.700 501.900 367.950 ;
        RECT 502.950 366.150 504.750 367.950 ;
        RECT 509.550 367.050 510.450 370.950 ;
        RECT 518.100 370.050 519.300 383.400 ;
        RECT 536.100 377.400 537.900 390.000 ;
        RECT 540.600 377.400 543.900 389.400 ;
        RECT 546.600 377.400 548.400 390.000 ;
        RECT 563.100 383.400 564.900 390.000 ;
        RECT 566.100 383.400 567.900 389.400 ;
        RECT 536.100 370.050 537.900 371.850 ;
        RECT 541.950 370.050 543.000 377.400 ;
        RECT 547.950 370.050 549.750 371.850 ;
        RECT 563.100 370.050 564.900 371.850 ;
        RECT 566.100 370.050 567.300 383.400 ;
        RECT 581.100 377.400 582.900 389.400 ;
        RECT 584.100 378.000 585.900 390.000 ;
        RECT 587.100 383.400 588.900 389.400 ;
        RECT 590.100 383.400 591.900 390.000 ;
        RECT 568.950 372.450 573.000 373.050 ;
        RECT 568.950 370.950 573.450 372.450 ;
        RECT 514.950 367.950 517.050 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 509.550 365.550 514.050 367.050 ;
        RECT 515.250 366.150 517.050 367.950 ;
        RECT 510.000 364.950 514.050 365.550 ;
        RECT 481.950 361.950 486.000 362.550 ;
        RECT 497.700 361.800 501.900 362.700 ;
        RECT 518.100 362.700 519.300 367.950 ;
        RECT 521.100 366.150 522.900 367.950 ;
        RECT 539.250 366.150 541.050 367.950 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 541.950 363.300 543.000 367.950 ;
        RECT 544.950 366.150 546.750 367.950 ;
        RECT 518.100 361.800 522.300 362.700 ;
        RECT 541.950 362.100 546.300 363.300 ;
        RECT 449.100 354.600 450.900 359.700 ;
        RECT 452.100 354.000 453.900 358.800 ;
        RECT 455.100 354.600 456.900 359.700 ;
        RECT 472.500 354.000 474.300 360.600 ;
        RECT 477.000 354.600 478.800 360.600 ;
        RECT 481.500 354.000 483.300 360.600 ;
        RECT 497.700 354.600 499.500 361.800 ;
        RECT 502.800 354.000 504.600 360.600 ;
        RECT 515.400 354.000 517.200 360.600 ;
        RECT 520.500 354.600 522.300 361.800 ;
        RECT 536.100 360.000 543.900 360.900 ;
        RECT 545.400 360.600 546.300 362.100 ;
        RECT 536.100 354.600 537.900 360.000 ;
        RECT 539.100 354.000 540.900 359.100 ;
        RECT 542.100 355.500 543.900 360.000 ;
        RECT 545.100 356.400 546.900 360.600 ;
        RECT 548.100 355.500 549.900 360.600 ;
        RECT 566.100 357.600 567.300 367.950 ;
        RECT 572.550 361.050 573.450 370.950 ;
        RECT 581.700 370.050 582.600 377.400 ;
        RECT 585.000 370.050 586.800 371.850 ;
        RECT 581.100 367.950 583.200 370.050 ;
        RECT 584.400 367.950 586.500 370.050 ;
        RECT 572.550 360.900 576.000 361.050 ;
        RECT 572.550 359.550 577.050 360.900 ;
        RECT 573.000 358.950 577.050 359.550 ;
        RECT 574.950 358.800 577.050 358.950 ;
        RECT 581.700 360.600 582.600 367.950 ;
        RECT 588.000 363.300 588.900 383.400 ;
        RECT 603.000 378.600 604.800 389.400 ;
        RECT 603.000 377.400 606.600 378.600 ;
        RECT 608.100 377.400 609.900 390.000 ;
        RECT 623.400 377.400 625.200 390.000 ;
        RECT 628.500 378.900 630.300 389.400 ;
        RECT 631.500 383.400 633.300 390.000 ;
        RECT 647.100 383.400 648.900 390.000 ;
        RECT 650.100 383.400 651.900 389.400 ;
        RECT 653.100 383.400 654.900 390.000 ;
        RECT 631.200 380.100 633.000 381.900 ;
        RECT 628.500 377.400 630.900 378.900 ;
        RECT 602.100 370.050 603.900 371.850 ;
        RECT 605.700 370.050 606.600 377.400 ;
        RECT 610.950 375.450 613.050 376.050 ;
        RECT 625.950 375.450 628.050 376.050 ;
        RECT 610.950 374.550 628.050 375.450 ;
        RECT 610.950 373.950 613.050 374.550 ;
        RECT 625.950 373.950 628.050 374.550 ;
        RECT 607.950 370.050 609.750 371.850 ;
        RECT 623.100 370.050 624.900 371.850 ;
        RECT 629.700 370.050 630.900 377.400 ;
        RECT 650.100 370.050 651.300 383.400 ;
        RECT 665.100 377.400 666.900 389.400 ;
        RECT 669.600 377.400 671.400 390.000 ;
        RECT 672.600 378.900 674.400 389.400 ;
        RECT 672.600 377.400 675.000 378.900 ;
        RECT 689.100 378.300 690.900 389.400 ;
        RECT 692.100 379.200 693.900 390.000 ;
        RECT 695.100 378.300 696.900 389.400 ;
        RECT 689.100 377.400 696.900 378.300 ;
        RECT 698.100 377.400 699.900 389.400 ;
        RECT 713.100 383.400 714.900 390.000 ;
        RECT 716.100 383.400 717.900 389.400 ;
        RECT 665.100 375.900 666.300 377.400 ;
        RECT 665.100 374.700 672.900 375.900 ;
        RECT 671.100 374.100 672.900 374.700 ;
        RECT 669.000 370.050 670.800 371.850 ;
        RECT 589.800 367.950 591.900 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 665.100 367.950 667.200 370.050 ;
        RECT 668.400 367.950 670.500 370.050 ;
        RECT 589.950 366.150 591.750 367.950 ;
        RECT 583.500 362.400 591.900 363.300 ;
        RECT 583.500 361.500 585.300 362.400 ;
        RECT 581.700 358.800 584.400 360.600 ;
        RECT 542.100 354.600 549.900 355.500 ;
        RECT 563.100 354.000 564.900 357.600 ;
        RECT 566.100 354.600 567.900 357.600 ;
        RECT 582.600 354.600 584.400 358.800 ;
        RECT 585.600 354.000 587.400 360.600 ;
        RECT 590.100 354.600 591.900 362.400 ;
        RECT 605.700 357.600 606.600 367.950 ;
        RECT 626.100 366.150 627.900 367.950 ;
        RECT 629.700 363.600 630.900 367.950 ;
        RECT 632.100 366.150 633.900 367.950 ;
        RECT 647.250 366.150 649.050 367.950 ;
        RECT 629.700 362.700 633.300 363.600 ;
        RECT 623.100 359.700 630.900 361.050 ;
        RECT 602.100 354.000 603.900 357.600 ;
        RECT 605.100 354.600 606.900 357.600 ;
        RECT 608.100 354.000 609.900 357.600 ;
        RECT 623.100 354.600 624.900 359.700 ;
        RECT 626.100 354.000 627.900 358.800 ;
        RECT 629.100 354.600 630.900 359.700 ;
        RECT 632.100 360.600 633.300 362.700 ;
        RECT 650.100 362.700 651.300 367.950 ;
        RECT 653.100 366.150 654.900 367.950 ;
        RECT 665.400 366.150 667.200 367.950 ;
        RECT 671.700 363.600 672.600 374.100 ;
        RECT 673.800 370.050 675.000 377.400 ;
        RECT 692.250 370.050 694.050 371.850 ;
        RECT 698.700 370.050 699.600 377.400 ;
        RECT 673.800 367.950 675.900 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 713.100 367.950 715.200 370.050 ;
        RECT 671.700 362.700 673.800 363.600 ;
        RECT 650.100 361.800 654.300 362.700 ;
        RECT 632.100 354.600 633.900 360.600 ;
        RECT 647.400 354.000 649.200 360.600 ;
        RECT 652.500 354.600 654.300 361.800 ;
        RECT 668.400 361.800 673.800 362.700 ;
        RECT 668.400 357.600 669.300 361.800 ;
        RECT 675.000 360.600 675.900 367.950 ;
        RECT 689.100 366.150 690.900 367.950 ;
        RECT 695.250 366.150 697.050 367.950 ;
        RECT 698.700 360.600 699.600 367.950 ;
        RECT 713.250 366.150 715.050 367.950 ;
        RECT 716.100 363.300 717.000 383.400 ;
        RECT 719.100 378.000 720.900 390.000 ;
        RECT 722.100 377.400 723.900 389.400 ;
        RECT 737.100 378.600 738.900 389.400 ;
        RECT 740.100 379.500 741.900 390.000 ;
        RECT 743.100 388.500 750.900 389.400 ;
        RECT 743.100 378.600 744.900 388.500 ;
        RECT 737.100 377.700 744.900 378.600 ;
        RECT 718.200 370.050 720.000 371.850 ;
        RECT 722.400 370.050 723.300 377.400 ;
        RECT 746.100 376.500 747.900 387.600 ;
        RECT 749.100 377.400 750.900 388.500 ;
        RECT 764.100 383.400 765.900 390.000 ;
        RECT 767.100 383.400 768.900 389.400 ;
        RECT 770.100 384.000 771.900 390.000 ;
        RECT 767.400 383.100 768.900 383.400 ;
        RECT 773.100 383.400 774.900 389.400 ;
        RECT 773.100 383.100 774.000 383.400 ;
        RECT 767.400 382.200 774.000 383.100 ;
        RECT 743.100 375.600 747.900 376.500 ;
        RECT 740.250 370.050 742.050 371.850 ;
        RECT 743.100 370.050 744.000 375.600 ;
        RECT 746.100 370.050 747.900 371.850 ;
        RECT 767.100 370.050 768.900 371.850 ;
        RECT 773.100 370.050 774.000 382.200 ;
        RECT 788.100 378.300 789.900 389.400 ;
        RECT 791.100 379.200 792.900 390.000 ;
        RECT 794.100 378.300 795.900 389.400 ;
        RECT 788.100 377.400 795.900 378.300 ;
        RECT 797.100 377.400 798.900 389.400 ;
        RECT 809.400 377.400 811.200 390.000 ;
        RECT 814.500 378.900 816.300 389.400 ;
        RECT 817.500 383.400 819.300 390.000 ;
        RECT 817.200 380.100 819.000 381.900 ;
        RECT 814.500 377.400 816.900 378.900 ;
        RECT 830.400 377.400 832.200 390.000 ;
        RECT 835.500 378.900 837.300 389.400 ;
        RECT 838.500 383.400 840.300 390.000 ;
        RECT 854.100 383.400 855.900 389.400 ;
        RECT 857.100 383.400 858.900 390.000 ;
        RECT 872.100 383.400 873.900 390.000 ;
        RECT 875.100 383.400 876.900 389.400 ;
        RECT 878.100 384.000 879.900 390.000 ;
        RECT 838.200 380.100 840.000 381.900 ;
        RECT 835.500 377.400 837.900 378.900 ;
        RECT 791.250 370.050 793.050 371.850 ;
        RECT 797.700 370.050 798.600 377.400 ;
        RECT 809.100 370.050 810.900 371.850 ;
        RECT 815.700 370.050 816.900 377.400 ;
        RECT 830.100 370.050 831.900 371.850 ;
        RECT 836.700 370.050 837.900 377.400 ;
        RECT 838.950 375.450 841.050 376.050 ;
        RECT 847.950 375.450 850.050 376.050 ;
        RECT 838.950 374.550 850.050 375.450 ;
        RECT 838.950 373.950 841.050 374.550 ;
        RECT 847.950 373.950 850.050 374.550 ;
        RECT 854.700 370.050 855.900 383.400 ;
        RECT 875.400 383.100 876.900 383.400 ;
        RECT 881.100 383.400 882.900 389.400 ;
        RECT 896.100 383.400 897.900 390.000 ;
        RECT 899.100 383.400 900.900 389.400 ;
        RECT 902.100 384.000 903.900 390.000 ;
        RECT 881.100 383.100 882.000 383.400 ;
        RECT 875.400 382.200 882.000 383.100 ;
        RECT 899.400 383.100 900.900 383.400 ;
        RECT 905.100 383.400 906.900 389.400 ;
        RECT 920.100 383.400 921.900 389.400 ;
        RECT 923.100 384.000 924.900 390.000 ;
        RECT 905.100 383.100 906.000 383.400 ;
        RECT 899.400 382.200 906.000 383.100 ;
        RECT 867.000 372.450 871.050 373.050 ;
        RECT 857.100 370.050 858.900 371.850 ;
        RECT 866.550 370.950 871.050 372.450 ;
        RECT 718.500 367.950 720.600 370.050 ;
        RECT 721.800 367.950 723.900 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 739.950 367.950 742.050 370.050 ;
        RECT 742.950 367.950 745.050 370.050 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 769.950 367.950 772.050 370.050 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 790.950 367.950 793.050 370.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 835.950 367.950 838.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 665.100 354.600 666.900 357.600 ;
        RECT 668.100 354.600 669.900 357.600 ;
        RECT 665.100 354.000 666.300 354.600 ;
        RECT 671.100 354.000 672.900 360.000 ;
        RECT 674.100 354.600 675.900 360.600 ;
        RECT 690.000 354.000 691.800 360.600 ;
        RECT 694.500 359.400 699.600 360.600 ;
        RECT 713.100 362.400 721.500 363.300 ;
        RECT 694.500 354.600 696.300 359.400 ;
        RECT 697.500 354.000 699.300 357.600 ;
        RECT 713.100 354.600 714.900 362.400 ;
        RECT 719.700 361.500 721.500 362.400 ;
        RECT 722.400 360.600 723.300 367.950 ;
        RECT 737.250 366.150 739.050 367.950 ;
        RECT 743.100 360.600 744.300 367.950 ;
        RECT 749.100 366.150 750.900 367.950 ;
        RECT 764.100 366.150 765.900 367.950 ;
        RECT 770.100 366.150 771.900 367.950 ;
        RECT 773.100 364.200 774.000 367.950 ;
        RECT 788.100 366.150 789.900 367.950 ;
        RECT 794.250 366.150 796.050 367.950 ;
        RECT 717.600 354.000 719.400 360.600 ;
        RECT 720.600 358.800 723.300 360.600 ;
        RECT 720.600 354.600 722.400 358.800 ;
        RECT 737.700 354.000 739.500 360.600 ;
        RECT 742.200 354.600 744.000 360.600 ;
        RECT 746.700 354.000 748.500 360.600 ;
        RECT 764.100 354.000 765.900 363.600 ;
        RECT 770.700 363.000 774.000 364.200 ;
        RECT 770.700 354.600 772.500 363.000 ;
        RECT 797.700 360.600 798.600 367.950 ;
        RECT 812.100 366.150 813.900 367.950 ;
        RECT 815.700 363.600 816.900 367.950 ;
        RECT 818.100 366.150 819.900 367.950 ;
        RECT 833.100 366.150 834.900 367.950 ;
        RECT 836.700 363.600 837.900 367.950 ;
        RECT 839.100 366.150 840.900 367.950 ;
        RECT 815.700 362.700 819.300 363.600 ;
        RECT 836.700 362.700 840.300 363.600 ;
        RECT 789.000 354.000 790.800 360.600 ;
        RECT 793.500 359.400 798.600 360.600 ;
        RECT 809.100 359.700 816.900 361.050 ;
        RECT 793.500 354.600 795.300 359.400 ;
        RECT 796.500 354.000 798.300 357.600 ;
        RECT 809.100 354.600 810.900 359.700 ;
        RECT 812.100 354.000 813.900 358.800 ;
        RECT 815.100 354.600 816.900 359.700 ;
        RECT 818.100 360.600 819.300 362.700 ;
        RECT 818.100 354.600 819.900 360.600 ;
        RECT 830.100 359.700 837.900 361.050 ;
        RECT 830.100 354.600 831.900 359.700 ;
        RECT 833.100 354.000 834.900 358.800 ;
        RECT 836.100 354.600 837.900 359.700 ;
        RECT 839.100 360.600 840.300 362.700 ;
        RECT 839.100 354.600 840.900 360.600 ;
        RECT 854.700 357.600 855.900 367.950 ;
        RECT 859.950 366.450 862.050 367.050 ;
        RECT 866.550 366.450 867.450 370.950 ;
        RECT 875.100 370.050 876.900 371.850 ;
        RECT 881.100 370.050 882.000 382.200 ;
        RECT 891.000 372.450 895.050 373.050 ;
        RECT 890.550 370.950 895.050 372.450 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 880.950 367.950 883.050 370.050 ;
        RECT 859.950 365.550 867.450 366.450 ;
        RECT 872.100 366.150 873.900 367.950 ;
        RECT 878.100 366.150 879.900 367.950 ;
        RECT 859.950 364.950 862.050 365.550 ;
        RECT 881.100 364.200 882.000 367.950 ;
        RECT 890.550 367.050 891.450 370.950 ;
        RECT 899.100 370.050 900.900 371.850 ;
        RECT 905.100 370.050 906.000 382.200 ;
        RECT 921.000 383.100 921.900 383.400 ;
        RECT 926.100 383.400 927.900 389.400 ;
        RECT 929.100 383.400 930.900 390.000 ;
        RECT 926.100 383.100 927.600 383.400 ;
        RECT 921.000 382.200 927.600 383.100 ;
        RECT 907.950 372.450 912.000 373.050 ;
        RECT 907.950 370.950 912.450 372.450 ;
        RECT 895.950 367.950 898.050 370.050 ;
        RECT 898.950 367.950 901.050 370.050 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 890.550 365.550 895.050 367.050 ;
        RECT 896.100 366.150 897.900 367.950 ;
        RECT 902.100 366.150 903.900 367.950 ;
        RECT 891.000 364.950 895.050 365.550 ;
        RECT 905.100 364.200 906.000 367.950 ;
        RECT 911.550 366.450 912.450 370.950 ;
        RECT 921.000 370.050 921.900 382.200 ;
        RECT 922.950 375.450 925.050 375.900 ;
        RECT 934.950 375.450 937.050 376.050 ;
        RECT 922.950 374.550 937.050 375.450 ;
        RECT 922.950 373.800 925.050 374.550 ;
        RECT 934.950 373.950 937.050 374.550 ;
        RECT 926.100 370.050 927.900 371.850 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 922.950 367.950 925.050 370.050 ;
        RECT 925.950 367.950 928.050 370.050 ;
        RECT 928.950 367.950 931.050 370.050 ;
        RECT 916.950 366.450 919.050 367.050 ;
        RECT 911.550 365.550 919.050 366.450 ;
        RECT 916.950 364.950 919.050 365.550 ;
        RECT 854.100 354.600 855.900 357.600 ;
        RECT 857.100 354.000 858.900 357.600 ;
        RECT 872.100 354.000 873.900 363.600 ;
        RECT 878.700 363.000 882.000 364.200 ;
        RECT 878.700 354.600 880.500 363.000 ;
        RECT 896.100 354.000 897.900 363.600 ;
        RECT 902.700 363.000 906.000 364.200 ;
        RECT 921.000 364.200 921.900 367.950 ;
        RECT 923.100 366.150 924.900 367.950 ;
        RECT 929.100 366.150 930.900 367.950 ;
        RECT 921.000 363.000 924.300 364.200 ;
        RECT 902.700 354.600 904.500 363.000 ;
        RECT 922.500 354.600 924.300 363.000 ;
        RECT 929.100 354.000 930.900 363.600 ;
        RECT 937.950 360.450 940.050 361.050 ;
        RECT 943.950 360.450 946.050 360.900 ;
        RECT 937.950 359.550 946.050 360.450 ;
        RECT 937.950 358.950 940.050 359.550 ;
        RECT 943.950 358.800 946.050 359.550 ;
        RECT 14.100 342.600 15.900 350.400 ;
        RECT 18.600 344.400 20.400 351.000 ;
        RECT 21.600 346.200 23.400 350.400 ;
        RECT 21.600 344.400 24.300 346.200 ;
        RECT 38.100 344.400 39.900 350.400 ;
        RECT 20.700 342.600 22.500 343.500 ;
        RECT 14.100 341.700 22.500 342.600 ;
        RECT 14.250 337.050 16.050 338.850 ;
        RECT 14.100 334.950 16.200 337.050 ;
        RECT 17.100 321.600 18.000 341.700 ;
        RECT 23.400 337.050 24.300 344.400 ;
        RECT 38.700 342.300 39.900 344.400 ;
        RECT 41.100 345.300 42.900 350.400 ;
        RECT 44.100 346.200 45.900 351.000 ;
        RECT 47.100 345.300 48.900 350.400 ;
        RECT 59.100 347.400 60.900 351.000 ;
        RECT 62.100 347.400 63.900 350.400 ;
        RECT 41.100 343.950 48.900 345.300 ;
        RECT 38.700 341.400 42.300 342.300 ;
        RECT 38.100 337.050 39.900 338.850 ;
        RECT 41.100 337.050 42.300 341.400 ;
        RECT 44.100 337.050 45.900 338.850 ;
        RECT 62.100 337.050 63.300 347.400 ;
        RECT 77.400 344.400 79.200 351.000 ;
        RECT 82.500 343.200 84.300 350.400 ;
        RECT 95.100 347.400 96.900 350.400 ;
        RECT 98.100 347.400 99.900 351.000 ;
        RECT 80.100 342.300 84.300 343.200 ;
        RECT 77.250 337.050 79.050 338.850 ;
        RECT 80.100 337.050 81.300 342.300 ;
        RECT 83.100 337.050 84.900 338.850 ;
        RECT 95.700 337.050 96.900 347.400 ;
        RECT 113.100 344.400 114.900 350.400 ;
        RECT 113.700 342.300 114.900 344.400 ;
        RECT 116.100 345.300 117.900 350.400 ;
        RECT 119.100 346.200 120.900 351.000 ;
        RECT 122.100 345.300 123.900 350.400 ;
        RECT 116.100 343.950 123.900 345.300 ;
        RECT 137.400 344.400 139.200 351.000 ;
        RECT 142.500 343.200 144.300 350.400 ;
        RECT 140.100 342.300 144.300 343.200 ;
        RECT 113.700 341.400 117.300 342.300 ;
        RECT 113.100 337.050 114.900 338.850 ;
        RECT 116.100 337.050 117.300 341.400 ;
        RECT 119.100 337.050 120.900 338.850 ;
        RECT 137.250 337.050 139.050 338.850 ;
        RECT 140.100 337.050 141.300 342.300 ;
        RECT 158.100 341.400 159.900 351.000 ;
        RECT 164.700 342.000 166.500 350.400 ;
        RECT 179.100 345.300 180.900 350.400 ;
        RECT 182.100 346.200 183.900 351.000 ;
        RECT 185.100 345.300 186.900 350.400 ;
        RECT 179.100 343.950 186.900 345.300 ;
        RECT 188.100 344.400 189.900 350.400 ;
        RECT 202.800 347.400 204.900 351.000 ;
        RECT 206.100 347.400 207.900 350.400 ;
        RECT 209.100 347.400 210.900 351.000 ;
        RECT 212.100 347.400 214.800 350.400 ;
        RECT 206.700 346.500 207.600 347.400 ;
        RECT 213.900 346.500 214.800 347.400 ;
        RECT 206.700 345.600 219.300 346.500 ;
        RECT 188.100 342.300 189.300 344.400 ;
        RECT 164.700 340.800 168.000 342.000 ;
        RECT 143.100 337.050 144.900 338.850 ;
        RECT 158.100 337.050 159.900 338.850 ;
        RECT 164.100 337.050 165.900 338.850 ;
        RECT 167.100 337.050 168.000 340.800 ;
        RECT 185.700 341.400 189.300 342.300 ;
        RECT 190.950 342.450 193.050 343.050 ;
        RECT 202.950 342.450 205.050 343.050 ;
        RECT 190.950 341.550 205.050 342.450 ;
        RECT 182.100 337.050 183.900 338.850 ;
        RECT 185.700 337.050 186.900 341.400 ;
        RECT 190.950 340.950 193.050 341.550 ;
        RECT 202.950 340.950 205.050 341.550 ;
        RECT 188.100 337.050 189.900 338.850 ;
        RECT 208.950 337.050 210.750 338.850 ;
        RECT 218.100 337.050 219.300 345.600 ;
        RECT 236.400 344.400 238.200 351.000 ;
        RECT 241.500 343.200 243.300 350.400 ;
        RECT 257.100 347.400 258.900 351.000 ;
        RECT 260.100 347.400 261.900 350.400 ;
        RECT 239.100 342.300 243.300 343.200 ;
        RECT 236.250 337.050 238.050 338.850 ;
        RECT 239.100 337.050 240.300 342.300 ;
        RECT 242.100 337.050 243.900 338.850 ;
        RECT 260.100 337.050 261.300 347.400 ;
        RECT 275.100 341.400 276.900 351.000 ;
        RECT 281.700 342.000 283.500 350.400 ;
        RECT 300.000 344.400 301.800 351.000 ;
        RECT 304.500 345.600 306.300 350.400 ;
        RECT 307.500 347.400 309.300 351.000 ;
        RECT 304.500 344.400 309.600 345.600 ;
        RECT 323.400 344.400 325.200 351.000 ;
        RECT 281.700 340.800 285.000 342.000 ;
        RECT 275.100 337.050 276.900 338.850 ;
        RECT 281.100 337.050 282.900 338.850 ;
        RECT 284.100 337.050 285.000 340.800 ;
        RECT 299.100 337.050 300.900 338.850 ;
        RECT 305.250 337.050 307.050 338.850 ;
        RECT 308.700 337.050 309.600 344.400 ;
        RECT 328.500 343.200 330.300 350.400 ;
        RECT 345.000 344.400 346.800 351.000 ;
        RECT 349.500 345.600 351.300 350.400 ;
        RECT 352.500 347.400 354.300 351.000 ;
        RECT 365.100 347.400 366.900 350.400 ;
        RECT 349.500 344.400 354.600 345.600 ;
        RECT 326.100 342.300 330.300 343.200 ;
        RECT 337.950 342.450 340.050 343.050 ;
        RECT 346.950 342.450 349.050 343.200 ;
        RECT 323.250 337.050 325.050 338.850 ;
        RECT 326.100 337.050 327.300 342.300 ;
        RECT 337.950 341.550 349.050 342.450 ;
        RECT 337.950 340.950 340.050 341.550 ;
        RECT 346.950 341.100 349.050 341.550 ;
        RECT 329.100 337.050 330.900 338.850 ;
        RECT 344.100 337.050 345.900 338.850 ;
        RECT 350.250 337.050 352.050 338.850 ;
        RECT 353.700 337.050 354.600 344.400 ;
        RECT 365.100 343.500 366.300 347.400 ;
        RECT 368.100 344.400 369.900 351.000 ;
        RECT 371.100 344.400 372.900 350.400 ;
        RECT 365.100 342.600 370.800 343.500 ;
        RECT 369.000 341.700 370.800 342.600 ;
        RECT 19.500 334.950 21.600 337.050 ;
        RECT 22.800 334.950 24.900 337.050 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 94.950 334.950 97.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 115.950 334.950 118.050 337.050 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 121.950 334.950 124.050 337.050 ;
        RECT 136.950 334.950 139.050 337.050 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 202.800 334.950 204.900 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 217.500 334.950 219.600 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 304.950 334.950 307.050 337.050 ;
        RECT 307.950 334.950 310.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 365.400 334.950 367.500 337.050 ;
        RECT 19.200 333.150 21.000 334.950 ;
        RECT 23.400 327.600 24.300 334.950 ;
        RECT 41.100 327.600 42.300 334.950 ;
        RECT 47.100 333.150 48.900 334.950 ;
        RECT 59.100 333.150 60.900 334.950 ;
        RECT 14.100 315.000 15.900 321.600 ;
        RECT 17.100 315.600 18.900 321.600 ;
        RECT 20.100 315.000 21.900 327.000 ;
        RECT 23.100 315.600 24.900 327.600 ;
        RECT 41.100 326.100 43.500 327.600 ;
        RECT 39.000 323.100 40.800 324.900 ;
        RECT 38.700 315.000 40.500 321.600 ;
        RECT 41.700 315.600 43.500 326.100 ;
        RECT 46.800 315.000 48.600 327.600 ;
        RECT 62.100 321.600 63.300 334.950 ;
        RECT 80.100 321.600 81.300 334.950 ;
        RECT 95.700 321.600 96.900 334.950 ;
        RECT 98.100 333.150 99.900 334.950 ;
        RECT 116.100 327.600 117.300 334.950 ;
        RECT 122.100 333.150 123.900 334.950 ;
        RECT 116.100 326.100 118.500 327.600 ;
        RECT 114.000 323.100 115.800 324.900 ;
        RECT 59.100 315.000 60.900 321.600 ;
        RECT 62.100 315.600 63.900 321.600 ;
        RECT 77.100 315.000 78.900 321.600 ;
        RECT 80.100 315.600 81.900 321.600 ;
        RECT 83.100 315.000 84.900 321.600 ;
        RECT 95.100 315.600 96.900 321.600 ;
        RECT 98.100 315.000 99.900 321.600 ;
        RECT 113.700 315.000 115.500 321.600 ;
        RECT 116.700 315.600 118.500 326.100 ;
        RECT 121.800 315.000 123.600 327.600 ;
        RECT 140.100 321.600 141.300 334.950 ;
        RECT 161.100 333.150 162.900 334.950 ;
        RECT 142.950 327.450 145.050 328.050 ;
        RECT 151.950 327.450 154.050 328.050 ;
        RECT 163.950 327.450 166.050 328.050 ;
        RECT 142.950 326.550 166.050 327.450 ;
        RECT 142.950 325.950 145.050 326.550 ;
        RECT 151.950 325.950 154.050 326.550 ;
        RECT 163.950 325.950 166.050 326.550 ;
        RECT 167.100 322.800 168.000 334.950 ;
        RECT 179.100 333.150 180.900 334.950 ;
        RECT 185.700 327.600 186.900 334.950 ;
        RECT 203.100 333.150 204.900 334.950 ;
        RECT 212.250 333.150 214.050 334.950 ;
        RECT 161.400 321.900 168.000 322.800 ;
        RECT 161.400 321.600 162.900 321.900 ;
        RECT 137.100 315.000 138.900 321.600 ;
        RECT 140.100 315.600 141.900 321.600 ;
        RECT 143.100 315.000 144.900 321.600 ;
        RECT 158.100 315.000 159.900 321.600 ;
        RECT 161.100 315.600 162.900 321.600 ;
        RECT 167.100 321.600 168.000 321.900 ;
        RECT 164.100 315.000 165.900 321.000 ;
        RECT 167.100 315.600 168.900 321.600 ;
        RECT 179.400 315.000 181.200 327.600 ;
        RECT 184.500 326.100 186.900 327.600 ;
        RECT 184.500 315.600 186.300 326.100 ;
        RECT 200.100 325.500 207.900 326.400 ;
        RECT 187.200 323.100 189.000 324.900 ;
        RECT 187.500 315.000 189.300 321.600 ;
        RECT 200.100 315.600 201.900 325.500 ;
        RECT 203.100 315.000 204.900 324.600 ;
        RECT 206.100 316.500 207.900 325.500 ;
        RECT 209.100 325.200 216.900 326.100 ;
        RECT 209.100 317.400 210.900 325.200 ;
        RECT 212.100 316.500 213.900 324.300 ;
        RECT 206.100 315.600 213.900 316.500 ;
        RECT 215.100 316.500 216.900 325.200 ;
        RECT 218.100 325.200 219.300 334.950 ;
        RECT 218.100 317.400 219.900 325.200 ;
        RECT 221.100 316.500 222.900 325.800 ;
        RECT 239.100 321.600 240.300 334.950 ;
        RECT 257.100 333.150 258.900 334.950 ;
        RECT 260.100 321.600 261.300 334.950 ;
        RECT 278.100 333.150 279.900 334.950 ;
        RECT 284.100 322.800 285.000 334.950 ;
        RECT 302.250 333.150 304.050 334.950 ;
        RECT 295.950 330.450 298.050 331.050 ;
        RECT 301.950 330.450 304.050 331.050 ;
        RECT 295.950 329.550 304.050 330.450 ;
        RECT 295.950 328.950 298.050 329.550 ;
        RECT 301.950 328.950 304.050 329.550 ;
        RECT 308.700 327.600 309.600 334.950 ;
        RECT 278.400 321.900 285.000 322.800 ;
        RECT 278.400 321.600 279.900 321.900 ;
        RECT 215.100 315.600 222.900 316.500 ;
        RECT 236.100 315.000 237.900 321.600 ;
        RECT 239.100 315.600 240.900 321.600 ;
        RECT 242.100 315.000 243.900 321.600 ;
        RECT 257.100 315.000 258.900 321.600 ;
        RECT 260.100 315.600 261.900 321.600 ;
        RECT 275.100 315.000 276.900 321.600 ;
        RECT 278.100 315.600 279.900 321.600 ;
        RECT 284.100 321.600 285.000 321.900 ;
        RECT 299.100 326.700 306.900 327.600 ;
        RECT 281.100 315.000 282.900 321.000 ;
        RECT 284.100 315.600 285.900 321.600 ;
        RECT 299.100 315.600 300.900 326.700 ;
        RECT 302.100 315.000 303.900 325.800 ;
        RECT 305.100 315.600 306.900 326.700 ;
        RECT 308.100 315.600 309.900 327.600 ;
        RECT 326.100 321.600 327.300 334.950 ;
        RECT 347.250 333.150 349.050 334.950 ;
        RECT 328.950 330.450 331.050 331.050 ;
        RECT 334.950 330.450 337.050 331.050 ;
        RECT 340.950 330.450 343.050 331.050 ;
        RECT 328.950 329.550 343.050 330.450 ;
        RECT 328.950 328.950 331.050 329.550 ;
        RECT 334.950 328.950 337.050 329.550 ;
        RECT 340.950 328.950 343.050 329.550 ;
        RECT 353.700 327.600 354.600 334.950 ;
        RECT 365.400 333.150 367.200 334.950 ;
        RECT 369.000 330.300 369.900 341.700 ;
        RECT 371.700 337.050 372.900 344.400 ;
        RECT 383.100 347.400 384.900 350.400 ;
        RECT 383.100 343.500 384.300 347.400 ;
        RECT 386.100 344.400 387.900 351.000 ;
        RECT 389.100 344.400 390.900 350.400 ;
        RECT 383.100 342.600 388.800 343.500 ;
        RECT 387.000 341.700 388.800 342.600 ;
        RECT 370.800 334.950 372.900 337.050 ;
        RECT 369.000 329.400 370.800 330.300 ;
        RECT 365.100 328.500 370.800 329.400 ;
        RECT 344.100 326.700 351.900 327.600 ;
        RECT 323.100 315.000 324.900 321.600 ;
        RECT 326.100 315.600 327.900 321.600 ;
        RECT 329.100 315.000 330.900 321.600 ;
        RECT 344.100 315.600 345.900 326.700 ;
        RECT 347.100 315.000 348.900 325.800 ;
        RECT 350.100 315.600 351.900 326.700 ;
        RECT 353.100 315.600 354.900 327.600 ;
        RECT 365.100 321.600 366.300 328.500 ;
        RECT 371.700 327.600 372.900 334.950 ;
        RECT 383.400 334.950 385.500 337.050 ;
        RECT 383.400 333.150 385.200 334.950 ;
        RECT 387.000 330.300 387.900 341.700 ;
        RECT 389.700 337.050 390.900 344.400 ;
        RECT 404.100 344.400 405.900 350.400 ;
        RECT 407.100 345.300 408.900 351.000 ;
        RECT 411.300 345.000 413.100 350.400 ;
        RECT 415.800 345.300 417.600 351.000 ;
        RECT 404.100 343.500 405.600 344.400 ;
        RECT 404.100 342.000 408.600 343.500 ;
        RECT 406.500 341.400 408.600 342.000 ;
        RECT 412.200 342.900 413.100 345.000 ;
        RECT 419.100 344.400 420.900 350.400 ;
        RECT 431.100 344.400 432.900 350.400 ;
        RECT 416.400 343.500 420.900 344.400 ;
        RECT 409.500 339.900 411.300 341.700 ;
        RECT 412.200 340.800 415.200 342.900 ;
        RECT 416.400 341.100 418.500 343.500 ;
        RECT 431.700 342.300 432.900 344.400 ;
        RECT 434.100 345.300 435.900 350.400 ;
        RECT 437.100 346.200 438.900 351.000 ;
        RECT 440.100 345.300 441.900 350.400 ;
        RECT 453.600 346.200 455.400 350.400 ;
        RECT 434.100 343.950 441.900 345.300 ;
        RECT 452.700 344.400 455.400 346.200 ;
        RECT 456.600 344.400 458.400 351.000 ;
        RECT 431.700 341.400 435.300 342.300 ;
        RECT 408.900 339.000 411.000 339.900 ;
        RECT 404.400 337.800 411.000 339.000 ;
        RECT 404.400 337.200 406.200 337.800 ;
        RECT 388.800 334.950 390.900 337.050 ;
        RECT 404.100 334.950 406.200 337.200 ;
        RECT 387.000 329.400 388.800 330.300 ;
        RECT 365.100 315.600 366.900 321.600 ;
        RECT 368.100 315.000 369.900 325.800 ;
        RECT 371.100 315.600 372.900 327.600 ;
        RECT 383.100 328.500 388.800 329.400 ;
        RECT 383.100 321.600 384.300 328.500 ;
        RECT 389.700 327.600 390.900 334.950 ;
        RECT 408.900 334.800 411.000 336.900 ;
        RECT 408.900 333.000 410.700 334.800 ;
        RECT 412.200 334.050 413.100 340.800 ;
        RECT 414.000 336.900 416.100 339.000 ;
        RECT 431.100 337.050 432.900 338.850 ;
        RECT 434.100 337.050 435.300 341.400 ;
        RECT 442.950 339.450 445.050 340.050 ;
        RECT 437.100 337.050 438.900 338.850 ;
        RECT 442.950 338.550 450.450 339.450 ;
        RECT 442.950 337.950 445.050 338.550 ;
        RECT 414.000 335.100 415.800 336.900 ;
        RECT 418.800 334.950 420.900 337.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 412.200 332.700 415.200 334.050 ;
        RECT 418.800 333.150 420.600 334.950 ;
        RECT 413.100 331.950 415.200 332.700 ;
        RECT 410.400 329.700 412.200 331.500 ;
        RECT 406.800 328.800 412.200 329.700 ;
        RECT 406.800 327.900 408.900 328.800 ;
        RECT 383.100 315.600 384.900 321.600 ;
        RECT 386.100 315.000 387.900 325.800 ;
        RECT 389.100 315.600 390.900 327.600 ;
        RECT 404.100 326.700 408.900 327.900 ;
        RECT 413.700 327.600 414.900 331.950 ;
        RECT 411.600 326.700 414.900 327.600 ;
        RECT 415.800 327.600 417.900 328.500 ;
        RECT 434.100 327.600 435.300 334.950 ;
        RECT 440.100 333.150 441.900 334.950 ;
        RECT 449.550 333.900 450.450 338.550 ;
        RECT 452.700 337.050 453.600 344.400 ;
        RECT 454.500 342.600 456.300 343.500 ;
        RECT 461.100 342.600 462.900 350.400 ;
        RECT 476.100 345.300 477.900 350.400 ;
        RECT 479.100 346.200 480.900 351.000 ;
        RECT 482.100 345.300 483.900 350.400 ;
        RECT 476.100 343.950 483.900 345.300 ;
        RECT 485.100 344.400 486.900 350.400 ;
        RECT 454.500 341.700 462.900 342.600 ;
        RECT 485.100 342.300 486.300 344.400 ;
        RECT 497.700 343.200 499.500 350.400 ;
        RECT 502.800 344.400 504.600 351.000 ;
        RECT 515.100 344.400 516.900 350.400 ;
        RECT 452.100 334.950 454.200 337.050 ;
        RECT 455.400 334.950 457.500 337.050 ;
        RECT 448.950 331.800 451.050 333.900 ;
        RECT 452.700 327.600 453.600 334.950 ;
        RECT 456.000 333.150 457.800 334.950 ;
        RECT 404.100 315.600 405.900 326.700 ;
        RECT 407.100 315.000 408.900 325.500 ;
        RECT 411.600 315.600 413.400 326.700 ;
        RECT 415.800 326.400 420.900 327.600 ;
        RECT 415.800 315.000 417.900 325.500 ;
        RECT 419.100 315.600 420.900 326.400 ;
        RECT 434.100 326.100 436.500 327.600 ;
        RECT 432.000 323.100 433.800 324.900 ;
        RECT 431.700 315.000 433.500 321.600 ;
        RECT 434.700 315.600 436.500 326.100 ;
        RECT 439.800 315.000 441.600 327.600 ;
        RECT 442.950 324.450 445.050 324.900 ;
        RECT 448.950 324.450 451.050 325.050 ;
        RECT 442.950 323.550 451.050 324.450 ;
        RECT 442.950 322.800 445.050 323.550 ;
        RECT 448.950 322.950 451.050 323.550 ;
        RECT 452.100 315.600 453.900 327.600 ;
        RECT 455.100 315.000 456.900 327.000 ;
        RECT 459.000 321.600 459.900 341.700 ;
        RECT 482.700 341.400 486.300 342.300 ;
        RECT 466.950 339.450 469.050 339.900 ;
        RECT 472.950 339.450 475.050 340.050 ;
        RECT 460.950 337.050 462.750 338.850 ;
        RECT 466.950 338.550 475.050 339.450 ;
        RECT 466.950 337.800 469.050 338.550 ;
        RECT 472.950 337.950 475.050 338.550 ;
        RECT 479.100 337.050 480.900 338.850 ;
        RECT 482.700 337.050 483.900 341.400 ;
        RECT 487.950 339.450 490.050 343.050 ;
        RECT 497.700 342.300 501.900 343.200 ;
        RECT 493.950 339.450 496.050 340.050 ;
        RECT 487.950 339.000 496.050 339.450 ;
        RECT 485.100 337.050 486.900 338.850 ;
        RECT 488.550 338.550 496.050 339.000 ;
        RECT 493.950 337.950 496.050 338.550 ;
        RECT 497.100 337.050 498.900 338.850 ;
        RECT 500.700 337.050 501.900 342.300 ;
        RECT 515.700 342.300 516.900 344.400 ;
        RECT 518.100 345.300 519.900 350.400 ;
        RECT 521.100 346.200 522.900 351.000 ;
        RECT 524.100 345.300 525.900 350.400 ;
        RECT 518.100 343.950 525.900 345.300 ;
        RECT 515.700 341.400 519.300 342.300 ;
        RECT 502.950 337.050 504.750 338.850 ;
        RECT 515.100 337.050 516.900 338.850 ;
        RECT 518.100 337.050 519.300 341.400 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 536.100 341.400 537.900 351.000 ;
        RECT 542.700 342.000 544.500 350.400 ;
        RECT 557.400 344.400 559.200 351.000 ;
        RECT 562.500 343.200 564.300 350.400 ;
        RECT 575.100 347.400 576.900 351.000 ;
        RECT 578.100 347.400 579.900 350.400 ;
        RECT 581.100 347.400 582.900 351.000 ;
        RECT 596.100 347.400 597.900 351.000 ;
        RECT 599.100 347.400 600.900 350.400 ;
        RECT 560.100 342.300 564.300 343.200 ;
        RECT 574.950 343.050 577.050 343.200 ;
        RECT 573.000 342.450 577.050 343.050 ;
        RECT 521.100 337.050 522.900 338.850 ;
        RECT 460.800 334.950 462.900 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 476.100 333.150 477.900 334.950 ;
        RECT 482.700 327.600 483.900 334.950 ;
        RECT 458.100 315.600 459.900 321.600 ;
        RECT 461.100 315.000 462.900 321.600 ;
        RECT 476.400 315.000 478.200 327.600 ;
        RECT 481.500 326.100 483.900 327.600 ;
        RECT 481.500 315.600 483.300 326.100 ;
        RECT 484.200 323.100 486.000 324.900 ;
        RECT 500.700 321.600 501.900 334.950 ;
        RECT 502.950 330.450 505.050 331.050 ;
        RECT 514.950 330.450 517.050 331.050 ;
        RECT 502.950 329.550 517.050 330.450 ;
        RECT 502.950 328.950 505.050 329.550 ;
        RECT 514.950 328.950 517.050 329.550 ;
        RECT 518.100 327.600 519.300 334.950 ;
        RECT 524.100 333.150 525.900 334.950 ;
        RECT 530.550 333.450 531.450 340.950 ;
        RECT 542.700 340.800 546.000 342.000 ;
        RECT 536.100 337.050 537.900 338.850 ;
        RECT 542.100 337.050 543.900 338.850 ;
        RECT 545.100 337.050 546.000 340.800 ;
        RECT 557.250 337.050 559.050 338.850 ;
        RECT 560.100 337.050 561.300 342.300 ;
        RECT 572.550 341.100 577.050 342.450 ;
        RECT 572.550 340.950 576.000 341.100 ;
        RECT 572.550 339.450 573.450 340.950 ;
        RECT 563.100 337.050 564.900 338.850 ;
        RECT 569.550 338.550 573.450 339.450 ;
        RECT 535.950 334.950 538.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 530.550 332.550 534.450 333.450 ;
        RECT 539.100 333.150 540.900 334.950 ;
        RECT 533.550 330.450 534.450 332.550 ;
        RECT 538.950 330.450 541.050 331.050 ;
        RECT 533.550 329.550 541.050 330.450 ;
        RECT 538.950 328.950 541.050 329.550 ;
        RECT 518.100 326.100 520.500 327.600 ;
        RECT 516.000 323.100 517.800 324.900 ;
        RECT 484.500 315.000 486.300 321.600 ;
        RECT 497.100 315.000 498.900 321.600 ;
        RECT 500.100 315.600 501.900 321.600 ;
        RECT 503.100 315.000 504.900 321.600 ;
        RECT 515.700 315.000 517.500 321.600 ;
        RECT 518.700 315.600 520.500 326.100 ;
        RECT 523.800 315.000 525.600 327.600 ;
        RECT 545.100 322.800 546.000 334.950 ;
        RECT 539.400 321.900 546.000 322.800 ;
        RECT 539.400 321.600 540.900 321.900 ;
        RECT 536.100 315.000 537.900 321.600 ;
        RECT 539.100 315.600 540.900 321.600 ;
        RECT 545.100 321.600 546.000 321.900 ;
        RECT 560.100 321.600 561.300 334.950 ;
        RECT 569.550 334.050 570.450 338.550 ;
        RECT 578.400 337.050 579.300 347.400 ;
        RECT 580.950 345.450 583.050 346.050 ;
        RECT 592.950 345.450 595.050 346.050 ;
        RECT 580.950 344.550 595.050 345.450 ;
        RECT 580.950 343.950 583.050 344.550 ;
        RECT 592.950 343.950 595.050 344.550 ;
        RECT 599.100 337.050 600.300 347.400 ;
        RECT 611.100 341.400 612.900 351.000 ;
        RECT 617.700 342.000 619.500 350.400 ;
        RECT 635.100 347.400 636.900 350.400 ;
        RECT 638.100 347.400 639.900 351.000 ;
        RECT 617.700 340.800 621.000 342.000 ;
        RECT 611.100 337.050 612.900 338.850 ;
        RECT 617.100 337.050 618.900 338.850 ;
        RECT 620.100 337.050 621.000 340.800 ;
        RECT 635.700 337.050 636.900 347.400 ;
        RECT 650.700 343.200 652.500 350.400 ;
        RECT 655.800 344.400 657.600 351.000 ;
        RECT 668.700 343.200 670.500 350.400 ;
        RECT 673.800 344.400 675.600 351.000 ;
        RECT 650.700 342.300 654.900 343.200 ;
        RECT 668.700 342.300 672.900 343.200 ;
        RECT 650.100 337.050 651.900 338.850 ;
        RECT 653.700 337.050 654.900 342.300 ;
        RECT 655.950 337.050 657.750 338.850 ;
        RECT 668.100 337.050 669.900 338.850 ;
        RECT 671.700 337.050 672.900 342.300 ;
        RECT 689.100 341.400 690.900 351.000 ;
        RECT 695.700 342.000 697.500 350.400 ;
        RECT 714.000 344.400 715.800 351.000 ;
        RECT 718.500 345.600 720.300 350.400 ;
        RECT 721.500 347.400 723.300 351.000 ;
        RECT 734.100 347.400 735.900 351.000 ;
        RECT 737.100 347.400 738.900 350.400 ;
        RECT 718.500 344.400 723.600 345.600 ;
        RECT 695.700 340.800 699.000 342.000 ;
        RECT 673.950 337.050 675.750 338.850 ;
        RECT 689.100 337.050 690.900 338.850 ;
        RECT 695.100 337.050 696.900 338.850 ;
        RECT 698.100 337.050 699.000 340.800 ;
        RECT 713.100 337.050 714.900 338.850 ;
        RECT 719.250 337.050 721.050 338.850 ;
        RECT 722.700 337.050 723.600 344.400 ;
        RECT 737.100 337.050 738.300 347.400 ;
        RECT 752.100 345.300 753.900 350.400 ;
        RECT 755.100 346.200 756.900 351.000 ;
        RECT 758.100 345.300 759.900 350.400 ;
        RECT 752.100 343.950 759.900 345.300 ;
        RECT 761.100 344.400 762.900 350.400 ;
        RECT 776.100 345.300 777.900 350.400 ;
        RECT 779.100 346.200 780.900 351.000 ;
        RECT 782.100 345.300 783.900 350.400 ;
        RECT 761.100 342.300 762.300 344.400 ;
        RECT 776.100 343.950 783.900 345.300 ;
        RECT 785.100 344.400 786.900 350.400 ;
        RECT 798.000 344.400 799.800 351.000 ;
        RECT 802.500 345.600 804.300 350.400 ;
        RECT 805.500 347.400 807.300 351.000 ;
        RECT 802.500 344.400 807.600 345.600 ;
        RECT 785.100 342.300 786.300 344.400 ;
        RECT 758.700 341.400 762.300 342.300 ;
        RECT 782.700 341.400 786.300 342.300 ;
        RECT 755.100 337.050 756.900 338.850 ;
        RECT 758.700 337.050 759.900 341.400 ;
        RECT 761.100 337.050 762.900 338.850 ;
        RECT 779.100 337.050 780.900 338.850 ;
        RECT 782.700 337.050 783.900 341.400 ;
        RECT 792.000 339.450 796.050 340.050 ;
        RECT 785.100 337.050 786.900 338.850 ;
        RECT 791.550 337.950 796.050 339.450 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 757.950 334.950 760.050 337.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 569.550 332.550 574.050 334.050 ;
        RECT 575.250 333.150 577.050 334.950 ;
        RECT 570.000 331.950 574.050 332.550 ;
        RECT 578.400 327.600 579.300 334.950 ;
        RECT 581.100 333.150 582.900 334.950 ;
        RECT 596.100 333.150 597.900 334.950 ;
        RECT 542.100 315.000 543.900 321.000 ;
        RECT 545.100 315.600 546.900 321.600 ;
        RECT 557.100 315.000 558.900 321.600 ;
        RECT 560.100 315.600 561.900 321.600 ;
        RECT 563.100 315.000 564.900 321.600 ;
        RECT 575.100 315.000 576.900 327.600 ;
        RECT 578.400 326.400 582.000 327.600 ;
        RECT 580.200 315.600 582.000 326.400 ;
        RECT 599.100 321.600 600.300 334.950 ;
        RECT 614.100 333.150 615.900 334.950 ;
        RECT 620.100 322.800 621.000 334.950 ;
        RECT 614.400 321.900 621.000 322.800 ;
        RECT 614.400 321.600 615.900 321.900 ;
        RECT 596.100 315.000 597.900 321.600 ;
        RECT 599.100 315.600 600.900 321.600 ;
        RECT 611.100 315.000 612.900 321.600 ;
        RECT 614.100 315.600 615.900 321.600 ;
        RECT 620.100 321.600 621.000 321.900 ;
        RECT 635.700 321.600 636.900 334.950 ;
        RECT 638.100 333.150 639.900 334.950 ;
        RECT 653.700 321.600 654.900 334.950 ;
        RECT 671.700 321.600 672.900 334.950 ;
        RECT 692.100 333.150 693.900 334.950 ;
        RECT 673.950 330.450 676.050 331.050 ;
        RECT 688.950 330.450 691.050 331.050 ;
        RECT 673.950 329.550 691.050 330.450 ;
        RECT 673.950 328.950 676.050 329.550 ;
        RECT 688.950 328.950 691.050 329.550 ;
        RECT 698.100 322.800 699.000 334.950 ;
        RECT 716.250 333.150 718.050 334.950 ;
        RECT 722.700 327.600 723.600 334.950 ;
        RECT 734.100 333.150 735.900 334.950 ;
        RECT 692.400 321.900 699.000 322.800 ;
        RECT 692.400 321.600 693.900 321.900 ;
        RECT 617.100 315.000 618.900 321.000 ;
        RECT 620.100 315.600 621.900 321.600 ;
        RECT 635.100 315.600 636.900 321.600 ;
        RECT 638.100 315.000 639.900 321.600 ;
        RECT 650.100 315.000 651.900 321.600 ;
        RECT 653.100 315.600 654.900 321.600 ;
        RECT 656.100 315.000 657.900 321.600 ;
        RECT 668.100 315.000 669.900 321.600 ;
        RECT 671.100 315.600 672.900 321.600 ;
        RECT 674.100 315.000 675.900 321.600 ;
        RECT 689.100 315.000 690.900 321.600 ;
        RECT 692.100 315.600 693.900 321.600 ;
        RECT 698.100 321.600 699.000 321.900 ;
        RECT 713.100 326.700 720.900 327.600 ;
        RECT 695.100 315.000 696.900 321.000 ;
        RECT 698.100 315.600 699.900 321.600 ;
        RECT 713.100 315.600 714.900 326.700 ;
        RECT 716.100 315.000 717.900 325.800 ;
        RECT 719.100 315.600 720.900 326.700 ;
        RECT 722.100 315.600 723.900 327.600 ;
        RECT 737.100 321.600 738.300 334.950 ;
        RECT 752.100 333.150 753.900 334.950 ;
        RECT 758.700 327.600 759.900 334.950 ;
        RECT 776.100 333.150 777.900 334.950 ;
        RECT 760.950 330.450 763.050 330.750 ;
        RECT 778.950 330.450 781.050 331.050 ;
        RECT 760.950 329.550 781.050 330.450 ;
        RECT 760.950 328.650 763.050 329.550 ;
        RECT 778.950 328.950 781.050 329.550 ;
        RECT 782.700 327.600 783.900 334.950 ;
        RECT 791.550 334.050 792.450 337.950 ;
        RECT 797.100 337.050 798.900 338.850 ;
        RECT 803.250 337.050 805.050 338.850 ;
        RECT 806.700 337.050 807.600 344.400 ;
        RECT 821.100 341.400 822.900 351.000 ;
        RECT 827.700 342.000 829.500 350.400 ;
        RECT 827.700 340.800 831.000 342.000 ;
        RECT 845.100 341.400 846.900 351.000 ;
        RECT 851.700 342.000 853.500 350.400 ;
        RECT 870.000 344.400 871.800 351.000 ;
        RECT 874.500 345.600 876.300 350.400 ;
        RECT 877.500 347.400 879.300 351.000 ;
        RECT 874.500 344.400 879.600 345.600 ;
        RECT 851.700 340.800 855.000 342.000 ;
        RECT 821.100 337.050 822.900 338.850 ;
        RECT 827.100 337.050 828.900 338.850 ;
        RECT 830.100 337.050 831.000 340.800 ;
        RECT 845.100 337.050 846.900 338.850 ;
        RECT 851.100 337.050 852.900 338.850 ;
        RECT 854.100 337.050 855.000 340.800 ;
        RECT 869.100 337.050 870.900 338.850 ;
        RECT 875.250 337.050 877.050 338.850 ;
        RECT 878.700 337.050 879.600 344.400 ;
        RECT 895.500 342.000 897.300 350.400 ;
        RECT 894.000 340.800 897.300 342.000 ;
        RECT 902.100 341.400 903.900 351.000 ;
        RECT 914.400 344.400 916.200 351.000 ;
        RECT 919.500 343.200 921.300 350.400 ;
        RECT 917.100 342.300 921.300 343.200 ;
        RECT 894.000 337.050 894.900 340.800 ;
        RECT 909.000 339.450 913.050 340.050 ;
        RECT 896.100 337.050 897.900 338.850 ;
        RECT 902.100 337.050 903.900 338.850 ;
        RECT 908.550 337.950 913.050 339.450 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 787.950 332.550 792.450 334.050 ;
        RECT 800.250 333.150 802.050 334.950 ;
        RECT 787.950 331.950 792.000 332.550 ;
        RECT 806.700 327.600 807.600 334.950 ;
        RECT 824.100 333.150 825.900 334.950 ;
        RECT 808.950 330.450 811.050 331.050 ;
        RECT 826.950 330.450 829.050 331.050 ;
        RECT 808.950 329.550 829.050 330.450 ;
        RECT 808.950 328.950 811.050 329.550 ;
        RECT 826.950 328.950 829.050 329.550 ;
        RECT 734.100 315.000 735.900 321.600 ;
        RECT 737.100 315.600 738.900 321.600 ;
        RECT 752.400 315.000 754.200 327.600 ;
        RECT 757.500 326.100 759.900 327.600 ;
        RECT 757.500 315.600 759.300 326.100 ;
        RECT 760.200 323.100 762.000 324.900 ;
        RECT 760.500 315.000 762.300 321.600 ;
        RECT 776.400 315.000 778.200 327.600 ;
        RECT 781.500 326.100 783.900 327.600 ;
        RECT 797.100 326.700 804.900 327.600 ;
        RECT 781.500 315.600 783.300 326.100 ;
        RECT 784.200 323.100 786.000 324.900 ;
        RECT 784.500 315.000 786.300 321.600 ;
        RECT 797.100 315.600 798.900 326.700 ;
        RECT 800.100 315.000 801.900 325.800 ;
        RECT 803.100 315.600 804.900 326.700 ;
        RECT 806.100 315.600 807.900 327.600 ;
        RECT 830.100 322.800 831.000 334.950 ;
        RECT 848.100 333.150 849.900 334.950 ;
        RECT 838.950 327.450 841.050 328.050 ;
        RECT 850.950 327.450 853.050 328.050 ;
        RECT 838.950 326.550 853.050 327.450 ;
        RECT 838.950 325.950 841.050 326.550 ;
        RECT 850.950 325.950 853.050 326.550 ;
        RECT 854.100 322.800 855.000 334.950 ;
        RECT 872.250 333.150 874.050 334.950 ;
        RECT 878.700 327.600 879.600 334.950 ;
        RECT 824.400 321.900 831.000 322.800 ;
        RECT 824.400 321.600 825.900 321.900 ;
        RECT 821.100 315.000 822.900 321.600 ;
        RECT 824.100 315.600 825.900 321.600 ;
        RECT 830.100 321.600 831.000 321.900 ;
        RECT 848.400 321.900 855.000 322.800 ;
        RECT 848.400 321.600 849.900 321.900 ;
        RECT 827.100 315.000 828.900 321.000 ;
        RECT 830.100 315.600 831.900 321.600 ;
        RECT 845.100 315.000 846.900 321.600 ;
        RECT 848.100 315.600 849.900 321.600 ;
        RECT 854.100 321.600 855.000 321.900 ;
        RECT 869.100 326.700 876.900 327.600 ;
        RECT 851.100 315.000 852.900 321.000 ;
        RECT 854.100 315.600 855.900 321.600 ;
        RECT 869.100 315.600 870.900 326.700 ;
        RECT 872.100 315.000 873.900 325.800 ;
        RECT 875.100 315.600 876.900 326.700 ;
        RECT 878.100 315.600 879.900 327.600 ;
        RECT 894.000 322.800 894.900 334.950 ;
        RECT 899.100 333.150 900.900 334.950 ;
        RECT 908.550 334.050 909.450 337.950 ;
        RECT 914.250 337.050 916.050 338.850 ;
        RECT 917.100 337.050 918.300 342.300 ;
        RECT 935.100 341.400 936.900 351.000 ;
        RECT 941.700 342.000 943.500 350.400 ;
        RECT 941.700 340.800 945.000 342.000 ;
        RECT 930.000 339.450 934.050 340.050 ;
        RECT 920.100 337.050 921.900 338.850 ;
        RECT 929.550 337.950 934.050 339.450 ;
        RECT 913.950 334.950 916.050 337.050 ;
        RECT 916.950 334.950 919.050 337.050 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 908.550 332.550 913.050 334.050 ;
        RECT 909.000 331.950 913.050 332.550 ;
        RECT 901.950 330.450 904.050 331.050 ;
        RECT 913.950 330.450 916.050 331.050 ;
        RECT 901.950 329.550 916.050 330.450 ;
        RECT 901.950 328.950 904.050 329.550 ;
        RECT 913.950 328.950 916.050 329.550 ;
        RECT 894.000 321.900 900.600 322.800 ;
        RECT 894.000 321.600 894.900 321.900 ;
        RECT 893.100 315.600 894.900 321.600 ;
        RECT 899.100 321.600 900.600 321.900 ;
        RECT 917.100 321.600 918.300 334.950 ;
        RECT 922.950 333.450 925.050 334.050 ;
        RECT 929.550 333.450 930.450 337.950 ;
        RECT 935.100 337.050 936.900 338.850 ;
        RECT 941.100 337.050 942.900 338.850 ;
        RECT 944.100 337.050 945.000 340.800 ;
        RECT 934.950 334.950 937.050 337.050 ;
        RECT 937.950 334.950 940.050 337.050 ;
        RECT 940.950 334.950 943.050 337.050 ;
        RECT 943.950 334.950 946.050 337.050 ;
        RECT 922.950 332.550 930.450 333.450 ;
        RECT 938.100 333.150 939.900 334.950 ;
        RECT 922.950 331.950 925.050 332.550 ;
        RECT 944.100 322.800 945.000 334.950 ;
        RECT 938.400 321.900 945.000 322.800 ;
        RECT 938.400 321.600 939.900 321.900 ;
        RECT 896.100 315.000 897.900 321.000 ;
        RECT 899.100 315.600 900.900 321.600 ;
        RECT 902.100 315.000 903.900 321.600 ;
        RECT 914.100 315.000 915.900 321.600 ;
        RECT 917.100 315.600 918.900 321.600 ;
        RECT 920.100 315.000 921.900 321.600 ;
        RECT 935.100 315.000 936.900 321.600 ;
        RECT 938.100 315.600 939.900 321.600 ;
        RECT 944.100 321.600 945.000 321.900 ;
        RECT 941.100 315.000 942.900 321.000 ;
        RECT 944.100 315.600 945.900 321.600 ;
        RECT 14.100 299.400 15.900 312.000 ;
        RECT 19.200 300.600 21.000 311.400 ;
        RECT 17.400 299.400 21.000 300.600 ;
        RECT 35.400 299.400 37.200 312.000 ;
        RECT 40.500 300.900 42.300 311.400 ;
        RECT 43.500 305.400 45.300 312.000 ;
        RECT 56.100 305.400 57.900 312.000 ;
        RECT 59.100 305.400 60.900 311.400 ;
        RECT 62.100 306.000 63.900 312.000 ;
        RECT 59.400 305.100 60.900 305.400 ;
        RECT 65.100 305.400 66.900 311.400 ;
        RECT 65.100 305.100 66.000 305.400 ;
        RECT 59.400 304.200 66.000 305.100 ;
        RECT 43.200 302.100 45.000 303.900 ;
        RECT 40.500 299.400 42.900 300.900 ;
        RECT 14.250 292.050 16.050 293.850 ;
        RECT 17.400 292.050 18.300 299.400 ;
        RECT 37.950 297.450 40.050 298.050 ;
        RECT 29.550 296.550 40.050 297.450 ;
        RECT 20.100 292.050 21.900 293.850 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 17.400 279.600 18.300 289.950 ;
        RECT 29.550 279.900 30.450 296.550 ;
        RECT 37.950 295.950 40.050 296.550 ;
        RECT 35.100 292.050 36.900 293.850 ;
        RECT 41.700 292.050 42.900 299.400 ;
        RECT 59.100 292.050 60.900 293.850 ;
        RECT 65.100 292.050 66.000 304.200 ;
        RECT 80.100 300.300 81.900 311.400 ;
        RECT 83.100 301.200 84.900 312.000 ;
        RECT 86.100 300.300 87.900 311.400 ;
        RECT 80.100 299.400 87.900 300.300 ;
        RECT 89.100 299.400 90.900 311.400 ;
        RECT 101.100 305.400 102.900 312.000 ;
        RECT 104.100 305.400 105.900 311.400 ;
        RECT 107.100 305.400 108.900 312.000 ;
        RECT 119.100 310.500 126.900 311.400 ;
        RECT 67.950 297.450 70.050 298.050 ;
        RECT 73.950 297.450 76.050 298.050 ;
        RECT 85.950 297.450 88.050 298.050 ;
        RECT 67.950 296.550 88.050 297.450 ;
        RECT 67.950 295.950 70.050 296.550 ;
        RECT 73.950 295.950 76.050 296.550 ;
        RECT 85.950 295.950 88.050 296.550 ;
        RECT 83.250 292.050 85.050 293.850 ;
        RECT 89.700 292.050 90.600 299.400 ;
        RECT 104.700 292.050 105.900 305.400 ;
        RECT 119.100 299.400 120.900 310.500 ;
        RECT 122.100 298.500 123.900 309.600 ;
        RECT 125.100 300.600 126.900 310.500 ;
        RECT 128.100 301.500 129.900 312.000 ;
        RECT 131.100 300.600 132.900 311.400 ;
        RECT 143.100 305.400 144.900 312.000 ;
        RECT 146.100 305.400 147.900 311.400 ;
        RECT 161.100 305.400 162.900 312.000 ;
        RECT 164.100 305.400 165.900 311.400 ;
        RECT 179.100 305.400 180.900 311.400 ;
        RECT 182.100 306.000 183.900 312.000 ;
        RECT 125.100 299.700 132.900 300.600 ;
        RECT 122.100 297.600 126.900 298.500 ;
        RECT 114.000 294.450 118.050 295.050 ;
        RECT 113.550 292.950 118.050 294.450 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 38.100 288.150 39.900 289.950 ;
        RECT 41.700 285.600 42.900 289.950 ;
        RECT 44.100 288.150 45.900 289.950 ;
        RECT 56.100 288.150 57.900 289.950 ;
        RECT 62.100 288.150 63.900 289.950 ;
        RECT 65.100 286.200 66.000 289.950 ;
        RECT 80.100 288.150 81.900 289.950 ;
        RECT 86.250 288.150 88.050 289.950 ;
        RECT 41.700 284.700 45.300 285.600 ;
        RECT 35.100 281.700 42.900 283.050 ;
        RECT 14.100 276.000 15.900 279.600 ;
        RECT 17.100 276.600 18.900 279.600 ;
        RECT 20.100 276.000 21.900 279.600 ;
        RECT 28.950 277.800 31.050 279.900 ;
        RECT 35.100 276.600 36.900 281.700 ;
        RECT 38.100 276.000 39.900 280.800 ;
        RECT 41.100 276.600 42.900 281.700 ;
        RECT 44.100 282.600 45.300 284.700 ;
        RECT 44.100 276.600 45.900 282.600 ;
        RECT 56.100 276.000 57.900 285.600 ;
        RECT 62.700 285.000 66.000 286.200 ;
        RECT 62.700 276.600 64.500 285.000 ;
        RECT 89.700 282.600 90.600 289.950 ;
        RECT 94.950 289.050 97.050 292.050 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 91.950 288.000 97.050 289.050 ;
        RECT 101.100 288.150 102.900 289.950 ;
        RECT 91.950 287.550 96.450 288.000 ;
        RECT 91.950 286.950 96.000 287.550 ;
        RECT 104.700 284.700 105.900 289.950 ;
        RECT 106.950 288.150 108.750 289.950 ;
        RECT 113.550 289.050 114.450 292.950 ;
        RECT 122.100 292.050 123.900 293.850 ;
        RECT 126.000 292.050 126.900 297.600 ;
        RECT 133.950 294.450 138.000 295.050 ;
        RECT 127.950 292.050 129.750 293.850 ;
        RECT 133.950 292.950 138.450 294.450 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 113.550 287.550 118.050 289.050 ;
        RECT 119.100 288.150 120.900 289.950 ;
        RECT 114.000 286.950 118.050 287.550 ;
        RECT 81.000 276.000 82.800 282.600 ;
        RECT 85.500 281.400 90.600 282.600 ;
        RECT 101.700 283.800 105.900 284.700 ;
        RECT 85.500 276.600 87.300 281.400 ;
        RECT 88.500 276.000 90.300 279.600 ;
        RECT 101.700 276.600 103.500 283.800 ;
        RECT 125.700 282.600 126.900 289.950 ;
        RECT 130.950 288.150 132.750 289.950 ;
        RECT 137.550 289.050 138.450 292.950 ;
        RECT 143.100 292.050 144.900 293.850 ;
        RECT 146.100 292.050 147.300 305.400 ;
        RECT 161.100 292.050 162.900 293.850 ;
        RECT 164.100 292.050 165.300 305.400 ;
        RECT 180.000 305.100 180.900 305.400 ;
        RECT 185.100 305.400 186.900 311.400 ;
        RECT 188.100 305.400 189.900 312.000 ;
        RECT 185.100 305.100 186.600 305.400 ;
        RECT 180.000 304.200 186.600 305.100 ;
        RECT 180.000 292.050 180.900 304.200 ;
        RECT 203.100 299.400 204.900 311.400 ;
        RECT 206.100 299.400 207.900 312.000 ;
        RECT 218.100 305.400 219.900 311.400 ;
        RECT 185.100 292.050 186.900 293.850 ;
        RECT 203.700 292.050 204.900 299.400 ;
        RECT 218.100 298.500 219.300 305.400 ;
        RECT 221.100 301.200 222.900 312.000 ;
        RECT 224.100 299.400 225.900 311.400 ;
        RECT 236.100 305.400 237.900 312.000 ;
        RECT 239.100 305.400 240.900 311.400 ;
        RECT 242.100 306.000 243.900 312.000 ;
        RECT 239.400 305.100 240.900 305.400 ;
        RECT 245.100 305.400 246.900 311.400 ;
        RECT 245.100 305.100 246.000 305.400 ;
        RECT 239.400 304.200 246.000 305.100 ;
        RECT 218.100 297.600 223.800 298.500 ;
        RECT 222.000 296.700 223.800 297.600 ;
        RECT 218.400 292.050 220.200 293.850 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 160.950 289.950 163.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 218.400 289.950 220.500 292.050 ;
        RECT 133.950 287.550 138.450 289.050 ;
        RECT 133.950 286.950 138.000 287.550 ;
        RECT 106.800 276.000 108.600 282.600 ;
        RECT 121.500 276.000 123.300 282.600 ;
        RECT 126.000 276.600 127.800 282.600 ;
        RECT 130.500 276.000 132.300 282.600 ;
        RECT 146.100 279.600 147.300 289.950 ;
        RECT 164.100 279.600 165.300 289.950 ;
        RECT 180.000 286.200 180.900 289.950 ;
        RECT 182.100 288.150 183.900 289.950 ;
        RECT 188.100 288.150 189.900 289.950 ;
        RECT 193.950 288.450 196.050 289.050 ;
        RECT 199.950 288.450 202.050 289.050 ;
        RECT 193.950 287.550 202.050 288.450 ;
        RECT 193.950 286.950 196.050 287.550 ;
        RECT 199.950 286.950 202.050 287.550 ;
        RECT 180.000 285.000 183.300 286.200 ;
        RECT 143.100 276.000 144.900 279.600 ;
        RECT 146.100 276.600 147.900 279.600 ;
        RECT 161.100 276.000 162.900 279.600 ;
        RECT 164.100 276.600 165.900 279.600 ;
        RECT 181.500 276.600 183.300 285.000 ;
        RECT 188.100 276.000 189.900 285.600 ;
        RECT 203.700 282.600 204.900 289.950 ;
        RECT 206.100 288.150 207.900 289.950 ;
        RECT 222.000 285.300 222.900 296.700 ;
        RECT 224.700 292.050 225.900 299.400 ;
        RECT 239.100 292.050 240.900 293.850 ;
        RECT 245.100 292.050 246.000 304.200 ;
        RECT 257.100 299.400 258.900 311.400 ;
        RECT 260.100 299.400 261.900 312.000 ;
        RECT 272.100 301.500 273.900 311.400 ;
        RECT 275.100 302.400 276.900 312.000 ;
        RECT 278.100 310.500 285.900 311.400 ;
        RECT 278.100 301.500 279.900 310.500 ;
        RECT 272.100 300.600 279.900 301.500 ;
        RECT 281.100 301.800 282.900 309.600 ;
        RECT 284.100 302.700 285.900 310.500 ;
        RECT 287.100 310.500 294.900 311.400 ;
        RECT 287.100 301.800 288.900 310.500 ;
        RECT 281.100 300.900 288.900 301.800 ;
        RECT 290.100 301.800 291.900 309.600 ;
        RECT 257.700 292.050 258.900 299.400 ;
        RECT 262.950 294.450 267.000 295.050 ;
        RECT 262.950 292.950 267.450 294.450 ;
        RECT 223.800 289.950 225.900 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 222.000 284.400 223.800 285.300 ;
        RECT 218.100 283.500 223.800 284.400 ;
        RECT 203.100 276.600 204.900 282.600 ;
        RECT 206.100 276.000 207.900 282.600 ;
        RECT 218.100 279.600 219.300 283.500 ;
        RECT 224.700 282.600 225.900 289.950 ;
        RECT 236.100 288.150 237.900 289.950 ;
        RECT 242.100 288.150 243.900 289.950 ;
        RECT 245.100 286.200 246.000 289.950 ;
        RECT 218.100 276.600 219.900 279.600 ;
        RECT 221.100 276.000 222.900 282.600 ;
        RECT 224.100 276.600 225.900 282.600 ;
        RECT 236.100 276.000 237.900 285.600 ;
        RECT 242.700 285.000 246.000 286.200 ;
        RECT 242.700 276.600 244.500 285.000 ;
        RECT 257.700 282.600 258.900 289.950 ;
        RECT 260.100 288.150 261.900 289.950 ;
        RECT 266.550 289.050 267.450 292.950 ;
        RECT 275.100 292.050 276.900 293.850 ;
        RECT 284.250 292.050 286.050 293.850 ;
        RECT 290.100 292.050 291.300 301.800 ;
        RECT 293.100 301.200 294.900 310.500 ;
        RECT 308.700 305.400 310.500 312.000 ;
        RECT 309.000 302.100 310.800 303.900 ;
        RECT 311.700 300.900 313.500 311.400 ;
        RECT 311.100 299.400 313.500 300.900 ;
        RECT 316.800 299.400 318.600 312.000 ;
        RECT 332.400 299.400 334.200 312.000 ;
        RECT 337.500 300.900 339.300 311.400 ;
        RECT 340.500 305.400 342.300 312.000 ;
        RECT 340.200 302.100 342.000 303.900 ;
        RECT 337.500 299.400 339.900 300.900 ;
        RECT 356.100 300.300 357.900 311.400 ;
        RECT 359.100 301.200 360.900 312.000 ;
        RECT 362.100 300.300 363.900 311.400 ;
        RECT 356.100 299.400 363.900 300.300 ;
        RECT 365.100 299.400 366.900 311.400 ;
        RECT 380.100 305.400 381.900 312.000 ;
        RECT 383.100 305.400 384.900 311.400 ;
        RECT 398.100 305.400 399.900 312.000 ;
        RECT 401.100 305.400 402.900 311.400 ;
        RECT 404.100 305.400 405.900 312.000 ;
        RECT 419.100 305.400 420.900 312.000 ;
        RECT 422.100 305.400 423.900 311.400 ;
        RECT 425.100 305.400 426.900 312.000 ;
        RECT 440.100 305.400 441.900 312.000 ;
        RECT 443.100 305.400 444.900 311.400 ;
        RECT 446.100 305.400 447.900 312.000 ;
        RECT 458.700 305.400 460.500 312.000 ;
        RECT 311.100 292.050 312.300 299.400 ;
        RECT 328.950 294.450 331.050 295.050 ;
        RECT 317.100 292.050 318.900 293.850 ;
        RECT 323.550 293.550 331.050 294.450 ;
        RECT 274.800 289.950 276.900 292.050 ;
        RECT 280.950 289.950 283.050 292.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 289.500 289.950 291.600 292.050 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 262.950 287.550 267.450 289.050 ;
        RECT 280.950 288.150 282.750 289.950 ;
        RECT 262.950 286.950 267.000 287.550 ;
        RECT 257.100 276.600 258.900 282.600 ;
        RECT 260.100 276.000 261.900 282.600 ;
        RECT 290.100 281.400 291.300 289.950 ;
        RECT 308.100 288.150 309.900 289.950 ;
        RECT 311.100 285.600 312.300 289.950 ;
        RECT 314.100 288.150 315.900 289.950 ;
        RECT 323.550 289.050 324.450 293.550 ;
        RECT 328.950 292.950 331.050 293.550 ;
        RECT 332.100 292.050 333.900 293.850 ;
        RECT 338.700 292.050 339.900 299.400 ;
        RECT 349.950 297.450 352.050 298.050 ;
        RECT 355.950 297.450 358.050 298.050 ;
        RECT 349.950 296.550 358.050 297.450 ;
        RECT 349.950 295.950 352.050 296.550 ;
        RECT 355.950 295.950 358.050 296.550 ;
        RECT 359.250 292.050 361.050 293.850 ;
        RECT 365.700 292.050 366.600 299.400 ;
        RECT 379.950 297.450 382.050 298.050 ;
        RECT 371.550 296.550 382.050 297.450 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 319.950 287.550 324.450 289.050 ;
        RECT 335.100 288.150 336.900 289.950 ;
        RECT 319.950 286.950 324.000 287.550 ;
        RECT 308.700 284.700 312.300 285.600 ;
        RECT 338.700 285.600 339.900 289.950 ;
        RECT 341.100 288.150 342.900 289.950 ;
        RECT 356.100 288.150 357.900 289.950 ;
        RECT 362.250 288.150 364.050 289.950 ;
        RECT 338.700 284.700 342.300 285.600 ;
        RECT 308.700 282.600 309.900 284.700 ;
        RECT 278.700 280.500 291.300 281.400 ;
        RECT 278.700 279.600 279.600 280.500 ;
        RECT 285.900 279.600 286.800 280.500 ;
        RECT 274.800 276.000 276.900 279.600 ;
        RECT 278.100 276.600 279.900 279.600 ;
        RECT 281.100 276.000 282.900 279.600 ;
        RECT 284.100 276.600 286.800 279.600 ;
        RECT 308.100 276.600 309.900 282.600 ;
        RECT 311.100 281.700 318.900 283.050 ;
        RECT 311.100 276.600 312.900 281.700 ;
        RECT 314.100 276.000 315.900 280.800 ;
        RECT 317.100 276.600 318.900 281.700 ;
        RECT 332.100 281.700 339.900 283.050 ;
        RECT 332.100 276.600 333.900 281.700 ;
        RECT 335.100 276.000 336.900 280.800 ;
        RECT 338.100 276.600 339.900 281.700 ;
        RECT 341.100 282.600 342.300 284.700 ;
        RECT 365.700 282.600 366.600 289.950 ;
        RECT 371.550 285.900 372.450 296.550 ;
        RECT 379.950 295.950 382.050 296.550 ;
        RECT 380.100 292.050 381.900 293.850 ;
        RECT 383.100 292.050 384.300 305.400 ;
        RECT 401.100 292.050 402.300 305.400 ;
        RECT 422.100 292.050 423.300 305.400 ;
        RECT 424.950 303.450 427.050 304.050 ;
        RECT 433.950 303.450 436.050 304.050 ;
        RECT 424.950 302.550 436.050 303.450 ;
        RECT 424.950 301.950 427.050 302.550 ;
        RECT 433.950 301.950 436.050 302.550 ;
        RECT 443.700 292.050 444.900 305.400 ;
        RECT 459.000 302.100 460.800 303.900 ;
        RECT 461.700 300.900 463.500 311.400 ;
        RECT 461.100 299.400 463.500 300.900 ;
        RECT 466.800 299.400 468.600 312.000 ;
        RECT 479.100 305.400 480.900 311.400 ;
        RECT 482.100 305.400 483.900 312.000 ;
        RECT 494.100 310.500 501.900 311.400 ;
        RECT 461.100 292.050 462.300 299.400 ;
        RECT 467.100 292.050 468.900 293.850 ;
        RECT 479.700 292.050 480.900 305.400 ;
        RECT 494.100 299.400 495.900 310.500 ;
        RECT 497.100 298.500 498.900 309.600 ;
        RECT 500.100 300.600 501.900 310.500 ;
        RECT 503.100 301.500 504.900 312.000 ;
        RECT 506.100 300.600 507.900 311.400 ;
        RECT 518.100 305.400 519.900 311.400 ;
        RECT 521.100 306.000 522.900 312.000 ;
        RECT 500.100 299.700 507.900 300.600 ;
        RECT 519.000 305.100 519.900 305.400 ;
        RECT 524.100 305.400 525.900 311.400 ;
        RECT 527.100 305.400 528.900 312.000 ;
        RECT 524.100 305.100 525.600 305.400 ;
        RECT 519.000 304.200 525.600 305.100 ;
        RECT 497.100 297.600 501.900 298.500 ;
        RECT 482.100 292.050 483.900 293.850 ;
        RECT 497.100 292.050 498.900 293.850 ;
        RECT 501.000 292.050 501.900 297.600 ;
        RECT 502.950 292.050 504.750 293.850 ;
        RECT 519.000 292.050 519.900 304.200 ;
        RECT 542.100 300.600 543.900 311.400 ;
        RECT 545.100 301.500 546.900 312.000 ;
        RECT 548.100 310.500 555.900 311.400 ;
        RECT 548.100 300.600 549.900 310.500 ;
        RECT 542.100 299.700 549.900 300.600 ;
        RECT 551.100 298.500 552.900 309.600 ;
        RECT 554.100 299.400 555.900 310.500 ;
        RECT 569.100 305.400 570.900 312.000 ;
        RECT 572.100 305.400 573.900 311.400 ;
        RECT 575.100 305.400 576.900 312.000 ;
        RECT 587.100 305.400 588.900 312.000 ;
        RECT 590.100 305.400 591.900 311.400 ;
        RECT 593.100 305.400 594.900 312.000 ;
        RECT 548.100 297.600 552.900 298.500 ;
        RECT 524.100 292.050 525.900 293.850 ;
        RECT 545.250 292.050 547.050 293.850 ;
        RECT 548.100 292.050 549.000 297.600 ;
        RECT 564.000 294.450 568.050 295.050 ;
        RECT 551.100 292.050 552.900 293.850 ;
        RECT 563.550 292.950 568.050 294.450 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 493.950 289.950 496.050 292.050 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 499.950 289.950 502.050 292.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 517.950 289.950 520.050 292.050 ;
        RECT 520.950 289.950 523.050 292.050 ;
        RECT 523.950 289.950 526.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 370.950 283.800 373.050 285.900 ;
        RECT 341.100 276.600 342.900 282.600 ;
        RECT 357.000 276.000 358.800 282.600 ;
        RECT 361.500 281.400 366.600 282.600 ;
        RECT 361.500 276.600 363.300 281.400 ;
        RECT 383.100 279.600 384.300 289.950 ;
        RECT 398.250 288.150 400.050 289.950 ;
        RECT 401.100 284.700 402.300 289.950 ;
        RECT 404.100 288.150 405.900 289.950 ;
        RECT 419.250 288.150 421.050 289.950 ;
        RECT 422.100 284.700 423.300 289.950 ;
        RECT 425.100 288.150 426.900 289.950 ;
        RECT 440.100 288.150 441.900 289.950 ;
        RECT 443.700 284.700 444.900 289.950 ;
        RECT 445.950 288.150 447.750 289.950 ;
        RECT 458.100 288.150 459.900 289.950 ;
        RECT 461.100 285.600 462.300 289.950 ;
        RECT 464.100 288.150 465.900 289.950 ;
        RECT 401.100 283.800 405.300 284.700 ;
        RECT 422.100 283.800 426.300 284.700 ;
        RECT 364.500 276.000 366.300 279.600 ;
        RECT 380.100 276.000 381.900 279.600 ;
        RECT 383.100 276.600 384.900 279.600 ;
        RECT 398.400 276.000 400.200 282.600 ;
        RECT 403.500 276.600 405.300 283.800 ;
        RECT 419.400 276.000 421.200 282.600 ;
        RECT 424.500 276.600 426.300 283.800 ;
        RECT 440.700 283.800 444.900 284.700 ;
        RECT 458.700 284.700 462.300 285.600 ;
        RECT 440.700 276.600 442.500 283.800 ;
        RECT 458.700 282.600 459.900 284.700 ;
        RECT 445.800 276.000 447.600 282.600 ;
        RECT 458.100 276.600 459.900 282.600 ;
        RECT 461.100 281.700 468.900 283.050 ;
        RECT 461.100 276.600 462.900 281.700 ;
        RECT 464.100 276.000 465.900 280.800 ;
        RECT 467.100 276.600 468.900 281.700 ;
        RECT 479.700 279.600 480.900 289.950 ;
        RECT 494.100 288.150 495.900 289.950 ;
        RECT 500.700 282.600 501.900 289.950 ;
        RECT 505.950 288.150 507.750 289.950 ;
        RECT 519.000 286.200 519.900 289.950 ;
        RECT 521.100 288.150 522.900 289.950 ;
        RECT 527.100 288.150 528.900 289.950 ;
        RECT 542.250 288.150 544.050 289.950 ;
        RECT 519.000 285.000 522.300 286.200 ;
        RECT 479.100 276.600 480.900 279.600 ;
        RECT 482.100 276.000 483.900 279.600 ;
        RECT 496.500 276.000 498.300 282.600 ;
        RECT 501.000 276.600 502.800 282.600 ;
        RECT 505.500 276.000 507.300 282.600 ;
        RECT 520.500 276.600 522.300 285.000 ;
        RECT 527.100 276.000 528.900 285.600 ;
        RECT 548.100 282.600 549.300 289.950 ;
        RECT 554.100 288.150 555.900 289.950 ;
        RECT 556.950 288.450 559.050 289.050 ;
        RECT 563.550 288.450 564.450 292.950 ;
        RECT 572.100 292.050 573.300 305.400 ;
        RECT 590.700 292.050 591.900 305.400 ;
        RECT 608.100 300.300 609.900 311.400 ;
        RECT 611.100 301.500 612.900 312.000 ;
        RECT 615.600 300.300 617.400 311.400 ;
        RECT 619.800 301.500 621.900 312.000 ;
        RECT 623.100 300.600 624.900 311.400 ;
        RECT 635.100 305.400 636.900 312.000 ;
        RECT 638.100 305.400 639.900 311.400 ;
        RECT 641.100 305.400 642.900 312.000 ;
        RECT 608.100 299.100 612.900 300.300 ;
        RECT 615.600 299.400 618.900 300.300 ;
        RECT 610.800 298.200 612.900 299.100 ;
        RECT 610.800 297.300 616.200 298.200 ;
        RECT 614.400 295.500 616.200 297.300 ;
        RECT 617.700 295.050 618.900 299.400 ;
        RECT 619.800 299.400 624.900 300.600 ;
        RECT 619.800 298.500 621.900 299.400 ;
        RECT 617.100 294.300 619.200 295.050 ;
        RECT 612.900 292.200 614.700 294.000 ;
        RECT 616.200 292.950 619.200 294.300 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 586.950 289.950 589.050 292.050 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 556.950 287.550 564.450 288.450 ;
        RECT 569.250 288.150 571.050 289.950 ;
        RECT 556.950 286.950 559.050 287.550 ;
        RECT 572.100 284.700 573.300 289.950 ;
        RECT 575.100 288.150 576.900 289.950 ;
        RECT 587.100 288.150 588.900 289.950 ;
        RECT 590.700 284.700 591.900 289.950 ;
        RECT 592.950 288.150 594.750 289.950 ;
        RECT 608.100 289.800 610.200 292.050 ;
        RECT 612.900 290.100 615.000 292.200 ;
        RECT 608.400 289.200 610.200 289.800 ;
        RECT 608.400 288.000 615.000 289.200 ;
        RECT 612.900 287.100 615.000 288.000 ;
        RECT 610.500 285.000 612.600 285.600 ;
        RECT 613.500 285.300 615.300 287.100 ;
        RECT 616.200 286.200 617.100 292.950 ;
        RECT 622.800 292.050 624.600 293.850 ;
        RECT 638.100 292.050 639.300 305.400 ;
        RECT 656.100 299.400 657.900 311.400 ;
        RECT 660.600 299.400 662.400 312.000 ;
        RECT 663.600 300.900 665.400 311.400 ;
        RECT 663.600 299.400 666.000 300.900 ;
        RECT 680.100 299.400 681.900 312.000 ;
        RECT 685.200 300.600 687.000 311.400 ;
        RECT 701.100 305.400 702.900 312.000 ;
        RECT 704.100 305.400 705.900 311.400 ;
        RECT 707.100 305.400 708.900 312.000 ;
        RECT 683.400 299.400 687.000 300.600 ;
        RECT 656.100 297.900 657.300 299.400 ;
        RECT 656.100 296.700 663.900 297.900 ;
        RECT 662.100 296.100 663.900 296.700 ;
        RECT 660.000 292.050 661.800 293.850 ;
        RECT 618.000 290.100 619.800 291.900 ;
        RECT 618.000 288.000 620.100 290.100 ;
        RECT 622.800 289.950 624.900 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 656.100 289.950 658.200 292.050 ;
        RECT 659.400 289.950 661.500 292.050 ;
        RECT 635.250 288.150 637.050 289.950 ;
        RECT 572.100 283.800 576.300 284.700 ;
        RECT 542.700 276.000 544.500 282.600 ;
        RECT 547.200 276.600 549.000 282.600 ;
        RECT 551.700 276.000 553.500 282.600 ;
        RECT 569.400 276.000 571.200 282.600 ;
        RECT 574.500 276.600 576.300 283.800 ;
        RECT 587.700 283.800 591.900 284.700 ;
        RECT 587.700 276.600 589.500 283.800 ;
        RECT 608.100 283.500 612.600 285.000 ;
        RECT 616.200 284.100 619.200 286.200 ;
        RECT 608.100 282.600 609.600 283.500 ;
        RECT 592.800 276.000 594.600 282.600 ;
        RECT 608.100 276.600 609.900 282.600 ;
        RECT 616.200 282.000 617.100 284.100 ;
        RECT 620.400 283.500 622.500 285.900 ;
        RECT 638.100 284.700 639.300 289.950 ;
        RECT 641.100 288.150 642.900 289.950 ;
        RECT 656.400 288.150 658.200 289.950 ;
        RECT 662.700 285.600 663.600 296.100 ;
        RECT 664.800 292.050 666.000 299.400 ;
        RECT 680.250 292.050 682.050 293.850 ;
        RECT 683.400 292.050 684.300 299.400 ;
        RECT 686.100 292.050 687.900 293.850 ;
        RECT 704.700 292.050 705.900 305.400 ;
        RECT 722.100 299.400 723.900 311.400 ;
        RECT 725.100 300.000 726.900 312.000 ;
        RECT 728.100 305.400 729.900 311.400 ;
        RECT 731.100 305.400 732.900 312.000 ;
        RECT 746.100 305.400 747.900 312.000 ;
        RECT 749.100 305.400 750.900 311.400 ;
        RECT 752.100 305.400 753.900 312.000 ;
        RECT 722.700 292.050 723.600 299.400 ;
        RECT 726.000 292.050 727.800 293.850 ;
        RECT 664.800 289.950 666.900 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 722.100 289.950 724.200 292.050 ;
        RECT 725.400 289.950 727.500 292.050 ;
        RECT 662.700 284.700 664.800 285.600 ;
        RECT 638.100 283.800 642.300 284.700 ;
        RECT 620.400 282.600 624.900 283.500 ;
        RECT 611.100 276.000 612.900 281.700 ;
        RECT 615.300 276.600 617.100 282.000 ;
        RECT 619.800 276.000 621.600 281.700 ;
        RECT 623.100 276.600 624.900 282.600 ;
        RECT 635.400 276.000 637.200 282.600 ;
        RECT 640.500 276.600 642.300 283.800 ;
        RECT 659.400 283.800 664.800 284.700 ;
        RECT 659.400 279.600 660.300 283.800 ;
        RECT 666.000 282.600 666.900 289.950 ;
        RECT 656.100 276.600 657.900 279.600 ;
        RECT 659.100 276.600 660.900 279.600 ;
        RECT 656.100 276.000 657.300 276.600 ;
        RECT 662.100 276.000 663.900 282.000 ;
        RECT 665.100 276.600 666.900 282.600 ;
        RECT 683.400 279.600 684.300 289.950 ;
        RECT 701.100 288.150 702.900 289.950 ;
        RECT 685.950 285.450 688.050 286.050 ;
        RECT 691.950 285.450 694.050 286.050 ;
        RECT 685.950 284.550 694.050 285.450 ;
        RECT 704.700 284.700 705.900 289.950 ;
        RECT 706.950 288.150 708.750 289.950 ;
        RECT 685.950 283.950 688.050 284.550 ;
        RECT 691.950 283.950 694.050 284.550 ;
        RECT 701.700 283.800 705.900 284.700 ;
        RECT 680.100 276.000 681.900 279.600 ;
        RECT 683.100 276.600 684.900 279.600 ;
        RECT 686.100 276.000 687.900 279.600 ;
        RECT 701.700 276.600 703.500 283.800 ;
        RECT 722.700 282.600 723.600 289.950 ;
        RECT 729.000 285.300 729.900 305.400 ;
        RECT 749.700 292.050 750.900 305.400 ;
        RECT 764.100 300.300 765.900 311.400 ;
        RECT 767.100 301.500 768.900 312.000 ;
        RECT 771.600 300.300 773.400 311.400 ;
        RECT 775.800 301.500 777.900 312.000 ;
        RECT 779.100 300.600 780.900 311.400 ;
        RECT 791.700 305.400 793.500 312.000 ;
        RECT 792.000 302.100 793.800 303.900 ;
        RECT 794.700 300.900 796.500 311.400 ;
        RECT 764.100 299.100 768.900 300.300 ;
        RECT 771.600 299.400 774.900 300.300 ;
        RECT 766.800 298.200 768.900 299.100 ;
        RECT 766.800 297.300 772.200 298.200 ;
        RECT 770.400 295.500 772.200 297.300 ;
        RECT 773.700 295.050 774.900 299.400 ;
        RECT 775.800 299.400 780.900 300.600 ;
        RECT 794.100 299.400 796.500 300.900 ;
        RECT 799.800 299.400 801.600 312.000 ;
        RECT 815.100 300.300 816.900 311.400 ;
        RECT 818.100 301.500 819.900 312.000 ;
        RECT 822.600 300.300 824.400 311.400 ;
        RECT 826.800 301.500 828.900 312.000 ;
        RECT 830.100 300.600 831.900 311.400 ;
        RECT 775.800 298.500 777.900 299.400 ;
        RECT 773.100 294.300 775.200 295.050 ;
        RECT 768.900 292.200 770.700 294.000 ;
        RECT 772.200 292.950 775.200 294.300 ;
        RECT 730.800 289.950 732.900 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 748.950 289.950 751.050 292.050 ;
        RECT 751.950 289.950 754.050 292.050 ;
        RECT 730.950 288.150 732.750 289.950 ;
        RECT 746.100 288.150 747.900 289.950 ;
        RECT 724.500 284.400 732.900 285.300 ;
        RECT 749.700 284.700 750.900 289.950 ;
        RECT 751.950 288.150 753.750 289.950 ;
        RECT 764.100 289.800 766.200 292.050 ;
        RECT 768.900 290.100 771.000 292.200 ;
        RECT 764.400 289.200 766.200 289.800 ;
        RECT 764.400 288.000 771.000 289.200 ;
        RECT 768.900 287.100 771.000 288.000 ;
        RECT 766.500 285.000 768.600 285.600 ;
        RECT 769.500 285.300 771.300 287.100 ;
        RECT 772.200 286.200 773.100 292.950 ;
        RECT 778.800 292.050 780.600 293.850 ;
        RECT 794.100 292.050 795.300 299.400 ;
        RECT 815.100 299.100 819.900 300.300 ;
        RECT 822.600 299.400 825.900 300.300 ;
        RECT 817.800 298.200 819.900 299.100 ;
        RECT 817.800 297.300 823.200 298.200 ;
        RECT 821.400 295.500 823.200 297.300 ;
        RECT 824.700 295.050 825.900 299.400 ;
        RECT 826.800 299.400 831.900 300.600 ;
        RECT 845.100 300.600 846.900 311.400 ;
        RECT 848.100 301.500 849.900 312.000 ;
        RECT 845.100 299.400 849.900 300.600 ;
        RECT 826.800 298.500 828.900 299.400 ;
        RECT 847.800 298.500 849.900 299.400 ;
        RECT 852.600 299.400 854.400 311.400 ;
        RECT 857.100 301.500 858.900 312.000 ;
        RECT 860.100 300.300 861.900 311.400 ;
        RECT 857.400 299.400 861.900 300.300 ;
        RECT 875.100 299.400 876.900 311.400 ;
        RECT 878.100 300.300 879.900 311.400 ;
        RECT 881.100 301.200 882.900 312.000 ;
        RECT 884.100 300.300 885.900 311.400 ;
        RECT 878.100 299.400 885.900 300.300 ;
        RECT 897.000 300.600 898.800 311.400 ;
        RECT 897.000 299.400 900.600 300.600 ;
        RECT 902.100 299.400 903.900 312.000 ;
        RECT 914.700 305.400 916.500 312.000 ;
        RECT 915.000 302.100 916.800 303.900 ;
        RECT 917.700 300.900 919.500 311.400 ;
        RECT 917.100 299.400 919.500 300.900 ;
        RECT 922.800 299.400 924.600 312.000 ;
        RECT 935.100 305.400 936.900 312.000 ;
        RECT 938.100 305.400 939.900 311.400 ;
        RECT 941.100 305.400 942.900 312.000 ;
        RECT 852.600 298.050 853.800 299.400 ;
        RECT 852.300 297.000 853.800 298.050 ;
        RECT 857.400 297.300 859.500 299.400 ;
        RECT 852.300 295.050 853.200 297.000 ;
        RECT 824.100 294.300 826.200 295.050 ;
        RECT 800.100 292.050 801.900 293.850 ;
        RECT 819.900 292.200 821.700 294.000 ;
        RECT 823.200 292.950 826.200 294.300 ;
        RECT 774.000 290.100 775.800 291.900 ;
        RECT 774.000 288.000 776.100 290.100 ;
        RECT 778.800 289.950 780.900 292.050 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 791.100 288.150 792.900 289.950 ;
        RECT 724.500 283.500 726.300 284.400 ;
        RECT 706.800 276.000 708.600 282.600 ;
        RECT 722.700 280.800 725.400 282.600 ;
        RECT 723.600 276.600 725.400 280.800 ;
        RECT 726.600 276.000 728.400 282.600 ;
        RECT 731.100 276.600 732.900 284.400 ;
        RECT 746.700 283.800 750.900 284.700 ;
        RECT 746.700 276.600 748.500 283.800 ;
        RECT 764.100 283.500 768.600 285.000 ;
        RECT 772.200 284.100 775.200 286.200 ;
        RECT 764.100 282.600 765.600 283.500 ;
        RECT 751.800 276.000 753.600 282.600 ;
        RECT 764.100 276.600 765.900 282.600 ;
        RECT 772.200 282.000 773.100 284.100 ;
        RECT 776.400 283.500 778.500 285.900 ;
        RECT 794.100 285.600 795.300 289.950 ;
        RECT 797.100 288.150 798.900 289.950 ;
        RECT 815.100 289.800 817.200 292.050 ;
        RECT 819.900 290.100 822.000 292.200 ;
        RECT 815.400 289.200 817.200 289.800 ;
        RECT 802.950 288.450 805.050 289.050 ;
        RECT 808.950 288.450 811.050 289.050 ;
        RECT 802.950 287.550 811.050 288.450 ;
        RECT 815.400 288.000 822.000 289.200 ;
        RECT 802.950 286.950 805.050 287.550 ;
        RECT 808.950 286.950 811.050 287.550 ;
        RECT 819.900 287.100 822.000 288.000 ;
        RECT 791.700 284.700 795.300 285.600 ;
        RECT 817.500 285.000 819.600 285.600 ;
        RECT 820.500 285.300 822.300 287.100 ;
        RECT 823.200 286.200 824.100 292.950 ;
        RECT 829.800 292.050 831.600 293.850 ;
        RECT 845.400 292.050 847.200 293.850 ;
        RECT 851.100 292.950 853.200 295.050 ;
        RECT 854.100 295.500 856.200 295.800 ;
        RECT 854.100 293.700 858.000 295.500 ;
        RECT 825.000 290.100 826.800 291.900 ;
        RECT 825.000 288.000 827.100 290.100 ;
        RECT 829.800 289.950 831.900 292.050 ;
        RECT 845.100 289.950 847.200 292.050 ;
        RECT 851.700 292.800 853.200 292.950 ;
        RECT 851.700 291.900 854.100 292.800 ;
        RECT 849.900 289.200 851.700 291.000 ;
        RECT 849.900 287.100 852.000 289.200 ;
        RECT 852.900 286.200 854.100 291.900 ;
        RECT 855.000 292.050 856.800 292.500 ;
        RECT 875.400 292.050 876.300 299.400 ;
        RECT 877.950 297.450 880.050 298.050 ;
        RECT 889.950 297.450 892.050 298.050 ;
        RECT 895.950 297.450 898.050 298.050 ;
        RECT 877.950 296.550 898.050 297.450 ;
        RECT 877.950 295.950 880.050 296.550 ;
        RECT 889.950 295.950 892.050 296.550 ;
        RECT 895.950 295.950 898.050 296.550 ;
        RECT 880.950 292.050 882.750 293.850 ;
        RECT 896.100 292.050 897.900 293.850 ;
        RECT 899.700 292.050 900.600 299.400 ;
        RECT 912.000 297.450 916.050 298.050 ;
        RECT 911.550 295.950 916.050 297.450 ;
        RECT 911.550 294.450 912.450 295.950 ;
        RECT 901.950 292.050 903.750 293.850 ;
        RECT 908.550 293.550 912.450 294.450 ;
        RECT 855.000 290.700 861.900 292.050 ;
        RECT 859.800 289.950 861.900 290.700 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 898.950 289.950 901.050 292.050 ;
        RECT 901.950 289.950 904.050 292.050 ;
        RECT 776.400 282.600 780.900 283.500 ;
        RECT 791.700 282.600 792.900 284.700 ;
        RECT 815.100 283.500 819.600 285.000 ;
        RECT 823.200 284.100 826.200 286.200 ;
        RECT 767.100 276.000 768.900 281.700 ;
        RECT 771.300 276.600 773.100 282.000 ;
        RECT 775.800 276.000 777.600 281.700 ;
        RECT 779.100 276.600 780.900 282.600 ;
        RECT 791.100 276.600 792.900 282.600 ;
        RECT 794.100 281.700 801.900 283.050 ;
        RECT 794.100 276.600 795.900 281.700 ;
        RECT 797.100 276.000 798.900 280.800 ;
        RECT 800.100 276.600 801.900 281.700 ;
        RECT 815.100 282.600 816.600 283.500 ;
        RECT 815.100 276.600 816.900 282.600 ;
        RECT 823.200 282.000 824.100 284.100 ;
        RECT 827.400 283.500 829.500 285.900 ;
        RECT 847.800 283.500 849.900 284.700 ;
        RECT 851.100 284.100 854.100 286.200 ;
        RECT 855.000 287.400 856.800 289.200 ;
        RECT 859.800 288.150 861.600 289.950 ;
        RECT 855.000 285.300 857.100 287.400 ;
        RECT 855.000 284.400 861.300 285.300 ;
        RECT 827.400 282.600 831.900 283.500 ;
        RECT 818.100 276.000 819.900 281.700 ;
        RECT 822.300 276.600 824.100 282.000 ;
        RECT 826.800 276.000 828.600 281.700 ;
        RECT 830.100 276.600 831.900 282.600 ;
        RECT 845.100 282.600 849.900 283.500 ;
        RECT 852.900 282.600 854.100 284.100 ;
        RECT 860.100 282.600 861.300 284.400 ;
        RECT 875.400 282.600 876.300 289.950 ;
        RECT 877.950 288.150 879.750 289.950 ;
        RECT 884.100 288.150 885.900 289.950 ;
        RECT 845.100 276.600 846.900 282.600 ;
        RECT 848.100 276.000 849.900 281.700 ;
        RECT 852.600 276.600 854.400 282.600 ;
        RECT 857.100 276.000 858.900 281.700 ;
        RECT 860.100 276.600 861.900 282.600 ;
        RECT 875.400 281.400 880.500 282.600 ;
        RECT 875.700 276.000 877.500 279.600 ;
        RECT 878.700 276.600 880.500 281.400 ;
        RECT 883.200 276.000 885.000 282.600 ;
        RECT 899.700 279.600 900.600 289.950 ;
        RECT 908.550 289.050 909.450 293.550 ;
        RECT 917.100 292.050 918.300 299.400 ;
        RECT 919.950 297.450 922.050 298.200 ;
        RECT 919.950 296.550 927.450 297.450 ;
        RECT 919.950 296.100 922.050 296.550 ;
        RECT 926.550 294.450 927.450 296.550 ;
        RECT 923.100 292.050 924.900 293.850 ;
        RECT 926.550 293.550 930.450 294.450 ;
        RECT 913.950 289.950 916.050 292.050 ;
        RECT 916.950 289.950 919.050 292.050 ;
        RECT 919.950 289.950 922.050 292.050 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 904.950 287.550 909.450 289.050 ;
        RECT 914.100 288.150 915.900 289.950 ;
        RECT 904.950 286.950 909.000 287.550 ;
        RECT 917.100 285.600 918.300 289.950 ;
        RECT 920.100 288.150 921.900 289.950 ;
        RECT 929.550 289.050 930.450 293.550 ;
        RECT 938.700 292.050 939.900 305.400 ;
        RECT 934.950 289.950 937.050 292.050 ;
        RECT 937.950 289.950 940.050 292.050 ;
        RECT 940.950 289.950 943.050 292.050 ;
        RECT 925.950 287.550 930.450 289.050 ;
        RECT 935.100 288.150 936.900 289.950 ;
        RECT 925.950 286.950 930.000 287.550 ;
        RECT 914.700 284.700 918.300 285.600 ;
        RECT 938.700 284.700 939.900 289.950 ;
        RECT 940.950 288.150 942.750 289.950 ;
        RECT 914.700 282.600 915.900 284.700 ;
        RECT 935.700 283.800 939.900 284.700 ;
        RECT 896.100 276.000 897.900 279.600 ;
        RECT 899.100 276.600 900.900 279.600 ;
        RECT 902.100 276.000 903.900 279.600 ;
        RECT 914.100 276.600 915.900 282.600 ;
        RECT 917.100 281.700 924.900 283.050 ;
        RECT 917.100 276.600 918.900 281.700 ;
        RECT 920.100 276.000 921.900 280.800 ;
        RECT 923.100 276.600 924.900 281.700 ;
        RECT 935.700 276.600 937.500 283.800 ;
        RECT 940.800 276.000 942.600 282.600 ;
        RECT 15.000 266.400 16.800 273.000 ;
        RECT 19.500 267.600 21.300 272.400 ;
        RECT 22.500 269.400 24.300 273.000 ;
        RECT 19.500 266.400 24.600 267.600 ;
        RECT 14.100 259.050 15.900 260.850 ;
        RECT 20.250 259.050 22.050 260.850 ;
        RECT 23.700 259.050 24.600 266.400 ;
        RECT 35.100 267.300 36.900 272.400 ;
        RECT 38.100 268.200 39.900 273.000 ;
        RECT 41.100 267.300 42.900 272.400 ;
        RECT 35.100 265.950 42.900 267.300 ;
        RECT 44.100 266.400 45.900 272.400 ;
        RECT 44.100 264.300 45.300 266.400 ;
        RECT 41.700 263.400 45.300 264.300 ;
        RECT 59.100 263.400 60.900 273.000 ;
        RECT 65.700 264.000 67.500 272.400 ;
        RECT 80.100 266.400 81.900 272.400 ;
        RECT 83.100 267.000 84.900 273.000 ;
        RECT 89.700 272.400 90.900 273.000 ;
        RECT 86.100 269.400 87.900 272.400 ;
        RECT 89.100 269.400 90.900 272.400 ;
        RECT 25.950 261.450 30.000 262.050 ;
        RECT 25.950 259.950 30.450 261.450 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 17.250 255.150 19.050 256.950 ;
        RECT 23.700 249.600 24.600 256.950 ;
        RECT 29.550 256.050 30.450 259.950 ;
        RECT 38.100 259.050 39.900 260.850 ;
        RECT 41.700 259.050 42.900 263.400 ;
        RECT 65.700 262.800 69.000 264.000 ;
        RECT 44.100 259.050 45.900 260.850 ;
        RECT 59.100 259.050 60.900 260.850 ;
        RECT 65.100 259.050 66.900 260.850 ;
        RECT 68.100 259.050 69.000 262.800 ;
        RECT 80.100 259.050 81.000 266.400 ;
        RECT 86.700 265.200 87.600 269.400 ;
        RECT 104.100 266.400 105.900 272.400 ;
        RECT 82.200 264.300 87.600 265.200 ;
        RECT 104.700 264.300 105.900 266.400 ;
        RECT 107.100 267.300 108.900 272.400 ;
        RECT 110.100 268.200 111.900 273.000 ;
        RECT 113.100 267.300 114.900 272.400 ;
        RECT 128.100 269.400 129.900 272.400 ;
        RECT 131.100 269.400 132.900 273.000 ;
        RECT 146.100 269.400 147.900 273.000 ;
        RECT 149.100 269.400 150.900 272.400 ;
        RECT 107.100 265.950 114.900 267.300 ;
        RECT 82.200 263.400 84.300 264.300 ;
        RECT 104.700 263.400 108.300 264.300 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 80.100 256.950 82.200 259.050 ;
        RECT 25.950 254.550 30.450 256.050 ;
        RECT 35.100 255.150 36.900 256.950 ;
        RECT 25.950 253.950 30.000 254.550 ;
        RECT 41.700 249.600 42.900 256.950 ;
        RECT 62.100 255.150 63.900 256.950 ;
        RECT 58.950 252.450 61.050 253.050 ;
        RECT 64.950 252.450 67.050 252.750 ;
        RECT 58.950 251.550 67.050 252.450 ;
        RECT 58.950 250.950 61.050 251.550 ;
        RECT 64.950 250.650 67.050 251.550 ;
        RECT 14.100 248.700 21.900 249.600 ;
        RECT 14.100 237.600 15.900 248.700 ;
        RECT 17.100 237.000 18.900 247.800 ;
        RECT 20.100 237.600 21.900 248.700 ;
        RECT 23.100 237.600 24.900 249.600 ;
        RECT 35.400 237.000 37.200 249.600 ;
        RECT 40.500 248.100 42.900 249.600 ;
        RECT 40.500 237.600 42.300 248.100 ;
        RECT 43.200 245.100 45.000 246.900 ;
        RECT 68.100 244.800 69.000 256.950 ;
        RECT 81.000 249.600 82.200 256.950 ;
        RECT 83.400 252.900 84.300 263.400 ;
        RECT 88.800 259.050 90.600 260.850 ;
        RECT 104.100 259.050 105.900 260.850 ;
        RECT 107.100 259.050 108.300 263.400 ;
        RECT 110.100 259.050 111.900 260.850 ;
        RECT 128.700 259.050 129.900 269.400 ;
        RECT 149.100 259.050 150.300 269.400 ;
        RECT 161.100 267.300 162.900 272.400 ;
        RECT 164.100 268.200 165.900 273.000 ;
        RECT 167.100 267.300 168.900 272.400 ;
        RECT 161.100 265.950 168.900 267.300 ;
        RECT 170.100 266.400 171.900 272.400 ;
        RECT 182.100 266.400 183.900 272.400 ;
        RECT 170.100 264.300 171.300 266.400 ;
        RECT 167.700 263.400 171.300 264.300 ;
        RECT 182.700 264.300 183.900 266.400 ;
        RECT 185.100 267.300 186.900 272.400 ;
        RECT 188.100 268.200 189.900 273.000 ;
        RECT 191.100 267.300 192.900 272.400 ;
        RECT 206.100 269.400 207.900 273.000 ;
        RECT 209.100 269.400 210.900 272.400 ;
        RECT 185.100 265.950 192.900 267.300 ;
        RECT 182.700 263.400 186.300 264.300 ;
        RECT 164.100 259.050 165.900 260.850 ;
        RECT 167.700 259.050 168.900 263.400 ;
        RECT 170.100 259.050 171.900 260.850 ;
        RECT 182.100 259.050 183.900 260.850 ;
        RECT 185.100 259.050 186.300 263.400 ;
        RECT 193.950 261.450 198.000 262.050 ;
        RECT 188.100 259.050 189.900 260.850 ;
        RECT 193.950 259.950 198.450 261.450 ;
        RECT 85.500 256.950 87.600 259.050 ;
        RECT 88.800 256.950 90.900 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 85.200 255.150 87.000 256.950 ;
        RECT 83.100 252.300 84.900 252.900 ;
        RECT 83.100 251.100 90.900 252.300 ;
        RECT 89.700 249.600 90.900 251.100 ;
        RECT 81.000 248.100 83.400 249.600 ;
        RECT 62.400 243.900 69.000 244.800 ;
        RECT 62.400 243.600 63.900 243.900 ;
        RECT 43.500 237.000 45.300 243.600 ;
        RECT 59.100 237.000 60.900 243.600 ;
        RECT 62.100 237.600 63.900 243.600 ;
        RECT 68.100 243.600 69.000 243.900 ;
        RECT 65.100 237.000 66.900 243.000 ;
        RECT 68.100 237.600 69.900 243.600 ;
        RECT 81.600 237.600 83.400 248.100 ;
        RECT 84.600 237.000 86.400 249.600 ;
        RECT 89.100 237.600 90.900 249.600 ;
        RECT 107.100 249.600 108.300 256.950 ;
        RECT 113.100 255.150 114.900 256.950 ;
        RECT 107.100 248.100 109.500 249.600 ;
        RECT 105.000 245.100 106.800 246.900 ;
        RECT 104.700 237.000 106.500 243.600 ;
        RECT 107.700 237.600 109.500 248.100 ;
        RECT 112.800 237.000 114.600 249.600 ;
        RECT 128.700 243.600 129.900 256.950 ;
        RECT 131.100 255.150 132.900 256.950 ;
        RECT 146.100 255.150 147.900 256.950 ;
        RECT 149.100 243.600 150.300 256.950 ;
        RECT 161.100 255.150 162.900 256.950 ;
        RECT 167.700 249.600 168.900 256.950 ;
        RECT 128.100 237.600 129.900 243.600 ;
        RECT 131.100 237.000 132.900 243.600 ;
        RECT 146.100 237.000 147.900 243.600 ;
        RECT 149.100 237.600 150.900 243.600 ;
        RECT 161.400 237.000 163.200 249.600 ;
        RECT 166.500 248.100 168.900 249.600 ;
        RECT 185.100 249.600 186.300 256.950 ;
        RECT 191.100 255.150 192.900 256.950 ;
        RECT 197.550 255.450 198.450 259.950 ;
        RECT 209.100 259.050 210.300 269.400 ;
        RECT 224.400 266.400 226.200 273.000 ;
        RECT 229.500 265.200 231.300 272.400 ;
        RECT 242.100 269.400 243.900 273.000 ;
        RECT 245.100 269.400 246.900 272.400 ;
        RECT 248.100 269.400 249.900 273.000 ;
        RECT 227.100 264.300 231.300 265.200 ;
        RECT 219.000 261.450 223.050 262.050 ;
        RECT 218.550 259.950 223.050 261.450 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 194.550 254.550 198.450 255.450 ;
        RECT 206.100 255.150 207.900 256.950 ;
        RECT 194.550 253.050 195.450 254.550 ;
        RECT 190.950 251.550 195.450 253.050 ;
        RECT 190.950 250.950 195.000 251.550 ;
        RECT 185.100 248.100 187.500 249.600 ;
        RECT 166.500 237.600 168.300 248.100 ;
        RECT 169.200 245.100 171.000 246.900 ;
        RECT 183.000 245.100 184.800 246.900 ;
        RECT 169.500 237.000 171.300 243.600 ;
        RECT 182.700 237.000 184.500 243.600 ;
        RECT 185.700 237.600 187.500 248.100 ;
        RECT 190.800 237.000 192.600 249.600 ;
        RECT 209.100 243.600 210.300 256.950 ;
        RECT 218.550 256.050 219.450 259.950 ;
        RECT 224.250 259.050 226.050 260.850 ;
        RECT 227.100 259.050 228.300 264.300 ;
        RECT 230.100 259.050 231.900 260.850 ;
        RECT 245.400 259.050 246.300 269.400 ;
        RECT 263.700 265.200 265.500 272.400 ;
        RECT 268.800 266.400 270.600 273.000 ;
        RECT 285.600 268.200 287.400 272.400 ;
        RECT 284.700 266.400 287.400 268.200 ;
        RECT 288.600 266.400 290.400 273.000 ;
        RECT 247.950 264.450 250.050 265.050 ;
        RECT 256.950 264.450 259.050 265.050 ;
        RECT 247.950 263.550 259.050 264.450 ;
        RECT 263.700 264.300 267.900 265.200 ;
        RECT 247.950 262.950 250.050 263.550 ;
        RECT 256.950 262.950 259.050 263.550 ;
        RECT 258.000 261.450 262.050 262.050 ;
        RECT 257.550 259.950 262.050 261.450 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 241.950 256.950 244.050 259.050 ;
        RECT 244.950 256.950 247.050 259.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 218.550 254.550 223.050 256.050 ;
        RECT 219.000 253.950 223.050 254.550 ;
        RECT 227.100 243.600 228.300 256.950 ;
        RECT 242.250 255.150 244.050 256.950 ;
        RECT 245.400 249.600 246.300 256.950 ;
        RECT 248.100 255.150 249.900 256.950 ;
        RECT 257.550 256.050 258.450 259.950 ;
        RECT 263.100 259.050 264.900 260.850 ;
        RECT 266.700 259.050 267.900 264.300 ;
        RECT 268.950 259.050 270.750 260.850 ;
        RECT 284.700 259.050 285.600 266.400 ;
        RECT 286.500 264.600 288.300 265.500 ;
        RECT 293.100 264.600 294.900 272.400 ;
        RECT 308.100 269.400 309.900 273.000 ;
        RECT 311.100 269.400 312.900 272.400 ;
        RECT 323.700 269.400 325.500 273.000 ;
        RECT 286.500 263.700 294.900 264.600 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 265.950 256.950 268.050 259.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 284.100 256.950 286.200 259.050 ;
        RECT 287.400 256.950 289.500 259.050 ;
        RECT 257.550 254.550 262.050 256.050 ;
        RECT 258.000 253.950 262.050 254.550 ;
        RECT 206.100 237.000 207.900 243.600 ;
        RECT 209.100 237.600 210.900 243.600 ;
        RECT 224.100 237.000 225.900 243.600 ;
        RECT 227.100 237.600 228.900 243.600 ;
        RECT 230.100 237.000 231.900 243.600 ;
        RECT 242.100 237.000 243.900 249.600 ;
        RECT 245.400 248.400 249.000 249.600 ;
        RECT 247.200 237.600 249.000 248.400 ;
        RECT 266.700 243.600 267.900 256.950 ;
        RECT 284.700 249.600 285.600 256.950 ;
        RECT 288.000 255.150 289.800 256.950 ;
        RECT 263.100 237.000 264.900 243.600 ;
        RECT 266.100 237.600 267.900 243.600 ;
        RECT 269.100 237.000 270.900 243.600 ;
        RECT 284.100 237.600 285.900 249.600 ;
        RECT 287.100 237.000 288.900 249.000 ;
        RECT 291.000 243.600 291.900 263.700 ;
        RECT 292.950 259.050 294.750 260.850 ;
        RECT 311.100 259.050 312.300 269.400 ;
        RECT 326.700 267.600 328.500 272.400 ;
        RECT 323.400 266.400 328.500 267.600 ;
        RECT 331.200 266.400 333.000 273.000 ;
        RECT 323.400 259.050 324.300 266.400 ;
        RECT 349.500 264.000 351.300 272.400 ;
        RECT 348.000 262.800 351.300 264.000 ;
        RECT 356.100 263.400 357.900 273.000 ;
        RECT 371.100 269.400 372.900 272.400 ;
        RECT 371.100 265.500 372.300 269.400 ;
        RECT 374.100 266.400 375.900 273.000 ;
        RECT 377.100 266.400 378.900 272.400 ;
        RECT 393.600 268.200 395.400 272.400 ;
        RECT 371.100 264.600 376.800 265.500 ;
        RECT 375.000 263.700 376.800 264.600 ;
        RECT 325.950 259.050 327.750 260.850 ;
        RECT 332.100 259.050 333.900 260.850 ;
        RECT 348.000 259.050 348.900 262.800 ;
        RECT 350.100 259.050 351.900 260.850 ;
        RECT 356.100 259.050 357.900 260.850 ;
        RECT 292.800 256.950 294.900 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 371.400 256.950 373.500 259.050 ;
        RECT 308.100 255.150 309.900 256.950 ;
        RECT 311.100 243.600 312.300 256.950 ;
        RECT 323.400 249.600 324.300 256.950 ;
        RECT 328.950 255.150 330.750 256.950 ;
        RECT 325.950 252.450 328.050 253.050 ;
        RECT 340.950 252.450 343.050 253.050 ;
        RECT 325.950 251.550 343.050 252.450 ;
        RECT 325.950 250.950 328.050 251.550 ;
        RECT 340.950 250.950 343.050 251.550 ;
        RECT 290.100 237.600 291.900 243.600 ;
        RECT 293.100 237.000 294.900 243.600 ;
        RECT 298.950 240.450 301.050 240.900 ;
        RECT 304.950 240.450 307.050 241.050 ;
        RECT 298.950 239.550 307.050 240.450 ;
        RECT 298.950 238.800 301.050 239.550 ;
        RECT 304.950 238.950 307.050 239.550 ;
        RECT 308.100 237.000 309.900 243.600 ;
        RECT 311.100 237.600 312.900 243.600 ;
        RECT 323.100 237.600 324.900 249.600 ;
        RECT 326.100 248.700 333.900 249.600 ;
        RECT 326.100 237.600 327.900 248.700 ;
        RECT 329.100 237.000 330.900 247.800 ;
        RECT 332.100 237.600 333.900 248.700 ;
        RECT 348.000 244.800 348.900 256.950 ;
        RECT 353.100 255.150 354.900 256.950 ;
        RECT 371.400 255.150 373.200 256.950 ;
        RECT 375.000 252.300 375.900 263.700 ;
        RECT 377.700 259.050 378.900 266.400 ;
        RECT 392.700 266.400 395.400 268.200 ;
        RECT 396.600 266.400 398.400 273.000 ;
        RECT 392.700 259.050 393.600 266.400 ;
        RECT 394.500 264.600 396.300 265.500 ;
        RECT 401.100 264.600 402.900 272.400 ;
        RECT 416.100 269.400 417.900 272.400 ;
        RECT 419.100 269.400 420.900 273.000 ;
        RECT 394.500 263.700 402.900 264.600 ;
        RECT 376.800 256.950 378.900 259.050 ;
        RECT 392.100 256.950 394.200 259.050 ;
        RECT 395.400 256.950 397.500 259.050 ;
        RECT 375.000 251.400 376.800 252.300 ;
        RECT 371.100 250.500 376.800 251.400 ;
        RECT 348.000 243.900 354.600 244.800 ;
        RECT 348.000 243.600 348.900 243.900 ;
        RECT 347.100 237.600 348.900 243.600 ;
        RECT 353.100 243.600 354.600 243.900 ;
        RECT 371.100 243.600 372.300 250.500 ;
        RECT 377.700 249.600 378.900 256.950 ;
        RECT 392.700 249.600 393.600 256.950 ;
        RECT 396.000 255.150 397.800 256.950 ;
        RECT 350.100 237.000 351.900 243.000 ;
        RECT 353.100 237.600 354.900 243.600 ;
        RECT 356.100 237.000 357.900 243.600 ;
        RECT 371.100 237.600 372.900 243.600 ;
        RECT 374.100 237.000 375.900 247.800 ;
        RECT 377.100 237.600 378.900 249.600 ;
        RECT 392.100 237.600 393.900 249.600 ;
        RECT 395.100 237.000 396.900 249.000 ;
        RECT 399.000 243.600 399.900 263.700 ;
        RECT 400.950 259.050 402.750 260.850 ;
        RECT 416.700 259.050 417.900 269.400 ;
        RECT 435.600 268.200 437.400 272.400 ;
        RECT 434.700 266.400 437.400 268.200 ;
        RECT 438.600 266.400 440.400 273.000 ;
        RECT 434.700 259.050 435.600 266.400 ;
        RECT 436.500 264.600 438.300 265.500 ;
        RECT 443.100 264.600 444.900 272.400 ;
        RECT 458.100 269.400 459.900 273.000 ;
        RECT 461.100 269.400 462.900 272.400 ;
        RECT 464.100 269.400 465.900 273.000 ;
        RECT 436.500 263.700 444.900 264.600 ;
        RECT 400.800 256.950 402.900 259.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 434.100 256.950 436.200 259.050 ;
        RECT 437.400 256.950 439.500 259.050 ;
        RECT 416.700 243.600 417.900 256.950 ;
        RECT 419.100 255.150 420.900 256.950 ;
        RECT 434.700 249.600 435.600 256.950 ;
        RECT 438.000 255.150 439.800 256.950 ;
        RECT 398.100 237.600 399.900 243.600 ;
        RECT 401.100 237.000 402.900 243.600 ;
        RECT 416.100 237.600 417.900 243.600 ;
        RECT 419.100 237.000 420.900 243.600 ;
        RECT 434.100 237.600 435.900 249.600 ;
        RECT 437.100 237.000 438.900 249.000 ;
        RECT 441.000 243.600 441.900 263.700 ;
        RECT 442.950 259.050 444.750 260.850 ;
        RECT 461.400 259.050 462.300 269.400 ;
        RECT 476.700 266.400 478.500 273.000 ;
        RECT 481.200 266.400 483.000 272.400 ;
        RECT 485.700 266.400 487.500 273.000 ;
        RECT 500.400 266.400 502.200 273.000 ;
        RECT 476.250 259.050 478.050 260.850 ;
        RECT 482.100 259.050 483.300 266.400 ;
        RECT 505.500 265.200 507.300 272.400 ;
        RECT 503.100 264.300 507.300 265.200 ;
        RECT 521.700 265.200 523.500 272.400 ;
        RECT 526.800 266.400 528.600 273.000 ;
        RECT 542.100 269.400 543.900 273.000 ;
        RECT 545.100 269.400 546.900 272.400 ;
        RECT 521.700 264.300 525.900 265.200 ;
        RECT 488.100 259.050 489.900 260.850 ;
        RECT 500.250 259.050 502.050 260.850 ;
        RECT 503.100 259.050 504.300 264.300 ;
        RECT 506.100 259.050 507.900 260.850 ;
        RECT 521.100 259.050 522.900 260.850 ;
        RECT 524.700 259.050 525.900 264.300 ;
        RECT 526.950 259.050 528.750 260.850 ;
        RECT 545.100 259.050 546.300 269.400 ;
        RECT 560.700 265.200 562.500 272.400 ;
        RECT 565.800 266.400 567.600 273.000 ;
        RECT 581.100 269.400 582.900 273.000 ;
        RECT 584.100 269.400 585.900 272.400 ;
        RECT 587.100 269.400 588.900 273.000 ;
        RECT 560.700 264.300 564.900 265.200 ;
        RECT 560.100 259.050 561.900 260.850 ;
        RECT 563.700 259.050 564.900 264.300 ;
        RECT 576.000 261.450 580.050 262.050 ;
        RECT 565.950 259.050 567.750 260.850 ;
        RECT 575.550 259.950 580.050 261.450 ;
        RECT 575.550 259.050 576.450 259.950 ;
        RECT 584.400 259.050 585.300 269.400 ;
        RECT 602.100 267.300 603.900 272.400 ;
        RECT 605.100 268.200 606.900 273.000 ;
        RECT 608.100 267.300 609.900 272.400 ;
        RECT 602.100 265.950 609.900 267.300 ;
        RECT 611.100 266.400 612.900 272.400 ;
        RECT 626.100 266.400 627.900 272.400 ;
        RECT 629.100 267.300 630.900 273.000 ;
        RECT 633.600 266.400 635.400 272.400 ;
        RECT 638.100 267.300 639.900 273.000 ;
        RECT 641.100 266.400 642.900 272.400 ;
        RECT 611.100 264.300 612.300 266.400 ;
        RECT 608.700 263.400 612.300 264.300 ;
        RECT 626.700 264.600 627.900 266.400 ;
        RECT 633.900 264.900 635.100 266.400 ;
        RECT 638.100 265.500 642.900 266.400 ;
        RECT 626.700 263.700 633.000 264.600 ;
        RECT 605.100 259.050 606.900 260.850 ;
        RECT 608.700 259.050 609.900 263.400 ;
        RECT 630.900 261.600 633.000 263.700 ;
        RECT 611.100 259.050 612.900 260.850 ;
        RECT 626.400 259.050 628.200 260.850 ;
        RECT 631.200 259.800 633.000 261.600 ;
        RECT 633.900 262.800 636.900 264.900 ;
        RECT 638.100 264.300 640.200 265.500 ;
        RECT 653.700 265.200 655.500 272.400 ;
        RECT 658.800 266.400 660.600 273.000 ;
        RECT 674.100 269.400 675.900 273.000 ;
        RECT 677.100 269.400 678.900 272.400 ;
        RECT 680.100 269.400 681.900 273.000 ;
        RECT 653.700 264.300 657.900 265.200 ;
        RECT 442.800 256.950 444.900 259.050 ;
        RECT 457.950 256.950 460.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 565.950 256.950 568.050 259.050 ;
        RECT 573.000 258.900 576.450 259.050 ;
        RECT 571.950 257.550 576.450 258.900 ;
        RECT 571.950 256.950 576.000 257.550 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 626.100 258.300 628.200 259.050 ;
        RECT 626.100 256.950 633.000 258.300 ;
        RECT 458.250 255.150 460.050 256.950 ;
        RECT 461.400 249.600 462.300 256.950 ;
        RECT 464.100 255.150 465.900 256.950 ;
        RECT 479.250 255.150 481.050 256.950 ;
        RECT 482.100 251.400 483.000 256.950 ;
        RECT 485.100 255.150 486.900 256.950 ;
        RECT 482.100 250.500 486.900 251.400 ;
        RECT 440.100 237.600 441.900 243.600 ;
        RECT 443.100 237.000 444.900 243.600 ;
        RECT 458.100 237.000 459.900 249.600 ;
        RECT 461.400 248.400 465.000 249.600 ;
        RECT 463.200 237.600 465.000 248.400 ;
        RECT 476.100 248.400 483.900 249.300 ;
        RECT 476.100 237.600 477.900 248.400 ;
        RECT 479.100 237.000 480.900 247.500 ;
        RECT 482.100 238.500 483.900 248.400 ;
        RECT 485.100 239.400 486.900 250.500 ;
        RECT 488.100 238.500 489.900 249.600 ;
        RECT 503.100 243.600 504.300 256.950 ;
        RECT 524.700 243.600 525.900 256.950 ;
        RECT 542.100 255.150 543.900 256.950 ;
        RECT 545.100 243.600 546.300 256.950 ;
        RECT 547.950 252.450 550.050 253.050 ;
        RECT 559.950 252.450 562.050 253.050 ;
        RECT 547.950 251.550 562.050 252.450 ;
        RECT 547.950 250.950 550.050 251.550 ;
        RECT 559.950 250.950 562.050 251.550 ;
        RECT 563.700 243.600 564.900 256.950 ;
        RECT 571.950 256.800 574.050 256.950 ;
        RECT 581.250 255.150 583.050 256.950 ;
        RECT 584.400 249.600 585.300 256.950 ;
        RECT 587.100 255.150 588.900 256.950 ;
        RECT 602.100 255.150 603.900 256.950 ;
        RECT 608.700 249.600 609.900 256.950 ;
        RECT 631.200 256.500 633.000 256.950 ;
        RECT 633.900 257.100 635.100 262.800 ;
        RECT 636.000 259.800 638.100 261.900 ;
        RECT 636.300 258.000 638.100 259.800 ;
        RECT 653.100 259.050 654.900 260.850 ;
        RECT 656.700 259.050 657.900 264.300 ;
        RECT 664.950 264.450 667.050 265.050 ;
        RECT 673.950 264.450 676.050 265.050 ;
        RECT 664.950 263.550 676.050 264.450 ;
        RECT 664.950 262.950 667.050 263.550 ;
        RECT 673.950 262.950 676.050 263.550 ;
        RECT 658.950 259.050 660.750 260.850 ;
        RECT 677.700 259.050 678.600 269.400 ;
        RECT 692.400 266.400 694.200 273.000 ;
        RECT 697.500 265.200 699.300 272.400 ;
        RECT 713.100 267.300 714.900 272.400 ;
        RECT 716.100 268.200 717.900 273.000 ;
        RECT 719.100 267.300 720.900 272.400 ;
        RECT 713.100 265.950 720.900 267.300 ;
        RECT 722.100 266.400 723.900 272.400 ;
        RECT 734.700 266.400 736.500 273.000 ;
        RECT 739.200 266.400 741.000 272.400 ;
        RECT 743.700 266.400 745.500 273.000 ;
        RECT 695.100 264.300 699.300 265.200 ;
        RECT 722.100 264.300 723.300 266.400 ;
        RECT 692.250 259.050 694.050 260.850 ;
        RECT 695.100 259.050 696.300 264.300 ;
        RECT 719.700 263.400 723.300 264.300 ;
        RECT 724.950 264.450 727.050 265.050 ;
        RECT 736.950 264.450 739.050 265.050 ;
        RECT 724.950 263.550 739.050 264.450 ;
        RECT 698.100 259.050 699.900 260.850 ;
        RECT 716.100 259.050 717.900 260.850 ;
        RECT 719.700 259.050 720.900 263.400 ;
        RECT 724.950 262.950 727.050 263.550 ;
        RECT 736.950 262.950 739.050 263.550 ;
        RECT 722.100 259.050 723.900 260.850 ;
        RECT 734.250 259.050 736.050 260.850 ;
        RECT 740.100 259.050 741.300 266.400 ;
        RECT 758.100 263.400 759.900 273.000 ;
        RECT 764.700 264.000 766.500 272.400 ;
        RECT 780.000 266.400 781.800 273.000 ;
        RECT 784.500 267.600 786.300 272.400 ;
        RECT 787.500 269.400 789.300 273.000 ;
        RECT 784.500 266.400 789.600 267.600 ;
        RECT 800.100 266.400 801.900 272.400 ;
        RECT 764.700 262.800 768.000 264.000 ;
        RECT 746.100 259.050 747.900 260.850 ;
        RECT 758.100 259.050 759.900 260.850 ;
        RECT 764.100 259.050 765.900 260.850 ;
        RECT 767.100 259.050 768.000 262.800 ;
        RECT 779.100 259.050 780.900 260.850 ;
        RECT 785.250 259.050 787.050 260.850 ;
        RECT 788.700 259.050 789.600 266.400 ;
        RECT 800.700 264.300 801.900 266.400 ;
        RECT 803.100 267.300 804.900 272.400 ;
        RECT 806.100 268.200 807.900 273.000 ;
        RECT 809.100 267.300 810.900 272.400 ;
        RECT 803.100 265.950 810.900 267.300 ;
        RECT 824.100 267.300 825.900 272.400 ;
        RECT 827.100 268.200 828.900 273.000 ;
        RECT 830.100 267.300 831.900 272.400 ;
        RECT 824.100 265.950 831.900 267.300 ;
        RECT 833.100 266.400 834.900 272.400 ;
        RECT 848.700 269.400 850.500 273.000 ;
        RECT 851.700 267.600 853.500 272.400 ;
        RECT 848.400 266.400 853.500 267.600 ;
        RECT 856.200 266.400 858.000 273.000 ;
        RECT 873.000 266.400 874.800 273.000 ;
        RECT 877.500 267.600 879.300 272.400 ;
        RECT 880.500 269.400 882.300 273.000 ;
        RECT 877.500 266.400 882.600 267.600 ;
        RECT 833.100 264.300 834.300 266.400 ;
        RECT 800.700 263.400 804.300 264.300 ;
        RECT 800.100 259.050 801.900 260.850 ;
        RECT 803.100 259.050 804.300 263.400 ;
        RECT 830.700 263.400 834.300 264.300 ;
        RECT 814.950 261.450 817.050 262.050 ;
        RECT 820.950 261.450 823.050 262.050 ;
        RECT 806.100 259.050 807.900 260.850 ;
        RECT 814.950 260.550 823.050 261.450 ;
        RECT 814.950 259.950 817.050 260.550 ;
        RECT 820.950 259.950 823.050 260.550 ;
        RECT 827.100 259.050 828.900 260.850 ;
        RECT 830.700 259.050 831.900 263.400 ;
        RECT 833.100 259.050 834.900 260.850 ;
        RECT 848.400 259.050 849.300 266.400 ;
        RECT 853.950 264.450 856.050 265.050 ;
        RECT 862.950 264.450 865.050 265.050 ;
        RECT 853.950 263.550 865.050 264.450 ;
        RECT 853.950 262.950 856.050 263.550 ;
        RECT 862.950 262.950 865.050 263.550 ;
        RECT 850.950 259.050 852.750 260.850 ;
        RECT 857.100 259.050 858.900 260.850 ;
        RECT 872.100 259.050 873.900 260.850 ;
        RECT 878.250 259.050 880.050 260.850 ;
        RECT 881.700 259.050 882.600 266.400 ;
        RECT 896.100 263.400 897.900 273.000 ;
        RECT 902.700 264.000 904.500 272.400 ;
        RECT 922.500 264.000 924.300 272.400 ;
        RECT 902.700 262.800 906.000 264.000 ;
        RECT 896.100 259.050 897.900 260.850 ;
        RECT 902.100 259.050 903.900 260.850 ;
        RECT 905.100 259.050 906.000 262.800 ;
        RECT 921.000 262.800 924.300 264.000 ;
        RECT 929.100 263.400 930.900 273.000 ;
        RECT 941.100 269.400 942.900 272.400 ;
        RECT 944.100 269.400 945.900 273.000 ;
        RECT 910.950 259.950 913.050 262.050 ;
        RECT 915.000 261.450 919.050 262.050 ;
        RECT 914.550 259.950 919.050 261.450 ;
        RECT 633.900 256.200 636.300 257.100 ;
        RECT 634.800 256.050 636.300 256.200 ;
        RECT 640.800 256.950 642.900 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 736.950 256.950 739.050 259.050 ;
        RECT 739.950 256.950 742.050 259.050 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 745.950 256.950 748.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 880.950 256.950 883.050 259.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 901.950 256.950 904.050 259.050 ;
        RECT 904.950 256.950 907.050 259.050 ;
        RECT 630.000 253.500 633.900 255.300 ;
        RECT 631.800 253.200 633.900 253.500 ;
        RECT 634.800 253.950 636.900 256.050 ;
        RECT 640.800 255.150 642.600 256.950 ;
        RECT 634.800 252.000 635.700 253.950 ;
        RECT 628.500 249.600 630.600 251.700 ;
        RECT 634.200 250.950 635.700 252.000 ;
        RECT 634.200 249.600 635.400 250.950 ;
        RECT 482.100 237.600 489.900 238.500 ;
        RECT 500.100 237.000 501.900 243.600 ;
        RECT 503.100 237.600 504.900 243.600 ;
        RECT 506.100 237.000 507.900 243.600 ;
        RECT 521.100 237.000 522.900 243.600 ;
        RECT 524.100 237.600 525.900 243.600 ;
        RECT 527.100 237.000 528.900 243.600 ;
        RECT 542.100 237.000 543.900 243.600 ;
        RECT 545.100 237.600 546.900 243.600 ;
        RECT 560.100 237.000 561.900 243.600 ;
        RECT 563.100 237.600 564.900 243.600 ;
        RECT 566.100 237.000 567.900 243.600 ;
        RECT 581.100 237.000 582.900 249.600 ;
        RECT 584.400 248.400 588.000 249.600 ;
        RECT 586.200 237.600 588.000 248.400 ;
        RECT 602.400 237.000 604.200 249.600 ;
        RECT 607.500 248.100 609.900 249.600 ;
        RECT 626.100 248.700 630.600 249.600 ;
        RECT 607.500 237.600 609.300 248.100 ;
        RECT 610.200 245.100 612.000 246.900 ;
        RECT 610.500 237.000 612.300 243.600 ;
        RECT 626.100 237.600 627.900 248.700 ;
        RECT 629.100 237.000 630.900 247.500 ;
        RECT 633.600 237.600 635.400 249.600 ;
        RECT 638.100 249.600 640.200 250.500 ;
        RECT 638.100 248.400 642.900 249.600 ;
        RECT 638.100 237.000 639.900 247.500 ;
        RECT 641.100 237.600 642.900 248.400 ;
        RECT 656.700 243.600 657.900 256.950 ;
        RECT 674.100 255.150 675.900 256.950 ;
        RECT 677.700 249.600 678.600 256.950 ;
        RECT 679.950 255.150 681.750 256.950 ;
        RECT 685.950 252.450 688.050 253.050 ;
        RECT 691.950 252.450 694.050 253.050 ;
        RECT 685.950 251.550 694.050 252.450 ;
        RECT 685.950 250.950 688.050 251.550 ;
        RECT 691.950 250.950 694.050 251.550 ;
        RECT 675.000 248.400 678.600 249.600 ;
        RECT 653.100 237.000 654.900 243.600 ;
        RECT 656.100 237.600 657.900 243.600 ;
        RECT 659.100 237.000 660.900 243.600 ;
        RECT 675.000 237.600 676.800 248.400 ;
        RECT 680.100 237.000 681.900 249.600 ;
        RECT 695.100 243.600 696.300 256.950 ;
        RECT 713.100 255.150 714.900 256.950 ;
        RECT 719.700 249.600 720.900 256.950 ;
        RECT 737.250 255.150 739.050 256.950 ;
        RECT 740.100 251.400 741.000 256.950 ;
        RECT 743.100 255.150 744.900 256.950 ;
        RECT 761.100 255.150 762.900 256.950 ;
        RECT 740.100 250.500 744.900 251.400 ;
        RECT 692.100 237.000 693.900 243.600 ;
        RECT 695.100 237.600 696.900 243.600 ;
        RECT 698.100 237.000 699.900 243.600 ;
        RECT 713.400 237.000 715.200 249.600 ;
        RECT 718.500 248.100 720.900 249.600 ;
        RECT 734.100 248.400 741.900 249.300 ;
        RECT 718.500 237.600 720.300 248.100 ;
        RECT 721.200 245.100 723.000 246.900 ;
        RECT 721.500 237.000 723.300 243.600 ;
        RECT 734.100 237.600 735.900 248.400 ;
        RECT 737.100 237.000 738.900 247.500 ;
        RECT 740.100 238.500 741.900 248.400 ;
        RECT 743.100 239.400 744.900 250.500 ;
        RECT 746.100 238.500 747.900 249.600 ;
        RECT 767.100 244.800 768.000 256.950 ;
        RECT 782.250 255.150 784.050 256.950 ;
        RECT 788.700 249.600 789.600 256.950 ;
        RECT 803.100 249.600 804.300 256.950 ;
        RECT 809.100 255.150 810.900 256.950 ;
        RECT 824.100 255.150 825.900 256.950 ;
        RECT 830.700 249.600 831.900 256.950 ;
        RECT 832.950 252.450 835.050 252.750 ;
        RECT 841.950 252.450 844.050 253.050 ;
        RECT 832.950 251.550 844.050 252.450 ;
        RECT 832.950 250.650 835.050 251.550 ;
        RECT 841.950 250.950 844.050 251.550 ;
        RECT 848.400 249.600 849.300 256.950 ;
        RECT 853.950 255.150 855.750 256.950 ;
        RECT 875.250 255.150 877.050 256.950 ;
        RECT 881.700 249.600 882.600 256.950 ;
        RECT 899.100 255.150 900.900 256.950 ;
        RECT 761.400 243.900 768.000 244.800 ;
        RECT 761.400 243.600 762.900 243.900 ;
        RECT 740.100 237.600 747.900 238.500 ;
        RECT 758.100 237.000 759.900 243.600 ;
        RECT 761.100 237.600 762.900 243.600 ;
        RECT 767.100 243.600 768.000 243.900 ;
        RECT 779.100 248.700 786.900 249.600 ;
        RECT 764.100 237.000 765.900 243.000 ;
        RECT 767.100 237.600 768.900 243.600 ;
        RECT 779.100 237.600 780.900 248.700 ;
        RECT 782.100 237.000 783.900 247.800 ;
        RECT 785.100 237.600 786.900 248.700 ;
        RECT 788.100 237.600 789.900 249.600 ;
        RECT 803.100 248.100 805.500 249.600 ;
        RECT 801.000 245.100 802.800 246.900 ;
        RECT 800.700 237.000 802.500 243.600 ;
        RECT 803.700 237.600 805.500 248.100 ;
        RECT 808.800 237.000 810.600 249.600 ;
        RECT 824.400 237.000 826.200 249.600 ;
        RECT 829.500 248.100 831.900 249.600 ;
        RECT 829.500 237.600 831.300 248.100 ;
        RECT 832.200 245.100 834.000 246.900 ;
        RECT 832.500 237.000 834.300 243.600 ;
        RECT 848.100 237.600 849.900 249.600 ;
        RECT 851.100 248.700 858.900 249.600 ;
        RECT 851.100 237.600 852.900 248.700 ;
        RECT 854.100 237.000 855.900 247.800 ;
        RECT 857.100 237.600 858.900 248.700 ;
        RECT 872.100 248.700 879.900 249.600 ;
        RECT 872.100 237.600 873.900 248.700 ;
        RECT 875.100 237.000 876.900 247.800 ;
        RECT 878.100 237.600 879.900 248.700 ;
        RECT 881.100 237.600 882.900 249.600 ;
        RECT 883.950 249.450 886.050 250.050 ;
        RECT 901.950 249.450 904.050 250.050 ;
        RECT 883.950 248.550 904.050 249.450 ;
        RECT 883.950 247.950 886.050 248.550 ;
        RECT 901.950 247.950 904.050 248.550 ;
        RECT 905.100 244.800 906.000 256.950 ;
        RECT 911.550 256.050 912.450 259.950 ;
        RECT 907.950 254.550 912.450 256.050 ;
        RECT 914.550 256.050 915.450 259.950 ;
        RECT 921.000 259.050 921.900 262.800 ;
        RECT 936.000 261.450 940.050 262.050 ;
        RECT 923.100 259.050 924.900 260.850 ;
        RECT 929.100 259.050 930.900 260.850 ;
        RECT 935.550 259.950 940.050 261.450 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 922.950 256.950 925.050 259.050 ;
        RECT 925.950 256.950 928.050 259.050 ;
        RECT 928.950 256.950 931.050 259.050 ;
        RECT 914.550 254.550 919.050 256.050 ;
        RECT 907.950 253.950 912.000 254.550 ;
        RECT 915.000 253.950 919.050 254.550 ;
        RECT 899.400 243.900 906.000 244.800 ;
        RECT 899.400 243.600 900.900 243.900 ;
        RECT 896.100 237.000 897.900 243.600 ;
        RECT 899.100 237.600 900.900 243.600 ;
        RECT 905.100 243.600 906.000 243.900 ;
        RECT 921.000 244.800 921.900 256.950 ;
        RECT 926.100 255.150 927.900 256.950 ;
        RECT 935.550 256.050 936.450 259.950 ;
        RECT 941.700 259.050 942.900 269.400 ;
        RECT 940.950 256.950 943.050 259.050 ;
        RECT 943.950 256.950 946.050 259.050 ;
        RECT 935.550 254.550 940.050 256.050 ;
        RECT 936.000 253.950 940.050 254.550 ;
        RECT 921.000 243.900 927.600 244.800 ;
        RECT 921.000 243.600 921.900 243.900 ;
        RECT 902.100 237.000 903.900 243.000 ;
        RECT 905.100 237.600 906.900 243.600 ;
        RECT 920.100 237.600 921.900 243.600 ;
        RECT 926.100 243.600 927.600 243.900 ;
        RECT 941.700 243.600 942.900 256.950 ;
        RECT 944.100 255.150 945.900 256.950 ;
        RECT 923.100 237.000 924.900 243.000 ;
        RECT 926.100 237.600 927.900 243.600 ;
        RECT 929.100 237.000 930.900 243.600 ;
        RECT 941.100 237.600 942.900 243.600 ;
        RECT 944.100 237.000 945.900 243.600 ;
        RECT 11.100 227.400 12.900 233.400 ;
        RECT 14.100 227.400 15.900 234.000 ;
        RECT 29.100 227.400 30.900 234.000 ;
        RECT 32.100 227.400 33.900 233.400 ;
        RECT 35.100 227.400 36.900 234.000 ;
        RECT 50.100 227.400 51.900 234.000 ;
        RECT 53.100 227.400 54.900 233.400 ;
        RECT 56.100 227.400 57.900 234.000 ;
        RECT 11.700 214.050 12.900 227.400 ;
        RECT 14.100 214.050 15.900 215.850 ;
        RECT 32.700 214.050 33.900 227.400 ;
        RECT 53.700 214.050 54.900 227.400 ;
        RECT 68.400 221.400 70.200 234.000 ;
        RECT 73.500 222.900 75.300 233.400 ;
        RECT 76.500 227.400 78.300 234.000 ;
        RECT 89.100 227.400 90.900 234.000 ;
        RECT 92.100 227.400 93.900 233.400 ;
        RECT 95.100 227.400 96.900 234.000 ;
        RECT 110.100 227.400 111.900 234.000 ;
        RECT 113.100 227.400 114.900 233.400 ;
        RECT 116.100 227.400 117.900 234.000 ;
        RECT 76.200 224.100 78.000 225.900 ;
        RECT 73.500 221.400 75.900 222.900 ;
        RECT 68.100 214.050 69.900 215.850 ;
        RECT 74.700 214.050 75.900 221.400 ;
        RECT 92.100 214.050 93.300 227.400 ;
        RECT 113.100 214.050 114.300 227.400 ;
        RECT 131.100 222.300 132.900 233.400 ;
        RECT 134.100 223.200 135.900 234.000 ;
        RECT 137.100 222.300 138.900 233.400 ;
        RECT 131.100 221.400 138.900 222.300 ;
        RECT 140.100 221.400 141.900 233.400 ;
        RECT 155.100 227.400 156.900 234.000 ;
        RECT 158.100 227.400 159.900 233.400 ;
        RECT 161.100 227.400 162.900 234.000 ;
        RECT 173.100 227.400 174.900 233.400 ;
        RECT 176.100 227.400 177.900 234.000 ;
        RECT 191.100 227.400 192.900 234.000 ;
        RECT 194.100 227.400 195.900 233.400 ;
        RECT 197.100 228.000 198.900 234.000 ;
        RECT 115.950 219.450 118.050 220.050 ;
        RECT 133.950 219.450 136.050 220.050 ;
        RECT 115.950 218.550 136.050 219.450 ;
        RECT 115.950 217.950 118.050 218.550 ;
        RECT 133.950 217.950 136.050 218.550 ;
        RECT 134.250 214.050 136.050 215.850 ;
        RECT 140.700 214.050 141.600 221.400 ;
        RECT 158.100 214.050 159.300 227.400 ;
        RECT 173.700 214.050 174.900 227.400 ;
        RECT 194.400 227.100 195.900 227.400 ;
        RECT 200.100 227.400 201.900 233.400 ;
        RECT 215.700 227.400 217.500 234.000 ;
        RECT 200.100 227.100 201.000 227.400 ;
        RECT 194.400 226.200 201.000 227.100 ;
        RECT 176.100 214.050 177.900 215.850 ;
        RECT 194.100 214.050 195.900 215.850 ;
        RECT 200.100 214.050 201.000 226.200 ;
        RECT 216.000 224.100 217.800 225.900 ;
        RECT 218.700 222.900 220.500 233.400 ;
        RECT 218.100 221.400 220.500 222.900 ;
        RECT 223.800 221.400 225.600 234.000 ;
        RECT 236.100 227.400 237.900 234.000 ;
        RECT 239.100 227.400 240.900 233.400 ;
        RECT 251.100 227.400 252.900 234.000 ;
        RECT 254.100 227.400 255.900 233.400 ;
        RECT 257.100 228.000 258.900 234.000 ;
        RECT 210.000 216.450 214.050 217.050 ;
        RECT 209.550 214.950 214.050 216.450 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 28.950 211.950 31.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 160.950 211.950 163.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 11.700 201.600 12.900 211.950 ;
        RECT 29.100 210.150 30.900 211.950 ;
        RECT 32.700 206.700 33.900 211.950 ;
        RECT 34.950 210.150 36.750 211.950 ;
        RECT 50.100 210.150 51.900 211.950 ;
        RECT 53.700 206.700 54.900 211.950 ;
        RECT 55.950 210.150 57.750 211.950 ;
        RECT 71.100 210.150 72.900 211.950 ;
        RECT 74.700 207.600 75.900 211.950 ;
        RECT 77.100 210.150 78.900 211.950 ;
        RECT 89.250 210.150 91.050 211.950 ;
        RECT 74.700 206.700 78.300 207.600 ;
        RECT 29.700 205.800 33.900 206.700 ;
        RECT 50.700 205.800 54.900 206.700 ;
        RECT 11.100 198.600 12.900 201.600 ;
        RECT 14.100 198.000 15.900 201.600 ;
        RECT 29.700 198.600 31.500 205.800 ;
        RECT 34.800 198.000 36.600 204.600 ;
        RECT 50.700 198.600 52.500 205.800 ;
        RECT 55.800 198.000 57.600 204.600 ;
        RECT 68.100 203.700 75.900 205.050 ;
        RECT 68.100 198.600 69.900 203.700 ;
        RECT 71.100 198.000 72.900 202.800 ;
        RECT 74.100 198.600 75.900 203.700 ;
        RECT 77.100 204.600 78.300 206.700 ;
        RECT 92.100 206.700 93.300 211.950 ;
        RECT 95.100 210.150 96.900 211.950 ;
        RECT 110.250 210.150 112.050 211.950 ;
        RECT 113.100 206.700 114.300 211.950 ;
        RECT 116.100 210.150 117.900 211.950 ;
        RECT 131.100 210.150 132.900 211.950 ;
        RECT 137.250 210.150 139.050 211.950 ;
        RECT 92.100 205.800 96.300 206.700 ;
        RECT 113.100 205.800 117.300 206.700 ;
        RECT 77.100 198.600 78.900 204.600 ;
        RECT 89.400 198.000 91.200 204.600 ;
        RECT 94.500 198.600 96.300 205.800 ;
        RECT 110.400 198.000 112.200 204.600 ;
        RECT 115.500 198.600 117.300 205.800 ;
        RECT 140.700 204.600 141.600 211.950 ;
        RECT 155.250 210.150 157.050 211.950 ;
        RECT 158.100 206.700 159.300 211.950 ;
        RECT 161.100 210.150 162.900 211.950 ;
        RECT 158.100 205.800 162.300 206.700 ;
        RECT 132.000 198.000 133.800 204.600 ;
        RECT 136.500 203.400 141.600 204.600 ;
        RECT 136.500 198.600 138.300 203.400 ;
        RECT 139.500 198.000 141.300 201.600 ;
        RECT 155.400 198.000 157.200 204.600 ;
        RECT 160.500 198.600 162.300 205.800 ;
        RECT 173.700 201.600 174.900 211.950 ;
        RECT 191.100 210.150 192.900 211.950 ;
        RECT 197.100 210.150 198.900 211.950 ;
        RECT 200.100 208.200 201.000 211.950 ;
        RECT 209.550 211.050 210.450 214.950 ;
        RECT 218.100 214.050 219.300 221.400 ;
        RECT 231.000 216.450 235.050 217.050 ;
        RECT 224.100 214.050 225.900 215.850 ;
        RECT 230.550 214.950 235.050 216.450 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 209.550 209.550 214.050 211.050 ;
        RECT 215.100 210.150 216.900 211.950 ;
        RECT 210.000 208.950 214.050 209.550 ;
        RECT 173.100 198.600 174.900 201.600 ;
        RECT 176.100 198.000 177.900 201.600 ;
        RECT 191.100 198.000 192.900 207.600 ;
        RECT 197.700 207.000 201.000 208.200 ;
        RECT 218.100 207.600 219.300 211.950 ;
        RECT 221.100 210.150 222.900 211.950 ;
        RECT 230.550 211.050 231.450 214.950 ;
        RECT 236.100 214.050 237.900 215.850 ;
        RECT 239.100 214.050 240.300 227.400 ;
        RECT 254.400 227.100 255.900 227.400 ;
        RECT 260.100 227.400 261.900 233.400 ;
        RECT 272.100 227.400 273.900 234.000 ;
        RECT 275.100 227.400 276.900 233.400 ;
        RECT 278.100 227.400 279.900 234.000 ;
        RECT 293.700 227.400 295.500 234.000 ;
        RECT 260.100 227.100 261.000 227.400 ;
        RECT 254.400 226.200 261.000 227.100 ;
        RECT 254.100 214.050 255.900 215.850 ;
        RECT 260.100 214.050 261.000 226.200 ;
        RECT 265.950 220.050 268.050 223.050 ;
        RECT 265.950 219.000 271.050 220.050 ;
        RECT 266.550 218.550 271.050 219.000 ;
        RECT 267.000 217.950 271.050 218.550 ;
        RECT 275.100 214.050 276.300 227.400 ;
        RECT 294.000 224.100 295.800 225.900 ;
        RECT 296.700 222.900 298.500 233.400 ;
        RECT 296.100 221.400 298.500 222.900 ;
        RECT 301.800 221.400 303.600 234.000 ;
        RECT 304.950 231.450 307.050 232.050 ;
        RECT 313.950 231.450 316.050 232.050 ;
        RECT 304.950 230.550 316.050 231.450 ;
        RECT 304.950 229.950 307.050 230.550 ;
        RECT 313.950 229.950 316.050 230.550 ;
        RECT 317.100 227.400 318.900 234.000 ;
        RECT 320.100 227.400 321.900 233.400 ;
        RECT 277.950 219.450 280.050 220.050 ;
        RECT 292.950 219.450 295.050 220.050 ;
        RECT 277.950 218.550 295.050 219.450 ;
        RECT 277.950 217.950 280.050 218.550 ;
        RECT 292.950 217.950 295.050 218.550 ;
        RECT 296.100 214.050 297.300 221.400 ;
        RECT 304.950 216.450 309.000 217.050 ;
        RECT 302.100 214.050 303.900 215.850 ;
        RECT 304.950 214.950 309.450 216.450 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 256.950 211.950 259.050 214.050 ;
        RECT 259.950 211.950 262.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 226.950 209.550 231.450 211.050 ;
        RECT 226.950 208.950 231.000 209.550 ;
        RECT 197.700 198.600 199.500 207.000 ;
        RECT 215.700 206.700 219.300 207.600 ;
        RECT 215.700 204.600 216.900 206.700 ;
        RECT 215.100 198.600 216.900 204.600 ;
        RECT 218.100 203.700 225.900 205.050 ;
        RECT 218.100 198.600 219.900 203.700 ;
        RECT 221.100 198.000 222.900 202.800 ;
        RECT 224.100 198.600 225.900 203.700 ;
        RECT 239.100 201.600 240.300 211.950 ;
        RECT 251.100 210.150 252.900 211.950 ;
        RECT 257.100 210.150 258.900 211.950 ;
        RECT 260.100 208.200 261.000 211.950 ;
        RECT 272.250 210.150 274.050 211.950 ;
        RECT 236.100 198.000 237.900 201.600 ;
        RECT 239.100 198.600 240.900 201.600 ;
        RECT 251.100 198.000 252.900 207.600 ;
        RECT 257.700 207.000 261.000 208.200 ;
        RECT 257.700 198.600 259.500 207.000 ;
        RECT 275.100 206.700 276.300 211.950 ;
        RECT 278.100 210.150 279.900 211.950 ;
        RECT 293.100 210.150 294.900 211.950 ;
        RECT 296.100 207.600 297.300 211.950 ;
        RECT 299.100 210.150 300.900 211.950 ;
        RECT 308.550 211.050 309.450 214.950 ;
        RECT 317.100 211.950 319.200 214.050 ;
        RECT 304.950 209.550 309.450 211.050 ;
        RECT 317.250 210.150 319.050 211.950 ;
        RECT 304.950 208.950 309.000 209.550 ;
        RECT 293.700 206.700 297.300 207.600 ;
        RECT 320.100 207.300 321.000 227.400 ;
        RECT 323.100 222.000 324.900 234.000 ;
        RECT 326.100 221.400 327.900 233.400 ;
        RECT 338.100 227.400 339.900 234.000 ;
        RECT 341.100 227.400 342.900 233.400 ;
        RECT 344.100 227.400 345.900 234.000 ;
        RECT 322.200 214.050 324.000 215.850 ;
        RECT 326.400 214.050 327.300 221.400 ;
        RECT 341.100 214.050 342.300 227.400 ;
        RECT 356.400 221.400 358.200 234.000 ;
        RECT 361.500 222.900 363.300 233.400 ;
        RECT 364.500 227.400 366.300 234.000 ;
        RECT 380.700 227.400 382.500 234.000 ;
        RECT 364.200 224.100 366.000 225.900 ;
        RECT 381.000 224.100 382.800 225.900 ;
        RECT 383.700 222.900 385.500 233.400 ;
        RECT 361.500 221.400 363.900 222.900 ;
        RECT 356.100 214.050 357.900 215.850 ;
        RECT 362.700 214.050 363.900 221.400 ;
        RECT 383.100 221.400 385.500 222.900 ;
        RECT 388.800 221.400 390.600 234.000 ;
        RECT 404.100 227.400 405.900 234.000 ;
        RECT 407.100 227.400 408.900 233.400 ;
        RECT 383.100 214.050 384.300 221.400 ;
        RECT 385.950 219.450 388.050 220.050 ;
        RECT 394.950 219.450 397.050 220.050 ;
        RECT 385.950 218.550 397.050 219.450 ;
        RECT 385.950 217.950 388.050 218.550 ;
        RECT 394.950 217.950 397.050 218.550 ;
        RECT 389.100 214.050 390.900 215.850 ;
        RECT 322.500 211.950 324.600 214.050 ;
        RECT 325.800 211.950 327.900 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 404.100 211.950 406.200 214.050 ;
        RECT 275.100 205.800 279.300 206.700 ;
        RECT 272.400 198.000 274.200 204.600 ;
        RECT 277.500 198.600 279.300 205.800 ;
        RECT 293.700 204.600 294.900 206.700 ;
        RECT 317.100 206.400 325.500 207.300 ;
        RECT 293.100 198.600 294.900 204.600 ;
        RECT 296.100 203.700 303.900 205.050 ;
        RECT 296.100 198.600 297.900 203.700 ;
        RECT 299.100 198.000 300.900 202.800 ;
        RECT 302.100 198.600 303.900 203.700 ;
        RECT 317.100 198.600 318.900 206.400 ;
        RECT 323.700 205.500 325.500 206.400 ;
        RECT 326.400 204.600 327.300 211.950 ;
        RECT 338.250 210.150 340.050 211.950 ;
        RECT 341.100 206.700 342.300 211.950 ;
        RECT 344.100 210.150 345.900 211.950 ;
        RECT 359.100 210.150 360.900 211.950 ;
        RECT 362.700 207.600 363.900 211.950 ;
        RECT 365.100 210.150 366.900 211.950 ;
        RECT 380.100 210.150 381.900 211.950 ;
        RECT 383.100 207.600 384.300 211.950 ;
        RECT 386.100 210.150 387.900 211.950 ;
        RECT 404.250 210.150 406.050 211.950 ;
        RECT 362.700 206.700 366.300 207.600 ;
        RECT 341.100 205.800 345.300 206.700 ;
        RECT 321.600 198.000 323.400 204.600 ;
        RECT 324.600 202.800 327.300 204.600 ;
        RECT 324.600 198.600 326.400 202.800 ;
        RECT 338.400 198.000 340.200 204.600 ;
        RECT 343.500 198.600 345.300 205.800 ;
        RECT 356.100 203.700 363.900 205.050 ;
        RECT 356.100 198.600 357.900 203.700 ;
        RECT 359.100 198.000 360.900 202.800 ;
        RECT 362.100 198.600 363.900 203.700 ;
        RECT 365.100 204.600 366.300 206.700 ;
        RECT 380.700 206.700 384.300 207.600 ;
        RECT 407.100 207.300 408.000 227.400 ;
        RECT 410.100 222.000 411.900 234.000 ;
        RECT 413.100 221.400 414.900 233.400 ;
        RECT 428.100 227.400 429.900 234.000 ;
        RECT 431.100 227.400 432.900 233.400 ;
        RECT 434.100 227.400 435.900 234.000 ;
        RECT 446.100 227.400 447.900 234.000 ;
        RECT 449.100 227.400 450.900 233.400 ;
        RECT 409.200 214.050 411.000 215.850 ;
        RECT 413.400 214.050 414.300 221.400 ;
        RECT 431.100 214.050 432.300 227.400 ;
        RECT 409.500 211.950 411.600 214.050 ;
        RECT 412.800 211.950 414.900 214.050 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 430.950 211.950 433.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 446.100 211.950 448.200 214.050 ;
        RECT 380.700 204.600 381.900 206.700 ;
        RECT 404.100 206.400 412.500 207.300 ;
        RECT 365.100 198.600 366.900 204.600 ;
        RECT 380.100 198.600 381.900 204.600 ;
        RECT 383.100 203.700 390.900 205.050 ;
        RECT 383.100 198.600 384.900 203.700 ;
        RECT 386.100 198.000 387.900 202.800 ;
        RECT 389.100 198.600 390.900 203.700 ;
        RECT 404.100 198.600 405.900 206.400 ;
        RECT 410.700 205.500 412.500 206.400 ;
        RECT 413.400 204.600 414.300 211.950 ;
        RECT 428.250 210.150 430.050 211.950 ;
        RECT 431.100 206.700 432.300 211.950 ;
        RECT 434.100 210.150 435.900 211.950 ;
        RECT 446.250 210.150 448.050 211.950 ;
        RECT 449.100 207.300 450.000 227.400 ;
        RECT 452.100 222.000 453.900 234.000 ;
        RECT 455.100 221.400 456.900 233.400 ;
        RECT 470.100 227.400 471.900 234.000 ;
        RECT 473.100 227.400 474.900 233.400 ;
        RECT 476.100 227.400 477.900 234.000 ;
        RECT 488.700 227.400 490.500 234.000 ;
        RECT 451.200 214.050 453.000 215.850 ;
        RECT 455.400 214.050 456.300 221.400 ;
        RECT 473.700 214.050 474.900 227.400 ;
        RECT 489.000 224.100 490.800 225.900 ;
        RECT 491.700 222.900 493.500 233.400 ;
        RECT 491.100 221.400 493.500 222.900 ;
        RECT 496.800 221.400 498.600 234.000 ;
        RECT 509.100 227.400 510.900 234.000 ;
        RECT 512.100 227.400 513.900 233.400 ;
        RECT 491.100 214.050 492.300 221.400 ;
        RECT 497.100 214.050 498.900 215.850 ;
        RECT 509.100 214.050 510.900 215.850 ;
        RECT 512.100 214.050 513.300 227.400 ;
        RECT 527.400 221.400 529.200 234.000 ;
        RECT 532.500 222.900 534.300 233.400 ;
        RECT 535.500 227.400 537.300 234.000 ;
        RECT 551.100 227.400 552.900 234.000 ;
        RECT 554.100 227.400 555.900 233.400 ;
        RECT 569.100 227.400 570.900 233.400 ;
        RECT 572.100 227.400 573.900 234.000 ;
        RECT 587.100 227.400 588.900 234.000 ;
        RECT 590.100 227.400 591.900 233.400 ;
        RECT 535.200 224.100 537.000 225.900 ;
        RECT 532.500 221.400 534.900 222.900 ;
        RECT 522.000 216.450 526.050 217.050 ;
        RECT 521.550 214.950 526.050 216.450 ;
        RECT 451.500 211.950 453.600 214.050 ;
        RECT 454.800 211.950 456.900 214.050 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 472.950 211.950 475.050 214.050 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 431.100 205.800 435.300 206.700 ;
        RECT 408.600 198.000 410.400 204.600 ;
        RECT 411.600 202.800 414.300 204.600 ;
        RECT 411.600 198.600 413.400 202.800 ;
        RECT 428.400 198.000 430.200 204.600 ;
        RECT 433.500 198.600 435.300 205.800 ;
        RECT 446.100 206.400 454.500 207.300 ;
        RECT 446.100 198.600 447.900 206.400 ;
        RECT 452.700 205.500 454.500 206.400 ;
        RECT 455.400 204.600 456.300 211.950 ;
        RECT 470.100 210.150 471.900 211.950 ;
        RECT 473.700 206.700 474.900 211.950 ;
        RECT 475.950 210.150 477.750 211.950 ;
        RECT 488.100 210.150 489.900 211.950 ;
        RECT 491.100 207.600 492.300 211.950 ;
        RECT 494.100 210.150 495.900 211.950 ;
        RECT 450.600 198.000 452.400 204.600 ;
        RECT 453.600 202.800 456.300 204.600 ;
        RECT 470.700 205.800 474.900 206.700 ;
        RECT 488.700 206.700 492.300 207.600 ;
        RECT 453.600 198.600 455.400 202.800 ;
        RECT 470.700 198.600 472.500 205.800 ;
        RECT 488.700 204.600 489.900 206.700 ;
        RECT 475.800 198.000 477.600 204.600 ;
        RECT 488.100 198.600 489.900 204.600 ;
        RECT 491.100 203.700 498.900 205.050 ;
        RECT 491.100 198.600 492.900 203.700 ;
        RECT 494.100 198.000 495.900 202.800 ;
        RECT 497.100 198.600 498.900 203.700 ;
        RECT 512.100 201.600 513.300 211.950 ;
        RECT 514.950 210.450 517.050 211.050 ;
        RECT 521.550 210.450 522.450 214.950 ;
        RECT 527.100 214.050 528.900 215.850 ;
        RECT 533.700 214.050 534.900 221.400 ;
        RECT 551.100 214.050 552.900 215.850 ;
        RECT 554.100 214.050 555.300 227.400 ;
        RECT 569.700 214.050 570.900 227.400 ;
        RECT 572.100 214.050 573.900 215.850 ;
        RECT 587.100 214.050 588.900 215.850 ;
        RECT 590.100 214.050 591.300 227.400 ;
        RECT 605.100 222.300 606.900 233.400 ;
        RECT 608.100 223.200 609.900 234.000 ;
        RECT 611.100 222.300 612.900 233.400 ;
        RECT 605.100 221.400 612.900 222.300 ;
        RECT 614.100 221.400 615.900 233.400 ;
        RECT 629.100 227.400 630.900 234.000 ;
        RECT 632.100 227.400 633.900 233.400 ;
        RECT 635.100 227.400 636.900 234.000 ;
        RECT 608.250 214.050 610.050 215.850 ;
        RECT 614.700 214.050 615.600 221.400 ;
        RECT 624.000 216.450 628.050 217.050 ;
        RECT 623.550 214.950 628.050 216.450 ;
        RECT 526.950 211.950 529.050 214.050 ;
        RECT 529.950 211.950 532.050 214.050 ;
        RECT 532.950 211.950 535.050 214.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 550.950 211.950 553.050 214.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 514.950 209.550 522.450 210.450 ;
        RECT 530.100 210.150 531.900 211.950 ;
        RECT 514.950 208.950 517.050 209.550 ;
        RECT 533.700 207.600 534.900 211.950 ;
        RECT 536.100 210.150 537.900 211.950 ;
        RECT 533.700 206.700 537.300 207.600 ;
        RECT 527.100 203.700 534.900 205.050 ;
        RECT 509.100 198.000 510.900 201.600 ;
        RECT 512.100 198.600 513.900 201.600 ;
        RECT 527.100 198.600 528.900 203.700 ;
        RECT 530.100 198.000 531.900 202.800 ;
        RECT 533.100 198.600 534.900 203.700 ;
        RECT 536.100 204.600 537.300 206.700 ;
        RECT 536.100 198.600 537.900 204.600 ;
        RECT 554.100 201.600 555.300 211.950 ;
        RECT 569.700 201.600 570.900 211.950 ;
        RECT 571.950 207.450 574.050 208.050 ;
        RECT 577.950 207.450 580.050 208.050 ;
        RECT 571.950 206.550 580.050 207.450 ;
        RECT 571.950 205.950 574.050 206.550 ;
        RECT 577.950 205.950 580.050 206.550 ;
        RECT 590.100 201.600 591.300 211.950 ;
        RECT 605.100 210.150 606.900 211.950 ;
        RECT 611.250 210.150 613.050 211.950 ;
        RECT 598.950 207.450 601.050 208.050 ;
        RECT 607.950 207.450 610.050 208.050 ;
        RECT 598.950 206.550 610.050 207.450 ;
        RECT 598.950 205.950 601.050 206.550 ;
        RECT 607.950 205.950 610.050 206.550 ;
        RECT 614.700 204.600 615.600 211.950 ;
        RECT 623.550 211.050 624.450 214.950 ;
        RECT 632.700 214.050 633.900 227.400 ;
        RECT 648.000 222.600 649.800 233.400 ;
        RECT 648.000 221.400 651.600 222.600 ;
        RECT 653.100 221.400 654.900 234.000 ;
        RECT 665.100 227.400 666.900 234.000 ;
        RECT 668.100 227.400 669.900 233.400 ;
        RECT 671.100 227.400 672.900 234.000 ;
        RECT 637.950 216.450 642.000 217.050 ;
        RECT 637.950 214.950 642.450 216.450 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 623.550 209.550 628.050 211.050 ;
        RECT 629.100 210.150 630.900 211.950 ;
        RECT 624.000 208.950 628.050 209.550 ;
        RECT 632.700 206.700 633.900 211.950 ;
        RECT 634.950 210.150 636.750 211.950 ;
        RECT 641.550 210.450 642.450 214.950 ;
        RECT 647.100 214.050 648.900 215.850 ;
        RECT 650.700 214.050 651.600 221.400 ;
        RECT 652.950 214.050 654.750 215.850 ;
        RECT 668.700 214.050 669.900 227.400 ;
        RECT 686.100 222.300 687.900 233.400 ;
        RECT 689.100 223.200 690.900 234.000 ;
        RECT 692.100 222.300 693.900 233.400 ;
        RECT 686.100 221.400 693.900 222.300 ;
        RECT 695.100 221.400 696.900 233.400 ;
        RECT 710.100 227.400 711.900 234.000 ;
        RECT 713.100 227.400 714.900 233.400 ;
        RECT 716.100 228.000 717.900 234.000 ;
        RECT 713.400 227.100 714.900 227.400 ;
        RECT 719.100 227.400 720.900 233.400 ;
        RECT 731.100 227.400 732.900 234.000 ;
        RECT 734.100 227.400 735.900 233.400 ;
        RECT 737.100 228.000 738.900 234.000 ;
        RECT 719.100 227.100 720.000 227.400 ;
        RECT 713.400 226.200 720.000 227.100 ;
        RECT 734.400 227.100 735.900 227.400 ;
        RECT 740.100 227.400 741.900 233.400 ;
        RECT 740.100 227.100 741.000 227.400 ;
        RECT 734.400 226.200 741.000 227.100 ;
        RECT 681.000 216.450 685.050 217.050 ;
        RECT 680.550 214.950 685.050 216.450 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 649.950 211.950 652.050 214.050 ;
        RECT 652.950 211.950 655.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 670.950 211.950 673.050 214.050 ;
        RECT 641.550 210.000 645.450 210.450 ;
        RECT 641.550 209.550 646.050 210.000 ;
        RECT 551.100 198.000 552.900 201.600 ;
        RECT 554.100 198.600 555.900 201.600 ;
        RECT 569.100 198.600 570.900 201.600 ;
        RECT 572.100 198.000 573.900 201.600 ;
        RECT 587.100 198.000 588.900 201.600 ;
        RECT 590.100 198.600 591.900 201.600 ;
        RECT 606.000 198.000 607.800 204.600 ;
        RECT 610.500 203.400 615.600 204.600 ;
        RECT 629.700 205.800 633.900 206.700 ;
        RECT 643.950 205.950 646.050 209.550 ;
        RECT 610.500 198.600 612.300 203.400 ;
        RECT 613.500 198.000 615.300 201.600 ;
        RECT 629.700 198.600 631.500 205.800 ;
        RECT 634.800 198.000 636.600 204.600 ;
        RECT 650.700 201.600 651.600 211.950 ;
        RECT 665.100 210.150 666.900 211.950 ;
        RECT 668.700 206.700 669.900 211.950 ;
        RECT 670.950 210.150 672.750 211.950 ;
        RECT 680.550 210.450 681.450 214.950 ;
        RECT 689.250 214.050 691.050 215.850 ;
        RECT 695.700 214.050 696.600 221.400 ;
        RECT 697.950 219.450 700.050 220.050 ;
        RECT 715.950 219.450 718.050 220.050 ;
        RECT 697.950 218.550 718.050 219.450 ;
        RECT 697.950 217.950 700.050 218.550 ;
        RECT 715.950 217.950 718.050 218.550 ;
        RECT 700.950 216.450 703.050 217.050 ;
        RECT 706.950 216.450 709.050 217.050 ;
        RECT 700.950 215.550 709.050 216.450 ;
        RECT 700.950 214.950 703.050 215.550 ;
        RECT 706.950 214.950 709.050 215.550 ;
        RECT 713.100 214.050 714.900 215.850 ;
        RECT 719.100 214.050 720.000 226.200 ;
        RECT 724.950 219.450 727.050 220.050 ;
        RECT 730.950 219.450 733.050 220.050 ;
        RECT 724.950 218.550 733.050 219.450 ;
        RECT 724.950 217.950 727.050 218.550 ;
        RECT 730.950 217.950 733.050 218.550 ;
        RECT 734.100 214.050 735.900 215.850 ;
        RECT 740.100 214.050 741.000 226.200 ;
        RECT 755.100 222.300 756.900 233.400 ;
        RECT 758.100 223.200 759.900 234.000 ;
        RECT 761.100 222.300 762.900 233.400 ;
        RECT 755.100 221.400 762.900 222.300 ;
        RECT 764.100 221.400 765.900 233.400 ;
        RECT 779.100 227.400 780.900 234.000 ;
        RECT 782.100 227.400 783.900 233.400 ;
        RECT 785.100 227.400 786.900 234.000 ;
        RECT 800.100 227.400 801.900 234.000 ;
        RECT 803.100 227.400 804.900 233.400 ;
        RECT 806.100 228.000 807.900 234.000 ;
        RECT 748.950 219.450 751.050 220.050 ;
        RECT 760.950 219.450 763.050 220.050 ;
        RECT 748.950 218.550 763.050 219.450 ;
        RECT 748.950 217.950 751.050 218.550 ;
        RECT 760.950 217.950 763.050 218.550 ;
        RECT 758.250 214.050 760.050 215.850 ;
        RECT 764.700 214.050 765.600 221.400 ;
        RECT 782.700 214.050 783.900 227.400 ;
        RECT 803.400 227.100 804.900 227.400 ;
        RECT 809.100 227.400 810.900 233.400 ;
        RECT 809.100 227.100 810.000 227.400 ;
        RECT 803.400 226.200 810.000 227.100 ;
        RECT 803.100 214.050 804.900 215.850 ;
        RECT 809.100 214.050 810.000 226.200 ;
        RECT 822.000 222.600 823.800 233.400 ;
        RECT 822.000 221.400 825.600 222.600 ;
        RECT 827.100 221.400 828.900 234.000 ;
        RECT 842.100 222.300 843.900 233.400 ;
        RECT 845.100 223.200 846.900 234.000 ;
        RECT 848.100 222.300 849.900 233.400 ;
        RECT 842.100 221.400 849.900 222.300 ;
        RECT 851.100 221.400 852.900 233.400 ;
        RECT 863.100 227.400 864.900 234.000 ;
        RECT 866.100 227.400 867.900 233.400 ;
        RECT 869.100 228.000 870.900 234.000 ;
        RECT 866.400 227.100 867.900 227.400 ;
        RECT 872.100 227.400 873.900 233.400 ;
        RECT 887.100 227.400 888.900 234.000 ;
        RECT 890.100 227.400 891.900 233.400 ;
        RECT 893.100 228.000 894.900 234.000 ;
        RECT 872.100 227.100 873.000 227.400 ;
        RECT 866.400 226.200 873.000 227.100 ;
        RECT 890.400 227.100 891.900 227.400 ;
        RECT 896.100 227.400 897.900 233.400 ;
        RECT 908.100 227.400 909.900 233.400 ;
        RECT 911.100 228.000 912.900 234.000 ;
        RECT 896.100 227.100 897.000 227.400 ;
        RECT 890.400 226.200 897.000 227.100 ;
        RECT 821.100 214.050 822.900 215.850 ;
        RECT 824.700 214.050 825.600 221.400 ;
        RECT 826.950 214.050 828.750 215.850 ;
        RECT 845.250 214.050 847.050 215.850 ;
        RECT 851.700 214.050 852.600 221.400 ;
        RECT 858.000 216.450 862.050 217.050 ;
        RECT 857.550 214.950 862.050 216.450 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 694.950 211.950 697.050 214.050 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 680.550 209.550 684.450 210.450 ;
        RECT 686.100 210.150 687.900 211.950 ;
        RECT 692.250 210.150 694.050 211.950 ;
        RECT 665.700 205.800 669.900 206.700 ;
        RECT 683.550 207.450 684.450 209.550 ;
        RECT 688.950 207.450 691.050 208.050 ;
        RECT 683.550 206.550 691.050 207.450 ;
        RECT 688.950 205.950 691.050 206.550 ;
        RECT 647.100 198.000 648.900 201.600 ;
        RECT 650.100 198.600 651.900 201.600 ;
        RECT 653.100 198.000 654.900 201.600 ;
        RECT 665.700 198.600 667.500 205.800 ;
        RECT 695.700 204.600 696.600 211.950 ;
        RECT 710.100 210.150 711.900 211.950 ;
        RECT 716.100 210.150 717.900 211.950 ;
        RECT 719.100 208.200 720.000 211.950 ;
        RECT 731.100 210.150 732.900 211.950 ;
        RECT 737.100 210.150 738.900 211.950 ;
        RECT 740.100 208.200 741.000 211.950 ;
        RECT 755.100 210.150 756.900 211.950 ;
        RECT 761.250 210.150 763.050 211.950 ;
        RECT 670.800 198.000 672.600 204.600 ;
        RECT 687.000 198.000 688.800 204.600 ;
        RECT 691.500 203.400 696.600 204.600 ;
        RECT 691.500 198.600 693.300 203.400 ;
        RECT 694.500 198.000 696.300 201.600 ;
        RECT 710.100 198.000 711.900 207.600 ;
        RECT 716.700 207.000 720.000 208.200 ;
        RECT 716.700 198.600 718.500 207.000 ;
        RECT 731.100 198.000 732.900 207.600 ;
        RECT 737.700 207.000 741.000 208.200 ;
        RECT 737.700 198.600 739.500 207.000 ;
        RECT 764.700 204.600 765.600 211.950 ;
        RECT 779.100 210.150 780.900 211.950 ;
        RECT 782.700 206.700 783.900 211.950 ;
        RECT 784.950 210.150 786.750 211.950 ;
        RECT 800.100 210.150 801.900 211.950 ;
        RECT 806.100 210.150 807.900 211.950 ;
        RECT 809.100 208.200 810.000 211.950 ;
        RECT 756.000 198.000 757.800 204.600 ;
        RECT 760.500 203.400 765.600 204.600 ;
        RECT 779.700 205.800 783.900 206.700 ;
        RECT 760.500 198.600 762.300 203.400 ;
        RECT 763.500 198.000 765.300 201.600 ;
        RECT 779.700 198.600 781.500 205.800 ;
        RECT 784.800 198.000 786.600 204.600 ;
        RECT 800.100 198.000 801.900 207.600 ;
        RECT 806.700 207.000 810.000 208.200 ;
        RECT 806.700 198.600 808.500 207.000 ;
        RECT 824.700 201.600 825.600 211.950 ;
        RECT 842.100 210.150 843.900 211.950 ;
        RECT 848.250 210.150 850.050 211.950 ;
        RECT 851.700 204.600 852.600 211.950 ;
        RECT 857.550 211.050 858.450 214.950 ;
        RECT 866.100 214.050 867.900 215.850 ;
        RECT 872.100 214.050 873.000 226.200 ;
        RECT 874.950 216.450 879.000 217.050 ;
        RECT 882.000 216.450 886.050 217.050 ;
        RECT 874.950 214.950 879.450 216.450 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 857.550 209.550 862.050 211.050 ;
        RECT 863.100 210.150 864.900 211.950 ;
        RECT 869.100 210.150 870.900 211.950 ;
        RECT 858.000 208.950 862.050 209.550 ;
        RECT 872.100 208.200 873.000 211.950 ;
        RECT 878.550 211.050 879.450 214.950 ;
        RECT 874.950 209.550 879.450 211.050 ;
        RECT 881.550 214.950 886.050 216.450 ;
        RECT 881.550 210.450 882.450 214.950 ;
        RECT 890.100 214.050 891.900 215.850 ;
        RECT 896.100 214.050 897.000 226.200 ;
        RECT 909.000 227.100 909.900 227.400 ;
        RECT 914.100 227.400 915.900 233.400 ;
        RECT 917.100 227.400 918.900 234.000 ;
        RECT 932.100 227.400 933.900 234.000 ;
        RECT 935.100 227.400 936.900 233.400 ;
        RECT 938.100 228.000 939.900 234.000 ;
        RECT 914.100 227.100 915.600 227.400 ;
        RECT 909.000 226.200 915.600 227.100 ;
        RECT 935.400 227.100 936.900 227.400 ;
        RECT 941.100 227.400 942.900 233.400 ;
        RECT 941.100 227.100 942.000 227.400 ;
        RECT 935.400 226.200 942.000 227.100 ;
        RECT 903.000 216.450 907.050 217.050 ;
        RECT 902.550 214.950 907.050 216.450 ;
        RECT 886.950 211.950 889.050 214.050 ;
        RECT 889.950 211.950 892.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 895.950 211.950 898.050 214.050 ;
        RECT 881.550 209.550 885.450 210.450 ;
        RECT 887.100 210.150 888.900 211.950 ;
        RECT 893.100 210.150 894.900 211.950 ;
        RECT 874.950 208.950 879.000 209.550 ;
        RECT 821.100 198.000 822.900 201.600 ;
        RECT 824.100 198.600 825.900 201.600 ;
        RECT 827.100 198.000 828.900 201.600 ;
        RECT 843.000 198.000 844.800 204.600 ;
        RECT 847.500 203.400 852.600 204.600 ;
        RECT 847.500 198.600 849.300 203.400 ;
        RECT 850.500 198.000 852.300 201.600 ;
        RECT 863.100 198.000 864.900 207.600 ;
        RECT 869.700 207.000 873.000 208.200 ;
        RECT 869.700 198.600 871.500 207.000 ;
        RECT 877.950 204.450 880.050 205.050 ;
        RECT 884.550 204.450 885.450 209.550 ;
        RECT 896.100 208.200 897.000 211.950 ;
        RECT 902.550 211.050 903.450 214.950 ;
        RECT 909.000 214.050 909.900 226.200 ;
        RECT 922.950 220.950 925.050 223.050 ;
        RECT 914.100 214.050 915.900 215.850 ;
        RECT 907.950 211.950 910.050 214.050 ;
        RECT 910.950 211.950 913.050 214.050 ;
        RECT 913.950 211.950 916.050 214.050 ;
        RECT 916.950 211.950 919.050 214.050 ;
        RECT 902.550 209.550 907.050 211.050 ;
        RECT 903.000 208.950 907.050 209.550 ;
        RECT 877.950 203.550 885.450 204.450 ;
        RECT 877.950 202.950 880.050 203.550 ;
        RECT 887.100 198.000 888.900 207.600 ;
        RECT 893.700 207.000 897.000 208.200 ;
        RECT 909.000 208.200 909.900 211.950 ;
        RECT 911.100 210.150 912.900 211.950 ;
        RECT 917.100 210.150 918.900 211.950 ;
        RECT 909.000 207.000 912.300 208.200 ;
        RECT 923.550 208.050 924.450 220.950 ;
        RECT 935.100 214.050 936.900 215.850 ;
        RECT 941.100 214.050 942.000 226.200 ;
        RECT 931.950 211.950 934.050 214.050 ;
        RECT 934.950 211.950 937.050 214.050 ;
        RECT 937.950 211.950 940.050 214.050 ;
        RECT 940.950 211.950 943.050 214.050 ;
        RECT 932.100 210.150 933.900 211.950 ;
        RECT 938.100 210.150 939.900 211.950 ;
        RECT 941.100 208.200 942.000 211.950 ;
        RECT 893.700 198.600 895.500 207.000 ;
        RECT 910.500 198.600 912.300 207.000 ;
        RECT 917.100 198.000 918.900 207.600 ;
        RECT 919.950 206.550 924.450 208.050 ;
        RECT 919.950 205.950 924.000 206.550 ;
        RECT 932.100 198.000 933.900 207.600 ;
        RECT 938.700 207.000 942.000 208.200 ;
        RECT 938.700 198.600 940.500 207.000 ;
        RECT 14.100 185.400 15.900 195.000 ;
        RECT 20.700 186.000 22.500 194.400 ;
        RECT 39.000 188.400 40.800 195.000 ;
        RECT 43.500 189.600 45.300 194.400 ;
        RECT 46.500 191.400 48.300 195.000 ;
        RECT 43.500 188.400 48.600 189.600 ;
        RECT 28.950 186.450 31.050 187.050 ;
        RECT 40.950 186.450 43.050 187.050 ;
        RECT 20.700 184.800 24.000 186.000 ;
        RECT 28.950 185.550 43.050 186.450 ;
        RECT 28.950 184.950 31.050 185.550 ;
        RECT 40.950 184.950 43.050 185.550 ;
        RECT 14.100 181.050 15.900 182.850 ;
        RECT 20.100 181.050 21.900 182.850 ;
        RECT 23.100 181.050 24.000 184.800 ;
        RECT 38.100 181.050 39.900 182.850 ;
        RECT 44.250 181.050 46.050 182.850 ;
        RECT 47.700 181.050 48.600 188.400 ;
        RECT 59.100 185.400 60.900 195.000 ;
        RECT 65.700 186.000 67.500 194.400 ;
        RECT 83.100 189.300 84.900 194.400 ;
        RECT 86.100 190.200 87.900 195.000 ;
        RECT 89.100 189.300 90.900 194.400 ;
        RECT 83.100 187.950 90.900 189.300 ;
        RECT 92.100 188.400 93.900 194.400 ;
        RECT 104.100 189.300 105.900 194.400 ;
        RECT 107.100 190.200 108.900 195.000 ;
        RECT 110.100 189.300 111.900 194.400 ;
        RECT 92.100 186.300 93.300 188.400 ;
        RECT 104.100 187.950 111.900 189.300 ;
        RECT 113.100 188.400 114.900 194.400 ;
        RECT 113.100 186.300 114.300 188.400 ;
        RECT 65.700 184.800 69.000 186.000 ;
        RECT 49.950 183.450 54.000 184.050 ;
        RECT 49.950 181.950 54.450 183.450 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 17.100 177.150 18.900 178.950 ;
        RECT 23.100 166.800 24.000 178.950 ;
        RECT 41.250 177.150 43.050 178.950 ;
        RECT 28.950 174.450 31.050 175.050 ;
        RECT 40.950 174.450 43.050 175.050 ;
        RECT 28.950 173.550 43.050 174.450 ;
        RECT 28.950 172.950 31.050 173.550 ;
        RECT 40.950 172.950 43.050 173.550 ;
        RECT 47.700 171.600 48.600 178.950 ;
        RECT 53.550 178.050 54.450 181.950 ;
        RECT 59.100 181.050 60.900 182.850 ;
        RECT 65.100 181.050 66.900 182.850 ;
        RECT 68.100 181.050 69.000 184.800 ;
        RECT 89.700 185.400 93.300 186.300 ;
        RECT 110.700 185.400 114.300 186.300 ;
        RECT 128.100 185.400 129.900 195.000 ;
        RECT 134.700 186.000 136.500 194.400 ;
        RECT 149.100 188.400 150.900 194.400 ;
        RECT 149.700 186.300 150.900 188.400 ;
        RECT 152.100 189.300 153.900 194.400 ;
        RECT 155.100 190.200 156.900 195.000 ;
        RECT 158.100 189.300 159.900 194.400 ;
        RECT 152.100 187.950 159.900 189.300 ;
        RECT 173.700 187.200 175.500 194.400 ;
        RECT 178.800 188.400 180.600 195.000 ;
        RECT 194.100 189.300 195.900 194.400 ;
        RECT 197.100 190.200 198.900 195.000 ;
        RECT 200.100 189.300 201.900 194.400 ;
        RECT 194.100 187.950 201.900 189.300 ;
        RECT 203.100 188.400 204.900 194.400 ;
        RECT 218.100 188.400 219.900 194.400 ;
        RECT 173.700 186.300 177.900 187.200 ;
        RECT 203.100 186.300 204.300 188.400 ;
        RECT 86.100 181.050 87.900 182.850 ;
        RECT 89.700 181.050 90.900 185.400 ;
        RECT 92.100 181.050 93.900 182.850 ;
        RECT 107.100 181.050 108.900 182.850 ;
        RECT 110.700 181.050 111.900 185.400 ;
        RECT 134.700 184.800 138.000 186.000 ;
        RECT 149.700 185.400 153.300 186.300 ;
        RECT 113.100 181.050 114.900 182.850 ;
        RECT 128.100 181.050 129.900 182.850 ;
        RECT 134.100 181.050 135.900 182.850 ;
        RECT 137.100 181.050 138.000 184.800 ;
        RECT 149.100 181.050 150.900 182.850 ;
        RECT 152.100 181.050 153.300 185.400 ;
        RECT 155.100 181.050 156.900 182.850 ;
        RECT 173.100 181.050 174.900 182.850 ;
        RECT 176.700 181.050 177.900 186.300 ;
        RECT 200.700 185.400 204.300 186.300 ;
        RECT 218.700 186.300 219.900 188.400 ;
        RECT 221.100 189.300 222.900 194.400 ;
        RECT 224.100 190.200 225.900 195.000 ;
        RECT 227.100 189.300 228.900 194.400 ;
        RECT 221.100 187.950 228.900 189.300 ;
        RECT 218.700 185.400 222.300 186.300 ;
        RECT 239.100 185.400 240.900 195.000 ;
        RECT 245.700 186.000 247.500 194.400 ;
        RECT 260.100 188.400 261.900 194.400 ;
        RECT 260.700 186.300 261.900 188.400 ;
        RECT 263.100 189.300 264.900 194.400 ;
        RECT 266.100 190.200 267.900 195.000 ;
        RECT 269.100 189.300 270.900 194.400 ;
        RECT 263.100 187.950 270.900 189.300 ;
        RECT 284.700 187.200 286.500 194.400 ;
        RECT 289.800 188.400 291.600 195.000 ;
        RECT 302.400 188.400 304.200 195.000 ;
        RECT 307.500 187.200 309.300 194.400 ;
        RECT 323.100 188.400 324.900 194.400 ;
        RECT 284.700 186.300 288.900 187.200 ;
        RECT 181.950 183.450 186.000 184.050 ;
        RECT 178.950 181.050 180.750 182.850 ;
        RECT 181.950 181.950 186.450 183.450 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 109.950 178.950 112.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 148.950 178.950 151.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 49.950 176.550 54.450 178.050 ;
        RECT 62.100 177.150 63.900 178.950 ;
        RECT 49.950 175.950 54.000 176.550 ;
        RECT 17.400 165.900 24.000 166.800 ;
        RECT 17.400 165.600 18.900 165.900 ;
        RECT 14.100 159.000 15.900 165.600 ;
        RECT 17.100 159.600 18.900 165.600 ;
        RECT 23.100 165.600 24.000 165.900 ;
        RECT 38.100 170.700 45.900 171.600 ;
        RECT 20.100 159.000 21.900 165.000 ;
        RECT 23.100 159.600 24.900 165.600 ;
        RECT 38.100 159.600 39.900 170.700 ;
        RECT 41.100 159.000 42.900 169.800 ;
        RECT 44.100 159.600 45.900 170.700 ;
        RECT 47.100 159.600 48.900 171.600 ;
        RECT 68.100 166.800 69.000 178.950 ;
        RECT 83.100 177.150 84.900 178.950 ;
        RECT 89.700 171.600 90.900 178.950 ;
        RECT 104.100 177.150 105.900 178.950 ;
        RECT 110.700 171.600 111.900 178.950 ;
        RECT 131.100 177.150 132.900 178.950 ;
        RECT 62.400 165.900 69.000 166.800 ;
        RECT 62.400 165.600 63.900 165.900 ;
        RECT 59.100 159.000 60.900 165.600 ;
        RECT 62.100 159.600 63.900 165.600 ;
        RECT 68.100 165.600 69.000 165.900 ;
        RECT 65.100 159.000 66.900 165.000 ;
        RECT 68.100 159.600 69.900 165.600 ;
        RECT 83.400 159.000 85.200 171.600 ;
        RECT 88.500 170.100 90.900 171.600 ;
        RECT 88.500 159.600 90.300 170.100 ;
        RECT 91.200 167.100 93.000 168.900 ;
        RECT 91.500 159.000 93.300 165.600 ;
        RECT 104.400 159.000 106.200 171.600 ;
        RECT 109.500 170.100 111.900 171.600 ;
        RECT 109.500 159.600 111.300 170.100 ;
        RECT 112.200 167.100 114.000 168.900 ;
        RECT 137.100 166.800 138.000 178.950 ;
        RECT 152.100 171.600 153.300 178.950 ;
        RECT 158.100 177.150 159.900 178.950 ;
        RECT 152.100 170.100 154.500 171.600 ;
        RECT 150.000 167.100 151.800 168.900 ;
        RECT 131.400 165.900 138.000 166.800 ;
        RECT 131.400 165.600 132.900 165.900 ;
        RECT 112.500 159.000 114.300 165.600 ;
        RECT 128.100 159.000 129.900 165.600 ;
        RECT 131.100 159.600 132.900 165.600 ;
        RECT 137.100 165.600 138.000 165.900 ;
        RECT 134.100 159.000 135.900 165.000 ;
        RECT 137.100 159.600 138.900 165.600 ;
        RECT 149.700 159.000 151.500 165.600 ;
        RECT 152.700 159.600 154.500 170.100 ;
        RECT 157.800 159.000 159.600 171.600 ;
        RECT 176.700 165.600 177.900 178.950 ;
        RECT 185.550 174.450 186.450 181.950 ;
        RECT 197.100 181.050 198.900 182.850 ;
        RECT 200.700 181.050 201.900 185.400 ;
        RECT 205.950 183.450 208.050 184.050 ;
        RECT 211.950 183.450 214.050 184.050 ;
        RECT 203.100 181.050 204.900 182.850 ;
        RECT 205.950 182.550 214.050 183.450 ;
        RECT 205.950 181.950 208.050 182.550 ;
        RECT 211.950 181.950 214.050 182.550 ;
        RECT 218.100 181.050 219.900 182.850 ;
        RECT 221.100 181.050 222.300 185.400 ;
        RECT 245.700 184.800 249.000 186.000 ;
        RECT 260.700 185.400 264.300 186.300 ;
        RECT 224.100 181.050 225.900 182.850 ;
        RECT 239.100 181.050 240.900 182.850 ;
        RECT 245.100 181.050 246.900 182.850 ;
        RECT 248.100 181.050 249.000 184.800 ;
        RECT 260.100 181.050 261.900 182.850 ;
        RECT 263.100 181.050 264.300 185.400 ;
        RECT 266.100 181.050 267.900 182.850 ;
        RECT 284.100 181.050 285.900 182.850 ;
        RECT 287.700 181.050 288.900 186.300 ;
        RECT 305.100 186.300 309.300 187.200 ;
        RECT 323.700 186.300 324.900 188.400 ;
        RECT 326.100 189.300 327.900 194.400 ;
        RECT 329.100 190.200 330.900 195.000 ;
        RECT 332.100 189.300 333.900 194.400 ;
        RECT 326.100 187.950 333.900 189.300 ;
        RECT 343.950 187.950 346.050 190.050 ;
        RECT 292.950 183.450 297.000 184.050 ;
        RECT 289.950 181.050 291.750 182.850 ;
        RECT 292.950 181.950 297.450 183.450 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 283.950 178.950 286.050 181.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 194.100 177.150 195.900 178.950 ;
        RECT 193.950 174.450 196.050 175.050 ;
        RECT 185.550 173.550 196.050 174.450 ;
        RECT 193.950 172.950 196.050 173.550 ;
        RECT 200.700 171.600 201.900 178.950 ;
        RECT 173.100 159.000 174.900 165.600 ;
        RECT 176.100 159.600 177.900 165.600 ;
        RECT 179.100 159.000 180.900 165.600 ;
        RECT 194.400 159.000 196.200 171.600 ;
        RECT 199.500 170.100 201.900 171.600 ;
        RECT 221.100 171.600 222.300 178.950 ;
        RECT 227.100 177.150 228.900 178.950 ;
        RECT 242.100 177.150 243.900 178.950 ;
        RECT 221.100 170.100 223.500 171.600 ;
        RECT 199.500 159.600 201.300 170.100 ;
        RECT 202.200 167.100 204.000 168.900 ;
        RECT 219.000 167.100 220.800 168.900 ;
        RECT 202.500 159.000 204.300 165.600 ;
        RECT 218.700 159.000 220.500 165.600 ;
        RECT 221.700 159.600 223.500 170.100 ;
        RECT 226.800 159.000 228.600 171.600 ;
        RECT 248.100 166.800 249.000 178.950 ;
        RECT 263.100 171.600 264.300 178.950 ;
        RECT 269.100 177.150 270.900 178.950 ;
        RECT 265.950 174.450 268.050 175.050 ;
        RECT 280.950 174.450 283.050 175.050 ;
        RECT 265.950 173.550 283.050 174.450 ;
        RECT 265.950 172.950 268.050 173.550 ;
        RECT 280.950 172.950 283.050 173.550 ;
        RECT 263.100 170.100 265.500 171.600 ;
        RECT 261.000 167.100 262.800 168.900 ;
        RECT 242.400 165.900 249.000 166.800 ;
        RECT 242.400 165.600 243.900 165.900 ;
        RECT 239.100 159.000 240.900 165.600 ;
        RECT 242.100 159.600 243.900 165.600 ;
        RECT 248.100 165.600 249.000 165.900 ;
        RECT 245.100 159.000 246.900 165.000 ;
        RECT 248.100 159.600 249.900 165.600 ;
        RECT 260.700 159.000 262.500 165.600 ;
        RECT 263.700 159.600 265.500 170.100 ;
        RECT 268.800 159.000 270.600 171.600 ;
        RECT 274.950 171.450 277.050 171.900 ;
        RECT 283.950 171.450 286.050 172.050 ;
        RECT 274.950 170.550 286.050 171.450 ;
        RECT 274.950 169.800 277.050 170.550 ;
        RECT 283.950 169.950 286.050 170.550 ;
        RECT 287.700 165.600 288.900 178.950 ;
        RECT 296.550 177.450 297.450 181.950 ;
        RECT 302.250 181.050 304.050 182.850 ;
        RECT 305.100 181.050 306.300 186.300 ;
        RECT 323.700 185.400 327.300 186.300 ;
        RECT 308.100 181.050 309.900 182.850 ;
        RECT 323.100 181.050 324.900 182.850 ;
        RECT 326.100 181.050 327.300 185.400 ;
        RECT 334.950 183.450 337.050 183.900 ;
        RECT 344.550 183.450 345.450 187.950 ;
        RECT 347.100 185.400 348.900 195.000 ;
        RECT 353.700 186.000 355.500 194.400 ;
        RECT 367.950 189.450 370.050 190.050 ;
        RECT 359.550 189.000 370.050 189.450 ;
        RECT 358.950 188.550 370.050 189.000 ;
        RECT 353.700 184.800 357.000 186.000 ;
        RECT 358.950 184.950 361.050 188.550 ;
        RECT 367.950 187.950 370.050 188.550 ;
        RECT 371.100 185.400 372.900 195.000 ;
        RECT 377.700 186.000 379.500 194.400 ;
        RECT 392.100 191.400 393.900 195.000 ;
        RECT 395.100 191.400 396.900 194.400 ;
        RECT 377.700 184.800 381.000 186.000 ;
        RECT 329.100 181.050 330.900 182.850 ;
        RECT 334.950 182.550 345.450 183.450 ;
        RECT 334.950 181.800 337.050 182.550 ;
        RECT 347.100 181.050 348.900 182.850 ;
        RECT 353.100 181.050 354.900 182.850 ;
        RECT 356.100 181.050 357.000 184.800 ;
        RECT 371.100 181.050 372.900 182.850 ;
        RECT 377.100 181.050 378.900 182.850 ;
        RECT 380.100 181.050 381.000 184.800 ;
        RECT 382.950 183.450 387.000 184.050 ;
        RECT 382.950 181.950 387.450 183.450 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 293.550 176.550 297.450 177.450 ;
        RECT 293.550 175.050 294.450 176.550 ;
        RECT 291.000 174.750 294.450 175.050 ;
        RECT 289.950 173.550 294.450 174.750 ;
        RECT 289.950 172.950 294.000 173.550 ;
        RECT 289.950 172.650 292.050 172.950 ;
        RECT 305.100 165.600 306.300 178.950 ;
        RECT 326.100 171.600 327.300 178.950 ;
        RECT 332.100 177.150 333.900 178.950 ;
        RECT 350.100 177.150 351.900 178.950 ;
        RECT 326.100 170.100 328.500 171.600 ;
        RECT 324.000 167.100 325.800 168.900 ;
        RECT 284.100 159.000 285.900 165.600 ;
        RECT 287.100 159.600 288.900 165.600 ;
        RECT 290.100 159.000 291.900 165.600 ;
        RECT 302.100 159.000 303.900 165.600 ;
        RECT 305.100 159.600 306.900 165.600 ;
        RECT 308.100 159.000 309.900 165.600 ;
        RECT 323.700 159.000 325.500 165.600 ;
        RECT 326.700 159.600 328.500 170.100 ;
        RECT 331.800 159.000 333.600 171.600 ;
        RECT 356.100 166.800 357.000 178.950 ;
        RECT 374.100 177.150 375.900 178.950 ;
        RECT 358.950 174.450 361.050 175.050 ;
        RECT 373.950 174.450 376.050 175.050 ;
        RECT 358.950 173.550 376.050 174.450 ;
        RECT 358.950 172.950 361.050 173.550 ;
        RECT 373.950 172.950 376.050 173.550 ;
        RECT 380.100 166.800 381.000 178.950 ;
        RECT 386.550 178.050 387.450 181.950 ;
        RECT 395.100 181.050 396.300 191.400 ;
        RECT 410.700 187.200 412.500 194.400 ;
        RECT 415.800 188.400 417.600 195.000 ;
        RECT 433.500 188.400 435.300 195.000 ;
        RECT 438.000 188.400 439.800 194.400 ;
        RECT 442.500 188.400 444.300 195.000 ;
        RECT 458.100 189.300 459.900 194.400 ;
        RECT 461.100 190.200 462.900 195.000 ;
        RECT 464.100 189.300 465.900 194.400 ;
        RECT 410.700 186.300 414.900 187.200 ;
        RECT 405.000 183.450 409.050 184.050 ;
        RECT 404.550 181.950 409.050 183.450 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 382.950 176.550 387.450 178.050 ;
        RECT 392.100 177.150 393.900 178.950 ;
        RECT 382.950 175.950 387.000 176.550 ;
        RECT 350.400 165.900 357.000 166.800 ;
        RECT 350.400 165.600 351.900 165.900 ;
        RECT 347.100 159.000 348.900 165.600 ;
        RECT 350.100 159.600 351.900 165.600 ;
        RECT 356.100 165.600 357.000 165.900 ;
        RECT 374.400 165.900 381.000 166.800 ;
        RECT 374.400 165.600 375.900 165.900 ;
        RECT 353.100 159.000 354.900 165.000 ;
        RECT 356.100 159.600 357.900 165.600 ;
        RECT 371.100 159.000 372.900 165.600 ;
        RECT 374.100 159.600 375.900 165.600 ;
        RECT 380.100 165.600 381.000 165.900 ;
        RECT 395.100 165.600 396.300 178.950 ;
        RECT 397.950 177.450 400.050 178.050 ;
        RECT 404.550 177.450 405.450 181.950 ;
        RECT 410.100 181.050 411.900 182.850 ;
        RECT 413.700 181.050 414.900 186.300 ;
        RECT 415.950 186.450 418.050 187.050 ;
        RECT 427.950 186.450 430.050 187.050 ;
        RECT 415.950 185.550 430.050 186.450 ;
        RECT 415.950 184.950 418.050 185.550 ;
        RECT 427.950 184.950 430.050 185.550 ;
        RECT 415.950 181.050 417.750 182.850 ;
        RECT 431.100 181.050 432.900 182.850 ;
        RECT 437.700 181.050 438.900 188.400 ;
        RECT 458.100 187.950 465.900 189.300 ;
        RECT 467.100 188.400 468.900 194.400 ;
        RECT 467.100 186.300 468.300 188.400 ;
        RECT 464.700 185.400 468.300 186.300 ;
        RECT 484.500 186.000 486.300 194.400 ;
        RECT 453.000 183.450 457.050 184.050 ;
        RECT 442.950 181.050 444.750 182.850 ;
        RECT 452.550 181.950 457.050 183.450 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 397.950 176.550 405.450 177.450 ;
        RECT 397.950 175.950 400.050 176.550 ;
        RECT 400.950 174.450 403.050 175.050 ;
        RECT 406.950 174.450 409.050 175.050 ;
        RECT 400.950 173.550 409.050 174.450 ;
        RECT 400.950 172.950 403.050 173.550 ;
        RECT 406.950 172.950 409.050 173.550 ;
        RECT 413.700 165.600 414.900 178.950 ;
        RECT 434.100 177.150 435.900 178.950 ;
        RECT 438.000 173.400 438.900 178.950 ;
        RECT 439.950 177.150 441.750 178.950 ;
        RECT 452.550 178.050 453.450 181.950 ;
        RECT 461.100 181.050 462.900 182.850 ;
        RECT 464.700 181.050 465.900 185.400 ;
        RECT 483.000 184.800 486.300 186.000 ;
        RECT 491.100 185.400 492.900 195.000 ;
        RECT 503.700 187.200 505.500 194.400 ;
        RECT 508.800 188.400 510.600 195.000 ;
        RECT 524.100 191.400 525.900 195.000 ;
        RECT 527.100 191.400 528.900 194.400 ;
        RECT 503.700 186.300 507.900 187.200 ;
        RECT 467.100 181.050 468.900 182.850 ;
        RECT 483.000 181.050 483.900 184.800 ;
        RECT 498.000 183.450 502.050 184.050 ;
        RECT 485.100 181.050 486.900 182.850 ;
        RECT 491.100 181.050 492.900 182.850 ;
        RECT 497.550 181.950 502.050 183.450 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 463.950 178.950 466.050 181.050 ;
        RECT 466.950 178.950 469.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 484.950 178.950 487.050 181.050 ;
        RECT 487.950 178.950 490.050 181.050 ;
        RECT 490.950 178.950 493.050 181.050 ;
        RECT 452.550 176.550 457.050 178.050 ;
        RECT 458.100 177.150 459.900 178.950 ;
        RECT 453.000 175.950 457.050 176.550 ;
        RECT 434.100 172.500 438.900 173.400 ;
        RECT 377.100 159.000 378.900 165.000 ;
        RECT 380.100 159.600 381.900 165.600 ;
        RECT 392.100 159.000 393.900 165.600 ;
        RECT 395.100 159.600 396.900 165.600 ;
        RECT 410.100 159.000 411.900 165.600 ;
        RECT 413.100 159.600 414.900 165.600 ;
        RECT 416.100 159.000 417.900 165.600 ;
        RECT 431.100 160.500 432.900 171.600 ;
        RECT 434.100 161.400 435.900 172.500 ;
        RECT 464.700 171.600 465.900 178.950 ;
        RECT 466.950 174.450 469.050 175.050 ;
        RECT 472.950 174.450 475.050 175.050 ;
        RECT 466.950 173.550 475.050 174.450 ;
        RECT 466.950 172.950 469.050 173.550 ;
        RECT 472.950 172.950 475.050 173.550 ;
        RECT 437.100 170.400 444.900 171.300 ;
        RECT 437.100 160.500 438.900 170.400 ;
        RECT 431.100 159.600 438.900 160.500 ;
        RECT 440.100 159.000 441.900 169.500 ;
        RECT 443.100 159.600 444.900 170.400 ;
        RECT 458.400 159.000 460.200 171.600 ;
        RECT 463.500 170.100 465.900 171.600 ;
        RECT 463.500 159.600 465.300 170.100 ;
        RECT 466.200 167.100 468.000 168.900 ;
        RECT 483.000 166.800 483.900 178.950 ;
        RECT 488.100 177.150 489.900 178.950 ;
        RECT 497.550 178.050 498.450 181.950 ;
        RECT 503.100 181.050 504.900 182.850 ;
        RECT 506.700 181.050 507.900 186.300 ;
        RECT 508.950 181.050 510.750 182.850 ;
        RECT 527.100 181.050 528.300 191.400 ;
        RECT 542.100 185.400 543.900 195.000 ;
        RECT 548.700 186.000 550.500 194.400 ;
        RECT 548.700 184.800 552.000 186.000 ;
        RECT 566.100 185.400 567.900 195.000 ;
        RECT 572.700 186.000 574.500 194.400 ;
        RECT 587.100 189.300 588.900 194.400 ;
        RECT 590.100 190.200 591.900 195.000 ;
        RECT 593.100 189.300 594.900 194.400 ;
        RECT 587.100 187.950 594.900 189.300 ;
        RECT 596.100 188.400 597.900 194.400 ;
        RECT 596.100 186.300 597.300 188.400 ;
        RECT 572.700 184.800 576.000 186.000 ;
        RECT 542.100 181.050 543.900 182.850 ;
        RECT 548.100 181.050 549.900 182.850 ;
        RECT 551.100 181.050 552.000 184.800 ;
        RECT 566.100 181.050 567.900 182.850 ;
        RECT 572.100 181.050 573.900 182.850 ;
        RECT 575.100 181.050 576.000 184.800 ;
        RECT 593.700 185.400 597.300 186.300 ;
        RECT 608.100 185.400 609.900 195.000 ;
        RECT 614.700 186.000 616.500 194.400 ;
        RECT 629.100 189.300 630.900 194.400 ;
        RECT 632.100 190.200 633.900 195.000 ;
        RECT 635.100 189.300 636.900 194.400 ;
        RECT 629.100 187.950 636.900 189.300 ;
        RECT 638.100 188.400 639.900 194.400 ;
        RECT 653.100 191.400 654.900 195.000 ;
        RECT 656.100 191.400 657.900 194.400 ;
        RECT 659.100 191.400 660.900 195.000 ;
        RECT 638.100 186.300 639.300 188.400 ;
        RECT 582.000 183.450 586.050 184.050 ;
        RECT 581.550 181.950 586.050 183.450 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 505.950 178.950 508.050 181.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 574.950 178.950 577.050 181.050 ;
        RECT 493.950 176.550 498.450 178.050 ;
        RECT 493.950 175.950 498.000 176.550 ;
        RECT 483.000 165.900 489.600 166.800 ;
        RECT 483.000 165.600 483.900 165.900 ;
        RECT 466.500 159.000 468.300 165.600 ;
        RECT 482.100 159.600 483.900 165.600 ;
        RECT 488.100 165.600 489.600 165.900 ;
        RECT 506.700 165.600 507.900 178.950 ;
        RECT 524.100 177.150 525.900 178.950 ;
        RECT 527.100 165.600 528.300 178.950 ;
        RECT 545.100 177.150 546.900 178.950 ;
        RECT 529.950 174.450 532.050 175.050 ;
        RECT 547.950 174.450 550.050 175.050 ;
        RECT 529.950 173.550 550.050 174.450 ;
        RECT 529.950 172.950 532.050 173.550 ;
        RECT 547.950 172.950 550.050 173.550 ;
        RECT 551.100 166.800 552.000 178.950 ;
        RECT 569.100 177.150 570.900 178.950 ;
        RECT 575.100 166.800 576.000 178.950 ;
        RECT 581.550 178.050 582.450 181.950 ;
        RECT 590.100 181.050 591.900 182.850 ;
        RECT 593.700 181.050 594.900 185.400 ;
        RECT 614.700 184.800 618.000 186.000 ;
        RECT 596.100 181.050 597.900 182.850 ;
        RECT 608.100 181.050 609.900 182.850 ;
        RECT 614.100 181.050 615.900 182.850 ;
        RECT 617.100 181.050 618.000 184.800 ;
        RECT 635.700 185.400 639.300 186.300 ;
        RECT 632.100 181.050 633.900 182.850 ;
        RECT 635.700 181.050 636.900 185.400 ;
        RECT 638.100 181.050 639.900 182.850 ;
        RECT 656.400 181.050 657.300 191.400 ;
        RECT 674.100 188.400 675.900 194.400 ;
        RECT 677.100 189.000 678.900 195.000 ;
        RECT 683.700 194.400 684.900 195.000 ;
        RECT 680.100 191.400 681.900 194.400 ;
        RECT 683.100 191.400 684.900 194.400 ;
        RECT 698.100 191.400 699.900 195.000 ;
        RECT 701.100 191.400 702.900 194.400 ;
        RECT 704.100 191.400 705.900 195.000 ;
        RECT 719.100 191.400 720.900 195.000 ;
        RECT 722.100 191.400 723.900 194.400 ;
        RECT 725.100 191.400 726.900 195.000 ;
        RECT 674.100 181.050 675.000 188.400 ;
        RECT 680.700 187.200 681.600 191.400 ;
        RECT 676.200 186.300 681.600 187.200 ;
        RECT 688.950 186.450 691.050 187.050 ;
        RECT 697.950 186.450 700.050 187.050 ;
        RECT 676.200 185.400 678.300 186.300 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 628.950 178.950 631.050 181.050 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 674.100 178.950 676.200 181.050 ;
        RECT 581.550 176.550 586.050 178.050 ;
        RECT 587.100 177.150 588.900 178.950 ;
        RECT 582.000 175.950 586.050 176.550 ;
        RECT 593.700 171.600 594.900 178.950 ;
        RECT 611.100 177.150 612.900 178.950 ;
        RECT 545.400 165.900 552.000 166.800 ;
        RECT 545.400 165.600 546.900 165.900 ;
        RECT 485.100 159.000 486.900 165.000 ;
        RECT 488.100 159.600 489.900 165.600 ;
        RECT 491.100 159.000 492.900 165.600 ;
        RECT 503.100 159.000 504.900 165.600 ;
        RECT 506.100 159.600 507.900 165.600 ;
        RECT 509.100 159.000 510.900 165.600 ;
        RECT 524.100 159.000 525.900 165.600 ;
        RECT 527.100 159.600 528.900 165.600 ;
        RECT 542.100 159.000 543.900 165.600 ;
        RECT 545.100 159.600 546.900 165.600 ;
        RECT 551.100 165.600 552.000 165.900 ;
        RECT 569.400 165.900 576.000 166.800 ;
        RECT 569.400 165.600 570.900 165.900 ;
        RECT 548.100 159.000 549.900 165.000 ;
        RECT 551.100 159.600 552.900 165.600 ;
        RECT 566.100 159.000 567.900 165.600 ;
        RECT 569.100 159.600 570.900 165.600 ;
        RECT 575.100 165.600 576.000 165.900 ;
        RECT 572.100 159.000 573.900 165.000 ;
        RECT 575.100 159.600 576.900 165.600 ;
        RECT 587.400 159.000 589.200 171.600 ;
        RECT 592.500 170.100 594.900 171.600 ;
        RECT 592.500 159.600 594.300 170.100 ;
        RECT 595.200 167.100 597.000 168.900 ;
        RECT 617.100 166.800 618.000 178.950 ;
        RECT 629.100 177.150 630.900 178.950 ;
        RECT 635.700 171.600 636.900 178.950 ;
        RECT 653.250 177.150 655.050 178.950 ;
        RECT 656.400 171.600 657.300 178.950 ;
        RECT 659.100 177.150 660.900 178.950 ;
        RECT 675.000 171.600 676.200 178.950 ;
        RECT 677.400 174.900 678.300 185.400 ;
        RECT 688.950 185.550 700.050 186.450 ;
        RECT 688.950 184.950 691.050 185.550 ;
        RECT 697.950 184.950 700.050 185.550 ;
        RECT 682.800 181.050 684.600 182.850 ;
        RECT 701.700 181.050 702.600 191.400 ;
        RECT 722.700 181.050 723.600 191.400 ;
        RECT 737.700 187.200 739.500 194.400 ;
        RECT 742.800 188.400 744.600 195.000 ;
        RECT 737.700 186.300 741.900 187.200 ;
        RECT 737.100 181.050 738.900 182.850 ;
        RECT 740.700 181.050 741.900 186.300 ;
        RECT 742.950 186.450 745.050 187.050 ;
        RECT 751.950 186.450 754.050 187.050 ;
        RECT 742.950 185.550 754.050 186.450 ;
        RECT 758.100 186.600 759.900 194.400 ;
        RECT 762.600 188.400 764.400 195.000 ;
        RECT 765.600 190.200 767.400 194.400 ;
        RECT 765.600 188.400 768.300 190.200 ;
        RECT 764.700 186.600 766.500 187.500 ;
        RECT 758.100 185.700 766.500 186.600 ;
        RECT 742.950 184.950 745.050 185.550 ;
        RECT 751.950 184.950 754.050 185.550 ;
        RECT 742.950 181.050 744.750 182.850 ;
        RECT 758.250 181.050 760.050 182.850 ;
        RECT 679.500 178.950 681.600 181.050 ;
        RECT 682.800 178.950 684.900 181.050 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 718.950 178.950 721.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 758.100 178.950 760.200 181.050 ;
        RECT 679.200 177.150 681.000 178.950 ;
        RECT 698.100 177.150 699.900 178.950 ;
        RECT 677.100 174.300 678.900 174.900 ;
        RECT 677.100 173.100 684.900 174.300 ;
        RECT 683.700 171.600 684.900 173.100 ;
        RECT 701.700 171.600 702.600 178.950 ;
        RECT 703.950 177.150 705.750 178.950 ;
        RECT 719.100 177.150 720.900 178.950 ;
        RECT 722.700 171.600 723.600 178.950 ;
        RECT 724.950 177.150 726.750 178.950 ;
        RECT 724.950 174.450 727.050 175.050 ;
        RECT 736.950 174.450 739.050 174.750 ;
        RECT 724.950 173.550 739.050 174.450 ;
        RECT 724.950 172.950 727.050 173.550 ;
        RECT 736.950 172.650 739.050 173.550 ;
        RECT 611.400 165.900 618.000 166.800 ;
        RECT 611.400 165.600 612.900 165.900 ;
        RECT 595.500 159.000 597.300 165.600 ;
        RECT 608.100 159.000 609.900 165.600 ;
        RECT 611.100 159.600 612.900 165.600 ;
        RECT 617.100 165.600 618.000 165.900 ;
        RECT 614.100 159.000 615.900 165.000 ;
        RECT 617.100 159.600 618.900 165.600 ;
        RECT 629.400 159.000 631.200 171.600 ;
        RECT 634.500 170.100 636.900 171.600 ;
        RECT 634.500 159.600 636.300 170.100 ;
        RECT 637.200 167.100 639.000 168.900 ;
        RECT 637.500 159.000 639.300 165.600 ;
        RECT 653.100 159.000 654.900 171.600 ;
        RECT 656.400 170.400 660.000 171.600 ;
        RECT 658.200 159.600 660.000 170.400 ;
        RECT 675.000 170.100 677.400 171.600 ;
        RECT 675.600 159.600 677.400 170.100 ;
        RECT 678.600 159.000 680.400 171.600 ;
        RECT 683.100 159.600 684.900 171.600 ;
        RECT 699.000 170.400 702.600 171.600 ;
        RECT 699.000 159.600 700.800 170.400 ;
        RECT 704.100 159.000 705.900 171.600 ;
        RECT 720.000 170.400 723.600 171.600 ;
        RECT 720.000 159.600 721.800 170.400 ;
        RECT 725.100 159.000 726.900 171.600 ;
        RECT 740.700 165.600 741.900 178.950 ;
        RECT 745.950 177.450 748.050 178.050 ;
        RECT 754.950 177.450 757.050 178.050 ;
        RECT 745.950 176.550 757.050 177.450 ;
        RECT 745.950 175.950 748.050 176.550 ;
        RECT 754.950 175.950 757.050 176.550 ;
        RECT 751.950 174.450 754.050 174.900 ;
        RECT 757.950 174.450 760.050 175.050 ;
        RECT 751.950 173.550 760.050 174.450 ;
        RECT 751.950 172.800 754.050 173.550 ;
        RECT 757.950 172.950 760.050 173.550 ;
        RECT 742.950 171.450 745.050 172.050 ;
        RECT 754.950 171.450 757.050 171.900 ;
        RECT 742.950 170.550 757.050 171.450 ;
        RECT 742.950 169.950 745.050 170.550 ;
        RECT 754.950 169.800 757.050 170.550 ;
        RECT 761.100 165.600 762.000 185.700 ;
        RECT 767.400 181.050 768.300 188.400 ;
        RECT 779.100 189.300 780.900 194.400 ;
        RECT 782.100 190.200 783.900 195.000 ;
        RECT 785.100 189.300 786.900 194.400 ;
        RECT 779.100 187.950 786.900 189.300 ;
        RECT 788.100 188.400 789.900 194.400 ;
        RECT 803.100 189.300 804.900 194.400 ;
        RECT 806.100 190.200 807.900 195.000 ;
        RECT 809.100 189.300 810.900 194.400 ;
        RECT 788.100 186.300 789.300 188.400 ;
        RECT 803.100 187.950 810.900 189.300 ;
        RECT 812.100 188.400 813.900 194.400 ;
        RECT 812.100 186.300 813.300 188.400 ;
        RECT 827.700 187.200 829.500 194.400 ;
        RECT 832.800 188.400 834.600 195.000 ;
        RECT 845.100 189.300 846.900 194.400 ;
        RECT 848.100 190.200 849.900 195.000 ;
        RECT 851.100 189.300 852.900 194.400 ;
        RECT 845.100 187.950 852.900 189.300 ;
        RECT 854.100 188.400 855.900 194.400 ;
        RECT 869.700 191.400 871.500 195.000 ;
        RECT 872.700 189.600 874.500 194.400 ;
        RECT 869.400 188.400 874.500 189.600 ;
        RECT 877.200 188.400 879.000 195.000 ;
        RECT 890.100 188.400 891.900 194.400 ;
        RECT 827.700 186.300 831.900 187.200 ;
        RECT 854.100 186.300 855.300 188.400 ;
        RECT 785.700 185.400 789.300 186.300 ;
        RECT 809.700 185.400 813.300 186.300 ;
        RECT 782.100 181.050 783.900 182.850 ;
        RECT 785.700 181.050 786.900 185.400 ;
        RECT 790.950 183.450 793.050 184.050 ;
        RECT 788.100 181.050 789.900 182.850 ;
        RECT 790.950 182.550 798.450 183.450 ;
        RECT 790.950 181.950 793.050 182.550 ;
        RECT 763.500 178.950 765.600 181.050 ;
        RECT 766.800 178.950 768.900 181.050 ;
        RECT 778.950 178.950 781.050 181.050 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 763.200 177.150 765.000 178.950 ;
        RECT 767.400 171.600 768.300 178.950 ;
        RECT 779.100 177.150 780.900 178.950 ;
        RECT 785.700 171.600 786.900 178.950 ;
        RECT 797.550 177.450 798.450 182.550 ;
        RECT 806.100 181.050 807.900 182.850 ;
        RECT 809.700 181.050 810.900 185.400 ;
        RECT 812.100 181.050 813.900 182.850 ;
        RECT 827.100 181.050 828.900 182.850 ;
        RECT 830.700 181.050 831.900 186.300 ;
        RECT 851.700 185.400 855.300 186.300 ;
        RECT 840.000 183.450 844.050 184.050 ;
        RECT 832.950 181.050 834.750 182.850 ;
        RECT 839.550 181.950 844.050 183.450 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 797.550 177.000 801.450 177.450 ;
        RECT 803.100 177.150 804.900 178.950 ;
        RECT 797.550 176.550 802.050 177.000 ;
        RECT 799.950 172.950 802.050 176.550 ;
        RECT 809.700 171.600 810.900 178.950 ;
        RECT 737.100 159.000 738.900 165.600 ;
        RECT 740.100 159.600 741.900 165.600 ;
        RECT 743.100 159.000 744.900 165.600 ;
        RECT 758.100 159.000 759.900 165.600 ;
        RECT 761.100 159.600 762.900 165.600 ;
        RECT 764.100 159.000 765.900 171.000 ;
        RECT 767.100 159.600 768.900 171.600 ;
        RECT 779.400 159.000 781.200 171.600 ;
        RECT 784.500 170.100 786.900 171.600 ;
        RECT 784.500 159.600 786.300 170.100 ;
        RECT 787.200 167.100 789.000 168.900 ;
        RECT 787.500 159.000 789.300 165.600 ;
        RECT 803.400 159.000 805.200 171.600 ;
        RECT 808.500 170.100 810.900 171.600 ;
        RECT 808.500 159.600 810.300 170.100 ;
        RECT 811.200 167.100 813.000 168.900 ;
        RECT 830.700 165.600 831.900 178.950 ;
        RECT 839.550 178.050 840.450 181.950 ;
        RECT 848.100 181.050 849.900 182.850 ;
        RECT 851.700 181.050 852.900 185.400 ;
        RECT 864.000 183.450 868.050 184.050 ;
        RECT 854.100 181.050 855.900 182.850 ;
        RECT 863.550 181.950 868.050 183.450 ;
        RECT 844.950 178.950 847.050 181.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 835.950 176.550 840.450 178.050 ;
        RECT 845.100 177.150 846.900 178.950 ;
        RECT 835.950 175.950 840.000 176.550 ;
        RECT 851.700 171.600 852.900 178.950 ;
        RECT 863.550 178.050 864.450 181.950 ;
        RECT 869.400 181.050 870.300 188.400 ;
        RECT 890.700 186.300 891.900 188.400 ;
        RECT 893.100 189.300 894.900 194.400 ;
        RECT 896.100 190.200 897.900 195.000 ;
        RECT 899.100 189.300 900.900 194.400 ;
        RECT 893.100 187.950 900.900 189.300 ;
        RECT 911.100 189.300 912.900 194.400 ;
        RECT 914.100 190.200 915.900 195.000 ;
        RECT 917.100 189.300 918.900 194.400 ;
        RECT 911.100 187.950 918.900 189.300 ;
        RECT 920.100 188.400 921.900 194.400 ;
        RECT 890.700 185.400 894.300 186.300 ;
        RECT 871.950 181.050 873.750 182.850 ;
        RECT 878.100 181.050 879.900 182.850 ;
        RECT 890.100 181.050 891.900 182.850 ;
        RECT 893.100 181.050 894.300 185.400 ;
        RECT 904.950 184.950 907.050 187.050 ;
        RECT 920.100 186.300 921.300 188.400 ;
        RECT 917.700 185.400 921.300 186.300 ;
        RECT 937.500 186.000 939.300 194.400 ;
        RECT 896.100 181.050 897.900 182.850 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 889.950 178.950 892.050 181.050 ;
        RECT 892.950 178.950 895.050 181.050 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 863.550 176.550 868.050 178.050 ;
        RECT 864.000 175.950 868.050 176.550 ;
        RECT 869.400 171.600 870.300 178.950 ;
        RECT 874.950 177.150 876.750 178.950 ;
        RECT 871.950 174.450 874.050 174.750 ;
        RECT 883.950 174.450 886.050 175.050 ;
        RECT 871.950 173.550 886.050 174.450 ;
        RECT 871.950 172.650 874.050 173.550 ;
        RECT 883.950 172.950 886.050 173.550 ;
        RECT 893.100 171.600 894.300 178.950 ;
        RECT 899.100 177.150 900.900 178.950 ;
        RECT 905.550 178.050 906.450 184.950 ;
        RECT 914.100 181.050 915.900 182.850 ;
        RECT 917.700 181.050 918.900 185.400 ;
        RECT 936.000 184.800 939.300 186.000 ;
        RECT 944.100 185.400 945.900 195.000 ;
        RECT 930.000 183.450 934.050 184.050 ;
        RECT 920.100 181.050 921.900 182.850 ;
        RECT 929.550 181.950 934.050 183.450 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 913.950 178.950 916.050 181.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 905.550 176.550 910.050 178.050 ;
        RECT 911.100 177.150 912.900 178.950 ;
        RECT 906.000 175.950 910.050 176.550 ;
        RECT 917.700 171.600 918.900 178.950 ;
        RECT 929.550 178.050 930.450 181.950 ;
        RECT 936.000 181.050 936.900 184.800 ;
        RECT 938.100 181.050 939.900 182.850 ;
        RECT 944.100 181.050 945.900 182.850 ;
        RECT 934.950 178.950 937.050 181.050 ;
        RECT 937.950 178.950 940.050 181.050 ;
        RECT 940.950 178.950 943.050 181.050 ;
        RECT 943.950 178.950 946.050 181.050 ;
        RECT 929.550 176.550 934.050 178.050 ;
        RECT 930.000 175.950 934.050 176.550 ;
        RECT 811.500 159.000 813.300 165.600 ;
        RECT 827.100 159.000 828.900 165.600 ;
        RECT 830.100 159.600 831.900 165.600 ;
        RECT 833.100 159.000 834.900 165.600 ;
        RECT 845.400 159.000 847.200 171.600 ;
        RECT 850.500 170.100 852.900 171.600 ;
        RECT 850.500 159.600 852.300 170.100 ;
        RECT 853.200 167.100 855.000 168.900 ;
        RECT 853.500 159.000 855.300 165.600 ;
        RECT 869.100 159.600 870.900 171.600 ;
        RECT 872.100 170.700 879.900 171.600 ;
        RECT 872.100 159.600 873.900 170.700 ;
        RECT 875.100 159.000 876.900 169.800 ;
        RECT 878.100 159.600 879.900 170.700 ;
        RECT 893.100 170.100 895.500 171.600 ;
        RECT 891.000 167.100 892.800 168.900 ;
        RECT 890.700 159.000 892.500 165.600 ;
        RECT 893.700 159.600 895.500 170.100 ;
        RECT 898.800 159.000 900.600 171.600 ;
        RECT 911.400 159.000 913.200 171.600 ;
        RECT 916.500 170.100 918.900 171.600 ;
        RECT 916.500 159.600 918.300 170.100 ;
        RECT 919.200 167.100 921.000 168.900 ;
        RECT 936.000 166.800 936.900 178.950 ;
        RECT 941.100 177.150 942.900 178.950 ;
        RECT 936.000 165.900 942.600 166.800 ;
        RECT 936.000 165.600 936.900 165.900 ;
        RECT 919.500 159.000 921.300 165.600 ;
        RECT 935.100 159.600 936.900 165.600 ;
        RECT 941.100 165.600 942.600 165.900 ;
        RECT 938.100 159.000 939.900 165.000 ;
        RECT 941.100 159.600 942.900 165.600 ;
        RECT 944.100 159.000 945.900 165.600 ;
        RECT 14.100 144.300 15.900 155.400 ;
        RECT 17.100 145.200 18.900 156.000 ;
        RECT 20.100 144.300 21.900 155.400 ;
        RECT 14.100 143.400 21.900 144.300 ;
        RECT 23.100 143.400 24.900 155.400 ;
        RECT 38.100 149.400 39.900 156.000 ;
        RECT 41.100 149.400 42.900 155.400 ;
        RECT 44.100 150.000 45.900 156.000 ;
        RECT 41.400 149.100 42.900 149.400 ;
        RECT 47.100 149.400 48.900 155.400 ;
        RECT 62.100 149.400 63.900 155.400 ;
        RECT 65.100 150.000 66.900 156.000 ;
        RECT 47.100 149.100 48.000 149.400 ;
        RECT 41.400 148.200 48.000 149.100 ;
        RECT 17.250 136.050 19.050 137.850 ;
        RECT 23.700 136.050 24.600 143.400 ;
        RECT 28.950 141.450 31.050 142.050 ;
        RECT 43.950 141.450 46.050 142.050 ;
        RECT 28.950 140.550 46.050 141.450 ;
        RECT 28.950 139.950 31.050 140.550 ;
        RECT 43.950 139.950 46.050 140.550 ;
        RECT 33.000 138.450 37.050 139.050 ;
        RECT 32.550 136.950 37.050 138.450 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 14.100 132.150 15.900 133.950 ;
        RECT 20.250 132.150 22.050 133.950 ;
        RECT 23.700 126.600 24.600 133.950 ;
        RECT 25.950 132.450 28.050 133.050 ;
        RECT 32.550 132.450 33.450 136.950 ;
        RECT 41.100 136.050 42.900 137.850 ;
        RECT 47.100 136.050 48.000 148.200 ;
        RECT 63.000 149.100 63.900 149.400 ;
        RECT 68.100 149.400 69.900 155.400 ;
        RECT 71.100 149.400 72.900 156.000 ;
        RECT 68.100 149.100 69.600 149.400 ;
        RECT 63.000 148.200 69.600 149.100 ;
        RECT 57.000 138.450 61.050 139.050 ;
        RECT 56.550 136.950 61.050 138.450 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 43.950 133.950 46.050 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 25.950 131.550 33.450 132.450 ;
        RECT 38.100 132.150 39.900 133.950 ;
        RECT 44.100 132.150 45.900 133.950 ;
        RECT 25.950 130.950 28.050 131.550 ;
        RECT 47.100 130.200 48.000 133.950 ;
        RECT 56.550 133.050 57.450 136.950 ;
        RECT 63.000 136.050 63.900 148.200 ;
        RECT 84.600 144.900 86.400 155.400 ;
        RECT 84.000 143.400 86.400 144.900 ;
        RECT 87.600 143.400 89.400 156.000 ;
        RECT 92.100 143.400 93.900 155.400 ;
        RECT 104.100 143.400 105.900 155.400 ;
        RECT 107.100 144.300 108.900 155.400 ;
        RECT 110.100 145.200 111.900 156.000 ;
        RECT 113.100 144.300 114.900 155.400 ;
        RECT 125.100 149.400 126.900 156.000 ;
        RECT 128.100 149.400 129.900 155.400 ;
        RECT 131.100 150.000 132.900 156.000 ;
        RECT 128.400 149.100 129.900 149.400 ;
        RECT 134.100 149.400 135.900 155.400 ;
        RECT 134.100 149.100 135.000 149.400 ;
        RECT 128.400 148.200 135.000 149.100 ;
        RECT 107.100 143.400 114.900 144.300 ;
        RECT 64.950 141.450 67.050 142.050 ;
        RECT 79.950 141.450 82.050 142.050 ;
        RECT 64.950 140.550 82.050 141.450 ;
        RECT 64.950 139.950 67.050 140.550 ;
        RECT 79.950 139.950 82.050 140.550 ;
        RECT 68.100 136.050 69.900 137.850 ;
        RECT 84.000 136.050 85.200 143.400 ;
        RECT 92.700 141.900 93.900 143.400 ;
        RECT 86.100 140.700 93.900 141.900 ;
        RECT 86.100 140.100 87.900 140.700 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 83.100 133.950 85.200 136.050 ;
        RECT 56.550 131.550 61.050 133.050 ;
        RECT 57.000 130.950 61.050 131.550 ;
        RECT 15.000 120.000 16.800 126.600 ;
        RECT 19.500 125.400 24.600 126.600 ;
        RECT 19.500 120.600 21.300 125.400 ;
        RECT 22.500 120.000 24.300 123.600 ;
        RECT 38.100 120.000 39.900 129.600 ;
        RECT 44.700 129.000 48.000 130.200 ;
        RECT 63.000 130.200 63.900 133.950 ;
        RECT 65.100 132.150 66.900 133.950 ;
        RECT 71.100 132.150 72.900 133.950 ;
        RECT 63.000 129.000 66.300 130.200 ;
        RECT 44.700 120.600 46.500 129.000 ;
        RECT 64.500 120.600 66.300 129.000 ;
        RECT 71.100 120.000 72.900 129.600 ;
        RECT 83.100 126.600 84.000 133.950 ;
        RECT 86.400 129.600 87.300 140.100 ;
        RECT 88.200 136.050 90.000 137.850 ;
        RECT 104.400 136.050 105.300 143.400 ;
        RECT 109.950 136.050 111.750 137.850 ;
        RECT 128.100 136.050 129.900 137.850 ;
        RECT 134.100 136.050 135.000 148.200 ;
        RECT 146.100 143.400 147.900 155.400 ;
        RECT 149.100 144.000 150.900 156.000 ;
        RECT 152.100 149.400 153.900 155.400 ;
        RECT 155.100 149.400 156.900 156.000 ;
        RECT 170.100 149.400 171.900 156.000 ;
        RECT 173.100 149.400 174.900 155.400 ;
        RECT 176.100 149.400 177.900 156.000 ;
        RECT 146.700 136.050 147.600 143.400 ;
        RECT 150.000 136.050 151.800 137.850 ;
        RECT 88.500 133.950 90.600 136.050 ;
        RECT 91.800 133.950 93.900 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 146.100 133.950 148.200 136.050 ;
        RECT 149.400 133.950 151.500 136.050 ;
        RECT 91.800 132.150 93.600 133.950 ;
        RECT 85.200 128.700 87.300 129.600 ;
        RECT 85.200 127.800 90.600 128.700 ;
        RECT 83.100 120.600 84.900 126.600 ;
        RECT 86.100 120.000 87.900 126.000 ;
        RECT 89.700 123.600 90.600 127.800 ;
        RECT 104.400 126.600 105.300 133.950 ;
        RECT 106.950 132.150 108.750 133.950 ;
        RECT 113.100 132.150 114.900 133.950 ;
        RECT 125.100 132.150 126.900 133.950 ;
        RECT 131.100 132.150 132.900 133.950 ;
        RECT 134.100 130.200 135.000 133.950 ;
        RECT 104.400 125.400 109.500 126.600 ;
        RECT 89.100 120.600 90.900 123.600 ;
        RECT 92.100 120.600 93.900 123.600 ;
        RECT 92.700 120.000 93.900 120.600 ;
        RECT 104.700 120.000 106.500 123.600 ;
        RECT 107.700 120.600 109.500 125.400 ;
        RECT 112.200 120.000 114.000 126.600 ;
        RECT 125.100 120.000 126.900 129.600 ;
        RECT 131.700 129.000 135.000 130.200 ;
        RECT 131.700 120.600 133.500 129.000 ;
        RECT 146.700 126.600 147.600 133.950 ;
        RECT 153.000 129.300 153.900 149.400 ;
        RECT 173.700 136.050 174.900 149.400 ;
        RECT 188.100 143.400 189.900 155.400 ;
        RECT 191.100 144.000 192.900 156.000 ;
        RECT 194.100 149.400 195.900 155.400 ;
        RECT 197.100 149.400 198.900 156.000 ;
        RECT 212.100 149.400 213.900 156.000 ;
        RECT 215.100 149.400 216.900 155.400 ;
        RECT 218.100 150.000 219.900 156.000 ;
        RECT 188.700 136.050 189.600 143.400 ;
        RECT 192.000 136.050 193.800 137.850 ;
        RECT 154.800 133.950 156.900 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 188.100 133.950 190.200 136.050 ;
        RECT 191.400 133.950 193.500 136.050 ;
        RECT 154.950 132.150 156.750 133.950 ;
        RECT 170.100 132.150 171.900 133.950 ;
        RECT 148.500 128.400 156.900 129.300 ;
        RECT 173.700 128.700 174.900 133.950 ;
        RECT 175.950 132.150 177.750 133.950 ;
        RECT 148.500 127.500 150.300 128.400 ;
        RECT 146.700 124.800 149.400 126.600 ;
        RECT 147.600 120.600 149.400 124.800 ;
        RECT 150.600 120.000 152.400 126.600 ;
        RECT 155.100 120.600 156.900 128.400 ;
        RECT 170.700 127.800 174.900 128.700 ;
        RECT 170.700 120.600 172.500 127.800 ;
        RECT 188.700 126.600 189.600 133.950 ;
        RECT 195.000 129.300 195.900 149.400 ;
        RECT 215.400 149.100 216.900 149.400 ;
        RECT 221.100 149.400 222.900 155.400 ;
        RECT 221.100 149.100 222.000 149.400 ;
        RECT 215.400 148.200 222.000 149.100 ;
        RECT 215.100 136.050 216.900 137.850 ;
        RECT 221.100 136.050 222.000 148.200 ;
        RECT 236.400 143.400 238.200 156.000 ;
        RECT 241.500 144.900 243.300 155.400 ;
        RECT 244.500 149.400 246.300 156.000 ;
        RECT 257.100 149.400 258.900 156.000 ;
        RECT 260.100 149.400 261.900 155.400 ;
        RECT 263.100 150.000 264.900 156.000 ;
        RECT 260.400 149.100 261.900 149.400 ;
        RECT 266.100 149.400 267.900 155.400 ;
        RECT 266.100 149.100 267.000 149.400 ;
        RECT 260.400 148.200 267.000 149.100 ;
        RECT 244.200 146.100 246.000 147.900 ;
        RECT 241.500 143.400 243.900 144.900 ;
        RECT 236.100 136.050 237.900 137.850 ;
        RECT 242.700 136.050 243.900 143.400 ;
        RECT 247.950 141.450 250.050 141.900 ;
        RECT 262.950 141.450 265.050 142.050 ;
        RECT 247.950 140.550 265.050 141.450 ;
        RECT 247.950 139.800 250.050 140.550 ;
        RECT 262.950 139.950 265.050 140.550 ;
        RECT 260.100 136.050 261.900 137.850 ;
        RECT 266.100 136.050 267.000 148.200 ;
        RECT 281.100 144.300 282.900 155.400 ;
        RECT 284.100 145.500 285.900 156.000 ;
        RECT 288.600 144.300 290.400 155.400 ;
        RECT 292.800 145.500 294.900 156.000 ;
        RECT 296.100 144.600 297.900 155.400 ;
        RECT 308.100 149.400 309.900 156.000 ;
        RECT 311.100 149.400 312.900 155.400 ;
        RECT 314.100 149.400 315.900 156.000 ;
        RECT 281.100 143.100 285.900 144.300 ;
        RECT 288.600 143.400 291.900 144.300 ;
        RECT 283.800 142.200 285.900 143.100 ;
        RECT 271.950 141.450 274.050 142.050 ;
        RECT 277.950 141.450 280.050 142.050 ;
        RECT 271.950 140.550 280.050 141.450 ;
        RECT 283.800 141.300 289.200 142.200 ;
        RECT 271.950 139.950 274.050 140.550 ;
        RECT 277.950 139.950 280.050 140.550 ;
        RECT 287.400 139.500 289.200 141.300 ;
        RECT 290.700 139.050 291.900 143.400 ;
        RECT 292.800 143.400 297.900 144.600 ;
        RECT 292.800 142.500 294.900 143.400 ;
        RECT 290.100 138.300 292.200 139.050 ;
        RECT 285.900 136.200 287.700 138.000 ;
        RECT 289.200 136.950 292.200 138.300 ;
        RECT 196.800 133.950 198.900 136.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 196.950 132.150 198.750 133.950 ;
        RECT 212.100 132.150 213.900 133.950 ;
        RECT 218.100 132.150 219.900 133.950 ;
        RECT 221.100 130.200 222.000 133.950 ;
        RECT 239.100 132.150 240.900 133.950 ;
        RECT 190.500 128.400 198.900 129.300 ;
        RECT 190.500 127.500 192.300 128.400 ;
        RECT 175.800 120.000 177.600 126.600 ;
        RECT 188.700 124.800 191.400 126.600 ;
        RECT 189.600 120.600 191.400 124.800 ;
        RECT 192.600 120.000 194.400 126.600 ;
        RECT 197.100 120.600 198.900 128.400 ;
        RECT 199.950 123.450 202.050 124.050 ;
        RECT 208.950 123.450 211.050 124.050 ;
        RECT 199.950 122.550 211.050 123.450 ;
        RECT 199.950 121.950 202.050 122.550 ;
        RECT 208.950 121.950 211.050 122.550 ;
        RECT 212.100 120.000 213.900 129.600 ;
        RECT 218.700 129.000 222.000 130.200 ;
        RECT 242.700 129.600 243.900 133.950 ;
        RECT 245.100 132.150 246.900 133.950 ;
        RECT 257.100 132.150 258.900 133.950 ;
        RECT 263.100 132.150 264.900 133.950 ;
        RECT 266.100 130.200 267.000 133.950 ;
        RECT 281.100 133.800 283.200 136.050 ;
        RECT 285.900 134.100 288.000 136.200 ;
        RECT 281.400 133.200 283.200 133.800 ;
        RECT 281.400 132.000 288.000 133.200 ;
        RECT 285.900 131.100 288.000 132.000 ;
        RECT 218.700 120.600 220.500 129.000 ;
        RECT 242.700 128.700 246.300 129.600 ;
        RECT 236.100 125.700 243.900 127.050 ;
        RECT 236.100 120.600 237.900 125.700 ;
        RECT 239.100 120.000 240.900 124.800 ;
        RECT 242.100 120.600 243.900 125.700 ;
        RECT 245.100 126.600 246.300 128.700 ;
        RECT 245.100 120.600 246.900 126.600 ;
        RECT 257.100 120.000 258.900 129.600 ;
        RECT 263.700 129.000 267.000 130.200 ;
        RECT 283.500 129.000 285.600 129.600 ;
        RECT 286.500 129.300 288.300 131.100 ;
        RECT 289.200 130.200 290.100 136.950 ;
        RECT 295.800 136.050 297.600 137.850 ;
        RECT 311.700 136.050 312.900 149.400 ;
        RECT 330.000 144.600 331.800 155.400 ;
        RECT 330.000 143.400 333.600 144.600 ;
        RECT 335.100 143.400 336.900 156.000 ;
        RECT 350.100 149.400 351.900 155.400 ;
        RECT 353.100 150.000 354.900 156.000 ;
        RECT 351.000 149.100 351.900 149.400 ;
        RECT 356.100 149.400 357.900 155.400 ;
        RECT 359.100 149.400 360.900 156.000 ;
        RECT 374.100 149.400 375.900 156.000 ;
        RECT 377.100 149.400 378.900 155.400 ;
        RECT 380.100 149.400 381.900 156.000 ;
        RECT 392.100 149.400 393.900 156.000 ;
        RECT 395.100 149.400 396.900 155.400 ;
        RECT 356.100 149.100 357.600 149.400 ;
        RECT 351.000 148.200 357.600 149.100 ;
        RECT 329.100 136.050 330.900 137.850 ;
        RECT 332.700 136.050 333.600 143.400 ;
        RECT 334.950 141.450 339.000 142.050 ;
        RECT 334.950 139.950 339.450 141.450 ;
        RECT 338.550 138.450 339.450 139.950 ;
        RECT 334.950 136.050 336.750 137.850 ;
        RECT 338.550 137.550 342.450 138.450 ;
        RECT 291.000 134.100 292.800 135.900 ;
        RECT 291.000 132.000 293.100 134.100 ;
        RECT 295.800 133.950 297.900 136.050 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 328.950 133.950 331.050 136.050 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 308.100 132.150 309.900 133.950 ;
        RECT 263.700 120.600 265.500 129.000 ;
        RECT 281.100 127.500 285.600 129.000 ;
        RECT 289.200 128.100 292.200 130.200 ;
        RECT 281.100 126.600 282.600 127.500 ;
        RECT 281.100 120.600 282.900 126.600 ;
        RECT 289.200 126.000 290.100 128.100 ;
        RECT 293.400 127.500 295.500 129.900 ;
        RECT 311.700 128.700 312.900 133.950 ;
        RECT 313.950 132.150 315.750 133.950 ;
        RECT 322.950 130.050 325.050 133.050 ;
        RECT 321.000 129.900 325.050 130.050 ;
        RECT 308.700 127.800 312.900 128.700 ;
        RECT 319.950 129.000 325.050 129.900 ;
        RECT 319.950 128.550 324.450 129.000 ;
        RECT 319.950 127.950 324.000 128.550 ;
        RECT 319.950 127.800 322.050 127.950 ;
        RECT 293.400 126.600 297.900 127.500 ;
        RECT 284.100 120.000 285.900 125.700 ;
        RECT 288.300 120.600 290.100 126.000 ;
        RECT 292.800 120.000 294.600 125.700 ;
        RECT 296.100 120.600 297.900 126.600 ;
        RECT 308.700 120.600 310.500 127.800 ;
        RECT 313.800 120.000 315.600 126.600 ;
        RECT 332.700 123.600 333.600 133.950 ;
        RECT 334.950 129.450 337.050 130.050 ;
        RECT 341.550 129.450 342.450 137.550 ;
        RECT 351.000 136.050 351.900 148.200 ;
        RECT 369.000 138.450 373.050 139.050 ;
        RECT 356.100 136.050 357.900 137.850 ;
        RECT 368.550 136.950 373.050 138.450 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 352.950 133.950 355.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 334.950 128.550 342.450 129.450 ;
        RECT 351.000 130.200 351.900 133.950 ;
        RECT 353.100 132.150 354.900 133.950 ;
        RECT 359.100 132.150 360.900 133.950 ;
        RECT 368.550 133.050 369.450 136.950 ;
        RECT 377.100 136.050 378.300 149.400 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 392.100 133.950 394.200 136.050 ;
        RECT 368.550 131.550 373.050 133.050 ;
        RECT 374.250 132.150 376.050 133.950 ;
        RECT 369.000 130.950 373.050 131.550 ;
        RECT 351.000 129.000 354.300 130.200 ;
        RECT 334.950 127.950 337.050 128.550 ;
        RECT 334.950 126.450 337.050 126.900 ;
        RECT 346.950 126.450 349.050 127.050 ;
        RECT 334.950 125.550 349.050 126.450 ;
        RECT 334.950 124.800 337.050 125.550 ;
        RECT 346.950 124.950 349.050 125.550 ;
        RECT 329.100 120.000 330.900 123.600 ;
        RECT 332.100 120.600 333.900 123.600 ;
        RECT 335.100 120.000 336.900 123.600 ;
        RECT 352.500 120.600 354.300 129.000 ;
        RECT 359.100 120.000 360.900 129.600 ;
        RECT 364.950 129.450 367.050 130.050 ;
        RECT 373.950 129.450 376.050 130.050 ;
        RECT 364.950 128.550 376.050 129.450 ;
        RECT 364.950 127.950 367.050 128.550 ;
        RECT 373.950 127.950 376.050 128.550 ;
        RECT 377.100 128.700 378.300 133.950 ;
        RECT 380.100 132.150 381.900 133.950 ;
        RECT 392.250 132.150 394.050 133.950 ;
        RECT 395.100 129.300 396.000 149.400 ;
        RECT 398.100 144.000 399.900 156.000 ;
        RECT 401.100 143.400 402.900 155.400 ;
        RECT 413.100 149.400 414.900 155.400 ;
        RECT 416.100 150.000 417.900 156.000 ;
        RECT 414.000 149.100 414.900 149.400 ;
        RECT 419.100 149.400 420.900 155.400 ;
        RECT 422.100 149.400 423.900 156.000 ;
        RECT 437.100 149.400 438.900 156.000 ;
        RECT 440.100 149.400 441.900 155.400 ;
        RECT 455.700 149.400 457.500 156.000 ;
        RECT 419.100 149.100 420.600 149.400 ;
        RECT 414.000 148.200 420.600 149.100 ;
        RECT 397.200 136.050 399.000 137.850 ;
        RECT 401.400 136.050 402.300 143.400 ;
        RECT 414.000 136.050 414.900 148.200 ;
        RECT 421.950 141.450 424.050 141.900 ;
        RECT 433.950 141.450 436.050 142.050 ;
        RECT 421.950 140.550 436.050 141.450 ;
        RECT 421.950 139.800 424.050 140.550 ;
        RECT 433.950 139.950 436.050 140.550 ;
        RECT 419.100 136.050 420.900 137.850 ;
        RECT 437.100 136.050 438.900 137.850 ;
        RECT 440.100 136.050 441.300 149.400 ;
        RECT 456.000 146.100 457.800 147.900 ;
        RECT 458.700 144.900 460.500 155.400 ;
        RECT 458.100 143.400 460.500 144.900 ;
        RECT 463.800 143.400 465.600 156.000 ;
        RECT 476.100 149.400 477.900 156.000 ;
        RECT 479.100 149.400 480.900 155.400 ;
        RECT 482.100 150.000 483.900 156.000 ;
        RECT 479.400 149.100 480.900 149.400 ;
        RECT 485.100 149.400 486.900 155.400 ;
        RECT 485.100 149.100 486.000 149.400 ;
        RECT 479.400 148.200 486.000 149.100 ;
        RECT 442.950 138.450 445.050 139.050 ;
        RECT 451.950 138.450 454.050 139.050 ;
        RECT 442.950 137.550 454.050 138.450 ;
        RECT 442.950 136.950 445.050 137.550 ;
        RECT 451.950 136.950 454.050 137.550 ;
        RECT 458.100 136.050 459.300 143.400 ;
        RECT 460.950 141.450 463.050 142.050 ;
        RECT 475.950 141.450 478.050 142.200 ;
        RECT 460.950 140.550 478.050 141.450 ;
        RECT 460.950 139.950 463.050 140.550 ;
        RECT 475.950 140.100 478.050 140.550 ;
        RECT 466.950 138.450 471.000 139.050 ;
        RECT 466.950 138.000 471.450 138.450 ;
        RECT 464.100 136.050 465.900 137.850 ;
        RECT 466.950 136.950 472.050 138.000 ;
        RECT 397.500 133.950 399.600 136.050 ;
        RECT 400.800 133.950 402.900 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 457.950 133.950 460.050 136.050 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 377.100 127.800 381.300 128.700 ;
        RECT 374.400 120.000 376.200 126.600 ;
        RECT 379.500 120.600 381.300 127.800 ;
        RECT 392.100 128.400 400.500 129.300 ;
        RECT 392.100 120.600 393.900 128.400 ;
        RECT 398.700 127.500 400.500 128.400 ;
        RECT 401.400 126.600 402.300 133.950 ;
        RECT 414.000 130.200 414.900 133.950 ;
        RECT 416.100 132.150 417.900 133.950 ;
        RECT 422.100 132.150 423.900 133.950 ;
        RECT 427.950 132.450 430.050 133.050 ;
        RECT 433.950 132.450 436.050 133.050 ;
        RECT 427.950 131.550 436.050 132.450 ;
        RECT 427.950 130.950 430.050 131.550 ;
        RECT 433.950 130.950 436.050 131.550 ;
        RECT 414.000 129.000 417.300 130.200 ;
        RECT 396.600 120.000 398.400 126.600 ;
        RECT 399.600 124.800 402.300 126.600 ;
        RECT 399.600 120.600 401.400 124.800 ;
        RECT 415.500 120.600 417.300 129.000 ;
        RECT 422.100 120.000 423.900 129.600 ;
        RECT 440.100 123.600 441.300 133.950 ;
        RECT 455.100 132.150 456.900 133.950 ;
        RECT 458.100 129.600 459.300 133.950 ;
        RECT 461.100 132.150 462.900 133.950 ;
        RECT 469.950 133.800 472.050 136.950 ;
        RECT 479.100 136.050 480.900 137.850 ;
        RECT 485.100 136.050 486.000 148.200 ;
        RECT 497.100 144.300 498.900 155.400 ;
        RECT 500.100 145.200 501.900 156.000 ;
        RECT 503.100 144.300 504.900 155.400 ;
        RECT 497.100 143.400 504.900 144.300 ;
        RECT 506.100 143.400 507.900 155.400 ;
        RECT 521.400 143.400 523.200 156.000 ;
        RECT 526.500 144.900 528.300 155.400 ;
        RECT 529.500 149.400 531.300 156.000 ;
        RECT 529.200 146.100 531.000 147.900 ;
        RECT 526.500 143.400 528.900 144.900 ;
        RECT 545.400 143.400 547.200 156.000 ;
        RECT 550.500 144.900 552.300 155.400 ;
        RECT 553.500 149.400 555.300 156.000 ;
        RECT 553.200 146.100 555.000 147.900 ;
        RECT 550.500 143.400 552.900 144.900 ;
        RECT 569.100 144.600 570.900 155.400 ;
        RECT 572.100 145.500 573.900 156.000 ;
        RECT 575.100 154.500 582.900 155.400 ;
        RECT 575.100 144.600 576.900 154.500 ;
        RECT 569.100 143.700 576.900 144.600 ;
        RECT 500.250 136.050 502.050 137.850 ;
        RECT 506.700 136.050 507.600 143.400 ;
        RECT 521.100 136.050 522.900 137.850 ;
        RECT 527.700 136.050 528.900 143.400 ;
        RECT 545.100 136.050 546.900 137.850 ;
        RECT 551.700 136.050 552.900 143.400 ;
        RECT 578.100 142.500 579.900 153.600 ;
        RECT 581.100 143.400 582.900 154.500 ;
        RECT 596.100 149.400 597.900 156.000 ;
        RECT 599.100 149.400 600.900 155.400 ;
        RECT 602.100 150.000 603.900 156.000 ;
        RECT 599.400 149.100 600.900 149.400 ;
        RECT 605.100 149.400 606.900 155.400 ;
        RECT 620.100 149.400 621.900 156.000 ;
        RECT 623.100 149.400 624.900 155.400 ;
        RECT 626.100 150.000 627.900 156.000 ;
        RECT 605.100 149.100 606.000 149.400 ;
        RECT 599.400 148.200 606.000 149.100 ;
        RECT 623.400 149.100 624.900 149.400 ;
        RECT 629.100 149.400 630.900 155.400 ;
        RECT 629.100 149.100 630.000 149.400 ;
        RECT 623.400 148.200 630.000 149.100 ;
        RECT 575.100 141.600 579.900 142.500 ;
        RECT 572.250 136.050 574.050 137.850 ;
        RECT 575.100 136.050 576.000 141.600 ;
        RECT 601.950 141.450 604.050 142.050 ;
        RECT 593.550 140.550 604.050 141.450 ;
        RECT 593.550 138.450 594.450 140.550 ;
        RECT 601.950 139.950 604.050 140.550 ;
        RECT 578.100 136.050 579.900 137.850 ;
        RECT 590.550 137.550 594.450 138.450 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 481.950 133.950 484.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 499.950 133.950 502.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 526.950 133.950 529.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 476.100 132.150 477.900 133.950 ;
        RECT 482.100 132.150 483.900 133.950 ;
        RECT 485.100 130.200 486.000 133.950 ;
        RECT 497.100 132.150 498.900 133.950 ;
        RECT 503.250 132.150 505.050 133.950 ;
        RECT 455.700 128.700 459.300 129.600 ;
        RECT 455.700 126.600 456.900 128.700 ;
        RECT 437.100 120.000 438.900 123.600 ;
        RECT 440.100 120.600 441.900 123.600 ;
        RECT 455.100 120.600 456.900 126.600 ;
        RECT 458.100 125.700 465.900 127.050 ;
        RECT 458.100 120.600 459.900 125.700 ;
        RECT 461.100 120.000 462.900 124.800 ;
        RECT 464.100 120.600 465.900 125.700 ;
        RECT 476.100 120.000 477.900 129.600 ;
        RECT 482.700 129.000 486.000 130.200 ;
        RECT 482.700 120.600 484.500 129.000 ;
        RECT 506.700 126.600 507.600 133.950 ;
        RECT 524.100 132.150 525.900 133.950 ;
        RECT 527.700 129.600 528.900 133.950 ;
        RECT 530.100 132.150 531.900 133.950 ;
        RECT 548.100 132.150 549.900 133.950 ;
        RECT 551.700 129.600 552.900 133.950 ;
        RECT 554.100 132.150 555.900 133.950 ;
        RECT 569.250 132.150 571.050 133.950 ;
        RECT 527.700 128.700 531.300 129.600 ;
        RECT 551.700 128.700 555.300 129.600 ;
        RECT 498.000 120.000 499.800 126.600 ;
        RECT 502.500 125.400 507.600 126.600 ;
        RECT 521.100 125.700 528.900 127.050 ;
        RECT 502.500 120.600 504.300 125.400 ;
        RECT 505.500 120.000 507.300 123.600 ;
        RECT 521.100 120.600 522.900 125.700 ;
        RECT 524.100 120.000 525.900 124.800 ;
        RECT 527.100 120.600 528.900 125.700 ;
        RECT 530.100 126.600 531.300 128.700 ;
        RECT 530.100 120.600 531.900 126.600 ;
        RECT 545.100 125.700 552.900 127.050 ;
        RECT 545.100 120.600 546.900 125.700 ;
        RECT 548.100 120.000 549.900 124.800 ;
        RECT 551.100 120.600 552.900 125.700 ;
        RECT 554.100 126.600 555.300 128.700 ;
        RECT 575.100 126.600 576.300 133.950 ;
        RECT 581.100 132.150 582.900 133.950 ;
        RECT 583.950 132.450 586.050 133.050 ;
        RECT 590.550 132.450 591.450 137.550 ;
        RECT 599.100 136.050 600.900 137.850 ;
        RECT 605.100 136.050 606.000 148.200 ;
        RECT 623.100 136.050 624.900 137.850 ;
        RECT 629.100 136.050 630.000 148.200 ;
        RECT 644.100 144.300 645.900 155.400 ;
        RECT 647.100 145.200 648.900 156.000 ;
        RECT 650.100 144.300 651.900 155.400 ;
        RECT 644.100 143.400 651.900 144.300 ;
        RECT 653.100 143.400 654.900 155.400 ;
        RECT 668.100 144.300 669.900 155.400 ;
        RECT 671.100 145.200 672.900 156.000 ;
        RECT 674.100 144.300 675.900 155.400 ;
        RECT 668.100 143.400 675.900 144.300 ;
        RECT 677.100 143.400 678.900 155.400 ;
        RECT 689.700 149.400 691.500 156.000 ;
        RECT 690.000 146.100 691.800 147.900 ;
        RECT 692.700 144.900 694.500 155.400 ;
        RECT 692.100 143.400 694.500 144.900 ;
        RECT 697.800 143.400 699.600 156.000 ;
        RECT 713.400 143.400 715.200 156.000 ;
        RECT 718.500 144.900 720.300 155.400 ;
        RECT 721.500 149.400 723.300 156.000 ;
        RECT 734.100 149.400 735.900 156.000 ;
        RECT 737.100 149.400 738.900 155.400 ;
        RECT 749.100 149.400 750.900 155.400 ;
        RECT 752.100 150.000 753.900 156.000 ;
        RECT 721.200 146.100 723.000 147.900 ;
        RECT 718.500 143.400 720.900 144.900 ;
        RECT 647.250 136.050 649.050 137.850 ;
        RECT 653.700 136.050 654.600 143.400 ;
        RECT 671.250 136.050 673.050 137.850 ;
        RECT 677.700 136.050 678.600 143.400 ;
        RECT 692.100 136.050 693.300 143.400 ;
        RECT 698.100 136.050 699.900 137.850 ;
        RECT 713.100 136.050 714.900 137.850 ;
        RECT 719.700 136.050 720.900 143.400 ;
        RECT 734.100 136.050 735.900 137.850 ;
        RECT 737.100 136.050 738.300 149.400 ;
        RECT 750.000 149.100 750.900 149.400 ;
        RECT 755.100 149.400 756.900 155.400 ;
        RECT 758.100 149.400 759.900 156.000 ;
        RECT 770.100 149.400 771.900 155.400 ;
        RECT 773.100 149.400 774.900 156.000 ;
        RECT 788.100 149.400 789.900 156.000 ;
        RECT 791.100 149.400 792.900 155.400 ;
        RECT 794.100 150.000 795.900 156.000 ;
        RECT 755.100 149.100 756.600 149.400 ;
        RECT 750.000 148.200 756.600 149.100 ;
        RECT 750.000 136.050 750.900 148.200 ;
        RECT 755.100 136.050 756.900 137.850 ;
        RECT 770.700 136.050 771.900 149.400 ;
        RECT 791.400 149.100 792.900 149.400 ;
        RECT 797.100 149.400 798.900 155.400 ;
        RECT 809.100 149.400 810.900 156.000 ;
        RECT 812.100 149.400 813.900 155.400 ;
        RECT 815.100 150.000 816.900 156.000 ;
        RECT 797.100 149.100 798.000 149.400 ;
        RECT 791.400 148.200 798.000 149.100 ;
        RECT 812.400 149.100 813.900 149.400 ;
        RECT 818.100 149.400 819.900 155.400 ;
        RECT 820.950 153.450 823.050 154.050 ;
        RECT 826.950 153.450 829.050 154.050 ;
        RECT 820.950 152.550 829.050 153.450 ;
        RECT 820.950 151.950 823.050 152.550 ;
        RECT 826.950 151.950 829.050 152.550 ;
        RECT 818.100 149.100 819.000 149.400 ;
        RECT 812.400 148.200 819.000 149.100 ;
        RECT 772.950 147.450 775.050 148.050 ;
        RECT 784.950 147.450 787.050 148.050 ;
        RECT 772.950 146.550 787.050 147.450 ;
        RECT 772.950 145.950 775.050 146.550 ;
        RECT 784.950 145.950 787.050 146.550 ;
        RECT 773.100 136.050 774.900 137.850 ;
        RECT 791.100 136.050 792.900 137.850 ;
        RECT 797.100 136.050 798.000 148.200 ;
        RECT 812.100 136.050 813.900 137.850 ;
        RECT 818.100 136.050 819.000 148.200 ;
        RECT 833.100 144.300 834.900 155.400 ;
        RECT 836.100 145.200 837.900 156.000 ;
        RECT 839.100 144.300 840.900 155.400 ;
        RECT 833.100 143.400 840.900 144.300 ;
        RECT 842.100 143.400 843.900 155.400 ;
        RECT 857.400 143.400 859.200 156.000 ;
        RECT 862.500 144.900 864.300 155.400 ;
        RECT 865.500 149.400 867.300 156.000 ;
        RECT 865.200 146.100 867.000 147.900 ;
        RECT 862.500 143.400 864.900 144.900 ;
        RECT 881.400 143.400 883.200 156.000 ;
        RECT 886.500 144.900 888.300 155.400 ;
        RECT 889.500 149.400 891.300 156.000 ;
        RECT 889.200 146.100 891.000 147.900 ;
        RECT 886.500 143.400 888.900 144.900 ;
        RECT 905.100 144.600 906.900 155.400 ;
        RECT 908.100 145.500 909.900 156.000 ;
        RECT 911.100 154.500 918.900 155.400 ;
        RECT 911.100 144.600 912.900 154.500 ;
        RECT 905.100 143.700 912.900 144.600 ;
        RECT 836.250 136.050 838.050 137.850 ;
        RECT 842.700 136.050 843.600 143.400 ;
        RECT 859.950 141.450 862.050 142.050 ;
        RECT 854.550 140.550 862.050 141.450 ;
        RECT 854.550 138.450 855.450 140.550 ;
        RECT 859.950 139.950 862.050 140.550 ;
        RECT 851.550 137.550 855.450 138.450 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 583.950 131.550 591.450 132.450 ;
        RECT 596.100 132.150 597.900 133.950 ;
        RECT 602.100 132.150 603.900 133.950 ;
        RECT 583.950 130.950 586.050 131.550 ;
        RECT 605.100 130.200 606.000 133.950 ;
        RECT 620.100 132.150 621.900 133.950 ;
        RECT 626.100 132.150 627.900 133.950 ;
        RECT 629.100 130.200 630.000 133.950 ;
        RECT 644.100 132.150 645.900 133.950 ;
        RECT 650.250 132.150 652.050 133.950 ;
        RECT 554.100 120.600 555.900 126.600 ;
        RECT 569.700 120.000 571.500 126.600 ;
        RECT 574.200 120.600 576.000 126.600 ;
        RECT 578.700 120.000 580.500 126.600 ;
        RECT 596.100 120.000 597.900 129.600 ;
        RECT 602.700 129.000 606.000 130.200 ;
        RECT 602.700 120.600 604.500 129.000 ;
        RECT 620.100 120.000 621.900 129.600 ;
        RECT 626.700 129.000 630.000 130.200 ;
        RECT 626.700 120.600 628.500 129.000 ;
        RECT 653.700 126.600 654.600 133.950 ;
        RECT 668.100 132.150 669.900 133.950 ;
        RECT 674.250 132.150 676.050 133.950 ;
        RECT 655.950 129.450 658.050 130.050 ;
        RECT 667.950 129.450 670.050 130.050 ;
        RECT 655.950 128.550 670.050 129.450 ;
        RECT 655.950 127.950 658.050 128.550 ;
        RECT 667.950 127.950 670.050 128.550 ;
        RECT 677.700 126.600 678.600 133.950 ;
        RECT 689.100 132.150 690.900 133.950 ;
        RECT 692.100 129.600 693.300 133.950 ;
        RECT 695.100 132.150 696.900 133.950 ;
        RECT 716.100 132.150 717.900 133.950 ;
        RECT 689.700 128.700 693.300 129.600 ;
        RECT 719.700 129.600 720.900 133.950 ;
        RECT 722.100 132.150 723.900 133.950 ;
        RECT 719.700 128.700 723.300 129.600 ;
        RECT 689.700 126.600 690.900 128.700 ;
        RECT 645.000 120.000 646.800 126.600 ;
        RECT 649.500 125.400 654.600 126.600 ;
        RECT 649.500 120.600 651.300 125.400 ;
        RECT 652.500 120.000 654.300 123.600 ;
        RECT 669.000 120.000 670.800 126.600 ;
        RECT 673.500 125.400 678.600 126.600 ;
        RECT 673.500 120.600 675.300 125.400 ;
        RECT 676.500 120.000 678.300 123.600 ;
        RECT 689.100 120.600 690.900 126.600 ;
        RECT 692.100 125.700 699.900 127.050 ;
        RECT 692.100 120.600 693.900 125.700 ;
        RECT 695.100 120.000 696.900 124.800 ;
        RECT 698.100 120.600 699.900 125.700 ;
        RECT 713.100 125.700 720.900 127.050 ;
        RECT 713.100 120.600 714.900 125.700 ;
        RECT 716.100 120.000 717.900 124.800 ;
        RECT 719.100 120.600 720.900 125.700 ;
        RECT 722.100 126.600 723.300 128.700 ;
        RECT 722.100 120.600 723.900 126.600 ;
        RECT 737.100 123.600 738.300 133.950 ;
        RECT 750.000 130.200 750.900 133.950 ;
        RECT 752.100 132.150 753.900 133.950 ;
        RECT 758.100 132.150 759.900 133.950 ;
        RECT 750.000 129.000 753.300 130.200 ;
        RECT 734.100 120.000 735.900 123.600 ;
        RECT 737.100 120.600 738.900 123.600 ;
        RECT 751.500 120.600 753.300 129.000 ;
        RECT 758.100 120.000 759.900 129.600 ;
        RECT 770.700 123.600 771.900 133.950 ;
        RECT 788.100 132.150 789.900 133.950 ;
        RECT 794.100 132.150 795.900 133.950 ;
        RECT 797.100 130.200 798.000 133.950 ;
        RECT 809.100 132.150 810.900 133.950 ;
        RECT 815.100 132.150 816.900 133.950 ;
        RECT 818.100 130.200 819.000 133.950 ;
        RECT 833.100 132.150 834.900 133.950 ;
        RECT 839.250 132.150 841.050 133.950 ;
        RECT 770.100 120.600 771.900 123.600 ;
        RECT 773.100 120.000 774.900 123.600 ;
        RECT 788.100 120.000 789.900 129.600 ;
        RECT 794.700 129.000 798.000 130.200 ;
        RECT 794.700 120.600 796.500 129.000 ;
        RECT 809.100 120.000 810.900 129.600 ;
        RECT 815.700 129.000 819.000 130.200 ;
        RECT 815.700 120.600 817.500 129.000 ;
        RECT 842.700 126.600 843.600 133.950 ;
        RECT 844.950 132.450 847.050 133.050 ;
        RECT 851.550 132.450 852.450 137.550 ;
        RECT 857.100 136.050 858.900 137.850 ;
        RECT 863.700 136.050 864.900 143.400 ;
        RECT 881.100 136.050 882.900 137.850 ;
        RECT 887.700 136.050 888.900 143.400 ;
        RECT 914.100 142.500 915.900 153.600 ;
        RECT 917.100 143.400 918.900 154.500 ;
        RECT 932.100 149.400 933.900 156.000 ;
        RECT 935.100 149.400 936.900 155.400 ;
        RECT 938.100 150.000 939.900 156.000 ;
        RECT 935.400 149.100 936.900 149.400 ;
        RECT 941.100 149.400 942.900 155.400 ;
        RECT 941.100 149.100 942.000 149.400 ;
        RECT 935.400 148.200 942.000 149.100 ;
        RECT 911.100 141.600 915.900 142.500 ;
        RECT 892.950 138.450 897.000 139.050 ;
        RECT 892.950 136.950 897.450 138.450 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 844.950 131.550 852.450 132.450 ;
        RECT 860.100 132.150 861.900 133.950 ;
        RECT 844.950 130.950 847.050 131.550 ;
        RECT 863.700 129.600 864.900 133.950 ;
        RECT 866.100 132.150 867.900 133.950 ;
        RECT 884.100 132.150 885.900 133.950 ;
        RECT 887.700 129.600 888.900 133.950 ;
        RECT 890.100 132.150 891.900 133.950 ;
        RECT 896.550 132.450 897.450 136.950 ;
        RECT 908.250 136.050 910.050 137.850 ;
        RECT 911.100 136.050 912.000 141.600 ;
        RECT 916.950 141.450 919.050 142.050 ;
        RECT 925.950 141.450 928.050 142.050 ;
        RECT 934.950 141.450 937.050 142.050 ;
        RECT 916.950 140.550 937.050 141.450 ;
        RECT 916.950 139.950 919.050 140.550 ;
        RECT 925.950 139.950 928.050 140.550 ;
        RECT 934.950 139.950 937.050 140.550 ;
        RECT 927.000 138.450 931.050 139.050 ;
        RECT 914.100 136.050 915.900 137.850 ;
        RECT 926.550 136.950 931.050 138.450 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 913.950 133.950 916.050 136.050 ;
        RECT 916.950 133.950 919.050 136.050 ;
        RECT 893.550 131.550 897.450 132.450 ;
        RECT 905.250 132.150 907.050 133.950 ;
        RECT 863.700 128.700 867.300 129.600 ;
        RECT 887.700 128.700 891.300 129.600 ;
        RECT 834.000 120.000 835.800 126.600 ;
        RECT 838.500 125.400 843.600 126.600 ;
        RECT 857.100 125.700 864.900 127.050 ;
        RECT 838.500 120.600 840.300 125.400 ;
        RECT 841.500 120.000 843.300 123.600 ;
        RECT 857.100 120.600 858.900 125.700 ;
        RECT 860.100 120.000 861.900 124.800 ;
        RECT 863.100 120.600 864.900 125.700 ;
        RECT 866.100 126.600 867.300 128.700 ;
        RECT 866.100 120.600 867.900 126.600 ;
        RECT 881.100 125.700 888.900 127.050 ;
        RECT 881.100 120.600 882.900 125.700 ;
        RECT 884.100 120.000 885.900 124.800 ;
        RECT 887.100 120.600 888.900 125.700 ;
        RECT 890.100 126.600 891.300 128.700 ;
        RECT 893.550 127.050 894.450 131.550 ;
        RECT 895.950 129.450 898.050 130.050 ;
        RECT 904.950 129.450 907.050 130.050 ;
        RECT 895.950 128.550 907.050 129.450 ;
        RECT 895.950 127.950 898.050 128.550 ;
        RECT 904.950 127.950 907.050 128.550 ;
        RECT 893.550 126.900 897.000 127.050 ;
        RECT 890.100 120.600 891.900 126.600 ;
        RECT 893.550 125.550 898.050 126.900 ;
        RECT 911.100 126.600 912.300 133.950 ;
        RECT 917.100 132.150 918.900 133.950 ;
        RECT 926.550 133.050 927.450 136.950 ;
        RECT 935.100 136.050 936.900 137.850 ;
        RECT 941.100 136.050 942.000 148.200 ;
        RECT 931.950 133.950 934.050 136.050 ;
        RECT 934.950 133.950 937.050 136.050 ;
        RECT 937.950 133.950 940.050 136.050 ;
        RECT 940.950 133.950 943.050 136.050 ;
        RECT 926.550 131.550 931.050 133.050 ;
        RECT 932.100 132.150 933.900 133.950 ;
        RECT 938.100 132.150 939.900 133.950 ;
        RECT 927.000 130.950 931.050 131.550 ;
        RECT 941.100 130.200 942.000 133.950 ;
        RECT 894.000 124.950 898.050 125.550 ;
        RECT 895.950 124.800 898.050 124.950 ;
        RECT 905.700 120.000 907.500 126.600 ;
        RECT 910.200 120.600 912.000 126.600 ;
        RECT 914.700 120.000 916.500 126.600 ;
        RECT 932.100 120.000 933.900 129.600 ;
        RECT 938.700 129.000 942.000 130.200 ;
        RECT 938.700 120.600 940.500 129.000 ;
        RECT 11.100 110.400 12.900 116.400 ;
        RECT 11.700 108.300 12.900 110.400 ;
        RECT 14.100 111.300 15.900 116.400 ;
        RECT 17.100 112.200 18.900 117.000 ;
        RECT 20.100 111.300 21.900 116.400 ;
        RECT 14.100 109.950 21.900 111.300 ;
        RECT 33.000 110.400 34.800 117.000 ;
        RECT 37.500 111.600 39.300 116.400 ;
        RECT 40.500 113.400 42.300 117.000 ;
        RECT 37.500 110.400 42.600 111.600 ;
        RECT 56.100 110.400 57.900 116.400 ;
        RECT 11.700 107.400 15.300 108.300 ;
        RECT 11.100 103.050 12.900 104.850 ;
        RECT 14.100 103.050 15.300 107.400 ;
        RECT 17.100 103.050 18.900 104.850 ;
        RECT 32.100 103.050 33.900 104.850 ;
        RECT 38.250 103.050 40.050 104.850 ;
        RECT 41.700 103.050 42.600 110.400 ;
        RECT 56.700 108.300 57.900 110.400 ;
        RECT 59.100 111.300 60.900 116.400 ;
        RECT 62.100 112.200 63.900 117.000 ;
        RECT 65.100 111.300 66.900 116.400 ;
        RECT 78.600 112.200 80.400 116.400 ;
        RECT 59.100 109.950 66.900 111.300 ;
        RECT 77.700 110.400 80.400 112.200 ;
        RECT 81.600 110.400 83.400 117.000 ;
        RECT 56.700 107.400 60.300 108.300 ;
        RECT 56.100 103.050 57.900 104.850 ;
        RECT 59.100 103.050 60.300 107.400 ;
        RECT 62.100 103.050 63.900 104.850 ;
        RECT 77.700 103.050 78.600 110.400 ;
        RECT 79.500 108.600 81.300 109.500 ;
        RECT 86.100 108.600 87.900 116.400 ;
        RECT 101.100 113.400 102.900 117.000 ;
        RECT 104.100 113.400 105.900 116.400 ;
        RECT 107.100 113.400 108.900 117.000 ;
        RECT 79.500 107.700 87.900 108.600 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 77.100 100.950 79.200 103.050 ;
        RECT 80.400 100.950 82.500 103.050 ;
        RECT 14.100 93.600 15.300 100.950 ;
        RECT 20.100 99.150 21.900 100.950 ;
        RECT 35.250 99.150 37.050 100.950 ;
        RECT 25.950 96.450 28.050 97.050 ;
        RECT 37.950 96.450 40.050 97.050 ;
        RECT 25.950 95.550 40.050 96.450 ;
        RECT 25.950 94.950 28.050 95.550 ;
        RECT 37.950 94.950 40.050 95.550 ;
        RECT 41.700 93.600 42.600 100.950 ;
        RECT 59.100 93.600 60.300 100.950 ;
        RECT 65.100 99.150 66.900 100.950 ;
        RECT 77.700 93.600 78.600 100.950 ;
        RECT 81.000 99.150 82.800 100.950 ;
        RECT 14.100 92.100 16.500 93.600 ;
        RECT 12.000 89.100 13.800 90.900 ;
        RECT 11.700 81.000 13.500 87.600 ;
        RECT 14.700 81.600 16.500 92.100 ;
        RECT 19.800 81.000 21.600 93.600 ;
        RECT 32.100 92.700 39.900 93.600 ;
        RECT 32.100 81.600 33.900 92.700 ;
        RECT 35.100 81.000 36.900 91.800 ;
        RECT 38.100 81.600 39.900 92.700 ;
        RECT 41.100 81.600 42.900 93.600 ;
        RECT 59.100 92.100 61.500 93.600 ;
        RECT 57.000 89.100 58.800 90.900 ;
        RECT 56.700 81.000 58.500 87.600 ;
        RECT 59.700 81.600 61.500 92.100 ;
        RECT 64.800 81.000 66.600 93.600 ;
        RECT 77.100 81.600 78.900 93.600 ;
        RECT 80.100 81.000 81.900 93.000 ;
        RECT 84.000 87.600 84.900 107.700 ;
        RECT 85.950 103.050 87.750 104.850 ;
        RECT 104.400 103.050 105.300 113.400 ;
        RECT 124.500 110.400 126.300 117.000 ;
        RECT 129.000 110.400 130.800 116.400 ;
        RECT 133.500 110.400 135.300 117.000 ;
        RECT 112.950 105.450 115.050 106.050 ;
        RECT 118.950 105.450 121.050 106.050 ;
        RECT 112.950 104.550 121.050 105.450 ;
        RECT 112.950 103.950 115.050 104.550 ;
        RECT 118.950 103.950 121.050 104.550 ;
        RECT 122.100 103.050 123.900 104.850 ;
        RECT 128.700 103.050 129.900 110.400 ;
        RECT 146.100 107.400 147.900 117.000 ;
        RECT 152.700 108.000 154.500 116.400 ;
        RECT 152.700 106.800 156.000 108.000 ;
        RECT 170.100 107.400 171.900 117.000 ;
        RECT 176.700 108.000 178.500 116.400 ;
        RECT 195.000 110.400 196.800 117.000 ;
        RECT 199.500 111.600 201.300 116.400 ;
        RECT 202.500 113.400 204.300 117.000 ;
        RECT 218.100 113.400 219.900 117.000 ;
        RECT 221.100 113.400 222.900 116.400 ;
        RECT 224.100 113.400 225.900 117.000 ;
        RECT 226.950 114.450 229.050 115.050 ;
        RECT 235.950 114.450 238.050 115.050 ;
        RECT 226.950 113.550 238.050 114.450 ;
        RECT 199.500 110.400 204.600 111.600 ;
        RECT 176.700 106.800 180.000 108.000 ;
        RECT 141.000 105.450 145.050 106.050 ;
        RECT 133.950 103.050 135.750 104.850 ;
        RECT 140.550 103.950 145.050 105.450 ;
        RECT 85.800 100.950 87.900 103.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 121.950 100.950 124.050 103.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 101.250 99.150 103.050 100.950 ;
        RECT 104.400 93.600 105.300 100.950 ;
        RECT 107.100 99.150 108.900 100.950 ;
        RECT 125.100 99.150 126.900 100.950 ;
        RECT 129.000 95.400 129.900 100.950 ;
        RECT 130.950 99.150 132.750 100.950 ;
        RECT 140.550 100.050 141.450 103.950 ;
        RECT 146.100 103.050 147.900 104.850 ;
        RECT 152.100 103.050 153.900 104.850 ;
        RECT 155.100 103.050 156.000 106.800 ;
        RECT 170.100 103.050 171.900 104.850 ;
        RECT 176.100 103.050 177.900 104.850 ;
        RECT 179.100 103.050 180.000 106.800 ;
        RECT 194.100 103.050 195.900 104.850 ;
        RECT 200.250 103.050 202.050 104.850 ;
        RECT 203.700 103.050 204.600 110.400 ;
        RECT 221.700 103.050 222.600 113.400 ;
        RECT 226.950 112.950 229.050 113.550 ;
        RECT 235.950 112.950 238.050 113.550 ;
        RECT 239.100 111.300 240.900 116.400 ;
        RECT 242.100 112.200 243.900 117.000 ;
        RECT 245.100 111.300 246.900 116.400 ;
        RECT 239.100 109.950 246.900 111.300 ;
        RECT 248.100 110.400 249.900 116.400 ;
        RECT 263.100 111.300 264.900 116.400 ;
        RECT 266.100 112.200 267.900 117.000 ;
        RECT 269.100 111.300 270.900 116.400 ;
        RECT 248.100 108.300 249.300 110.400 ;
        RECT 263.100 109.950 270.900 111.300 ;
        RECT 272.100 110.400 273.900 116.400 ;
        RECT 272.100 108.300 273.300 110.400 ;
        RECT 245.700 107.400 249.300 108.300 ;
        RECT 269.700 107.400 273.300 108.300 ;
        RECT 287.100 107.400 288.900 117.000 ;
        RECT 293.700 108.000 295.500 116.400 ;
        RECT 313.500 110.400 315.300 117.000 ;
        RECT 318.000 110.400 319.800 116.400 ;
        RECT 322.500 110.400 324.300 117.000 ;
        RECT 335.100 113.400 336.900 116.400 ;
        RECT 338.100 113.400 339.900 117.000 ;
        RECT 242.100 103.050 243.900 104.850 ;
        RECT 245.700 103.050 246.900 107.400 ;
        RECT 248.100 103.050 249.900 104.850 ;
        RECT 266.100 103.050 267.900 104.850 ;
        RECT 269.700 103.050 270.900 107.400 ;
        RECT 293.700 106.800 297.000 108.000 ;
        RECT 274.950 105.450 277.050 106.050 ;
        RECT 280.950 105.450 283.050 106.050 ;
        RECT 272.100 103.050 273.900 104.850 ;
        RECT 274.950 104.550 283.050 105.450 ;
        RECT 274.950 103.950 277.050 104.550 ;
        RECT 280.950 103.950 283.050 104.550 ;
        RECT 287.100 103.050 288.900 104.850 ;
        RECT 293.100 103.050 294.900 104.850 ;
        RECT 296.100 103.050 297.000 106.800 ;
        RECT 298.950 105.450 303.000 106.050 ;
        RECT 298.950 103.950 303.450 105.450 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 154.950 100.950 157.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 175.950 100.950 178.050 103.050 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 220.950 100.950 223.050 103.050 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 136.950 98.550 141.450 100.050 ;
        RECT 149.100 99.150 150.900 100.950 ;
        RECT 136.950 97.950 141.000 98.550 ;
        RECT 125.100 94.500 129.900 95.400 ;
        RECT 130.950 96.450 133.050 97.050 ;
        RECT 139.950 96.450 142.050 97.050 ;
        RECT 130.950 95.550 142.050 96.450 ;
        RECT 130.950 94.950 133.050 95.550 ;
        RECT 139.950 94.950 142.050 95.550 ;
        RECT 83.100 81.600 84.900 87.600 ;
        RECT 86.100 81.000 87.900 87.600 ;
        RECT 101.100 81.000 102.900 93.600 ;
        RECT 104.400 92.400 108.000 93.600 ;
        RECT 106.200 81.600 108.000 92.400 ;
        RECT 122.100 82.500 123.900 93.600 ;
        RECT 125.100 83.400 126.900 94.500 ;
        RECT 128.100 92.400 135.900 93.300 ;
        RECT 128.100 82.500 129.900 92.400 ;
        RECT 122.100 81.600 129.900 82.500 ;
        RECT 131.100 81.000 132.900 91.500 ;
        RECT 134.100 81.600 135.900 92.400 ;
        RECT 155.100 88.800 156.000 100.950 ;
        RECT 173.100 99.150 174.900 100.950 ;
        RECT 179.100 88.800 180.000 100.950 ;
        RECT 197.250 99.150 199.050 100.950 ;
        RECT 190.950 96.450 193.050 97.050 ;
        RECT 199.950 96.450 202.050 97.050 ;
        RECT 190.950 95.550 202.050 96.450 ;
        RECT 190.950 94.950 193.050 95.550 ;
        RECT 199.950 94.950 202.050 95.550 ;
        RECT 203.700 93.600 204.600 100.950 ;
        RECT 218.100 99.150 219.900 100.950 ;
        RECT 221.700 93.600 222.600 100.950 ;
        RECT 223.950 99.150 225.750 100.950 ;
        RECT 239.100 99.150 240.900 100.950 ;
        RECT 245.700 93.600 246.900 100.950 ;
        RECT 263.100 99.150 264.900 100.950 ;
        RECT 253.950 96.450 256.050 97.050 ;
        RECT 265.950 96.450 268.050 96.750 ;
        RECT 253.950 95.550 268.050 96.450 ;
        RECT 253.950 94.950 256.050 95.550 ;
        RECT 265.950 94.650 268.050 95.550 ;
        RECT 269.700 93.600 270.900 100.950 ;
        RECT 290.100 99.150 291.900 100.950 ;
        RECT 271.950 96.450 274.050 96.750 ;
        RECT 292.950 96.450 295.050 97.050 ;
        RECT 271.950 95.550 295.050 96.450 ;
        RECT 271.950 94.650 274.050 95.550 ;
        RECT 292.950 94.950 295.050 95.550 ;
        RECT 149.400 87.900 156.000 88.800 ;
        RECT 149.400 87.600 150.900 87.900 ;
        RECT 146.100 81.000 147.900 87.600 ;
        RECT 149.100 81.600 150.900 87.600 ;
        RECT 155.100 87.600 156.000 87.900 ;
        RECT 173.400 87.900 180.000 88.800 ;
        RECT 173.400 87.600 174.900 87.900 ;
        RECT 152.100 81.000 153.900 87.000 ;
        RECT 155.100 81.600 156.900 87.600 ;
        RECT 170.100 81.000 171.900 87.600 ;
        RECT 173.100 81.600 174.900 87.600 ;
        RECT 179.100 87.600 180.000 87.900 ;
        RECT 194.100 92.700 201.900 93.600 ;
        RECT 176.100 81.000 177.900 87.000 ;
        RECT 179.100 81.600 180.900 87.600 ;
        RECT 194.100 81.600 195.900 92.700 ;
        RECT 197.100 81.000 198.900 91.800 ;
        RECT 200.100 81.600 201.900 92.700 ;
        RECT 203.100 81.600 204.900 93.600 ;
        RECT 219.000 92.400 222.600 93.600 ;
        RECT 219.000 81.600 220.800 92.400 ;
        RECT 224.100 81.000 225.900 93.600 ;
        RECT 239.400 81.000 241.200 93.600 ;
        RECT 244.500 92.100 246.900 93.600 ;
        RECT 244.500 81.600 246.300 92.100 ;
        RECT 247.200 89.100 249.000 90.900 ;
        RECT 247.500 81.000 249.300 87.600 ;
        RECT 263.400 81.000 265.200 93.600 ;
        RECT 268.500 92.100 270.900 93.600 ;
        RECT 268.500 81.600 270.300 92.100 ;
        RECT 271.200 89.100 273.000 90.900 ;
        RECT 296.100 88.800 297.000 100.950 ;
        RECT 302.550 99.450 303.450 103.950 ;
        RECT 311.100 103.050 312.900 104.850 ;
        RECT 317.700 103.050 318.900 110.400 ;
        RECT 322.950 103.050 324.750 104.850 ;
        RECT 335.700 103.050 336.900 113.400 ;
        RECT 350.100 111.300 351.900 116.400 ;
        RECT 353.100 112.200 354.900 117.000 ;
        RECT 356.100 111.300 357.900 116.400 ;
        RECT 350.100 109.950 357.900 111.300 ;
        RECT 359.100 110.400 360.900 116.400 ;
        RECT 359.100 108.300 360.300 110.400 ;
        RECT 371.700 109.200 373.500 116.400 ;
        RECT 376.800 110.400 378.600 117.000 ;
        RECT 392.700 113.400 394.500 117.000 ;
        RECT 395.700 111.600 397.500 116.400 ;
        RECT 392.400 110.400 397.500 111.600 ;
        RECT 400.200 110.400 402.000 117.000 ;
        RECT 371.700 108.300 375.900 109.200 ;
        RECT 356.700 107.400 360.300 108.300 ;
        RECT 353.100 103.050 354.900 104.850 ;
        RECT 356.700 103.050 357.900 107.400 ;
        RECT 359.100 103.050 360.900 104.850 ;
        RECT 371.100 103.050 372.900 104.850 ;
        RECT 374.700 103.050 375.900 108.300 ;
        RECT 376.950 103.050 378.750 104.850 ;
        RECT 392.400 103.050 393.300 110.400 ;
        RECT 416.100 107.400 417.900 117.000 ;
        RECT 422.700 108.000 424.500 116.400 ;
        RECT 439.500 108.000 441.300 116.400 ;
        RECT 422.700 106.800 426.000 108.000 ;
        RECT 403.950 105.450 408.000 106.050 ;
        RECT 394.950 103.050 396.750 104.850 ;
        RECT 401.100 103.050 402.900 104.850 ;
        RECT 403.950 103.950 408.450 105.450 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 313.950 100.950 316.050 103.050 ;
        RECT 316.950 100.950 319.050 103.050 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 352.950 100.950 355.050 103.050 ;
        RECT 355.950 100.950 358.050 103.050 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 373.950 100.950 376.050 103.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 394.950 100.950 397.050 103.050 ;
        RECT 397.950 100.950 400.050 103.050 ;
        RECT 400.950 100.950 403.050 103.050 ;
        RECT 299.550 99.000 303.450 99.450 ;
        RECT 314.100 99.150 315.900 100.950 ;
        RECT 298.950 98.550 303.450 99.000 ;
        RECT 298.950 94.950 301.050 98.550 ;
        RECT 318.000 95.400 318.900 100.950 ;
        RECT 319.950 99.150 321.750 100.950 ;
        RECT 314.100 94.500 318.900 95.400 ;
        RECT 290.400 87.900 297.000 88.800 ;
        RECT 290.400 87.600 291.900 87.900 ;
        RECT 271.500 81.000 273.300 87.600 ;
        RECT 287.100 81.000 288.900 87.600 ;
        RECT 290.100 81.600 291.900 87.600 ;
        RECT 296.100 87.600 297.000 87.900 ;
        RECT 293.100 81.000 294.900 87.000 ;
        RECT 296.100 81.600 297.900 87.600 ;
        RECT 311.100 82.500 312.900 93.600 ;
        RECT 314.100 83.400 315.900 94.500 ;
        RECT 317.100 92.400 324.900 93.300 ;
        RECT 317.100 82.500 318.900 92.400 ;
        RECT 311.100 81.600 318.900 82.500 ;
        RECT 320.100 81.000 321.900 91.500 ;
        RECT 323.100 81.600 324.900 92.400 ;
        RECT 335.700 87.600 336.900 100.950 ;
        RECT 338.100 99.150 339.900 100.950 ;
        RECT 350.100 99.150 351.900 100.950 ;
        RECT 356.700 93.600 357.900 100.950 ;
        RECT 335.100 81.600 336.900 87.600 ;
        RECT 338.100 81.000 339.900 87.600 ;
        RECT 350.400 81.000 352.200 93.600 ;
        RECT 355.500 92.100 357.900 93.600 ;
        RECT 355.500 81.600 357.300 92.100 ;
        RECT 358.200 89.100 360.000 90.900 ;
        RECT 374.700 87.600 375.900 100.950 ;
        RECT 392.400 93.600 393.300 100.950 ;
        RECT 397.950 99.150 399.750 100.950 ;
        RECT 407.550 99.900 408.450 103.950 ;
        RECT 416.100 103.050 417.900 104.850 ;
        RECT 422.100 103.050 423.900 104.850 ;
        RECT 425.100 103.050 426.000 106.800 ;
        RECT 438.000 106.800 441.300 108.000 ;
        RECT 446.100 107.400 447.900 117.000 ;
        RECT 461.700 113.400 463.500 117.000 ;
        RECT 464.700 111.600 466.500 116.400 ;
        RECT 461.400 110.400 466.500 111.600 ;
        RECT 469.200 110.400 471.000 117.000 ;
        RECT 485.700 113.400 487.500 117.000 ;
        RECT 488.700 111.600 490.500 116.400 ;
        RECT 485.400 110.400 490.500 111.600 ;
        RECT 493.200 110.400 495.000 117.000 ;
        RECT 438.000 103.050 438.900 106.800 ;
        RECT 440.100 103.050 441.900 104.850 ;
        RECT 446.100 103.050 447.900 104.850 ;
        RECT 461.400 103.050 462.300 110.400 ;
        RECT 463.950 103.050 465.750 104.850 ;
        RECT 470.100 103.050 471.900 104.850 ;
        RECT 485.400 103.050 486.300 110.400 ;
        RECT 508.500 108.000 510.300 116.400 ;
        RECT 507.000 106.800 510.300 108.000 ;
        RECT 515.100 107.400 516.900 117.000 ;
        RECT 529.500 108.000 531.300 116.400 ;
        RECT 528.000 106.800 531.300 108.000 ;
        RECT 536.100 107.400 537.900 117.000 ;
        RECT 551.700 113.400 553.500 117.000 ;
        RECT 554.700 111.600 556.500 116.400 ;
        RECT 551.400 110.400 556.500 111.600 ;
        RECT 559.200 110.400 561.000 117.000 ;
        RECT 487.950 103.050 489.750 104.850 ;
        RECT 494.100 103.050 495.900 104.850 ;
        RECT 507.000 103.050 507.900 106.800 ;
        RECT 509.100 103.050 510.900 104.850 ;
        RECT 515.100 103.050 516.900 104.850 ;
        RECT 528.000 103.050 528.900 106.800 ;
        RECT 530.100 103.050 531.900 104.850 ;
        RECT 536.100 103.050 537.900 104.850 ;
        RECT 551.400 103.050 552.300 110.400 ;
        RECT 575.100 107.400 576.900 117.000 ;
        RECT 581.700 108.000 583.500 116.400 ;
        RECT 596.100 108.600 597.900 116.400 ;
        RECT 600.600 110.400 602.400 117.000 ;
        RECT 603.600 112.200 605.400 116.400 ;
        RECT 603.600 110.400 606.300 112.200 ;
        RECT 617.400 110.400 619.200 117.000 ;
        RECT 602.700 108.600 604.500 109.500 ;
        RECT 581.700 106.800 585.000 108.000 ;
        RECT 596.100 107.700 604.500 108.600 ;
        RECT 553.950 103.050 555.750 104.850 ;
        RECT 560.100 103.050 561.900 104.850 ;
        RECT 575.100 103.050 576.900 104.850 ;
        RECT 581.100 103.050 582.900 104.850 ;
        RECT 584.100 103.050 585.000 106.800 ;
        RECT 596.250 103.050 598.050 104.850 ;
        RECT 415.950 100.950 418.050 103.050 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 596.100 100.950 598.200 103.050 ;
        RECT 406.950 97.800 409.050 99.900 ;
        RECT 419.100 99.150 420.900 100.950 ;
        RECT 394.950 96.450 397.050 97.050 ;
        RECT 412.950 96.450 415.050 97.050 ;
        RECT 394.950 95.550 415.050 96.450 ;
        RECT 394.950 94.950 397.050 95.550 ;
        RECT 412.950 94.950 415.050 95.550 ;
        RECT 358.500 81.000 360.300 87.600 ;
        RECT 371.100 81.000 372.900 87.600 ;
        RECT 374.100 81.600 375.900 87.600 ;
        RECT 377.100 81.000 378.900 87.600 ;
        RECT 392.100 81.600 393.900 93.600 ;
        RECT 395.100 92.700 402.900 93.600 ;
        RECT 395.100 81.600 396.900 92.700 ;
        RECT 398.100 81.000 399.900 91.800 ;
        RECT 401.100 81.600 402.900 92.700 ;
        RECT 425.100 88.800 426.000 100.950 ;
        RECT 419.400 87.900 426.000 88.800 ;
        RECT 419.400 87.600 420.900 87.900 ;
        RECT 416.100 81.000 417.900 87.600 ;
        RECT 419.100 81.600 420.900 87.600 ;
        RECT 425.100 87.600 426.000 87.900 ;
        RECT 438.000 88.800 438.900 100.950 ;
        RECT 443.100 99.150 444.900 100.950 ;
        RECT 461.400 93.600 462.300 100.950 ;
        RECT 466.950 99.150 468.750 100.950 ;
        RECT 485.400 93.600 486.300 100.950 ;
        RECT 490.950 99.150 492.750 100.950 ;
        RECT 438.000 87.900 444.600 88.800 ;
        RECT 438.000 87.600 438.900 87.900 ;
        RECT 422.100 81.000 423.900 87.000 ;
        RECT 425.100 81.600 426.900 87.600 ;
        RECT 437.100 81.600 438.900 87.600 ;
        RECT 443.100 87.600 444.600 87.900 ;
        RECT 440.100 81.000 441.900 87.000 ;
        RECT 443.100 81.600 444.900 87.600 ;
        RECT 446.100 81.000 447.900 87.600 ;
        RECT 461.100 81.600 462.900 93.600 ;
        RECT 464.100 92.700 471.900 93.600 ;
        RECT 464.100 81.600 465.900 92.700 ;
        RECT 467.100 81.000 468.900 91.800 ;
        RECT 470.100 81.600 471.900 92.700 ;
        RECT 485.100 81.600 486.900 93.600 ;
        RECT 488.100 92.700 495.900 93.600 ;
        RECT 488.100 81.600 489.900 92.700 ;
        RECT 491.100 81.000 492.900 91.800 ;
        RECT 494.100 81.600 495.900 92.700 ;
        RECT 507.000 88.800 507.900 100.950 ;
        RECT 512.100 99.150 513.900 100.950 ;
        RECT 528.000 88.800 528.900 100.950 ;
        RECT 533.100 99.150 534.900 100.950 ;
        RECT 551.400 93.600 552.300 100.950 ;
        RECT 556.950 99.150 558.750 100.950 ;
        RECT 578.100 99.150 579.900 100.950 ;
        RECT 565.950 96.450 568.050 97.050 ;
        RECT 580.950 96.450 583.050 97.050 ;
        RECT 565.950 95.550 583.050 96.450 ;
        RECT 565.950 94.950 568.050 95.550 ;
        RECT 580.950 94.950 583.050 95.550 ;
        RECT 507.000 87.900 513.600 88.800 ;
        RECT 507.000 87.600 507.900 87.900 ;
        RECT 506.100 81.600 507.900 87.600 ;
        RECT 512.100 87.600 513.600 87.900 ;
        RECT 528.000 87.900 534.600 88.800 ;
        RECT 528.000 87.600 528.900 87.900 ;
        RECT 509.100 81.000 510.900 87.000 ;
        RECT 512.100 81.600 513.900 87.600 ;
        RECT 515.100 81.000 516.900 87.600 ;
        RECT 527.100 81.600 528.900 87.600 ;
        RECT 533.100 87.600 534.600 87.900 ;
        RECT 530.100 81.000 531.900 87.000 ;
        RECT 533.100 81.600 534.900 87.600 ;
        RECT 536.100 81.000 537.900 87.600 ;
        RECT 551.100 81.600 552.900 93.600 ;
        RECT 554.100 92.700 561.900 93.600 ;
        RECT 554.100 81.600 555.900 92.700 ;
        RECT 557.100 81.000 558.900 91.800 ;
        RECT 560.100 81.600 561.900 92.700 ;
        RECT 584.100 88.800 585.000 100.950 ;
        RECT 578.400 87.900 585.000 88.800 ;
        RECT 578.400 87.600 579.900 87.900 ;
        RECT 575.100 81.000 576.900 87.600 ;
        RECT 578.100 81.600 579.900 87.600 ;
        RECT 584.100 87.600 585.000 87.900 ;
        RECT 599.100 87.600 600.000 107.700 ;
        RECT 605.400 103.050 606.300 110.400 ;
        RECT 622.500 109.200 624.300 116.400 ;
        RECT 635.100 110.400 636.900 116.400 ;
        RECT 620.100 108.300 624.300 109.200 ;
        RECT 635.700 108.300 636.900 110.400 ;
        RECT 638.100 111.300 639.900 116.400 ;
        RECT 641.100 112.200 642.900 117.000 ;
        RECT 644.100 111.300 645.900 116.400 ;
        RECT 638.100 109.950 645.900 111.300 ;
        RECT 659.100 110.400 660.900 116.400 ;
        RECT 659.700 108.300 660.900 110.400 ;
        RECT 662.100 111.300 663.900 116.400 ;
        RECT 665.100 112.200 666.900 117.000 ;
        RECT 668.100 111.300 669.900 116.400 ;
        RECT 662.100 109.950 669.900 111.300 ;
        RECT 617.250 103.050 619.050 104.850 ;
        RECT 620.100 103.050 621.300 108.300 ;
        RECT 635.700 107.400 639.300 108.300 ;
        RECT 659.700 107.400 663.300 108.300 ;
        RECT 685.500 108.000 687.300 116.400 ;
        RECT 623.100 103.050 624.900 104.850 ;
        RECT 635.100 103.050 636.900 104.850 ;
        RECT 638.100 103.050 639.300 107.400 ;
        RECT 641.100 103.050 642.900 104.850 ;
        RECT 659.100 103.050 660.900 104.850 ;
        RECT 662.100 103.050 663.300 107.400 ;
        RECT 684.000 106.800 687.300 108.000 ;
        RECT 692.100 107.400 693.900 117.000 ;
        RECT 707.100 111.300 708.900 116.400 ;
        RECT 710.100 112.200 711.900 117.000 ;
        RECT 713.100 111.300 714.900 116.400 ;
        RECT 707.100 109.950 714.900 111.300 ;
        RECT 716.100 110.400 717.900 116.400 ;
        RECT 716.100 108.300 717.300 110.400 ;
        RECT 713.700 107.400 717.300 108.300 ;
        RECT 733.500 108.000 735.300 116.400 ;
        RECT 665.100 103.050 666.900 104.850 ;
        RECT 684.000 103.050 684.900 106.800 ;
        RECT 694.950 105.450 699.000 106.050 ;
        RECT 686.100 103.050 687.900 104.850 ;
        RECT 692.100 103.050 693.900 104.850 ;
        RECT 694.950 103.950 699.450 105.450 ;
        RECT 601.500 100.950 603.600 103.050 ;
        RECT 604.800 100.950 606.900 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 601.200 99.150 603.000 100.950 ;
        RECT 605.400 93.600 606.300 100.950 ;
        RECT 581.100 81.000 582.900 87.000 ;
        RECT 584.100 81.600 585.900 87.600 ;
        RECT 596.100 81.000 597.900 87.600 ;
        RECT 599.100 81.600 600.900 87.600 ;
        RECT 602.100 81.000 603.900 93.000 ;
        RECT 605.100 81.600 606.900 93.600 ;
        RECT 620.100 87.600 621.300 100.950 ;
        RECT 638.100 93.600 639.300 100.950 ;
        RECT 644.100 99.150 645.900 100.950 ;
        RECT 640.950 96.450 643.050 96.750 ;
        RECT 652.950 96.450 655.050 97.050 ;
        RECT 640.950 95.550 655.050 96.450 ;
        RECT 640.950 94.650 643.050 95.550 ;
        RECT 652.950 94.950 655.050 95.550 ;
        RECT 662.100 93.600 663.300 100.950 ;
        RECT 668.100 99.150 669.900 100.950 ;
        RECT 638.100 92.100 640.500 93.600 ;
        RECT 636.000 89.100 637.800 90.900 ;
        RECT 617.100 81.000 618.900 87.600 ;
        RECT 620.100 81.600 621.900 87.600 ;
        RECT 623.100 81.000 624.900 87.600 ;
        RECT 635.700 81.000 637.500 87.600 ;
        RECT 638.700 81.600 640.500 92.100 ;
        RECT 643.800 81.000 645.600 93.600 ;
        RECT 662.100 92.100 664.500 93.600 ;
        RECT 660.000 89.100 661.800 90.900 ;
        RECT 659.700 81.000 661.500 87.600 ;
        RECT 662.700 81.600 664.500 92.100 ;
        RECT 667.800 81.000 669.600 93.600 ;
        RECT 684.000 88.800 684.900 100.950 ;
        RECT 689.100 99.150 690.900 100.950 ;
        RECT 698.550 100.050 699.450 103.950 ;
        RECT 710.100 103.050 711.900 104.850 ;
        RECT 713.700 103.050 714.900 107.400 ;
        RECT 732.000 106.800 735.300 108.000 ;
        RECT 740.100 107.400 741.900 117.000 ;
        RECT 752.700 109.200 754.500 116.400 ;
        RECT 757.800 110.400 759.600 117.000 ;
        RECT 773.700 109.200 775.500 116.400 ;
        RECT 778.800 110.400 780.600 117.000 ;
        RECT 794.100 111.300 795.900 116.400 ;
        RECT 797.100 112.200 798.900 117.000 ;
        RECT 800.100 111.300 801.900 116.400 ;
        RECT 794.100 109.950 801.900 111.300 ;
        RECT 803.100 110.400 804.900 116.400 ;
        RECT 818.400 110.400 820.200 117.000 ;
        RECT 752.700 108.300 756.900 109.200 ;
        RECT 773.700 108.300 777.900 109.200 ;
        RECT 803.100 108.300 804.300 110.400 ;
        RECT 823.500 109.200 825.300 116.400 ;
        RECT 836.700 110.400 838.500 117.000 ;
        RECT 841.200 110.400 843.000 116.400 ;
        RECT 845.700 110.400 847.500 117.000 ;
        RECT 716.100 103.050 717.900 104.850 ;
        RECT 732.000 103.050 732.900 106.800 ;
        RECT 734.100 103.050 735.900 104.850 ;
        RECT 740.100 103.050 741.900 104.850 ;
        RECT 752.100 103.050 753.900 104.850 ;
        RECT 755.700 103.050 756.900 108.300 ;
        RECT 760.950 105.450 763.050 106.050 ;
        RECT 757.950 103.050 759.750 104.850 ;
        RECT 760.950 104.550 768.450 105.450 ;
        RECT 760.950 103.950 763.050 104.550 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 751.950 100.950 754.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 694.950 98.550 699.450 100.050 ;
        RECT 707.100 99.150 708.900 100.950 ;
        RECT 694.950 97.950 699.000 98.550 ;
        RECT 713.700 93.600 714.900 100.950 ;
        RECT 684.000 87.900 690.600 88.800 ;
        RECT 684.000 87.600 684.900 87.900 ;
        RECT 683.100 81.600 684.900 87.600 ;
        RECT 689.100 87.600 690.600 87.900 ;
        RECT 686.100 81.000 687.900 87.000 ;
        RECT 689.100 81.600 690.900 87.600 ;
        RECT 692.100 81.000 693.900 87.600 ;
        RECT 707.400 81.000 709.200 93.600 ;
        RECT 712.500 92.100 714.900 93.600 ;
        RECT 712.500 81.600 714.300 92.100 ;
        RECT 715.200 89.100 717.000 90.900 ;
        RECT 732.000 88.800 732.900 100.950 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 732.000 87.900 738.600 88.800 ;
        RECT 732.000 87.600 732.900 87.900 ;
        RECT 715.500 81.000 717.300 87.600 ;
        RECT 731.100 81.600 732.900 87.600 ;
        RECT 737.100 87.600 738.600 87.900 ;
        RECT 755.700 87.600 756.900 100.950 ;
        RECT 767.550 100.050 768.450 104.550 ;
        RECT 773.100 103.050 774.900 104.850 ;
        RECT 776.700 103.050 777.900 108.300 ;
        RECT 800.700 107.400 804.300 108.300 ;
        RECT 821.100 108.300 825.300 109.200 ;
        RECT 781.950 105.450 784.050 106.050 ;
        RECT 787.950 105.450 790.050 106.050 ;
        RECT 778.950 103.050 780.750 104.850 ;
        RECT 781.950 104.550 790.050 105.450 ;
        RECT 781.950 103.950 784.050 104.550 ;
        RECT 787.950 103.950 790.050 104.550 ;
        RECT 797.100 103.050 798.900 104.850 ;
        RECT 800.700 103.050 801.900 107.400 ;
        RECT 803.100 103.050 804.900 104.850 ;
        RECT 818.250 103.050 820.050 104.850 ;
        RECT 821.100 103.050 822.300 108.300 ;
        RECT 831.000 105.450 835.050 106.050 ;
        RECT 824.100 103.050 825.900 104.850 ;
        RECT 830.550 103.950 835.050 105.450 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 767.550 98.550 772.050 100.050 ;
        RECT 768.000 97.950 772.050 98.550 ;
        RECT 776.700 87.600 777.900 100.950 ;
        RECT 794.100 99.150 795.900 100.950 ;
        RECT 800.700 93.600 801.900 100.950 ;
        RECT 734.100 81.000 735.900 87.000 ;
        RECT 737.100 81.600 738.900 87.600 ;
        RECT 740.100 81.000 741.900 87.600 ;
        RECT 752.100 81.000 753.900 87.600 ;
        RECT 755.100 81.600 756.900 87.600 ;
        RECT 758.100 81.000 759.900 87.600 ;
        RECT 773.100 81.000 774.900 87.600 ;
        RECT 776.100 81.600 777.900 87.600 ;
        RECT 779.100 81.000 780.900 87.600 ;
        RECT 794.400 81.000 796.200 93.600 ;
        RECT 799.500 92.100 801.900 93.600 ;
        RECT 799.500 81.600 801.300 92.100 ;
        RECT 802.200 89.100 804.000 90.900 ;
        RECT 821.100 87.600 822.300 100.950 ;
        RECT 830.550 100.050 831.450 103.950 ;
        RECT 836.250 103.050 838.050 104.850 ;
        RECT 842.100 103.050 843.300 110.400 ;
        RECT 863.100 108.600 864.900 116.400 ;
        RECT 867.600 110.400 869.400 117.000 ;
        RECT 870.600 112.200 872.400 116.400 ;
        RECT 870.600 110.400 873.300 112.200 ;
        RECT 885.000 110.400 886.800 117.000 ;
        RECT 889.500 111.600 891.300 116.400 ;
        RECT 892.500 113.400 894.300 117.000 ;
        RECT 910.800 113.400 912.900 117.000 ;
        RECT 914.100 113.400 915.900 116.400 ;
        RECT 917.100 113.400 918.900 117.000 ;
        RECT 920.100 113.400 922.800 116.400 ;
        RECT 914.700 112.500 915.600 113.400 ;
        RECT 921.900 112.500 922.800 113.400 ;
        RECT 914.700 111.600 927.300 112.500 ;
        RECT 889.500 110.400 894.600 111.600 ;
        RECT 869.700 108.600 871.500 109.500 ;
        RECT 863.100 107.700 871.500 108.600 ;
        RECT 850.950 105.450 853.050 106.050 ;
        RECT 856.950 105.450 859.050 106.050 ;
        RECT 848.100 103.050 849.900 104.850 ;
        RECT 850.950 104.550 859.050 105.450 ;
        RECT 850.950 103.950 853.050 104.550 ;
        RECT 856.950 103.950 859.050 104.550 ;
        RECT 863.250 103.050 865.050 104.850 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 863.100 100.950 865.200 103.050 ;
        RECT 830.550 98.550 835.050 100.050 ;
        RECT 839.250 99.150 841.050 100.950 ;
        RECT 831.000 97.950 835.050 98.550 ;
        RECT 842.100 95.400 843.000 100.950 ;
        RECT 845.100 99.150 846.900 100.950 ;
        RECT 847.950 96.450 850.050 97.050 ;
        RECT 856.950 96.450 859.050 97.050 ;
        RECT 847.950 95.550 859.050 96.450 ;
        RECT 842.100 94.500 846.900 95.400 ;
        RECT 847.950 94.950 850.050 95.550 ;
        RECT 856.950 94.950 859.050 95.550 ;
        RECT 836.100 92.400 843.900 93.300 ;
        RECT 802.500 81.000 804.300 87.600 ;
        RECT 818.100 81.000 819.900 87.600 ;
        RECT 821.100 81.600 822.900 87.600 ;
        RECT 824.100 81.000 825.900 87.600 ;
        RECT 836.100 81.600 837.900 92.400 ;
        RECT 839.100 81.000 840.900 91.500 ;
        RECT 842.100 82.500 843.900 92.400 ;
        RECT 845.100 83.400 846.900 94.500 ;
        RECT 848.100 82.500 849.900 93.600 ;
        RECT 866.100 87.600 867.000 107.700 ;
        RECT 872.400 103.050 873.300 110.400 ;
        RECT 886.950 109.050 889.050 109.200 ;
        RECT 883.950 107.100 889.050 109.050 ;
        RECT 883.950 106.950 888.000 107.100 ;
        RECT 884.100 103.050 885.900 104.850 ;
        RECT 890.250 103.050 892.050 104.850 ;
        RECT 893.700 103.050 894.600 110.400 ;
        RECT 916.950 103.050 918.750 104.850 ;
        RECT 926.100 103.050 927.300 111.600 ;
        RECT 868.500 100.950 870.600 103.050 ;
        RECT 871.800 100.950 873.900 103.050 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 889.950 100.950 892.050 103.050 ;
        RECT 892.950 100.950 895.050 103.050 ;
        RECT 910.800 100.950 912.900 103.050 ;
        RECT 916.950 100.950 919.050 103.050 ;
        RECT 919.950 100.950 922.050 103.050 ;
        RECT 925.500 100.950 927.600 103.050 ;
        RECT 868.200 99.150 870.000 100.950 ;
        RECT 872.400 93.600 873.300 100.950 ;
        RECT 887.250 99.150 889.050 100.950 ;
        RECT 893.700 93.600 894.600 100.950 ;
        RECT 911.100 99.150 912.900 100.950 ;
        RECT 920.250 99.150 922.050 100.950 ;
        RECT 842.100 81.600 849.900 82.500 ;
        RECT 863.100 81.000 864.900 87.600 ;
        RECT 866.100 81.600 867.900 87.600 ;
        RECT 869.100 81.000 870.900 93.000 ;
        RECT 872.100 81.600 873.900 93.600 ;
        RECT 884.100 92.700 891.900 93.600 ;
        RECT 884.100 81.600 885.900 92.700 ;
        RECT 887.100 81.000 888.900 91.800 ;
        RECT 890.100 81.600 891.900 92.700 ;
        RECT 893.100 81.600 894.900 93.600 ;
        RECT 908.100 91.500 915.900 92.400 ;
        RECT 908.100 81.600 909.900 91.500 ;
        RECT 911.100 81.000 912.900 90.600 ;
        RECT 914.100 82.500 915.900 91.500 ;
        RECT 917.100 91.200 924.900 92.100 ;
        RECT 917.100 83.400 918.900 91.200 ;
        RECT 920.100 82.500 921.900 90.300 ;
        RECT 914.100 81.600 921.900 82.500 ;
        RECT 923.100 82.500 924.900 91.200 ;
        RECT 926.100 91.200 927.300 100.950 ;
        RECT 926.100 83.400 927.900 91.200 ;
        RECT 929.100 82.500 930.900 91.800 ;
        RECT 923.100 81.600 930.900 82.500 ;
        RECT 14.100 71.400 15.900 77.400 ;
        RECT 17.100 71.400 18.900 78.000 ;
        RECT 14.700 58.050 15.900 71.400 ;
        RECT 32.400 65.400 34.200 78.000 ;
        RECT 37.500 66.900 39.300 77.400 ;
        RECT 40.500 71.400 42.300 78.000 ;
        RECT 53.700 71.400 55.500 78.000 ;
        RECT 40.200 68.100 42.000 69.900 ;
        RECT 54.000 68.100 55.800 69.900 ;
        RECT 56.700 66.900 58.500 77.400 ;
        RECT 37.500 65.400 39.900 66.900 ;
        RECT 16.950 63.450 19.050 64.050 ;
        RECT 34.950 63.450 37.050 64.050 ;
        RECT 16.950 62.550 37.050 63.450 ;
        RECT 16.950 61.950 19.050 62.550 ;
        RECT 34.950 61.950 37.050 62.550 ;
        RECT 17.100 58.050 18.900 59.850 ;
        RECT 32.100 58.050 33.900 59.850 ;
        RECT 38.700 58.050 39.900 65.400 ;
        RECT 56.100 65.400 58.500 66.900 ;
        RECT 61.800 65.400 63.600 78.000 ;
        RECT 77.100 71.400 78.900 78.000 ;
        RECT 80.100 71.400 81.900 77.400 ;
        RECT 83.100 72.000 84.900 78.000 ;
        RECT 80.400 71.100 81.900 71.400 ;
        RECT 86.100 71.400 87.900 77.400 ;
        RECT 86.100 71.100 87.000 71.400 ;
        RECT 80.400 70.200 87.000 71.100 ;
        RECT 56.100 58.050 57.300 65.400 ;
        RECT 62.100 58.050 63.900 59.850 ;
        RECT 80.100 58.050 81.900 59.850 ;
        RECT 86.100 58.050 87.000 70.200 ;
        RECT 101.400 65.400 103.200 78.000 ;
        RECT 106.500 66.900 108.300 77.400 ;
        RECT 109.500 71.400 111.300 78.000 ;
        RECT 109.200 68.100 111.000 69.900 ;
        RECT 106.500 65.400 108.900 66.900 ;
        RECT 122.400 65.400 124.200 78.000 ;
        RECT 127.500 66.900 129.300 77.400 ;
        RECT 130.500 71.400 132.300 78.000 ;
        RECT 143.100 71.400 144.900 77.400 ;
        RECT 146.100 72.000 147.900 78.000 ;
        RECT 144.000 71.100 144.900 71.400 ;
        RECT 149.100 71.400 150.900 77.400 ;
        RECT 152.100 71.400 153.900 78.000 ;
        RECT 149.100 71.100 150.600 71.400 ;
        RECT 144.000 70.200 150.600 71.100 ;
        RECT 130.200 68.100 132.000 69.900 ;
        RECT 127.500 65.400 129.900 66.900 ;
        RECT 101.100 58.050 102.900 59.850 ;
        RECT 107.700 58.050 108.900 65.400 ;
        RECT 122.100 58.050 123.900 59.850 ;
        RECT 128.700 58.050 129.900 65.400 ;
        RECT 144.000 58.050 144.900 70.200 ;
        RECT 154.950 69.450 157.050 70.050 ;
        RECT 160.950 69.450 163.050 70.050 ;
        RECT 154.950 68.550 163.050 69.450 ;
        RECT 154.950 67.950 157.050 68.550 ;
        RECT 160.950 67.950 163.050 68.550 ;
        RECT 167.100 65.400 168.900 77.400 ;
        RECT 170.100 66.300 171.900 77.400 ;
        RECT 173.100 67.200 174.900 78.000 ;
        RECT 176.100 66.300 177.900 77.400 ;
        RECT 191.700 71.400 193.500 78.000 ;
        RECT 192.000 68.100 193.800 69.900 ;
        RECT 194.700 66.900 196.500 77.400 ;
        RECT 170.100 65.400 177.900 66.300 ;
        RECT 194.100 65.400 196.500 66.900 ;
        RECT 199.800 65.400 201.600 78.000 ;
        RECT 215.100 71.400 216.900 77.400 ;
        RECT 218.100 72.000 219.900 78.000 ;
        RECT 216.000 71.100 216.900 71.400 ;
        RECT 221.100 71.400 222.900 77.400 ;
        RECT 224.100 71.400 225.900 78.000 ;
        RECT 236.100 71.400 237.900 77.400 ;
        RECT 239.100 71.400 240.900 78.000 ;
        RECT 254.100 71.400 255.900 78.000 ;
        RECT 257.100 71.400 258.900 77.400 ;
        RECT 260.100 72.000 261.900 78.000 ;
        RECT 221.100 71.100 222.600 71.400 ;
        RECT 216.000 70.200 222.600 71.100 ;
        RECT 151.950 63.450 154.050 64.050 ;
        RECT 160.950 63.450 163.050 64.050 ;
        RECT 151.950 62.550 163.050 63.450 ;
        RECT 151.950 61.950 154.050 62.550 ;
        RECT 160.950 61.950 163.050 62.550 ;
        RECT 149.100 58.050 150.900 59.850 ;
        RECT 167.400 58.050 168.300 65.400 ;
        RECT 178.950 60.450 183.000 61.050 ;
        RECT 172.950 58.050 174.750 59.850 ;
        RECT 178.950 58.950 183.450 60.450 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 14.700 45.600 15.900 55.950 ;
        RECT 35.100 54.150 36.900 55.950 ;
        RECT 38.700 51.600 39.900 55.950 ;
        RECT 41.100 54.150 42.900 55.950 ;
        RECT 53.100 54.150 54.900 55.950 ;
        RECT 56.100 51.600 57.300 55.950 ;
        RECT 59.100 54.150 60.900 55.950 ;
        RECT 77.100 54.150 78.900 55.950 ;
        RECT 83.100 54.150 84.900 55.950 ;
        RECT 86.100 52.200 87.000 55.950 ;
        RECT 104.100 54.150 105.900 55.950 ;
        RECT 38.700 50.700 42.300 51.600 ;
        RECT 32.100 47.700 39.900 49.050 ;
        RECT 14.100 42.600 15.900 45.600 ;
        RECT 17.100 42.000 18.900 45.600 ;
        RECT 32.100 42.600 33.900 47.700 ;
        RECT 35.100 42.000 36.900 46.800 ;
        RECT 38.100 42.600 39.900 47.700 ;
        RECT 41.100 48.600 42.300 50.700 ;
        RECT 53.700 50.700 57.300 51.600 ;
        RECT 53.700 48.600 54.900 50.700 ;
        RECT 41.100 42.600 42.900 48.600 ;
        RECT 53.100 42.600 54.900 48.600 ;
        RECT 56.100 47.700 63.900 49.050 ;
        RECT 56.100 42.600 57.900 47.700 ;
        RECT 59.100 42.000 60.900 46.800 ;
        RECT 62.100 42.600 63.900 47.700 ;
        RECT 77.100 42.000 78.900 51.600 ;
        RECT 83.700 51.000 87.000 52.200 ;
        RECT 107.700 51.600 108.900 55.950 ;
        RECT 110.100 54.150 111.900 55.950 ;
        RECT 125.100 54.150 126.900 55.950 ;
        RECT 128.700 51.600 129.900 55.950 ;
        RECT 131.100 54.150 132.900 55.950 ;
        RECT 144.000 52.200 144.900 55.950 ;
        RECT 146.100 54.150 147.900 55.950 ;
        RECT 152.100 54.150 153.900 55.950 ;
        RECT 83.700 42.600 85.500 51.000 ;
        RECT 107.700 50.700 111.300 51.600 ;
        RECT 128.700 50.700 132.300 51.600 ;
        RECT 144.000 51.000 147.300 52.200 ;
        RECT 101.100 47.700 108.900 49.050 ;
        RECT 101.100 42.600 102.900 47.700 ;
        RECT 104.100 42.000 105.900 46.800 ;
        RECT 107.100 42.600 108.900 47.700 ;
        RECT 110.100 48.600 111.300 50.700 ;
        RECT 110.100 42.600 111.900 48.600 ;
        RECT 122.100 47.700 129.900 49.050 ;
        RECT 122.100 42.600 123.900 47.700 ;
        RECT 125.100 42.000 126.900 46.800 ;
        RECT 128.100 42.600 129.900 47.700 ;
        RECT 131.100 48.600 132.300 50.700 ;
        RECT 131.100 42.600 132.900 48.600 ;
        RECT 145.500 42.600 147.300 51.000 ;
        RECT 152.100 42.000 153.900 51.600 ;
        RECT 167.400 48.600 168.300 55.950 ;
        RECT 169.950 54.150 171.750 55.950 ;
        RECT 176.100 54.150 177.900 55.950 ;
        RECT 182.550 55.050 183.450 58.950 ;
        RECT 194.100 58.050 195.300 65.400 ;
        RECT 200.100 58.050 201.900 59.850 ;
        RECT 216.000 58.050 216.900 70.200 ;
        RECT 221.100 58.050 222.900 59.850 ;
        RECT 236.700 58.050 237.900 71.400 ;
        RECT 257.400 71.100 258.900 71.400 ;
        RECT 263.100 71.400 264.900 77.400 ;
        RECT 278.100 71.400 279.900 78.000 ;
        RECT 281.100 71.400 282.900 77.400 ;
        RECT 284.100 72.000 285.900 78.000 ;
        RECT 263.100 71.100 264.000 71.400 ;
        RECT 257.400 70.200 264.000 71.100 ;
        RECT 281.400 71.100 282.900 71.400 ;
        RECT 287.100 71.400 288.900 77.400 ;
        RECT 299.700 71.400 301.500 78.000 ;
        RECT 287.100 71.100 288.000 71.400 ;
        RECT 281.400 70.200 288.000 71.100 ;
        RECT 239.100 58.050 240.900 59.850 ;
        RECT 257.100 58.050 258.900 59.850 ;
        RECT 263.100 58.050 264.000 70.200 ;
        RECT 283.950 63.450 286.050 64.050 ;
        RECT 275.550 62.550 286.050 63.450 ;
        RECT 275.550 60.450 276.450 62.550 ;
        RECT 283.950 61.950 286.050 62.550 ;
        RECT 272.550 59.550 276.450 60.450 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 220.950 55.950 223.050 58.050 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 181.950 52.950 184.050 55.050 ;
        RECT 191.100 54.150 192.900 55.950 ;
        RECT 194.100 51.600 195.300 55.950 ;
        RECT 197.100 54.150 198.900 55.950 ;
        RECT 191.700 50.700 195.300 51.600 ;
        RECT 216.000 52.200 216.900 55.950 ;
        RECT 218.100 54.150 219.900 55.950 ;
        RECT 224.100 54.150 225.900 55.950 ;
        RECT 216.000 51.000 219.300 52.200 ;
        RECT 191.700 48.600 192.900 50.700 ;
        RECT 167.400 47.400 172.500 48.600 ;
        RECT 167.700 42.000 169.500 45.600 ;
        RECT 170.700 42.600 172.500 47.400 ;
        RECT 175.200 42.000 177.000 48.600 ;
        RECT 191.100 42.600 192.900 48.600 ;
        RECT 194.100 47.700 201.900 49.050 ;
        RECT 194.100 42.600 195.900 47.700 ;
        RECT 197.100 42.000 198.900 46.800 ;
        RECT 200.100 42.600 201.900 47.700 ;
        RECT 217.500 42.600 219.300 51.000 ;
        RECT 224.100 42.000 225.900 51.600 ;
        RECT 236.700 45.600 237.900 55.950 ;
        RECT 254.100 54.150 255.900 55.950 ;
        RECT 260.100 54.150 261.900 55.950 ;
        RECT 263.100 52.200 264.000 55.950 ;
        RECT 265.950 54.450 268.050 55.050 ;
        RECT 272.550 54.450 273.450 59.550 ;
        RECT 281.100 58.050 282.900 59.850 ;
        RECT 287.100 58.050 288.000 70.200 ;
        RECT 300.000 68.100 301.800 69.900 ;
        RECT 302.700 66.900 304.500 77.400 ;
        RECT 302.100 65.400 304.500 66.900 ;
        RECT 307.800 65.400 309.600 78.000 ;
        RECT 323.400 65.400 325.200 78.000 ;
        RECT 328.500 66.900 330.300 77.400 ;
        RECT 331.500 71.400 333.300 78.000 ;
        RECT 331.200 68.100 333.000 69.900 ;
        RECT 328.500 65.400 330.900 66.900 ;
        RECT 344.400 65.400 346.200 78.000 ;
        RECT 349.500 66.900 351.300 77.400 ;
        RECT 352.500 71.400 354.300 78.000 ;
        RECT 365.100 71.400 366.900 77.400 ;
        RECT 368.100 72.000 369.900 78.000 ;
        RECT 366.000 71.100 366.900 71.400 ;
        RECT 371.100 71.400 372.900 77.400 ;
        RECT 374.100 71.400 375.900 78.000 ;
        RECT 371.100 71.100 372.600 71.400 ;
        RECT 366.000 70.200 372.600 71.100 ;
        RECT 352.200 68.100 354.000 69.900 ;
        RECT 349.500 65.400 351.900 66.900 ;
        RECT 289.950 63.450 292.050 64.050 ;
        RECT 298.950 63.450 301.050 64.050 ;
        RECT 289.950 62.550 301.050 63.450 ;
        RECT 289.950 61.950 292.050 62.550 ;
        RECT 298.950 61.950 301.050 62.550 ;
        RECT 302.100 58.050 303.300 65.400 ;
        RECT 304.950 63.450 307.050 64.050 ;
        RECT 325.950 63.450 328.050 64.050 ;
        RECT 304.950 62.550 328.050 63.450 ;
        RECT 304.950 61.950 307.050 62.550 ;
        RECT 325.950 61.950 328.050 62.550 ;
        RECT 308.100 58.050 309.900 59.850 ;
        RECT 323.100 58.050 324.900 59.850 ;
        RECT 329.700 58.050 330.900 65.400 ;
        RECT 344.100 58.050 345.900 59.850 ;
        RECT 350.700 58.050 351.900 65.400 ;
        RECT 360.000 60.450 364.050 61.050 ;
        RECT 359.550 58.950 364.050 60.450 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 265.950 53.550 273.450 54.450 ;
        RECT 278.100 54.150 279.900 55.950 ;
        RECT 284.100 54.150 285.900 55.950 ;
        RECT 265.950 52.950 268.050 53.550 ;
        RECT 287.100 52.200 288.000 55.950 ;
        RECT 299.100 54.150 300.900 55.950 ;
        RECT 236.100 42.600 237.900 45.600 ;
        RECT 239.100 42.000 240.900 45.600 ;
        RECT 254.100 42.000 255.900 51.600 ;
        RECT 260.700 51.000 264.000 52.200 ;
        RECT 260.700 42.600 262.500 51.000 ;
        RECT 278.100 42.000 279.900 51.600 ;
        RECT 284.700 51.000 288.000 52.200 ;
        RECT 302.100 51.600 303.300 55.950 ;
        RECT 305.100 54.150 306.900 55.950 ;
        RECT 326.100 54.150 327.900 55.950 ;
        RECT 284.700 42.600 286.500 51.000 ;
        RECT 299.700 50.700 303.300 51.600 ;
        RECT 329.700 51.600 330.900 55.950 ;
        RECT 332.100 54.150 333.900 55.950 ;
        RECT 347.100 54.150 348.900 55.950 ;
        RECT 350.700 51.600 351.900 55.950 ;
        RECT 353.100 54.150 354.900 55.950 ;
        RECT 359.550 55.050 360.450 58.950 ;
        RECT 366.000 58.050 366.900 70.200 ;
        RECT 389.100 65.400 390.900 77.400 ;
        RECT 392.100 66.300 393.900 77.400 ;
        RECT 395.100 67.200 396.900 78.000 ;
        RECT 398.100 66.300 399.900 77.400 ;
        RECT 413.700 71.400 415.500 78.000 ;
        RECT 414.000 68.100 415.800 69.900 ;
        RECT 416.700 66.900 418.500 77.400 ;
        RECT 392.100 65.400 399.900 66.300 ;
        RECT 416.100 65.400 418.500 66.900 ;
        RECT 421.800 65.400 423.600 78.000 ;
        RECT 437.100 71.400 438.900 78.000 ;
        RECT 440.100 71.400 441.900 77.400 ;
        RECT 443.100 72.000 444.900 78.000 ;
        RECT 440.400 71.100 441.900 71.400 ;
        RECT 446.100 71.400 447.900 77.400 ;
        RECT 446.100 71.100 447.000 71.400 ;
        RECT 440.400 70.200 447.000 71.100 ;
        RECT 371.100 58.050 372.900 59.850 ;
        RECT 389.400 58.050 390.300 65.400 ;
        RECT 394.950 58.050 396.750 59.850 ;
        RECT 416.100 58.050 417.300 65.400 ;
        RECT 432.000 60.450 436.050 61.050 ;
        RECT 422.100 58.050 423.900 59.850 ;
        RECT 431.550 58.950 436.050 60.450 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 355.950 53.550 360.450 55.050 ;
        RECT 355.950 52.950 360.000 53.550 ;
        RECT 366.000 52.200 366.900 55.950 ;
        RECT 368.100 54.150 369.900 55.950 ;
        RECT 374.100 54.150 375.900 55.950 ;
        RECT 329.700 50.700 333.300 51.600 ;
        RECT 350.700 50.700 354.300 51.600 ;
        RECT 366.000 51.000 369.300 52.200 ;
        RECT 299.700 48.600 300.900 50.700 ;
        RECT 299.100 42.600 300.900 48.600 ;
        RECT 302.100 47.700 309.900 49.050 ;
        RECT 302.100 42.600 303.900 47.700 ;
        RECT 305.100 42.000 306.900 46.800 ;
        RECT 308.100 42.600 309.900 47.700 ;
        RECT 323.100 47.700 330.900 49.050 ;
        RECT 323.100 42.600 324.900 47.700 ;
        RECT 326.100 42.000 327.900 46.800 ;
        RECT 329.100 42.600 330.900 47.700 ;
        RECT 332.100 48.600 333.300 50.700 ;
        RECT 332.100 42.600 333.900 48.600 ;
        RECT 344.100 47.700 351.900 49.050 ;
        RECT 344.100 42.600 345.900 47.700 ;
        RECT 347.100 42.000 348.900 46.800 ;
        RECT 350.100 42.600 351.900 47.700 ;
        RECT 353.100 48.600 354.300 50.700 ;
        RECT 353.100 42.600 354.900 48.600 ;
        RECT 367.500 42.600 369.300 51.000 ;
        RECT 374.100 42.000 375.900 51.600 ;
        RECT 389.400 48.600 390.300 55.950 ;
        RECT 391.950 54.150 393.750 55.950 ;
        RECT 398.100 54.150 399.900 55.950 ;
        RECT 413.100 54.150 414.900 55.950 ;
        RECT 416.100 51.600 417.300 55.950 ;
        RECT 419.100 54.150 420.900 55.950 ;
        RECT 427.950 55.050 430.050 58.050 ;
        RECT 424.950 54.000 430.050 55.050 ;
        RECT 431.550 55.050 432.450 58.950 ;
        RECT 440.100 58.050 441.900 59.850 ;
        RECT 446.100 58.050 447.000 70.200 ;
        RECT 461.100 66.300 462.900 77.400 ;
        RECT 464.100 67.200 465.900 78.000 ;
        RECT 467.100 66.300 468.900 77.400 ;
        RECT 461.100 65.400 468.900 66.300 ;
        RECT 470.100 65.400 471.900 77.400 ;
        RECT 485.400 65.400 487.200 78.000 ;
        RECT 490.500 66.900 492.300 77.400 ;
        RECT 493.500 71.400 495.300 78.000 ;
        RECT 493.200 68.100 495.000 69.900 ;
        RECT 490.500 65.400 492.900 66.900 ;
        RECT 506.400 65.400 508.200 78.000 ;
        RECT 511.500 66.900 513.300 77.400 ;
        RECT 514.500 71.400 516.300 78.000 ;
        RECT 514.200 68.100 516.000 69.900 ;
        RECT 511.500 65.400 513.900 66.900 ;
        RECT 530.100 66.300 531.900 77.400 ;
        RECT 533.100 67.200 534.900 78.000 ;
        RECT 536.100 66.300 537.900 77.400 ;
        RECT 530.100 65.400 537.900 66.300 ;
        RECT 539.100 65.400 540.900 77.400 ;
        RECT 554.100 71.400 555.900 77.400 ;
        RECT 557.100 71.400 558.900 78.000 ;
        RECT 448.950 63.450 451.050 64.050 ;
        RECT 466.950 63.450 469.050 64.200 ;
        RECT 448.950 62.550 469.050 63.450 ;
        RECT 448.950 61.950 451.050 62.550 ;
        RECT 466.950 62.100 469.050 62.550 ;
        RECT 464.250 58.050 466.050 59.850 ;
        RECT 470.700 58.050 471.600 65.400 ;
        RECT 485.100 58.050 486.900 59.850 ;
        RECT 491.700 58.050 492.900 65.400 ;
        RECT 496.950 60.450 501.000 61.050 ;
        RECT 496.950 58.950 501.450 60.450 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 424.950 53.550 429.450 54.000 ;
        RECT 431.550 53.550 436.050 55.050 ;
        RECT 437.100 54.150 438.900 55.950 ;
        RECT 443.100 54.150 444.900 55.950 ;
        RECT 424.950 52.950 429.000 53.550 ;
        RECT 432.000 52.950 436.050 53.550 ;
        RECT 446.100 52.200 447.000 55.950 ;
        RECT 461.100 54.150 462.900 55.950 ;
        RECT 467.250 54.150 469.050 55.950 ;
        RECT 413.700 50.700 417.300 51.600 ;
        RECT 413.700 48.600 414.900 50.700 ;
        RECT 389.400 47.400 394.500 48.600 ;
        RECT 389.700 42.000 391.500 45.600 ;
        RECT 392.700 42.600 394.500 47.400 ;
        RECT 397.200 42.000 399.000 48.600 ;
        RECT 413.100 42.600 414.900 48.600 ;
        RECT 416.100 47.700 423.900 49.050 ;
        RECT 416.100 42.600 417.900 47.700 ;
        RECT 419.100 42.000 420.900 46.800 ;
        RECT 422.100 42.600 423.900 47.700 ;
        RECT 437.100 42.000 438.900 51.600 ;
        RECT 443.700 51.000 447.000 52.200 ;
        RECT 443.700 42.600 445.500 51.000 ;
        RECT 470.700 48.600 471.600 55.950 ;
        RECT 488.100 54.150 489.900 55.950 ;
        RECT 491.700 51.600 492.900 55.950 ;
        RECT 494.100 54.150 495.900 55.950 ;
        RECT 500.550 55.050 501.450 58.950 ;
        RECT 506.100 58.050 507.900 59.850 ;
        RECT 512.700 58.050 513.900 65.400 ;
        RECT 533.250 58.050 535.050 59.850 ;
        RECT 539.700 58.050 540.600 65.400 ;
        RECT 549.000 60.450 553.050 61.050 ;
        RECT 548.550 58.950 553.050 60.450 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 496.950 53.550 501.450 55.050 ;
        RECT 509.100 54.150 510.900 55.950 ;
        RECT 496.950 52.950 501.000 53.550 ;
        RECT 512.700 51.600 513.900 55.950 ;
        RECT 515.100 54.150 516.900 55.950 ;
        RECT 530.100 54.150 531.900 55.950 ;
        RECT 536.250 54.150 538.050 55.950 ;
        RECT 491.700 50.700 495.300 51.600 ;
        RECT 512.700 50.700 516.300 51.600 ;
        RECT 462.000 42.000 463.800 48.600 ;
        RECT 466.500 47.400 471.600 48.600 ;
        RECT 485.100 47.700 492.900 49.050 ;
        RECT 466.500 42.600 468.300 47.400 ;
        RECT 469.500 42.000 471.300 45.600 ;
        RECT 485.100 42.600 486.900 47.700 ;
        RECT 488.100 42.000 489.900 46.800 ;
        RECT 491.100 42.600 492.900 47.700 ;
        RECT 494.100 48.600 495.300 50.700 ;
        RECT 494.100 42.600 495.900 48.600 ;
        RECT 506.100 47.700 513.900 49.050 ;
        RECT 506.100 42.600 507.900 47.700 ;
        RECT 509.100 42.000 510.900 46.800 ;
        RECT 512.100 42.600 513.900 47.700 ;
        RECT 515.100 48.600 516.300 50.700 ;
        RECT 539.700 48.600 540.600 55.950 ;
        RECT 541.950 54.450 544.050 55.050 ;
        RECT 548.550 54.450 549.450 58.950 ;
        RECT 554.700 58.050 555.900 71.400 ;
        RECT 572.400 65.400 574.200 78.000 ;
        RECT 577.500 66.900 579.300 77.400 ;
        RECT 580.500 71.400 582.300 78.000 ;
        RECT 596.100 71.400 597.900 77.400 ;
        RECT 599.100 72.000 600.900 78.000 ;
        RECT 597.000 71.100 597.900 71.400 ;
        RECT 602.100 71.400 603.900 77.400 ;
        RECT 605.100 71.400 606.900 78.000 ;
        RECT 602.100 71.100 603.600 71.400 ;
        RECT 597.000 70.200 603.600 71.100 ;
        RECT 580.200 68.100 582.000 69.900 ;
        RECT 577.500 65.400 579.900 66.900 ;
        RECT 557.100 58.050 558.900 59.850 ;
        RECT 572.100 58.050 573.900 59.850 ;
        RECT 578.700 58.050 579.900 65.400 ;
        RECT 597.000 58.050 597.900 70.200 ;
        RECT 617.100 65.400 618.900 77.400 ;
        RECT 620.100 66.300 621.900 77.400 ;
        RECT 623.100 67.200 624.900 78.000 ;
        RECT 626.100 66.300 627.900 77.400 ;
        RECT 638.100 71.400 639.900 77.400 ;
        RECT 641.100 72.000 642.900 78.000 ;
        RECT 620.100 65.400 627.900 66.300 ;
        RECT 639.000 71.100 639.900 71.400 ;
        RECT 644.100 71.400 645.900 77.400 ;
        RECT 647.100 71.400 648.900 78.000 ;
        RECT 659.100 71.400 660.900 78.000 ;
        RECT 662.100 71.400 663.900 77.400 ;
        RECT 665.100 71.400 666.900 78.000 ;
        RECT 680.100 71.400 681.900 77.400 ;
        RECT 683.100 72.000 684.900 78.000 ;
        RECT 644.100 71.100 645.600 71.400 ;
        RECT 639.000 70.200 645.600 71.100 ;
        RECT 604.950 63.450 607.050 64.050 ;
        RECT 610.950 63.450 613.050 64.050 ;
        RECT 604.950 62.550 613.050 63.450 ;
        RECT 604.950 61.950 607.050 62.550 ;
        RECT 610.950 61.950 613.050 62.550 ;
        RECT 602.100 58.050 603.900 59.850 ;
        RECT 617.400 58.050 618.300 65.400 ;
        RECT 622.950 58.050 624.750 59.850 ;
        RECT 639.000 58.050 639.900 70.200 ;
        RECT 644.100 58.050 645.900 59.850 ;
        RECT 662.100 58.050 663.300 71.400 ;
        RECT 681.000 71.100 681.900 71.400 ;
        RECT 686.100 71.400 687.900 77.400 ;
        RECT 689.100 71.400 690.900 78.000 ;
        RECT 704.100 71.400 705.900 77.400 ;
        RECT 707.100 72.000 708.900 78.000 ;
        RECT 686.100 71.100 687.600 71.400 ;
        RECT 681.000 70.200 687.600 71.100 ;
        RECT 705.000 71.100 705.900 71.400 ;
        RECT 710.100 71.400 711.900 77.400 ;
        RECT 713.100 71.400 714.900 78.000 ;
        RECT 728.100 71.400 729.900 77.400 ;
        RECT 731.100 72.000 732.900 78.000 ;
        RECT 710.100 71.100 711.600 71.400 ;
        RECT 705.000 70.200 711.600 71.100 ;
        RECT 729.000 71.100 729.900 71.400 ;
        RECT 734.100 71.400 735.900 77.400 ;
        RECT 737.100 71.400 738.900 78.000 ;
        RECT 749.100 71.400 750.900 77.400 ;
        RECT 752.100 71.400 753.900 78.000 ;
        RECT 764.100 71.400 765.900 78.000 ;
        RECT 767.100 71.400 768.900 77.400 ;
        RECT 770.100 71.400 771.900 78.000 ;
        RECT 782.100 71.400 783.900 77.400 ;
        RECT 785.100 72.000 786.900 78.000 ;
        RECT 734.100 71.100 735.600 71.400 ;
        RECT 729.000 70.200 735.600 71.100 ;
        RECT 670.950 60.450 673.050 61.050 ;
        RECT 676.950 60.450 679.050 61.050 ;
        RECT 670.950 59.550 679.050 60.450 ;
        RECT 670.950 58.950 673.050 59.550 ;
        RECT 676.950 58.950 679.050 59.550 ;
        RECT 681.000 58.050 681.900 70.200 ;
        RECT 686.100 58.050 687.900 59.850 ;
        RECT 705.000 58.050 705.900 70.200 ;
        RECT 710.100 58.050 711.900 59.850 ;
        RECT 729.000 58.050 729.900 70.200 ;
        RECT 734.100 58.050 735.900 59.850 ;
        RECT 749.700 58.050 750.900 71.400 ;
        RECT 752.100 58.050 753.900 59.850 ;
        RECT 767.700 58.050 768.900 71.400 ;
        RECT 783.000 71.100 783.900 71.400 ;
        RECT 788.100 71.400 789.900 77.400 ;
        RECT 791.100 71.400 792.900 78.000 ;
        RECT 788.100 71.100 789.600 71.400 ;
        RECT 783.000 70.200 789.600 71.100 ;
        RECT 783.000 58.050 783.900 70.200 ;
        RECT 806.100 66.300 807.900 77.400 ;
        RECT 809.100 67.200 810.900 78.000 ;
        RECT 812.100 66.300 813.900 77.400 ;
        RECT 806.100 65.400 813.900 66.300 ;
        RECT 815.100 65.400 816.900 77.400 ;
        RECT 827.700 71.400 829.500 78.000 ;
        RECT 828.000 68.100 829.800 69.900 ;
        RECT 830.700 66.900 832.500 77.400 ;
        RECT 830.100 65.400 832.500 66.900 ;
        RECT 835.800 65.400 837.600 78.000 ;
        RECT 851.100 71.400 852.900 77.400 ;
        RECT 854.100 72.000 855.900 78.000 ;
        RECT 852.000 71.100 852.900 71.400 ;
        RECT 857.100 71.400 858.900 77.400 ;
        RECT 860.100 71.400 861.900 78.000 ;
        RECT 875.100 71.400 876.900 77.400 ;
        RECT 878.100 72.000 879.900 78.000 ;
        RECT 857.100 71.100 858.600 71.400 ;
        RECT 852.000 70.200 858.600 71.100 ;
        RECT 876.000 71.100 876.900 71.400 ;
        RECT 881.100 71.400 882.900 77.400 ;
        RECT 884.100 71.400 885.900 78.000 ;
        RECT 881.100 71.100 882.600 71.400 ;
        RECT 876.000 70.200 882.600 71.100 ;
        RECT 788.100 58.050 789.900 59.850 ;
        RECT 809.250 58.050 811.050 59.850 ;
        RECT 815.700 58.050 816.600 65.400 ;
        RECT 830.100 58.050 831.300 65.400 ;
        RECT 836.100 58.050 837.900 59.850 ;
        RECT 852.000 58.050 852.900 70.200 ;
        RECT 862.950 60.450 867.000 61.050 ;
        RECT 857.100 58.050 858.900 59.850 ;
        RECT 862.950 58.950 867.450 60.450 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 580.950 55.950 583.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 769.950 55.950 772.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 811.950 55.950 814.050 58.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 835.950 55.950 838.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 859.950 55.950 862.050 58.050 ;
        RECT 541.950 53.550 549.450 54.450 ;
        RECT 541.950 52.950 544.050 53.550 ;
        RECT 515.100 42.600 516.900 48.600 ;
        RECT 531.000 42.000 532.800 48.600 ;
        RECT 535.500 47.400 540.600 48.600 ;
        RECT 535.500 42.600 537.300 47.400 ;
        RECT 554.700 45.600 555.900 55.950 ;
        RECT 559.950 54.450 562.050 55.050 ;
        RECT 565.950 54.450 568.050 55.050 ;
        RECT 559.950 53.550 568.050 54.450 ;
        RECT 575.100 54.150 576.900 55.950 ;
        RECT 559.950 52.950 562.050 53.550 ;
        RECT 565.950 52.950 568.050 53.550 ;
        RECT 578.700 51.600 579.900 55.950 ;
        RECT 581.100 54.150 582.900 55.950 ;
        RECT 597.000 52.200 597.900 55.950 ;
        RECT 599.100 54.150 600.900 55.950 ;
        RECT 605.100 54.150 606.900 55.950 ;
        RECT 578.700 50.700 582.300 51.600 ;
        RECT 597.000 51.000 600.300 52.200 ;
        RECT 572.100 47.700 579.900 49.050 ;
        RECT 538.500 42.000 540.300 45.600 ;
        RECT 554.100 42.600 555.900 45.600 ;
        RECT 557.100 42.000 558.900 45.600 ;
        RECT 559.950 45.450 562.050 46.050 ;
        RECT 565.950 45.450 568.050 46.050 ;
        RECT 559.950 44.550 568.050 45.450 ;
        RECT 559.950 43.950 562.050 44.550 ;
        RECT 565.950 43.950 568.050 44.550 ;
        RECT 572.100 42.600 573.900 47.700 ;
        RECT 575.100 42.000 576.900 46.800 ;
        RECT 578.100 42.600 579.900 47.700 ;
        RECT 581.100 48.600 582.300 50.700 ;
        RECT 581.100 42.600 582.900 48.600 ;
        RECT 598.500 42.600 600.300 51.000 ;
        RECT 605.100 42.000 606.900 51.600 ;
        RECT 617.400 48.600 618.300 55.950 ;
        RECT 619.950 54.150 621.750 55.950 ;
        RECT 626.100 54.150 627.900 55.950 ;
        RECT 639.000 52.200 639.900 55.950 ;
        RECT 641.100 54.150 642.900 55.950 ;
        RECT 647.100 54.150 648.900 55.950 ;
        RECT 659.250 54.150 661.050 55.950 ;
        RECT 639.000 51.000 642.300 52.200 ;
        RECT 617.400 47.400 622.500 48.600 ;
        RECT 617.700 42.000 619.500 45.600 ;
        RECT 620.700 42.600 622.500 47.400 ;
        RECT 625.200 42.000 627.000 48.600 ;
        RECT 640.500 42.600 642.300 51.000 ;
        RECT 647.100 42.000 648.900 51.600 ;
        RECT 662.100 50.700 663.300 55.950 ;
        RECT 665.100 54.150 666.900 55.950 ;
        RECT 681.000 52.200 681.900 55.950 ;
        RECT 683.100 54.150 684.900 55.950 ;
        RECT 689.100 54.150 690.900 55.950 ;
        RECT 705.000 52.200 705.900 55.950 ;
        RECT 707.100 54.150 708.900 55.950 ;
        RECT 713.100 54.150 714.900 55.950 ;
        RECT 729.000 52.200 729.900 55.950 ;
        RECT 731.100 54.150 732.900 55.950 ;
        RECT 737.100 54.150 738.900 55.950 ;
        RECT 681.000 51.000 684.300 52.200 ;
        RECT 662.100 49.800 666.300 50.700 ;
        RECT 659.400 42.000 661.200 48.600 ;
        RECT 664.500 42.600 666.300 49.800 ;
        RECT 682.500 42.600 684.300 51.000 ;
        RECT 689.100 42.000 690.900 51.600 ;
        RECT 705.000 51.000 708.300 52.200 ;
        RECT 706.500 42.600 708.300 51.000 ;
        RECT 713.100 42.000 714.900 51.600 ;
        RECT 729.000 51.000 732.300 52.200 ;
        RECT 730.500 42.600 732.300 51.000 ;
        RECT 737.100 42.000 738.900 51.600 ;
        RECT 749.700 45.600 750.900 55.950 ;
        RECT 764.100 54.150 765.900 55.950 ;
        RECT 767.700 50.700 768.900 55.950 ;
        RECT 769.950 54.150 771.750 55.950 ;
        RECT 783.000 52.200 783.900 55.950 ;
        RECT 785.100 54.150 786.900 55.950 ;
        RECT 791.100 54.150 792.900 55.950 ;
        RECT 806.100 54.150 807.900 55.950 ;
        RECT 812.250 54.150 814.050 55.950 ;
        RECT 783.000 51.000 786.300 52.200 ;
        RECT 764.700 49.800 768.900 50.700 ;
        RECT 749.100 42.600 750.900 45.600 ;
        RECT 752.100 42.000 753.900 45.600 ;
        RECT 764.700 42.600 766.500 49.800 ;
        RECT 769.800 42.000 771.600 48.600 ;
        RECT 784.500 42.600 786.300 51.000 ;
        RECT 791.100 42.000 792.900 51.600 ;
        RECT 796.950 51.450 799.050 52.050 ;
        RECT 808.950 51.450 811.050 52.050 ;
        RECT 796.950 50.550 811.050 51.450 ;
        RECT 796.950 49.950 799.050 50.550 ;
        RECT 808.950 49.950 811.050 50.550 ;
        RECT 815.700 48.600 816.600 55.950 ;
        RECT 827.100 54.150 828.900 55.950 ;
        RECT 830.100 51.600 831.300 55.950 ;
        RECT 833.100 54.150 834.900 55.950 ;
        RECT 827.700 50.700 831.300 51.600 ;
        RECT 852.000 52.200 852.900 55.950 ;
        RECT 854.100 54.150 855.900 55.950 ;
        RECT 860.100 54.150 861.900 55.950 ;
        RECT 866.550 54.900 867.450 58.950 ;
        RECT 876.000 58.050 876.900 70.200 ;
        RECT 896.100 65.400 897.900 77.400 ;
        RECT 899.100 66.300 900.900 77.400 ;
        RECT 902.100 67.200 903.900 78.000 ;
        RECT 905.100 66.300 906.900 77.400 ;
        RECT 917.100 71.400 918.900 77.400 ;
        RECT 920.100 72.000 921.900 78.000 ;
        RECT 899.100 65.400 906.900 66.300 ;
        RECT 918.000 71.100 918.900 71.400 ;
        RECT 923.100 71.400 924.900 77.400 ;
        RECT 926.100 71.400 927.900 78.000 ;
        RECT 923.100 71.100 924.600 71.400 ;
        RECT 918.000 70.200 924.600 71.100 ;
        RECT 877.950 63.450 880.050 64.200 ;
        RECT 883.950 63.450 886.050 64.050 ;
        RECT 877.950 62.550 886.050 63.450 ;
        RECT 877.950 62.100 880.050 62.550 ;
        RECT 883.950 61.950 886.050 62.550 ;
        RECT 881.100 58.050 882.900 59.850 ;
        RECT 896.400 58.050 897.300 65.400 ;
        RECT 901.950 63.450 904.050 64.050 ;
        RECT 910.950 63.450 913.050 64.050 ;
        RECT 901.950 62.550 913.050 63.450 ;
        RECT 901.950 61.950 904.050 62.550 ;
        RECT 910.950 61.950 913.050 62.550 ;
        RECT 901.950 58.050 903.750 59.850 ;
        RECT 918.000 58.050 918.900 70.200 ;
        RECT 923.100 58.050 924.900 59.850 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 883.950 55.950 886.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 898.950 55.950 901.050 58.050 ;
        RECT 901.950 55.950 904.050 58.050 ;
        RECT 904.950 55.950 907.050 58.050 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 919.950 55.950 922.050 58.050 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 865.950 52.800 868.050 54.900 ;
        RECT 876.000 52.200 876.900 55.950 ;
        RECT 878.100 54.150 879.900 55.950 ;
        RECT 884.100 54.150 885.900 55.950 ;
        RECT 852.000 51.000 855.300 52.200 ;
        RECT 827.700 48.600 828.900 50.700 ;
        RECT 807.000 42.000 808.800 48.600 ;
        RECT 811.500 47.400 816.600 48.600 ;
        RECT 811.500 42.600 813.300 47.400 ;
        RECT 814.500 42.000 816.300 45.600 ;
        RECT 827.100 42.600 828.900 48.600 ;
        RECT 830.100 47.700 837.900 49.050 ;
        RECT 830.100 42.600 831.900 47.700 ;
        RECT 833.100 42.000 834.900 46.800 ;
        RECT 836.100 42.600 837.900 47.700 ;
        RECT 853.500 42.600 855.300 51.000 ;
        RECT 860.100 42.000 861.900 51.600 ;
        RECT 876.000 51.000 879.300 52.200 ;
        RECT 877.500 42.600 879.300 51.000 ;
        RECT 884.100 42.000 885.900 51.600 ;
        RECT 896.400 48.600 897.300 55.950 ;
        RECT 898.950 54.150 900.750 55.950 ;
        RECT 905.100 54.150 906.900 55.950 ;
        RECT 918.000 52.200 918.900 55.950 ;
        RECT 920.100 54.150 921.900 55.950 ;
        RECT 926.100 54.150 927.900 55.950 ;
        RECT 918.000 51.000 921.300 52.200 ;
        RECT 896.400 47.400 901.500 48.600 ;
        RECT 896.700 42.000 898.500 45.600 ;
        RECT 899.700 42.600 901.500 47.400 ;
        RECT 904.200 42.000 906.000 48.600 ;
        RECT 919.500 42.600 921.300 51.000 ;
        RECT 926.100 42.000 927.900 51.600 ;
        RECT 14.100 29.400 15.900 39.000 ;
        RECT 20.700 30.000 22.500 38.400 ;
        RECT 36.000 32.400 37.800 39.000 ;
        RECT 40.500 33.600 42.300 38.400 ;
        RECT 43.500 35.400 45.300 39.000 ;
        RECT 40.500 32.400 45.600 33.600 ;
        RECT 37.950 30.450 40.050 31.050 ;
        RECT 20.700 28.800 24.000 30.000 ;
        RECT 14.100 25.050 15.900 26.850 ;
        RECT 20.100 25.050 21.900 26.850 ;
        RECT 23.100 25.050 24.000 28.800 ;
        RECT 29.550 29.550 40.050 30.450 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 22.950 22.950 25.050 25.050 ;
        RECT 17.100 21.150 18.900 22.950 ;
        RECT 23.100 10.800 24.000 22.950 ;
        RECT 29.550 22.050 30.450 29.550 ;
        RECT 37.950 28.950 40.050 29.550 ;
        RECT 35.100 25.050 36.900 26.850 ;
        RECT 41.250 25.050 43.050 26.850 ;
        RECT 44.700 25.050 45.600 32.400 ;
        RECT 61.500 30.000 63.300 38.400 ;
        RECT 60.000 28.800 63.300 30.000 ;
        RECT 68.100 29.400 69.900 39.000 ;
        RECT 84.000 32.400 85.800 39.000 ;
        RECT 88.500 33.600 90.300 38.400 ;
        RECT 91.500 35.400 93.300 39.000 ;
        RECT 88.500 32.400 93.600 33.600 ;
        RECT 104.100 32.400 105.900 38.400 ;
        RECT 73.950 30.450 76.050 31.050 ;
        RECT 85.950 30.450 88.050 31.050 ;
        RECT 73.950 29.550 88.050 30.450 ;
        RECT 73.950 28.950 76.050 29.550 ;
        RECT 85.950 28.950 88.050 29.550 ;
        RECT 60.000 25.050 60.900 28.800 ;
        RECT 62.100 25.050 63.900 26.850 ;
        RECT 68.100 25.050 69.900 26.850 ;
        RECT 83.100 25.050 84.900 26.850 ;
        RECT 89.250 25.050 91.050 26.850 ;
        RECT 92.700 25.050 93.600 32.400 ;
        RECT 104.700 30.300 105.900 32.400 ;
        RECT 107.100 33.300 108.900 38.400 ;
        RECT 110.100 34.200 111.900 39.000 ;
        RECT 113.100 33.300 114.900 38.400 ;
        RECT 128.100 35.400 129.900 39.000 ;
        RECT 131.100 35.400 132.900 38.400 ;
        RECT 107.100 31.950 114.900 33.300 ;
        RECT 104.700 29.400 108.300 30.300 ;
        RECT 104.100 25.050 105.900 26.850 ;
        RECT 107.100 25.050 108.300 29.400 ;
        RECT 110.100 25.050 111.900 26.850 ;
        RECT 131.100 25.050 132.300 35.400 ;
        RECT 145.500 30.000 147.300 38.400 ;
        RECT 144.000 28.800 147.300 30.000 ;
        RECT 152.100 29.400 153.900 39.000 ;
        RECT 165.000 32.400 166.800 39.000 ;
        RECT 169.500 33.600 171.300 38.400 ;
        RECT 172.500 35.400 174.300 39.000 ;
        RECT 169.500 32.400 174.600 33.600 ;
        RECT 157.950 30.450 160.050 31.050 ;
        RECT 169.950 30.450 172.050 31.050 ;
        RECT 157.950 29.550 172.050 30.450 ;
        RECT 157.950 28.950 160.050 29.550 ;
        RECT 169.950 28.950 172.050 29.550 ;
        RECT 144.000 25.050 144.900 28.800 ;
        RECT 146.100 25.050 147.900 26.850 ;
        RECT 152.100 25.050 153.900 26.850 ;
        RECT 164.100 25.050 165.900 26.850 ;
        RECT 170.250 25.050 172.050 26.850 ;
        RECT 173.700 25.050 174.600 32.400 ;
        RECT 188.100 29.400 189.900 39.000 ;
        RECT 194.700 30.000 196.500 38.400 ;
        RECT 210.000 32.400 211.800 39.000 ;
        RECT 214.500 33.600 216.300 38.400 ;
        RECT 217.500 35.400 219.300 39.000 ;
        RECT 214.500 32.400 219.600 33.600 ;
        RECT 234.000 32.400 235.800 39.000 ;
        RECT 238.500 33.600 240.300 38.400 ;
        RECT 241.500 35.400 243.300 39.000 ;
        RECT 254.100 35.400 255.900 38.400 ;
        RECT 257.100 35.400 258.900 39.000 ;
        RECT 238.500 32.400 243.600 33.600 ;
        RECT 194.700 28.800 198.000 30.000 ;
        RECT 175.950 27.450 178.050 28.050 ;
        RECT 175.950 26.550 183.450 27.450 ;
        RECT 175.950 25.950 178.050 26.550 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 40.950 22.950 43.050 25.050 ;
        RECT 43.950 22.950 46.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 25.950 20.550 30.450 22.050 ;
        RECT 38.250 21.150 40.050 22.950 ;
        RECT 25.950 19.950 30.000 20.550 ;
        RECT 28.950 18.450 31.050 18.900 ;
        RECT 40.950 18.450 43.050 19.050 ;
        RECT 28.950 17.550 43.050 18.450 ;
        RECT 28.950 16.800 31.050 17.550 ;
        RECT 40.950 16.950 43.050 17.550 ;
        RECT 44.700 15.600 45.600 22.950 ;
        RECT 17.400 9.900 24.000 10.800 ;
        RECT 17.400 9.600 18.900 9.900 ;
        RECT 14.100 3.000 15.900 9.600 ;
        RECT 17.100 3.600 18.900 9.600 ;
        RECT 23.100 9.600 24.000 9.900 ;
        RECT 35.100 14.700 42.900 15.600 ;
        RECT 20.100 3.000 21.900 9.000 ;
        RECT 23.100 3.600 24.900 9.600 ;
        RECT 35.100 3.600 36.900 14.700 ;
        RECT 38.100 3.000 39.900 13.800 ;
        RECT 41.100 3.600 42.900 14.700 ;
        RECT 44.100 3.600 45.900 15.600 ;
        RECT 60.000 10.800 60.900 22.950 ;
        RECT 65.100 21.150 66.900 22.950 ;
        RECT 86.250 21.150 88.050 22.950 ;
        RECT 61.950 18.450 64.050 19.050 ;
        RECT 73.950 18.450 76.050 19.050 ;
        RECT 61.950 17.550 76.050 18.450 ;
        RECT 61.950 16.950 64.050 17.550 ;
        RECT 73.950 16.950 76.050 17.550 ;
        RECT 92.700 15.600 93.600 22.950 ;
        RECT 107.100 15.600 108.300 22.950 ;
        RECT 113.100 21.150 114.900 22.950 ;
        RECT 128.100 21.150 129.900 22.950 ;
        RECT 83.100 14.700 90.900 15.600 ;
        RECT 60.000 9.900 66.600 10.800 ;
        RECT 60.000 9.600 60.900 9.900 ;
        RECT 59.100 3.600 60.900 9.600 ;
        RECT 65.100 9.600 66.600 9.900 ;
        RECT 62.100 3.000 63.900 9.000 ;
        RECT 65.100 3.600 66.900 9.600 ;
        RECT 68.100 3.000 69.900 9.600 ;
        RECT 83.100 3.600 84.900 14.700 ;
        RECT 86.100 3.000 87.900 13.800 ;
        RECT 89.100 3.600 90.900 14.700 ;
        RECT 92.100 3.600 93.900 15.600 ;
        RECT 107.100 14.100 109.500 15.600 ;
        RECT 105.000 11.100 106.800 12.900 ;
        RECT 104.700 3.000 106.500 9.600 ;
        RECT 107.700 3.600 109.500 14.100 ;
        RECT 112.800 3.000 114.600 15.600 ;
        RECT 131.100 9.600 132.300 22.950 ;
        RECT 144.000 10.800 144.900 22.950 ;
        RECT 149.100 21.150 150.900 22.950 ;
        RECT 167.250 21.150 169.050 22.950 ;
        RECT 145.950 18.450 148.050 19.050 ;
        RECT 157.950 18.450 160.050 19.050 ;
        RECT 145.950 17.550 160.050 18.450 ;
        RECT 145.950 16.950 148.050 17.550 ;
        RECT 157.950 16.950 160.050 17.550 ;
        RECT 173.700 15.600 174.600 22.950 ;
        RECT 182.550 22.050 183.450 26.550 ;
        RECT 188.100 25.050 189.900 26.850 ;
        RECT 194.100 25.050 195.900 26.850 ;
        RECT 197.100 25.050 198.000 28.800 ;
        RECT 209.100 25.050 210.900 26.850 ;
        RECT 215.250 25.050 217.050 26.850 ;
        RECT 218.700 25.050 219.600 32.400 ;
        RECT 223.950 27.450 226.050 28.050 ;
        RECT 229.950 27.450 232.050 28.050 ;
        RECT 223.950 26.550 232.050 27.450 ;
        RECT 223.950 25.950 226.050 26.550 ;
        RECT 229.950 25.950 232.050 26.550 ;
        RECT 233.100 25.050 234.900 26.850 ;
        RECT 239.250 25.050 241.050 26.850 ;
        RECT 242.700 25.050 243.600 32.400 ;
        RECT 254.700 25.050 255.900 35.400 ;
        RECT 272.100 32.400 273.900 38.400 ;
        RECT 259.950 27.450 262.050 31.050 ;
        RECT 272.700 30.300 273.900 32.400 ;
        RECT 275.100 33.300 276.900 38.400 ;
        RECT 278.100 34.200 279.900 39.000 ;
        RECT 281.100 33.300 282.900 38.400 ;
        RECT 296.700 35.400 298.500 39.000 ;
        RECT 299.700 33.600 301.500 38.400 ;
        RECT 275.100 31.950 282.900 33.300 ;
        RECT 296.400 32.400 301.500 33.600 ;
        RECT 304.200 32.400 306.000 39.000 ;
        RECT 272.700 29.400 276.300 30.300 ;
        RECT 259.950 27.000 267.450 27.450 ;
        RECT 260.550 26.550 267.450 27.000 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 182.550 20.550 187.050 22.050 ;
        RECT 191.100 21.150 192.900 22.950 ;
        RECT 183.000 19.950 187.050 20.550 ;
        RECT 164.100 14.700 171.900 15.600 ;
        RECT 144.000 9.900 150.600 10.800 ;
        RECT 144.000 9.600 144.900 9.900 ;
        RECT 128.100 3.000 129.900 9.600 ;
        RECT 131.100 3.600 132.900 9.600 ;
        RECT 143.100 3.600 144.900 9.600 ;
        RECT 149.100 9.600 150.600 9.900 ;
        RECT 146.100 3.000 147.900 9.000 ;
        RECT 149.100 3.600 150.900 9.600 ;
        RECT 152.100 3.000 153.900 9.600 ;
        RECT 164.100 3.600 165.900 14.700 ;
        RECT 167.100 3.000 168.900 13.800 ;
        RECT 170.100 3.600 171.900 14.700 ;
        RECT 173.100 3.600 174.900 15.600 ;
        RECT 197.100 10.800 198.000 22.950 ;
        RECT 202.950 22.050 205.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 202.950 21.000 208.050 22.050 ;
        RECT 212.250 21.150 214.050 22.950 ;
        RECT 203.550 20.550 208.050 21.000 ;
        RECT 204.000 19.950 208.050 20.550 ;
        RECT 202.950 18.450 205.050 19.050 ;
        RECT 211.950 18.450 214.050 19.050 ;
        RECT 202.950 17.550 214.050 18.450 ;
        RECT 202.950 16.950 205.050 17.550 ;
        RECT 211.950 16.950 214.050 17.550 ;
        RECT 218.700 15.600 219.600 22.950 ;
        RECT 236.250 21.150 238.050 22.950 ;
        RECT 226.950 18.450 229.050 19.050 ;
        RECT 238.950 18.450 241.050 19.050 ;
        RECT 226.950 17.550 241.050 18.450 ;
        RECT 226.950 16.950 229.050 17.550 ;
        RECT 238.950 16.950 241.050 17.550 ;
        RECT 242.700 15.600 243.600 22.950 ;
        RECT 191.400 9.900 198.000 10.800 ;
        RECT 191.400 9.600 192.900 9.900 ;
        RECT 188.100 3.000 189.900 9.600 ;
        RECT 191.100 3.600 192.900 9.600 ;
        RECT 197.100 9.600 198.000 9.900 ;
        RECT 209.100 14.700 216.900 15.600 ;
        RECT 194.100 3.000 195.900 9.000 ;
        RECT 197.100 3.600 198.900 9.600 ;
        RECT 209.100 3.600 210.900 14.700 ;
        RECT 212.100 3.000 213.900 13.800 ;
        RECT 215.100 3.600 216.900 14.700 ;
        RECT 218.100 3.600 219.900 15.600 ;
        RECT 233.100 14.700 240.900 15.600 ;
        RECT 220.950 6.450 223.050 7.050 ;
        RECT 226.950 6.450 229.050 7.050 ;
        RECT 220.950 5.550 229.050 6.450 ;
        RECT 220.950 4.950 223.050 5.550 ;
        RECT 226.950 4.950 229.050 5.550 ;
        RECT 233.100 3.600 234.900 14.700 ;
        RECT 236.100 3.000 237.900 13.800 ;
        RECT 239.100 3.600 240.900 14.700 ;
        RECT 242.100 3.600 243.900 15.600 ;
        RECT 254.700 9.600 255.900 22.950 ;
        RECT 257.100 21.150 258.900 22.950 ;
        RECT 266.550 22.050 267.450 26.550 ;
        RECT 272.100 25.050 273.900 26.850 ;
        RECT 275.100 25.050 276.300 29.400 ;
        RECT 278.100 25.050 279.900 26.850 ;
        RECT 296.400 25.050 297.300 32.400 ;
        RECT 317.100 29.400 318.900 39.000 ;
        RECT 323.700 30.000 325.500 38.400 ;
        RECT 340.500 30.000 342.300 38.400 ;
        RECT 323.700 28.800 327.000 30.000 ;
        RECT 307.950 27.450 312.000 28.050 ;
        RECT 298.950 25.050 300.750 26.850 ;
        RECT 305.100 25.050 306.900 26.850 ;
        RECT 307.950 25.950 312.450 27.450 ;
        RECT 271.950 22.950 274.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 266.550 20.550 271.050 22.050 ;
        RECT 267.000 19.950 271.050 20.550 ;
        RECT 275.100 15.600 276.300 22.950 ;
        RECT 281.100 21.150 282.900 22.950 ;
        RECT 277.950 18.450 280.050 18.750 ;
        RECT 289.950 18.450 292.050 19.050 ;
        RECT 277.950 17.550 292.050 18.450 ;
        RECT 277.950 16.650 280.050 17.550 ;
        RECT 289.950 16.950 292.050 17.550 ;
        RECT 296.400 15.600 297.300 22.950 ;
        RECT 301.950 21.150 303.750 22.950 ;
        RECT 311.550 22.050 312.450 25.950 ;
        RECT 317.100 25.050 318.900 26.850 ;
        RECT 323.100 25.050 324.900 26.850 ;
        RECT 326.100 25.050 327.000 28.800 ;
        RECT 339.000 28.800 342.300 30.000 ;
        RECT 347.100 29.400 348.900 39.000 ;
        RECT 362.100 33.300 363.900 38.400 ;
        RECT 365.100 34.200 366.900 39.000 ;
        RECT 368.100 33.300 369.900 38.400 ;
        RECT 362.100 31.950 369.900 33.300 ;
        RECT 371.100 32.400 372.900 38.400 ;
        RECT 386.700 35.400 388.500 39.000 ;
        RECT 389.700 33.600 391.500 38.400 ;
        RECT 386.400 32.400 391.500 33.600 ;
        RECT 394.200 32.400 396.000 39.000 ;
        RECT 371.100 30.300 372.300 32.400 ;
        RECT 368.700 29.400 372.300 30.300 ;
        RECT 333.000 27.450 337.050 28.050 ;
        RECT 332.550 25.950 337.050 27.450 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 311.550 20.550 316.050 22.050 ;
        RECT 320.100 21.150 321.900 22.950 ;
        RECT 312.000 19.950 316.050 20.550 ;
        RECT 298.950 18.450 301.050 19.050 ;
        RECT 322.950 18.450 325.050 19.050 ;
        RECT 298.950 17.550 325.050 18.450 ;
        RECT 298.950 16.950 301.050 17.550 ;
        RECT 322.950 16.950 325.050 17.550 ;
        RECT 275.100 14.100 277.500 15.600 ;
        RECT 273.000 11.100 274.800 12.900 ;
        RECT 254.100 3.600 255.900 9.600 ;
        RECT 257.100 3.000 258.900 9.600 ;
        RECT 272.700 3.000 274.500 9.600 ;
        RECT 275.700 3.600 277.500 14.100 ;
        RECT 280.800 3.000 282.600 15.600 ;
        RECT 296.100 3.600 297.900 15.600 ;
        RECT 299.100 14.700 306.900 15.600 ;
        RECT 299.100 3.600 300.900 14.700 ;
        RECT 302.100 3.000 303.900 13.800 ;
        RECT 305.100 3.600 306.900 14.700 ;
        RECT 326.100 10.800 327.000 22.950 ;
        RECT 332.550 22.050 333.450 25.950 ;
        RECT 339.000 25.050 339.900 28.800 ;
        RECT 341.100 25.050 342.900 26.850 ;
        RECT 347.100 25.050 348.900 26.850 ;
        RECT 365.100 25.050 366.900 26.850 ;
        RECT 368.700 25.050 369.900 29.400 ;
        RECT 371.100 25.050 372.900 26.850 ;
        RECT 386.400 25.050 387.300 32.400 ;
        RECT 410.100 29.400 411.900 39.000 ;
        RECT 416.700 30.000 418.500 38.400 ;
        RECT 436.500 30.000 438.300 38.400 ;
        RECT 416.700 28.800 420.000 30.000 ;
        RECT 388.950 25.050 390.750 26.850 ;
        RECT 395.100 25.050 396.900 26.850 ;
        RECT 410.100 25.050 411.900 26.850 ;
        RECT 416.100 25.050 417.900 26.850 ;
        RECT 419.100 25.050 420.000 28.800 ;
        RECT 435.000 28.800 438.300 30.000 ;
        RECT 443.100 29.400 444.900 39.000 ;
        RECT 456.000 32.400 457.800 39.000 ;
        RECT 460.500 33.600 462.300 38.400 ;
        RECT 463.500 35.400 465.300 39.000 ;
        RECT 479.700 35.400 481.500 39.000 ;
        RECT 460.500 32.400 465.600 33.600 ;
        RECT 435.000 25.050 435.900 28.800 ;
        RECT 437.100 25.050 438.900 26.850 ;
        RECT 443.100 25.050 444.900 26.850 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 461.250 25.050 463.050 26.850 ;
        RECT 464.700 25.050 465.600 32.400 ;
        RECT 466.950 33.450 469.050 33.900 ;
        RECT 475.950 33.450 478.050 34.050 ;
        RECT 482.700 33.600 484.500 38.400 ;
        RECT 466.950 32.550 478.050 33.450 ;
        RECT 466.950 31.800 469.050 32.550 ;
        RECT 475.950 31.950 478.050 32.550 ;
        RECT 479.400 32.400 484.500 33.600 ;
        RECT 487.200 32.400 489.000 39.000 ;
        RECT 479.400 25.050 480.300 32.400 ;
        RECT 503.100 29.400 504.900 39.000 ;
        RECT 509.700 30.000 511.500 38.400 ;
        RECT 529.500 30.000 531.300 38.400 ;
        RECT 509.700 28.800 513.000 30.000 ;
        RECT 481.950 25.050 483.750 26.850 ;
        RECT 488.100 25.050 489.900 26.850 ;
        RECT 503.100 25.050 504.900 26.850 ;
        RECT 509.100 25.050 510.900 26.850 ;
        RECT 512.100 25.050 513.000 28.800 ;
        RECT 528.000 28.800 531.300 30.000 ;
        RECT 536.100 29.400 537.900 39.000 ;
        RECT 550.500 30.000 552.300 38.400 ;
        RECT 549.000 28.800 552.300 30.000 ;
        RECT 557.100 29.400 558.900 39.000 ;
        RECT 572.100 32.400 573.900 38.400 ;
        RECT 572.700 30.300 573.900 32.400 ;
        RECT 575.100 33.300 576.900 38.400 ;
        RECT 578.100 34.200 579.900 39.000 ;
        RECT 581.100 33.300 582.900 38.400 ;
        RECT 575.100 31.950 582.900 33.300 ;
        RECT 596.100 32.400 597.900 38.400 ;
        RECT 596.700 30.300 597.900 32.400 ;
        RECT 599.100 33.300 600.900 38.400 ;
        RECT 602.100 34.200 603.900 39.000 ;
        RECT 605.100 33.300 606.900 38.400 ;
        RECT 599.100 31.950 606.900 33.300 ;
        RECT 620.100 32.400 621.900 38.400 ;
        RECT 610.950 30.450 613.050 31.050 ;
        RECT 616.950 30.450 619.050 31.050 ;
        RECT 572.700 29.400 576.300 30.300 ;
        RECT 596.700 29.400 600.300 30.300 ;
        RECT 528.000 25.050 528.900 28.800 ;
        RECT 530.100 25.050 531.900 26.850 ;
        RECT 536.100 25.050 537.900 26.850 ;
        RECT 549.000 25.050 549.900 28.800 ;
        RECT 551.100 25.050 552.900 26.850 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 572.100 25.050 573.900 26.850 ;
        RECT 575.100 25.050 576.300 29.400 ;
        RECT 578.100 25.050 579.900 26.850 ;
        RECT 596.100 25.050 597.900 26.850 ;
        RECT 599.100 25.050 600.300 29.400 ;
        RECT 610.950 29.550 619.050 30.450 ;
        RECT 610.950 28.950 613.050 29.550 ;
        RECT 616.950 28.950 619.050 29.550 ;
        RECT 620.700 30.300 621.900 32.400 ;
        RECT 623.100 33.300 624.900 38.400 ;
        RECT 626.100 34.200 627.900 39.000 ;
        RECT 629.100 33.300 630.900 38.400 ;
        RECT 623.100 31.950 630.900 33.300 ;
        RECT 645.000 32.400 646.800 39.000 ;
        RECT 649.500 33.600 651.300 38.400 ;
        RECT 652.500 35.400 654.300 39.000 ;
        RECT 649.500 32.400 654.600 33.600 ;
        RECT 631.950 30.450 634.050 31.050 ;
        RECT 649.950 30.450 652.050 31.050 ;
        RECT 620.700 29.400 624.300 30.300 ;
        RECT 607.950 27.450 610.050 28.050 ;
        RECT 613.950 27.450 616.050 28.050 ;
        RECT 602.100 25.050 603.900 26.850 ;
        RECT 607.950 26.550 616.050 27.450 ;
        RECT 607.950 25.950 610.050 26.550 ;
        RECT 613.950 25.950 616.050 26.550 ;
        RECT 620.100 25.050 621.900 26.850 ;
        RECT 623.100 25.050 624.300 29.400 ;
        RECT 631.950 29.550 652.050 30.450 ;
        RECT 631.950 28.950 634.050 29.550 ;
        RECT 649.950 28.950 652.050 29.550 ;
        RECT 626.100 25.050 627.900 26.850 ;
        RECT 644.100 25.050 645.900 26.850 ;
        RECT 650.250 25.050 652.050 26.850 ;
        RECT 653.700 25.050 654.600 32.400 ;
        RECT 665.700 31.200 667.500 38.400 ;
        RECT 670.800 32.400 672.600 39.000 ;
        RECT 686.100 32.400 687.900 38.400 ;
        RECT 665.700 30.300 669.900 31.200 ;
        RECT 665.100 25.050 666.900 26.850 ;
        RECT 668.700 25.050 669.900 30.300 ;
        RECT 686.700 30.300 687.900 32.400 ;
        RECT 689.100 33.300 690.900 38.400 ;
        RECT 692.100 34.200 693.900 39.000 ;
        RECT 695.100 33.300 696.900 38.400 ;
        RECT 689.100 31.950 696.900 33.300 ;
        RECT 707.100 33.300 708.900 38.400 ;
        RECT 710.100 34.200 711.900 39.000 ;
        RECT 713.100 33.300 714.900 38.400 ;
        RECT 707.100 31.950 714.900 33.300 ;
        RECT 716.100 32.400 717.900 38.400 ;
        RECT 716.100 30.300 717.300 32.400 ;
        RECT 686.700 29.400 690.300 30.300 ;
        RECT 670.950 25.050 672.750 26.850 ;
        RECT 686.100 25.050 687.900 26.850 ;
        RECT 689.100 25.050 690.300 29.400 ;
        RECT 713.700 29.400 717.300 30.300 ;
        RECT 733.500 30.000 735.300 38.400 ;
        RECT 692.100 25.050 693.900 26.850 ;
        RECT 710.100 25.050 711.900 26.850 ;
        RECT 713.700 25.050 714.900 29.400 ;
        RECT 732.000 28.800 735.300 30.000 ;
        RECT 740.100 29.400 741.900 39.000 ;
        RECT 752.100 29.400 753.900 39.000 ;
        RECT 758.700 30.000 760.500 38.400 ;
        RECT 774.000 32.400 775.800 39.000 ;
        RECT 778.500 33.600 780.300 38.400 ;
        RECT 781.500 35.400 783.300 39.000 ;
        RECT 778.500 32.400 783.600 33.600 ;
        RECT 798.000 32.400 799.800 39.000 ;
        RECT 802.500 33.600 804.300 38.400 ;
        RECT 805.500 35.400 807.300 39.000 ;
        RECT 802.500 32.400 807.600 33.600 ;
        RECT 758.700 28.800 762.000 30.000 ;
        RECT 716.100 25.050 717.900 26.850 ;
        RECT 732.000 25.050 732.900 28.800 ;
        RECT 734.100 25.050 735.900 26.850 ;
        RECT 740.100 25.050 741.900 26.850 ;
        RECT 752.100 25.050 753.900 26.850 ;
        RECT 758.100 25.050 759.900 26.850 ;
        RECT 761.100 25.050 762.000 28.800 ;
        RECT 773.100 25.050 774.900 26.850 ;
        RECT 779.250 25.050 781.050 26.850 ;
        RECT 782.700 25.050 783.600 32.400 ;
        RECT 797.100 25.050 798.900 26.850 ;
        RECT 803.250 25.050 805.050 26.850 ;
        RECT 806.700 25.050 807.600 32.400 ;
        RECT 821.100 29.400 822.900 39.000 ;
        RECT 827.700 30.000 829.500 38.400 ;
        RECT 845.100 35.400 846.900 38.400 ;
        RECT 848.100 35.400 849.900 39.000 ;
        RECT 827.700 28.800 831.000 30.000 ;
        RECT 821.100 25.050 822.900 26.850 ;
        RECT 827.100 25.050 828.900 26.850 ;
        RECT 830.100 25.050 831.000 28.800 ;
        RECT 845.700 25.050 846.900 35.400 ;
        RECT 863.100 33.300 864.900 38.400 ;
        RECT 866.100 34.200 867.900 39.000 ;
        RECT 869.100 33.300 870.900 38.400 ;
        RECT 863.100 31.950 870.900 33.300 ;
        RECT 872.100 32.400 873.900 38.400 ;
        RECT 887.100 33.300 888.900 38.400 ;
        RECT 890.100 34.200 891.900 39.000 ;
        RECT 893.100 33.300 894.900 38.400 ;
        RECT 872.100 30.300 873.300 32.400 ;
        RECT 887.100 31.950 894.900 33.300 ;
        RECT 896.100 32.400 897.900 38.400 ;
        RECT 912.000 32.400 913.800 39.000 ;
        RECT 916.500 33.600 918.300 38.400 ;
        RECT 919.500 35.400 921.300 39.000 ;
        RECT 932.100 35.400 933.900 38.400 ;
        RECT 935.100 35.400 936.900 39.000 ;
        RECT 916.500 32.400 921.600 33.600 ;
        RECT 896.100 30.300 897.300 32.400 ;
        RECT 869.700 29.400 873.300 30.300 ;
        RECT 893.700 29.400 897.300 30.300 ;
        RECT 866.100 25.050 867.900 26.850 ;
        RECT 869.700 25.050 870.900 29.400 ;
        RECT 872.100 25.050 873.900 26.850 ;
        RECT 890.100 25.050 891.900 26.850 ;
        RECT 893.700 25.050 894.900 29.400 ;
        RECT 896.100 25.050 897.900 26.850 ;
        RECT 911.100 25.050 912.900 26.850 ;
        RECT 917.250 25.050 919.050 26.850 ;
        RECT 920.700 25.050 921.600 32.400 ;
        RECT 932.700 25.050 933.900 35.400 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 370.950 22.950 373.050 25.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 394.950 22.950 397.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 415.950 22.950 418.050 25.050 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 715.950 22.950 718.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 778.950 22.950 781.050 25.050 ;
        RECT 781.950 22.950 784.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 829.950 22.950 832.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 868.950 22.950 871.050 25.050 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 895.950 22.950 898.050 25.050 ;
        RECT 910.950 22.950 913.050 25.050 ;
        RECT 913.950 22.950 916.050 25.050 ;
        RECT 916.950 22.950 919.050 25.050 ;
        RECT 919.950 22.950 922.050 25.050 ;
        RECT 931.950 22.950 934.050 25.050 ;
        RECT 934.950 22.950 937.050 25.050 ;
        RECT 328.950 20.550 333.450 22.050 ;
        RECT 328.950 19.950 333.000 20.550 ;
        RECT 320.400 9.900 327.000 10.800 ;
        RECT 320.400 9.600 321.900 9.900 ;
        RECT 317.100 3.000 318.900 9.600 ;
        RECT 320.100 3.600 321.900 9.600 ;
        RECT 326.100 9.600 327.000 9.900 ;
        RECT 339.000 10.800 339.900 22.950 ;
        RECT 344.100 21.150 345.900 22.950 ;
        RECT 362.100 21.150 363.900 22.950 ;
        RECT 346.950 18.450 349.050 19.050 ;
        RECT 355.950 18.450 358.050 19.050 ;
        RECT 364.950 18.450 367.050 18.750 ;
        RECT 346.950 17.550 367.050 18.450 ;
        RECT 346.950 16.950 349.050 17.550 ;
        RECT 355.950 16.950 358.050 17.550 ;
        RECT 364.950 16.650 367.050 17.550 ;
        RECT 368.700 15.600 369.900 22.950 ;
        RECT 339.000 9.900 345.600 10.800 ;
        RECT 339.000 9.600 339.900 9.900 ;
        RECT 323.100 3.000 324.900 9.000 ;
        RECT 326.100 3.600 327.900 9.600 ;
        RECT 338.100 3.600 339.900 9.600 ;
        RECT 344.100 9.600 345.600 9.900 ;
        RECT 341.100 3.000 342.900 9.000 ;
        RECT 344.100 3.600 345.900 9.600 ;
        RECT 347.100 3.000 348.900 9.600 ;
        RECT 349.950 9.450 352.050 10.050 ;
        RECT 355.950 9.450 358.050 10.050 ;
        RECT 349.950 8.550 358.050 9.450 ;
        RECT 349.950 7.950 352.050 8.550 ;
        RECT 355.950 7.950 358.050 8.550 ;
        RECT 362.400 3.000 364.200 15.600 ;
        RECT 367.500 14.100 369.900 15.600 ;
        RECT 370.950 15.450 373.050 16.050 ;
        RECT 379.950 15.450 382.050 16.050 ;
        RECT 386.400 15.600 387.300 22.950 ;
        RECT 391.950 21.150 393.750 22.950 ;
        RECT 413.100 21.150 414.900 22.950 ;
        RECT 370.950 14.550 382.050 15.450 ;
        RECT 367.500 3.600 369.300 14.100 ;
        RECT 370.950 13.950 373.050 14.550 ;
        RECT 379.950 13.950 382.050 14.550 ;
        RECT 370.200 11.100 372.000 12.900 ;
        RECT 370.500 3.000 372.300 9.600 ;
        RECT 386.100 3.600 387.900 15.600 ;
        RECT 389.100 14.700 396.900 15.600 ;
        RECT 389.100 3.600 390.900 14.700 ;
        RECT 392.100 3.000 393.900 13.800 ;
        RECT 395.100 3.600 396.900 14.700 ;
        RECT 419.100 10.800 420.000 22.950 ;
        RECT 413.400 9.900 420.000 10.800 ;
        RECT 413.400 9.600 414.900 9.900 ;
        RECT 410.100 3.000 411.900 9.600 ;
        RECT 413.100 3.600 414.900 9.600 ;
        RECT 419.100 9.600 420.000 9.900 ;
        RECT 435.000 10.800 435.900 22.950 ;
        RECT 440.100 21.150 441.900 22.950 ;
        RECT 458.250 21.150 460.050 22.950 ;
        RECT 436.950 18.450 439.050 19.050 ;
        RECT 460.950 18.450 463.050 19.050 ;
        RECT 436.950 17.550 463.050 18.450 ;
        RECT 436.950 16.950 439.050 17.550 ;
        RECT 460.950 16.950 463.050 17.550 ;
        RECT 464.700 15.600 465.600 22.950 ;
        RECT 479.400 15.600 480.300 22.950 ;
        RECT 484.950 21.150 486.750 22.950 ;
        RECT 506.100 21.150 507.900 22.950 ;
        RECT 496.950 18.450 499.050 19.050 ;
        RECT 508.950 18.450 511.050 19.050 ;
        RECT 496.950 17.550 511.050 18.450 ;
        RECT 496.950 16.950 499.050 17.550 ;
        RECT 508.950 16.950 511.050 17.550 ;
        RECT 455.100 14.700 462.900 15.600 ;
        RECT 435.000 9.900 441.600 10.800 ;
        RECT 435.000 9.600 435.900 9.900 ;
        RECT 416.100 3.000 417.900 9.000 ;
        RECT 419.100 3.600 420.900 9.600 ;
        RECT 434.100 3.600 435.900 9.600 ;
        RECT 440.100 9.600 441.600 9.900 ;
        RECT 437.100 3.000 438.900 9.000 ;
        RECT 440.100 3.600 441.900 9.600 ;
        RECT 443.100 3.000 444.900 9.600 ;
        RECT 455.100 3.600 456.900 14.700 ;
        RECT 458.100 3.000 459.900 13.800 ;
        RECT 461.100 3.600 462.900 14.700 ;
        RECT 464.100 3.600 465.900 15.600 ;
        RECT 479.100 3.600 480.900 15.600 ;
        RECT 482.100 14.700 489.900 15.600 ;
        RECT 482.100 3.600 483.900 14.700 ;
        RECT 485.100 3.000 486.900 13.800 ;
        RECT 488.100 3.600 489.900 14.700 ;
        RECT 493.950 15.450 496.050 16.050 ;
        RECT 502.950 15.450 505.050 15.900 ;
        RECT 493.950 14.550 505.050 15.450 ;
        RECT 493.950 13.950 496.050 14.550 ;
        RECT 502.950 13.800 505.050 14.550 ;
        RECT 512.100 10.800 513.000 22.950 ;
        RECT 506.400 9.900 513.000 10.800 ;
        RECT 506.400 9.600 507.900 9.900 ;
        RECT 503.100 3.000 504.900 9.600 ;
        RECT 506.100 3.600 507.900 9.600 ;
        RECT 512.100 9.600 513.000 9.900 ;
        RECT 528.000 10.800 528.900 22.950 ;
        RECT 533.100 21.150 534.900 22.950 ;
        RECT 549.000 10.800 549.900 22.950 ;
        RECT 554.100 21.150 555.900 22.950 ;
        RECT 575.100 15.600 576.300 22.950 ;
        RECT 581.100 21.150 582.900 22.950 ;
        RECT 589.950 18.450 592.050 19.050 ;
        RECT 595.950 18.450 598.050 19.050 ;
        RECT 589.950 17.550 598.050 18.450 ;
        RECT 589.950 16.950 592.050 17.550 ;
        RECT 595.950 16.950 598.050 17.550 ;
        RECT 599.100 15.600 600.300 22.950 ;
        RECT 605.100 21.150 606.900 22.950 ;
        RECT 623.100 15.600 624.300 22.950 ;
        RECT 629.100 21.150 630.900 22.950 ;
        RECT 647.250 21.150 649.050 22.950 ;
        RECT 653.700 15.600 654.600 22.950 ;
        RECT 575.100 14.100 577.500 15.600 ;
        RECT 573.000 11.100 574.800 12.900 ;
        RECT 528.000 9.900 534.600 10.800 ;
        RECT 528.000 9.600 528.900 9.900 ;
        RECT 509.100 3.000 510.900 9.000 ;
        RECT 512.100 3.600 513.900 9.600 ;
        RECT 527.100 3.600 528.900 9.600 ;
        RECT 533.100 9.600 534.600 9.900 ;
        RECT 549.000 9.900 555.600 10.800 ;
        RECT 549.000 9.600 549.900 9.900 ;
        RECT 530.100 3.000 531.900 9.000 ;
        RECT 533.100 3.600 534.900 9.600 ;
        RECT 536.100 3.000 537.900 9.600 ;
        RECT 548.100 3.600 549.900 9.600 ;
        RECT 554.100 9.600 555.600 9.900 ;
        RECT 551.100 3.000 552.900 9.000 ;
        RECT 554.100 3.600 555.900 9.600 ;
        RECT 557.100 3.000 558.900 9.600 ;
        RECT 572.700 3.000 574.500 9.600 ;
        RECT 575.700 3.600 577.500 14.100 ;
        RECT 580.800 3.000 582.600 15.600 ;
        RECT 599.100 14.100 601.500 15.600 ;
        RECT 597.000 11.100 598.800 12.900 ;
        RECT 596.700 3.000 598.500 9.600 ;
        RECT 599.700 3.600 601.500 14.100 ;
        RECT 604.800 3.000 606.600 15.600 ;
        RECT 623.100 14.100 625.500 15.600 ;
        RECT 621.000 11.100 622.800 12.900 ;
        RECT 620.700 3.000 622.500 9.600 ;
        RECT 623.700 3.600 625.500 14.100 ;
        RECT 628.800 3.000 630.600 15.600 ;
        RECT 644.100 14.700 651.900 15.600 ;
        RECT 644.100 3.600 645.900 14.700 ;
        RECT 647.100 3.000 648.900 13.800 ;
        RECT 650.100 3.600 651.900 14.700 ;
        RECT 653.100 3.600 654.900 15.600 ;
        RECT 658.950 13.950 664.050 16.050 ;
        RECT 668.700 9.600 669.900 22.950 ;
        RECT 689.100 15.600 690.300 22.950 ;
        RECT 695.100 21.150 696.900 22.950 ;
        RECT 707.100 21.150 708.900 22.950 ;
        RECT 713.700 15.600 714.900 22.950 ;
        RECT 689.100 14.100 691.500 15.600 ;
        RECT 687.000 11.100 688.800 12.900 ;
        RECT 665.100 3.000 666.900 9.600 ;
        RECT 668.100 3.600 669.900 9.600 ;
        RECT 671.100 3.000 672.900 9.600 ;
        RECT 686.700 3.000 688.500 9.600 ;
        RECT 689.700 3.600 691.500 14.100 ;
        RECT 694.800 3.000 696.600 15.600 ;
        RECT 707.400 3.000 709.200 15.600 ;
        RECT 712.500 14.100 714.900 15.600 ;
        RECT 712.500 3.600 714.300 14.100 ;
        RECT 715.200 11.100 717.000 12.900 ;
        RECT 732.000 10.800 732.900 22.950 ;
        RECT 737.100 21.150 738.900 22.950 ;
        RECT 755.100 21.150 756.900 22.950 ;
        RECT 761.100 10.800 762.000 22.950 ;
        RECT 776.250 21.150 778.050 22.950 ;
        RECT 782.700 15.600 783.600 22.950 ;
        RECT 800.250 21.150 802.050 22.950 ;
        RECT 787.950 18.450 790.050 19.050 ;
        RECT 799.950 18.450 802.050 19.050 ;
        RECT 787.950 17.550 802.050 18.450 ;
        RECT 787.950 16.950 790.050 17.550 ;
        RECT 799.950 16.950 802.050 17.550 ;
        RECT 806.700 15.600 807.600 22.950 ;
        RECT 824.100 21.150 825.900 22.950 ;
        RECT 817.950 18.450 820.050 19.050 ;
        RECT 826.950 18.450 829.050 19.050 ;
        RECT 817.950 17.550 829.050 18.450 ;
        RECT 817.950 16.950 820.050 17.550 ;
        RECT 826.950 16.950 829.050 17.550 ;
        RECT 732.000 9.900 738.600 10.800 ;
        RECT 732.000 9.600 732.900 9.900 ;
        RECT 715.500 3.000 717.300 9.600 ;
        RECT 731.100 3.600 732.900 9.600 ;
        RECT 737.100 9.600 738.600 9.900 ;
        RECT 755.400 9.900 762.000 10.800 ;
        RECT 755.400 9.600 756.900 9.900 ;
        RECT 734.100 3.000 735.900 9.000 ;
        RECT 737.100 3.600 738.900 9.600 ;
        RECT 740.100 3.000 741.900 9.600 ;
        RECT 752.100 3.000 753.900 9.600 ;
        RECT 755.100 3.600 756.900 9.600 ;
        RECT 761.100 9.600 762.000 9.900 ;
        RECT 773.100 14.700 780.900 15.600 ;
        RECT 758.100 3.000 759.900 9.000 ;
        RECT 761.100 3.600 762.900 9.600 ;
        RECT 773.100 3.600 774.900 14.700 ;
        RECT 776.100 3.000 777.900 13.800 ;
        RECT 779.100 3.600 780.900 14.700 ;
        RECT 782.100 3.600 783.900 15.600 ;
        RECT 797.100 14.700 804.900 15.600 ;
        RECT 797.100 3.600 798.900 14.700 ;
        RECT 800.100 3.000 801.900 13.800 ;
        RECT 803.100 3.600 804.900 14.700 ;
        RECT 806.100 3.600 807.900 15.600 ;
        RECT 808.950 15.450 811.050 16.050 ;
        RECT 823.950 15.450 826.050 15.900 ;
        RECT 808.950 14.550 826.050 15.450 ;
        RECT 808.950 13.950 811.050 14.550 ;
        RECT 823.950 13.800 826.050 14.550 ;
        RECT 830.100 10.800 831.000 22.950 ;
        RECT 824.400 9.900 831.000 10.800 ;
        RECT 824.400 9.600 825.900 9.900 ;
        RECT 821.100 3.000 822.900 9.600 ;
        RECT 824.100 3.600 825.900 9.600 ;
        RECT 830.100 9.600 831.000 9.900 ;
        RECT 845.700 9.600 846.900 22.950 ;
        RECT 848.100 21.150 849.900 22.950 ;
        RECT 863.100 21.150 864.900 22.950 ;
        RECT 869.700 15.600 870.900 22.950 ;
        RECT 887.100 21.150 888.900 22.950 ;
        RECT 893.700 15.600 894.900 22.950 ;
        RECT 914.250 21.150 916.050 22.950 ;
        RECT 920.700 15.600 921.600 22.950 ;
        RECT 827.100 3.000 828.900 9.000 ;
        RECT 830.100 3.600 831.900 9.600 ;
        RECT 845.100 3.600 846.900 9.600 ;
        RECT 848.100 3.000 849.900 9.600 ;
        RECT 863.400 3.000 865.200 15.600 ;
        RECT 868.500 14.100 870.900 15.600 ;
        RECT 868.500 3.600 870.300 14.100 ;
        RECT 871.200 11.100 873.000 12.900 ;
        RECT 871.500 3.000 873.300 9.600 ;
        RECT 887.400 3.000 889.200 15.600 ;
        RECT 892.500 14.100 894.900 15.600 ;
        RECT 911.100 14.700 918.900 15.600 ;
        RECT 892.500 3.600 894.300 14.100 ;
        RECT 895.200 11.100 897.000 12.900 ;
        RECT 895.500 3.000 897.300 9.600 ;
        RECT 911.100 3.600 912.900 14.700 ;
        RECT 914.100 3.000 915.900 13.800 ;
        RECT 917.100 3.600 918.900 14.700 ;
        RECT 920.100 3.600 921.900 15.600 ;
        RECT 932.700 9.600 933.900 22.950 ;
        RECT 935.100 21.150 936.900 22.950 ;
        RECT 932.100 3.600 933.900 9.600 ;
        RECT 935.100 3.000 936.900 9.600 ;
      LAYER metal2 ;
        RECT 244.950 931.950 247.050 934.050 ;
        RECT 274.950 931.950 277.050 934.050 ;
        RECT 220.950 928.950 223.050 931.050 ;
        RECT 16.950 925.950 19.050 928.050 ;
        RECT 106.950 925.950 109.050 928.050 ;
        RECT 17.400 918.600 18.450 925.950 ;
        RECT 34.500 921.300 36.600 923.400 ;
        RECT 44.100 922.500 46.200 924.600 ;
        RECT 55.950 922.950 58.050 925.050 ;
        RECT 97.950 922.950 100.050 925.050 ;
        RECT 17.400 916.350 18.600 918.600 ;
        RECT 32.400 918.450 33.600 918.600 ;
        RECT 29.400 917.400 33.600 918.450 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 14.400 911.400 15.600 913.650 ;
        RECT 14.400 892.050 15.450 911.400 ;
        RECT 29.400 909.450 30.450 917.400 ;
        RECT 32.400 916.350 33.600 917.400 ;
        RECT 32.100 913.950 34.200 916.050 ;
        RECT 35.400 912.300 36.300 921.300 ;
        RECT 37.800 917.700 39.900 919.800 ;
        RECT 41.400 919.350 42.600 921.600 ;
        RECT 39.000 915.300 39.900 917.700 ;
        RECT 40.800 916.950 42.900 919.050 ;
        RECT 44.700 915.300 45.900 922.500 ;
        RECT 52.950 917.100 55.050 919.200 ;
        RECT 39.000 914.100 45.900 915.300 ;
        RECT 42.000 912.300 44.100 913.200 ;
        RECT 35.400 911.100 44.100 912.300 ;
        RECT 29.400 908.400 33.450 909.450 ;
        RECT 36.900 909.300 39.000 911.100 ;
        RECT 13.950 889.950 16.050 892.050 ;
        RECT 14.400 885.600 15.450 889.950 ;
        RECT 14.400 883.350 15.600 885.600 ;
        RECT 19.950 884.100 22.050 886.200 ;
        RECT 25.950 884.100 28.050 886.200 ;
        RECT 32.400 885.600 33.450 908.400 ;
        RECT 40.800 908.100 42.900 910.200 ;
        RECT 45.000 908.700 45.900 914.100 ;
        RECT 46.800 913.950 48.900 916.050 ;
        RECT 47.400 912.450 48.600 913.650 ;
        RECT 47.400 911.400 51.450 912.450 ;
        RECT 41.400 907.050 42.600 907.800 ;
        RECT 40.950 904.950 43.050 907.050 ;
        RECT 44.100 906.600 46.200 908.700 ;
        RECT 20.400 883.350 21.600 884.100 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 19.950 880.950 22.050 883.050 ;
        RECT 17.400 878.400 18.600 880.650 ;
        RECT 17.400 877.050 18.450 878.400 ;
        RECT 22.950 877.950 25.050 880.050 ;
        RECT 17.400 875.400 22.050 877.050 ;
        RECT 18.000 874.950 22.050 875.400 ;
        RECT 23.400 871.050 24.450 877.950 ;
        RECT 26.400 877.050 27.450 884.100 ;
        RECT 32.400 883.350 33.600 885.600 ;
        RECT 37.950 884.100 40.050 886.200 ;
        RECT 38.400 883.350 39.600 884.100 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 35.400 879.900 36.600 880.650 ;
        RECT 34.950 877.800 37.050 879.900 ;
        RECT 41.400 879.450 42.600 880.650 ;
        RECT 41.400 878.400 45.450 879.450 ;
        RECT 25.950 874.950 28.050 877.050 ;
        RECT 40.950 871.950 43.050 874.050 ;
        RECT 22.950 868.950 25.050 871.050 ;
        RECT 41.400 841.200 42.450 871.950 ;
        RECT 44.400 868.050 45.450 878.400 ;
        RECT 46.950 877.800 49.050 879.900 ;
        RECT 43.950 865.950 46.050 868.050 ;
        RECT 16.950 839.100 19.050 841.200 ;
        RECT 24.000 840.600 28.050 841.050 ;
        RECT 17.400 838.350 18.600 839.100 ;
        RECT 23.400 838.950 28.050 840.600 ;
        RECT 28.950 839.100 31.050 841.200 ;
        RECT 31.950 840.600 36.000 841.050 ;
        RECT 23.400 838.350 24.600 838.950 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 22.950 835.950 25.050 838.050 ;
        RECT 14.400 833.400 15.600 835.650 ;
        RECT 20.400 834.900 21.600 835.650 ;
        RECT 14.400 829.050 15.450 833.400 ;
        RECT 19.950 832.800 22.050 834.900 ;
        RECT 29.400 832.050 30.450 839.100 ;
        RECT 31.950 838.950 36.600 840.600 ;
        RECT 40.950 839.100 43.050 841.200 ;
        RECT 47.400 841.050 48.450 877.800 ;
        RECT 35.400 838.350 36.600 838.950 ;
        RECT 41.400 838.350 42.600 839.100 ;
        RECT 46.950 838.950 49.050 841.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 43.950 835.950 46.050 838.050 ;
        RECT 22.950 829.950 25.050 832.050 ;
        RECT 28.950 829.950 31.050 832.050 ;
        RECT 31.950 829.950 34.050 835.050 ;
        RECT 38.400 833.400 39.600 835.650 ;
        RECT 44.400 834.000 45.600 835.650 ;
        RECT 13.950 826.950 16.050 829.050 ;
        RECT 23.400 817.050 24.450 829.950 ;
        RECT 28.950 826.800 31.050 828.900 ;
        RECT 31.950 826.800 34.050 828.900 ;
        RECT 16.950 814.950 19.050 817.050 ;
        RECT 22.950 814.950 25.050 817.050 ;
        RECT 1.950 806.100 4.050 808.200 ;
        RECT 17.400 807.600 18.450 814.950 ;
        RECT 2.400 715.050 3.450 806.100 ;
        RECT 17.400 805.350 18.600 807.600 ;
        RECT 22.950 806.100 25.050 808.200 ;
        RECT 23.400 805.350 24.600 806.100 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 14.400 801.000 15.600 802.650 ;
        RECT 20.400 801.000 21.600 802.650 ;
        RECT 29.400 801.900 30.450 826.800 ;
        RECT 13.950 796.950 16.050 801.000 ;
        RECT 19.950 796.950 22.050 801.000 ;
        RECT 28.950 799.800 31.050 801.900 ;
        RECT 25.950 796.950 28.050 799.050 ;
        RECT 4.950 761.100 7.050 763.200 ;
        RECT 13.950 761.100 16.050 763.200 ;
        RECT 19.950 761.100 22.050 763.200 ;
        RECT 5.400 751.050 6.450 761.100 ;
        RECT 14.400 760.350 15.600 761.100 ;
        RECT 20.400 760.350 21.600 761.100 ;
        RECT 10.950 757.950 13.050 760.050 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 7.950 754.800 10.050 756.900 ;
        RECT 11.400 755.400 12.600 757.650 ;
        RECT 17.400 756.900 18.600 757.650 ;
        RECT 4.950 748.950 7.050 751.050 ;
        RECT 4.950 739.950 7.050 742.050 ;
        RECT 1.950 712.950 4.050 715.050 ;
        RECT 5.400 676.050 6.450 739.950 ;
        RECT 8.400 721.050 9.450 754.800 ;
        RECT 11.400 754.050 12.450 755.400 ;
        RECT 16.950 754.800 19.050 756.900 ;
        RECT 22.950 754.950 25.050 757.050 ;
        RECT 11.400 752.400 16.050 754.050 ;
        RECT 12.000 751.950 16.050 752.400 ;
        RECT 16.950 748.950 19.050 751.050 ;
        RECT 17.400 729.600 18.450 748.950 ;
        RECT 23.400 730.200 24.450 754.950 ;
        RECT 26.400 754.050 27.450 796.950 ;
        RECT 25.950 751.950 28.050 754.050 ;
        RECT 17.400 727.350 18.600 729.600 ;
        RECT 22.950 728.100 25.050 730.200 ;
        RECT 23.400 727.350 24.600 728.100 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 22.950 724.950 25.050 727.050 ;
        RECT 14.400 722.400 15.600 724.650 ;
        RECT 20.400 722.400 21.600 724.650 ;
        RECT 29.400 723.450 30.450 799.800 ;
        RECT 32.400 799.050 33.450 826.800 ;
        RECT 38.400 826.050 39.450 833.400 ;
        RECT 43.950 829.950 46.050 834.000 ;
        RECT 46.950 832.950 49.050 835.050 ;
        RECT 47.400 826.050 48.450 832.950 ;
        RECT 50.400 828.450 51.450 911.400 ;
        RECT 53.400 904.050 54.450 917.100 ;
        RECT 56.400 907.050 57.450 922.950 ;
        RECT 61.950 917.100 64.050 919.200 ;
        RECT 67.950 917.100 70.050 919.200 ;
        RECT 76.950 917.100 79.050 922.050 ;
        RECT 82.950 917.100 85.050 919.200 ;
        RECT 88.950 918.000 91.050 922.050 ;
        RECT 62.400 916.350 63.600 917.100 ;
        RECT 68.400 916.350 69.600 917.100 ;
        RECT 61.950 913.950 64.050 916.050 ;
        RECT 64.950 913.950 67.050 916.050 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 65.400 911.400 66.600 913.650 ;
        RECT 71.400 911.400 72.600 913.650 ;
        RECT 55.950 904.950 58.050 907.050 ;
        RECT 52.950 901.950 55.050 904.050 ;
        RECT 65.400 892.050 66.450 911.400 ;
        RECT 71.400 904.050 72.450 911.400 ;
        RECT 67.800 901.950 69.900 904.050 ;
        RECT 70.950 901.950 73.050 904.050 ;
        RECT 64.950 889.950 67.050 892.050 ;
        RECT 55.950 884.100 58.050 886.200 ;
        RECT 56.400 883.350 57.600 884.100 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 52.950 877.950 55.050 880.050 ;
        RECT 59.400 879.900 60.600 880.650 ;
        RECT 53.400 871.050 54.450 877.950 ;
        RECT 58.950 877.800 61.050 879.900 ;
        RECT 65.400 874.050 66.450 889.950 ;
        RECT 64.950 871.950 67.050 874.050 ;
        RECT 52.950 868.950 55.050 871.050 ;
        RECT 53.400 853.050 54.450 868.950 ;
        RECT 68.400 859.050 69.450 901.950 ;
        RECT 77.400 885.600 78.450 917.100 ;
        RECT 83.400 916.350 84.600 917.100 ;
        RECT 89.400 916.350 90.600 918.000 ;
        RECT 98.400 916.050 99.450 922.950 ;
        RECT 100.950 919.950 103.050 922.050 ;
        RECT 82.950 913.950 85.050 916.050 ;
        RECT 85.950 913.950 88.050 916.050 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 97.950 913.950 100.050 916.050 ;
        RECT 86.400 912.900 87.600 913.650 ;
        RECT 85.950 910.800 88.050 912.900 ;
        RECT 92.400 911.400 93.600 913.650 ;
        RECT 88.950 907.950 91.050 910.050 ;
        RECT 89.400 904.050 90.450 907.950 ;
        RECT 88.950 901.950 91.050 904.050 ;
        RECT 92.400 895.050 93.450 911.400 ;
        RECT 101.400 901.050 102.450 919.950 ;
        RECT 107.400 919.200 108.450 925.950 ;
        RECT 121.950 922.950 124.050 925.050 ;
        RECT 184.950 922.950 187.050 925.050 ;
        RECT 106.950 917.100 109.050 919.200 ;
        RECT 112.950 918.000 115.050 922.050 ;
        RECT 107.400 916.350 108.600 917.100 ;
        RECT 113.400 916.350 114.600 918.000 ;
        RECT 122.400 916.050 123.450 922.950 ;
        RECT 132.000 918.600 136.050 919.050 ;
        RECT 131.400 916.950 136.050 918.600 ;
        RECT 136.950 917.100 139.050 919.200 ;
        RECT 142.950 917.100 145.050 919.200 ;
        RECT 148.950 917.100 151.050 919.200 ;
        RECT 157.950 917.100 160.050 919.200 ;
        RECT 163.950 917.100 166.050 919.200 ;
        RECT 169.950 917.100 172.050 919.200 ;
        RECT 185.400 918.600 186.450 922.950 ;
        RECT 202.950 919.950 205.050 922.050 ;
        RECT 131.400 916.350 132.600 916.950 ;
        RECT 106.950 913.950 109.050 916.050 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 121.950 913.950 124.050 916.050 ;
        RECT 127.950 913.950 130.050 916.050 ;
        RECT 130.950 913.950 133.050 916.050 ;
        RECT 110.400 911.400 111.600 913.650 ;
        RECT 128.400 911.400 129.600 913.650 ;
        RECT 110.400 907.050 111.450 911.400 ;
        RECT 109.950 904.950 112.050 907.050 ;
        RECT 94.950 898.950 97.050 901.050 ;
        RECT 100.950 898.950 103.050 901.050 ;
        RECT 106.950 898.950 109.050 901.050 ;
        RECT 91.950 892.950 94.050 895.050 ;
        RECT 85.950 889.950 88.050 892.050 ;
        RECT 77.400 883.350 78.600 885.600 ;
        RECT 73.950 880.950 76.050 883.050 ;
        RECT 76.950 880.950 79.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 74.400 878.400 75.600 880.650 ;
        RECT 80.400 879.900 81.600 880.650 ;
        RECT 86.400 880.050 87.450 889.950 ;
        RECT 95.400 885.600 96.450 898.950 ;
        RECT 95.400 883.350 96.600 885.600 ;
        RECT 100.950 884.100 103.050 886.200 ;
        RECT 101.400 883.350 102.600 884.100 ;
        RECT 91.950 880.950 94.050 883.050 ;
        RECT 94.950 880.950 97.050 883.050 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 100.950 880.950 103.050 883.050 ;
        RECT 74.400 874.050 75.450 878.400 ;
        RECT 79.950 877.800 82.050 879.900 ;
        RECT 85.950 877.950 88.050 880.050 ;
        RECT 92.400 878.400 93.600 880.650 ;
        RECT 98.400 878.400 99.600 880.650 ;
        RECT 73.950 871.950 76.050 874.050 ;
        RECT 74.400 868.050 75.450 871.950 ;
        RECT 73.950 865.950 76.050 868.050 ;
        RECT 92.400 859.050 93.450 878.400 ;
        RECT 98.400 862.050 99.450 878.400 ;
        RECT 103.950 877.950 106.050 880.050 ;
        RECT 107.400 879.450 108.450 898.950 ;
        RECT 128.400 898.050 129.450 911.400 ;
        RECT 137.400 910.050 138.450 917.100 ;
        RECT 143.400 916.350 144.600 917.100 ;
        RECT 149.400 916.350 150.600 917.100 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 148.950 913.950 151.050 916.050 ;
        RECT 151.950 913.950 154.050 916.050 ;
        RECT 146.400 912.900 147.600 913.650 ;
        RECT 136.950 907.950 139.050 910.050 ;
        RECT 139.950 907.950 142.050 912.900 ;
        RECT 145.950 910.800 148.050 912.900 ;
        RECT 152.400 911.400 153.600 913.650 ;
        RECT 130.950 904.950 136.050 907.050 ;
        RECT 138.000 906.900 141.000 907.050 ;
        RECT 136.950 904.950 142.050 906.900 ;
        RECT 136.950 904.800 139.050 904.950 ;
        RECT 139.950 904.800 142.050 904.950 ;
        RECT 152.400 904.050 153.450 911.400 ;
        RECT 158.400 907.050 159.450 917.100 ;
        RECT 164.400 916.350 165.600 917.100 ;
        RECT 170.400 916.350 171.600 917.100 ;
        RECT 185.400 916.350 186.600 918.600 ;
        RECT 190.950 917.100 193.050 919.200 ;
        RECT 191.400 916.350 192.600 917.100 ;
        RECT 199.950 916.950 202.050 919.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 166.950 913.950 169.050 916.050 ;
        RECT 169.950 913.950 172.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 190.950 913.950 193.050 916.050 ;
        RECT 193.950 913.950 196.050 916.050 ;
        RECT 167.400 912.900 168.600 913.650 ;
        RECT 166.950 910.800 169.050 912.900 ;
        RECT 188.400 912.000 189.600 913.650 ;
        RECT 194.400 912.900 195.600 913.650 ;
        RECT 187.950 907.950 190.050 912.000 ;
        RECT 193.950 910.800 196.050 912.900 ;
        RECT 157.950 904.950 160.050 907.050 ;
        RECT 151.950 901.950 154.050 904.050 ;
        RECT 200.400 901.050 201.450 916.950 ;
        RECT 203.400 904.050 204.450 919.950 ;
        RECT 208.950 919.050 211.050 919.200 ;
        RECT 205.950 917.100 211.050 919.050 ;
        RECT 214.950 918.000 217.050 922.050 ;
        RECT 205.950 916.950 210.600 917.100 ;
        RECT 209.400 916.350 210.600 916.950 ;
        RECT 215.400 916.350 216.600 918.000 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 211.950 913.950 214.050 916.050 ;
        RECT 214.950 913.950 217.050 916.050 ;
        RECT 212.400 912.900 213.600 913.650 ;
        RECT 221.400 913.050 222.450 928.950 ;
        RECT 226.950 917.100 229.050 919.200 ;
        RECT 232.950 917.100 235.050 919.200 ;
        RECT 241.950 917.100 244.050 919.200 ;
        RECT 227.400 916.350 228.600 917.100 ;
        RECT 233.400 916.350 234.600 917.100 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 235.950 913.950 238.050 916.050 ;
        RECT 205.950 910.800 208.050 912.900 ;
        RECT 211.950 910.800 214.050 912.900 ;
        RECT 220.950 910.950 223.050 913.050 ;
        RECT 230.400 911.400 231.600 913.650 ;
        RECT 236.400 913.050 237.600 913.650 ;
        RECT 236.400 911.400 241.050 913.050 ;
        RECT 202.950 901.950 205.050 904.050 ;
        RECT 206.400 901.050 207.450 910.800 ;
        RECT 230.400 904.050 231.450 911.400 ;
        RECT 237.000 910.950 241.050 911.400 ;
        RECT 242.400 910.050 243.450 917.100 ;
        RECT 245.400 913.050 246.450 931.950 ;
        RECT 256.950 928.950 259.050 931.050 ;
        RECT 250.950 922.950 253.050 925.050 ;
        RECT 251.400 918.600 252.450 922.950 ;
        RECT 257.400 918.600 258.450 928.950 ;
        RECT 275.400 918.600 276.450 931.950 ;
        RECT 352.950 928.950 355.050 931.050 ;
        RECT 365.700 930.300 367.800 932.400 ;
        RECT 286.950 925.950 289.050 928.050 ;
        RECT 251.400 916.350 252.600 918.600 ;
        RECT 257.400 916.350 258.600 918.600 ;
        RECT 275.400 916.350 276.600 918.600 ;
        RECT 280.950 917.100 283.050 919.200 ;
        RECT 281.400 916.350 282.600 917.100 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 256.950 913.950 259.050 916.050 ;
        RECT 259.950 913.950 262.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 280.950 913.950 283.050 916.050 ;
        RECT 244.950 910.950 247.050 913.050 ;
        RECT 254.400 911.400 255.600 913.650 ;
        RECT 260.400 912.900 261.600 913.650 ;
        RECT 278.400 912.900 279.600 913.650 ;
        RECT 287.400 912.900 288.450 925.950 ;
        RECT 305.400 918.450 306.600 918.600 ;
        RECT 305.400 917.400 309.450 918.450 ;
        RECT 305.400 916.350 306.600 917.400 ;
        RECT 296.100 913.950 298.200 916.050 ;
        RECT 299.400 913.950 301.500 916.050 ;
        RECT 304.800 913.950 306.900 916.050 ;
        RECT 241.950 907.950 244.050 910.050 ;
        RECT 242.400 904.050 243.450 907.950 ;
        RECT 229.950 901.950 232.050 904.050 ;
        RECT 241.950 901.950 244.050 904.050 ;
        RECT 139.950 898.950 142.050 901.050 ;
        RECT 199.950 898.950 202.050 901.050 ;
        RECT 205.950 898.950 208.050 901.050 ;
        RECT 238.950 898.950 241.050 901.050 ;
        RECT 127.950 895.950 130.050 898.050 ;
        RECT 133.950 895.950 136.050 898.050 ;
        RECT 115.950 884.100 118.050 886.200 ;
        RECT 128.400 886.050 129.450 895.950 ;
        RECT 116.400 883.350 117.600 884.100 ;
        RECT 124.950 883.950 127.050 886.050 ;
        RECT 127.950 883.950 130.050 886.050 ;
        RECT 134.400 885.600 135.450 895.950 ;
        RECT 140.400 885.600 141.450 898.950 ;
        RECT 148.950 892.950 151.050 895.050 ;
        RECT 196.950 892.950 199.050 895.050 ;
        RECT 217.950 894.450 220.050 895.050 ;
        RECT 223.950 894.450 226.050 895.050 ;
        RECT 217.950 893.400 226.050 894.450 ;
        RECT 217.950 892.950 220.050 893.400 ;
        RECT 223.950 892.950 226.050 893.400 ;
        RECT 112.950 880.950 115.050 883.050 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 118.950 880.950 121.050 883.050 ;
        RECT 113.400 879.450 114.600 880.650 ;
        RECT 107.400 878.400 114.600 879.450 ;
        RECT 119.400 878.400 120.600 880.650 ;
        RECT 97.950 859.950 100.050 862.050 ;
        RECT 58.950 856.950 61.050 859.050 ;
        RECT 67.950 856.950 70.050 859.050 ;
        RECT 91.950 856.950 94.050 859.050 ;
        RECT 52.950 850.950 55.050 853.050 ;
        RECT 59.400 844.050 60.450 856.950 ;
        RECT 104.400 853.050 105.450 877.950 ;
        RECT 109.950 871.950 112.050 874.050 ;
        RECT 73.950 850.950 76.050 853.050 ;
        RECT 103.950 850.950 106.050 853.050 ;
        RECT 64.950 844.950 67.050 847.050 ;
        RECT 52.950 841.950 55.050 844.050 ;
        RECT 53.400 832.050 54.450 841.950 ;
        RECT 58.950 840.000 61.050 844.050 ;
        RECT 65.400 840.600 66.450 844.950 ;
        RECT 59.400 838.350 60.600 840.000 ;
        RECT 65.400 838.350 66.600 840.600 ;
        RECT 74.400 838.050 75.450 850.950 ;
        RECT 88.950 844.950 91.050 847.050 ;
        RECT 89.400 841.200 90.450 844.950 ;
        RECT 76.950 839.100 79.050 841.200 ;
        RECT 82.950 839.100 85.050 841.200 ;
        RECT 88.950 839.100 91.050 841.200 ;
        RECT 97.950 839.100 100.050 841.200 ;
        RECT 104.400 840.600 105.450 850.950 ;
        RECT 110.400 841.200 111.450 871.950 ;
        RECT 119.400 871.050 120.450 878.400 ;
        RECT 121.950 877.950 124.050 880.050 ;
        RECT 118.950 868.950 121.050 871.050 ;
        RECT 122.400 867.450 123.450 877.950 ;
        RECT 125.400 877.050 126.450 883.950 ;
        RECT 134.400 883.350 135.600 885.600 ;
        RECT 140.400 883.350 141.600 885.600 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 131.400 879.900 132.600 880.650 ;
        RECT 130.950 877.800 133.050 879.900 ;
        RECT 137.400 879.000 138.600 880.650 ;
        RECT 149.400 879.900 150.450 892.950 ;
        RECT 166.950 889.950 169.050 892.050 ;
        RECT 154.950 888.450 157.050 889.050 ;
        RECT 160.950 888.450 163.050 889.050 ;
        RECT 154.950 887.400 163.050 888.450 ;
        RECT 154.950 886.950 157.050 887.400 ;
        RECT 160.950 886.950 163.050 887.400 ;
        RECT 157.950 884.100 160.050 886.200 ;
        RECT 158.400 883.350 159.600 884.100 ;
        RECT 154.950 880.950 157.050 883.050 ;
        RECT 157.950 880.950 160.050 883.050 ;
        RECT 160.950 880.950 163.050 883.050 ;
        RECT 155.400 879.900 156.600 880.650 ;
        RECT 161.400 879.900 162.600 880.650 ;
        RECT 167.400 879.900 168.450 889.950 ;
        RECT 175.950 884.100 178.050 886.200 ;
        RECT 176.400 883.350 177.600 884.100 ;
        RECT 187.950 883.950 190.050 886.050 ;
        RECT 197.400 885.600 198.450 892.950 ;
        RECT 220.950 889.950 223.050 892.050 ;
        RECT 229.950 889.950 232.050 892.050 ;
        RECT 172.950 880.950 175.050 883.050 ;
        RECT 175.950 880.950 178.050 883.050 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 124.950 874.950 127.050 877.050 ;
        RECT 136.950 874.950 139.050 879.000 ;
        RECT 148.950 877.800 151.050 879.900 ;
        RECT 154.950 877.800 157.050 879.900 ;
        RECT 160.950 877.800 163.050 879.900 ;
        RECT 166.950 877.800 169.050 879.900 ;
        RECT 173.400 878.400 174.600 880.650 ;
        RECT 179.400 879.900 180.600 880.650 ;
        RECT 188.400 879.900 189.450 883.950 ;
        RECT 197.400 883.350 198.600 885.600 ;
        RECT 205.950 883.950 208.050 886.050 ;
        RECT 214.950 884.100 217.050 886.200 ;
        RECT 221.400 885.600 222.450 889.950 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 194.400 879.900 195.600 880.650 ;
        RECT 200.400 879.900 201.600 880.650 ;
        RECT 157.950 874.950 160.050 877.050 ;
        RECT 154.950 871.950 157.050 874.050 ;
        RECT 119.400 866.400 123.450 867.450 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 62.400 834.900 63.600 835.650 ;
        RECT 61.950 832.800 64.050 834.900 ;
        RECT 68.400 833.400 69.600 835.650 ;
        RECT 52.950 829.950 55.050 832.050 ;
        RECT 68.400 829.050 69.450 833.400 ;
        RECT 50.400 827.400 54.450 828.450 ;
        RECT 37.950 823.950 40.050 826.050 ;
        RECT 46.950 823.950 49.050 826.050 ;
        RECT 46.950 811.950 49.050 814.050 ;
        RECT 40.950 806.100 43.050 811.050 ;
        RECT 47.400 807.600 48.450 811.950 ;
        RECT 41.400 805.350 42.600 806.100 ;
        RECT 47.400 805.350 48.600 807.600 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 38.400 801.900 39.600 802.650 ;
        RECT 37.950 799.800 40.050 801.900 ;
        RECT 44.400 801.000 45.600 802.650 ;
        RECT 31.950 796.950 34.050 799.050 ;
        RECT 43.950 796.950 46.050 801.000 ;
        RECT 53.400 799.050 54.450 827.400 ;
        RECT 67.950 826.950 70.050 829.050 ;
        RECT 77.400 828.450 78.450 839.100 ;
        RECT 83.400 838.350 84.600 839.100 ;
        RECT 89.400 838.350 90.600 839.100 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 88.950 835.950 91.050 838.050 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 86.400 834.000 87.600 835.650 ;
        RECT 85.950 829.950 88.050 834.000 ;
        RECT 92.400 833.400 93.600 835.650 ;
        RECT 79.950 828.450 82.050 829.050 ;
        RECT 77.400 827.400 82.050 828.450 ;
        RECT 79.950 826.950 82.050 827.400 ;
        RECT 70.950 817.950 73.050 820.050 ;
        RECT 55.950 811.950 58.050 814.050 ;
        RECT 71.400 813.450 72.450 817.950 ;
        RECT 56.400 801.900 57.450 811.950 ;
        RECT 71.400 811.200 72.600 813.450 ;
        RECT 58.950 806.100 61.050 808.200 ;
        RECT 66.900 807.900 69.000 809.700 ;
        RECT 70.800 808.800 72.900 810.900 ;
        RECT 74.100 810.300 76.200 812.400 ;
        RECT 65.400 806.700 74.100 807.900 ;
        RECT 55.950 799.800 58.050 801.900 ;
        RECT 46.950 796.950 49.050 799.050 ;
        RECT 52.950 796.950 55.050 799.050 ;
        RECT 34.950 790.950 37.050 793.050 ;
        RECT 43.950 790.950 46.050 793.050 ;
        RECT 35.400 762.600 36.450 790.950 ;
        RECT 35.400 760.350 36.600 762.600 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 38.400 755.400 39.600 757.650 ;
        RECT 38.400 745.050 39.450 755.400 ;
        RECT 37.950 742.950 40.050 745.050 ;
        RECT 34.950 733.950 37.050 736.050 ;
        RECT 31.950 728.100 34.050 730.200 ;
        RECT 32.400 724.050 33.450 728.100 ;
        RECT 26.400 722.400 30.450 723.450 ;
        RECT 7.950 718.950 10.050 721.050 ;
        RECT 14.400 718.050 15.450 722.400 ;
        RECT 20.400 721.050 21.450 722.400 ;
        RECT 19.950 718.950 22.050 721.050 ;
        RECT 13.950 715.950 16.050 718.050 ;
        RECT 7.950 706.950 10.050 709.050 ;
        RECT 4.950 673.950 7.050 676.050 ;
        RECT 8.400 609.450 9.450 706.950 ;
        RECT 14.400 691.050 15.450 715.950 ;
        RECT 13.950 688.950 16.050 691.050 ;
        RECT 11.400 679.950 13.500 682.050 ;
        RECT 16.500 679.950 18.600 682.050 ;
        RECT 17.400 678.900 18.600 679.650 ;
        RECT 16.950 676.800 19.050 678.900 ;
        RECT 10.950 673.950 13.050 676.050 ;
        RECT 5.400 608.400 9.450 609.450 ;
        RECT 5.400 567.900 6.450 608.400 ;
        RECT 11.400 607.050 12.450 673.950 ;
        RECT 20.400 664.050 21.450 718.950 ;
        RECT 22.950 688.950 25.050 691.050 ;
        RECT 23.400 679.050 24.450 688.950 ;
        RECT 22.950 676.950 25.050 679.050 ;
        RECT 19.950 661.950 22.050 664.050 ;
        RECT 14.400 646.950 16.500 649.050 ;
        RECT 19.800 646.950 21.900 649.050 ;
        RECT 20.400 644.400 21.600 646.650 ;
        RECT 20.400 634.050 21.450 644.400 ;
        RECT 19.950 631.950 22.050 634.050 ;
        RECT 26.400 613.050 27.450 722.400 ;
        RECT 31.950 721.950 34.050 724.050 ;
        RECT 35.400 718.050 36.450 733.950 ;
        RECT 44.400 733.050 45.450 790.950 ;
        RECT 47.400 756.450 48.450 796.950 ;
        RECT 59.400 793.050 60.450 806.100 ;
        RECT 62.100 802.950 64.200 805.050 ;
        RECT 62.400 801.900 63.600 802.650 ;
        RECT 61.950 799.800 64.050 801.900 ;
        RECT 65.400 797.700 66.300 806.700 ;
        RECT 72.000 805.800 74.100 806.700 ;
        RECT 75.000 804.900 75.900 810.300 ;
        RECT 76.950 806.100 79.050 808.200 ;
        RECT 77.400 805.350 78.600 806.100 ;
        RECT 69.000 803.700 75.900 804.900 ;
        RECT 69.000 801.300 69.900 803.700 ;
        RECT 67.800 799.200 69.900 801.300 ;
        RECT 70.800 799.950 72.900 802.050 ;
        RECT 64.500 795.600 66.600 797.700 ;
        RECT 71.400 797.400 72.600 799.650 ;
        RECT 74.700 796.500 75.900 803.700 ;
        RECT 76.800 802.950 78.900 805.050 ;
        RECT 74.100 794.400 76.200 796.500 ;
        RECT 58.950 790.950 61.050 793.050 ;
        RECT 49.950 769.950 52.050 772.050 ;
        RECT 50.400 763.200 51.450 769.950 ;
        RECT 80.400 769.050 81.450 826.950 ;
        RECT 82.950 820.950 85.050 823.050 ;
        RECT 83.400 793.050 84.450 820.950 ;
        RECT 88.950 810.450 91.050 811.050 ;
        RECT 92.400 810.450 93.450 833.400 ;
        RECT 98.400 823.050 99.450 839.100 ;
        RECT 104.400 838.350 105.600 840.600 ;
        RECT 109.950 839.100 112.050 841.200 ;
        RECT 115.950 839.100 118.050 841.200 ;
        RECT 119.400 841.050 120.450 866.400 ;
        RECT 155.400 862.050 156.450 871.950 ;
        RECT 158.400 868.050 159.450 874.950 ;
        RECT 173.400 874.050 174.450 878.400 ;
        RECT 178.950 877.800 181.050 879.900 ;
        RECT 187.950 877.800 190.050 879.900 ;
        RECT 193.950 877.800 196.050 879.900 ;
        RECT 199.950 877.800 202.050 879.900 ;
        RECT 200.400 876.450 201.450 877.800 ;
        RECT 206.400 877.050 207.450 883.950 ;
        RECT 215.400 883.350 216.600 884.100 ;
        RECT 221.400 883.350 222.600 885.600 ;
        RECT 211.950 880.950 214.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 217.950 880.950 220.050 883.050 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 212.400 878.400 213.600 880.650 ;
        RECT 218.400 879.000 219.600 880.650 ;
        RECT 230.400 879.900 231.450 889.950 ;
        RECT 239.400 885.600 240.450 898.950 ;
        RECT 254.400 885.600 255.450 911.400 ;
        RECT 259.950 910.800 262.050 912.900 ;
        RECT 277.950 910.800 280.050 912.900 ;
        RECT 286.950 910.800 289.050 912.900 ;
        RECT 299.400 911.400 300.600 913.650 ;
        RECT 299.400 904.050 300.450 911.400 ;
        RECT 298.950 901.950 301.050 904.050 ;
        RECT 256.950 894.450 259.050 895.050 ;
        RECT 262.950 894.450 265.050 895.050 ;
        RECT 256.950 893.400 265.050 894.450 ;
        RECT 256.950 892.950 259.050 893.400 ;
        RECT 262.950 892.950 265.050 893.400 ;
        RECT 295.950 892.950 298.050 895.050 ;
        RECT 259.950 889.950 262.050 892.050 ;
        RECT 260.400 886.200 261.450 889.950 ;
        RECT 239.400 883.350 240.600 885.600 ;
        RECT 254.400 883.350 255.600 885.600 ;
        RECT 259.950 884.100 262.050 886.200 ;
        RECT 277.950 884.100 280.050 886.200 ;
        RECT 283.950 885.000 286.050 889.050 ;
        RECT 289.950 886.950 292.050 889.050 ;
        RECT 260.400 883.350 261.600 884.100 ;
        RECT 278.400 883.350 279.600 884.100 ;
        RECT 284.400 883.350 285.600 885.000 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 262.950 880.950 265.050 883.050 ;
        RECT 277.950 880.950 280.050 883.050 ;
        RECT 280.950 880.950 283.050 883.050 ;
        RECT 283.950 880.950 286.050 883.050 ;
        RECT 236.400 879.900 237.600 880.650 ;
        RECT 197.400 875.400 201.450 876.450 ;
        RECT 172.950 871.950 175.050 874.050 ;
        RECT 157.950 865.950 160.050 868.050 ;
        RECT 154.950 859.950 157.050 862.050 ;
        RECT 110.400 838.350 111.600 839.100 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 109.950 835.950 112.050 838.050 ;
        RECT 107.400 834.900 108.600 835.650 ;
        RECT 106.950 832.800 109.050 834.900 ;
        RECT 112.950 832.950 115.050 835.050 ;
        RECT 97.950 820.950 100.050 823.050 ;
        RECT 113.400 820.050 114.450 832.950 ;
        RECT 112.950 817.950 115.050 820.050 ;
        RECT 116.400 814.050 117.450 839.100 ;
        RECT 118.950 838.950 121.050 841.050 ;
        RECT 121.950 839.100 124.050 841.200 ;
        RECT 127.950 839.100 130.050 841.200 ;
        RECT 148.950 839.100 151.050 841.200 ;
        RECT 122.400 838.350 123.600 839.100 ;
        RECT 128.400 838.350 129.600 839.100 ;
        RECT 149.400 838.350 150.600 839.100 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 130.950 835.950 133.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 148.950 835.950 151.050 838.050 ;
        RECT 125.400 834.900 126.600 835.650 ;
        RECT 124.950 832.800 127.050 834.900 ;
        RECT 131.400 833.400 132.600 835.650 ;
        RECT 146.400 833.400 147.600 835.650 ;
        RECT 131.400 829.050 132.450 833.400 ;
        RECT 146.400 829.050 147.450 833.400 ;
        RECT 155.400 831.450 156.450 859.950 ;
        RECT 197.400 847.050 198.450 875.400 ;
        RECT 205.950 874.950 208.050 877.050 ;
        RECT 212.400 874.050 213.450 878.400 ;
        RECT 217.950 874.950 220.050 879.000 ;
        RECT 229.950 877.800 232.050 879.900 ;
        RECT 235.950 877.800 238.050 879.900 ;
        RECT 257.400 878.400 258.600 880.650 ;
        RECT 281.400 878.400 282.600 880.650 ;
        RECT 257.400 874.050 258.450 878.400 ;
        RECT 199.950 871.950 202.050 874.050 ;
        RECT 211.950 871.950 214.050 874.050 ;
        RECT 220.950 871.950 223.050 874.050 ;
        RECT 256.950 871.950 259.050 874.050 ;
        RECT 200.400 853.050 201.450 871.950 ;
        RECT 221.400 868.050 222.450 871.950 ;
        RECT 220.950 865.950 223.050 868.050 ;
        RECT 199.950 850.950 202.050 853.050 ;
        RECT 163.800 844.500 165.900 846.600 ;
        RECT 157.950 838.950 160.050 841.050 ;
        RECT 152.400 830.400 156.450 831.450 ;
        RECT 158.400 834.450 159.450 838.950 ;
        RECT 161.100 835.950 163.200 838.050 ;
        RECT 164.100 837.300 165.300 844.500 ;
        RECT 167.400 841.350 168.600 843.600 ;
        RECT 173.400 843.300 175.500 845.400 ;
        RECT 196.950 844.950 199.050 847.050 ;
        RECT 167.100 838.950 169.200 841.050 ;
        RECT 170.100 839.700 172.200 841.800 ;
        RECT 170.100 837.300 171.000 839.700 ;
        RECT 164.100 836.100 171.000 837.300 ;
        RECT 161.400 834.450 162.600 835.650 ;
        RECT 158.400 833.400 162.600 834.450 ;
        RECT 118.950 826.950 121.050 829.050 ;
        RECT 130.950 826.950 133.050 829.050 ;
        RECT 145.950 826.950 148.050 829.050 ;
        RECT 94.950 811.950 97.050 814.050 ;
        RECT 115.950 811.950 118.050 814.050 ;
        RECT 88.950 809.400 93.450 810.450 ;
        RECT 88.950 807.000 91.050 809.400 ;
        RECT 95.400 807.600 96.450 811.950 ;
        RECT 89.400 805.350 90.600 807.000 ;
        RECT 95.400 805.350 96.600 807.600 ;
        RECT 106.950 806.100 109.050 808.200 ;
        RECT 112.950 806.100 115.050 808.200 ;
        RECT 119.400 807.600 120.450 826.950 ;
        RECT 127.950 811.950 130.050 814.050 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 91.950 802.950 94.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 92.400 800.400 93.600 802.650 ;
        RECT 98.400 801.000 99.600 802.650 ;
        RECT 92.400 798.450 93.450 800.400 ;
        RECT 92.400 797.400 96.450 798.450 ;
        RECT 82.950 790.950 85.050 793.050 ;
        RECT 91.950 790.950 94.050 793.050 ;
        RECT 79.950 766.950 82.050 769.050 ;
        RECT 88.950 766.950 91.050 769.050 ;
        RECT 49.950 761.100 52.050 763.200 ;
        RECT 55.950 761.100 58.050 763.200 ;
        RECT 61.950 761.100 64.050 763.200 ;
        RECT 67.950 761.100 70.050 763.200 ;
        RECT 76.950 761.100 79.050 763.200 ;
        RECT 82.950 761.100 85.050 763.200 ;
        RECT 56.400 760.350 57.600 761.100 ;
        RECT 62.400 760.350 63.600 761.100 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 47.400 755.400 51.450 756.450 ;
        RECT 43.950 730.950 46.050 733.050 ;
        RECT 38.100 724.950 40.200 727.050 ;
        RECT 43.500 724.950 45.600 727.050 ;
        RECT 38.400 723.900 39.600 724.650 ;
        RECT 37.950 721.800 40.050 723.900 ;
        RECT 34.950 715.950 37.050 718.050 ;
        RECT 50.400 705.450 51.450 755.400 ;
        RECT 53.400 755.400 54.600 757.650 ;
        RECT 59.400 756.900 60.600 757.650 ;
        RECT 53.400 753.450 54.450 755.400 ;
        RECT 58.950 754.800 61.050 756.900 ;
        RECT 53.400 752.400 57.450 753.450 ;
        RECT 52.950 748.950 55.050 751.050 ;
        RECT 53.400 709.050 54.450 748.950 ;
        RECT 56.400 748.050 57.450 752.400 ;
        RECT 55.950 745.950 58.050 748.050 ;
        RECT 56.400 729.450 57.450 745.950 ;
        RECT 64.950 735.450 67.050 736.050 ;
        RECT 68.400 735.450 69.450 761.100 ;
        RECT 77.400 760.350 78.600 761.100 ;
        RECT 83.400 760.350 84.600 761.100 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 74.400 755.400 75.600 757.650 ;
        RECT 80.400 755.400 81.600 757.650 ;
        RECT 74.400 745.050 75.450 755.400 ;
        RECT 80.400 754.050 81.450 755.400 ;
        RECT 85.950 754.950 88.050 757.050 ;
        RECT 76.950 752.400 81.450 754.050 ;
        RECT 76.950 751.950 81.000 752.400 ;
        RECT 82.950 751.950 85.050 754.050 ;
        RECT 73.950 742.950 76.050 745.050 ;
        RECT 64.950 734.400 69.450 735.450 ;
        RECT 64.950 733.950 67.050 734.400 ;
        RECT 58.950 729.450 61.050 730.200 ;
        RECT 56.400 728.400 61.050 729.450 ;
        RECT 58.950 728.100 61.050 728.400 ;
        RECT 65.400 729.600 66.450 733.950 ;
        RECT 59.400 727.350 60.600 728.100 ;
        RECT 65.400 727.350 66.600 729.600 ;
        RECT 70.950 728.100 73.050 730.200 ;
        RECT 76.950 728.100 79.050 730.200 ;
        RECT 83.400 729.600 84.450 751.950 ;
        RECT 86.400 748.050 87.450 754.950 ;
        RECT 89.400 754.050 90.450 766.950 ;
        RECT 88.950 751.950 91.050 754.050 ;
        RECT 85.950 745.950 88.050 748.050 ;
        RECT 92.400 745.050 93.450 790.950 ;
        RECT 95.400 790.050 96.450 797.400 ;
        RECT 97.950 796.950 100.050 801.000 ;
        RECT 107.400 799.050 108.450 806.100 ;
        RECT 113.400 805.350 114.600 806.100 ;
        RECT 119.400 805.350 120.600 807.600 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 116.400 801.000 117.600 802.650 ;
        RECT 122.400 801.900 123.600 802.650 ;
        RECT 128.400 801.900 129.450 811.950 ;
        RECT 136.950 807.000 139.050 811.050 ;
        RECT 137.400 805.350 138.600 807.000 ;
        RECT 145.950 806.100 148.050 808.200 ;
        RECT 134.100 802.950 136.200 805.050 ;
        RECT 137.400 802.950 139.500 805.050 ;
        RECT 142.800 802.950 144.900 805.050 ;
        RECT 106.950 796.950 109.050 799.050 ;
        RECT 109.950 796.950 112.050 799.050 ;
        RECT 112.950 796.950 115.050 799.050 ;
        RECT 110.400 790.050 111.450 796.950 ;
        RECT 94.950 787.950 97.050 790.050 ;
        RECT 109.950 787.950 112.050 790.050 ;
        RECT 94.950 772.950 97.050 775.050 ;
        RECT 95.400 763.050 96.450 772.950 ;
        RECT 103.950 766.950 106.050 769.050 ;
        RECT 94.950 760.950 97.050 763.050 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 104.400 762.600 105.450 766.950 ;
        RECT 110.400 763.050 111.450 787.950 ;
        RECT 98.400 760.350 99.600 761.100 ;
        RECT 104.400 760.350 105.600 762.600 ;
        RECT 109.950 760.950 112.050 763.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 101.400 755.400 102.600 757.650 ;
        RECT 107.400 756.900 108.600 757.650 ;
        RECT 97.950 753.450 100.050 754.050 ;
        RECT 101.400 753.450 102.450 755.400 ;
        RECT 106.950 754.800 109.050 756.900 ;
        RECT 97.950 752.400 102.450 753.450 ;
        RECT 97.950 751.950 100.050 752.400 ;
        RECT 91.950 742.950 94.050 745.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 61.950 724.950 64.050 727.050 ;
        RECT 64.950 724.950 67.050 727.050 ;
        RECT 62.400 722.400 63.600 724.650 ;
        RECT 62.400 715.050 63.450 722.400 ;
        RECT 71.400 718.050 72.450 728.100 ;
        RECT 77.400 727.350 78.600 728.100 ;
        RECT 83.400 727.350 84.600 729.600 ;
        RECT 88.950 728.100 91.050 730.200 ;
        RECT 89.400 727.350 90.600 728.100 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 80.400 723.900 81.600 724.650 ;
        RECT 79.950 721.800 82.050 723.900 ;
        RECT 86.400 722.400 87.600 724.650 ;
        RECT 64.950 715.950 67.050 718.050 ;
        RECT 70.950 715.950 73.050 718.050 ;
        RECT 61.950 712.950 64.050 715.050 ;
        RECT 52.950 706.950 55.050 709.050 ;
        RECT 50.400 704.400 54.450 705.450 ;
        RECT 53.400 684.600 54.450 704.400 ;
        RECT 53.400 682.350 54.600 684.600 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 28.950 676.950 31.050 679.050 ;
        RECT 35.400 678.900 36.600 679.650 ;
        RECT 50.400 678.900 51.600 679.650 ;
        RECT 29.400 640.050 30.450 676.950 ;
        RECT 34.950 676.800 37.050 678.900 ;
        RECT 49.950 676.800 52.050 678.900 ;
        RECT 56.400 677.400 57.600 679.650 ;
        RECT 35.400 654.450 36.450 676.800 ;
        RECT 56.400 673.050 57.450 677.400 ;
        RECT 55.950 670.950 58.050 673.050 ;
        RECT 58.950 667.950 61.050 670.050 ;
        RECT 49.950 661.950 52.050 664.050 ;
        RECT 40.950 658.950 43.050 661.050 ;
        RECT 41.400 654.450 42.450 658.950 ;
        RECT 32.400 653.400 36.450 654.450 ;
        RECT 38.400 653.400 42.450 654.450 ;
        RECT 28.950 637.950 31.050 640.050 ;
        RECT 32.400 619.050 33.450 653.400 ;
        RECT 38.400 651.600 39.450 653.400 ;
        RECT 38.400 649.350 39.600 651.600 ;
        RECT 35.100 646.950 37.200 649.050 ;
        RECT 38.400 646.950 40.500 649.050 ;
        RECT 43.800 646.950 45.900 649.050 ;
        RECT 35.400 644.400 36.600 646.650 ;
        RECT 44.400 645.000 45.600 646.650 ;
        RECT 31.950 616.950 34.050 619.050 ;
        RECT 22.950 610.950 25.050 613.050 ;
        RECT 25.950 610.950 28.050 613.050 ;
        RECT 31.950 610.950 34.050 613.050 ;
        RECT 23.400 607.050 24.450 610.950 ;
        RECT 10.950 604.950 13.050 607.050 ;
        RECT 22.950 604.950 25.050 607.050 ;
        RECT 32.400 606.600 33.450 610.950 ;
        RECT 35.400 610.050 36.450 644.400 ;
        RECT 43.950 640.950 46.050 645.000 ;
        RECT 50.400 631.050 51.450 661.950 ;
        RECT 59.400 651.600 60.450 667.950 ;
        RECT 62.400 658.050 63.450 712.950 ;
        RECT 65.400 679.050 66.450 715.950 ;
        RECT 86.400 715.050 87.450 722.400 ;
        RECT 76.950 712.950 79.050 715.050 ;
        RECT 85.950 712.950 88.050 715.050 ;
        RECT 73.950 700.950 76.050 703.050 ;
        RECT 74.400 687.450 75.450 700.950 ;
        RECT 71.400 686.400 75.450 687.450 ;
        RECT 71.400 684.600 72.450 686.400 ;
        RECT 77.400 684.600 78.450 712.950 ;
        RECT 98.400 709.050 99.450 751.950 ;
        RECT 113.400 750.450 114.450 796.950 ;
        RECT 115.950 793.950 118.050 801.000 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 127.950 799.800 130.050 801.900 ;
        RECT 134.400 800.400 135.600 802.650 ;
        RECT 143.400 801.450 144.600 802.650 ;
        RECT 146.400 801.450 147.450 806.100 ;
        RECT 152.400 802.050 153.450 830.400 ;
        RECT 158.400 814.050 159.450 833.400 ;
        RECT 164.100 830.700 165.000 836.100 ;
        RECT 165.900 834.300 168.000 835.200 ;
        RECT 173.700 834.300 174.600 843.300 ;
        RECT 176.400 840.450 177.600 840.600 ;
        RECT 176.400 839.400 180.450 840.450 ;
        RECT 176.400 838.350 177.600 839.400 ;
        RECT 175.800 835.950 177.900 838.050 ;
        RECT 179.400 835.050 180.450 839.400 ;
        RECT 190.950 839.100 193.050 841.200 ;
        RECT 191.400 838.350 192.600 839.100 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 165.900 833.100 174.600 834.300 ;
        RECT 163.800 828.600 165.900 830.700 ;
        RECT 167.100 830.100 169.200 832.200 ;
        RECT 171.000 831.300 173.100 833.100 ;
        RECT 178.950 832.950 181.050 835.050 ;
        RECT 188.400 833.400 189.600 835.650 ;
        RECT 188.400 831.450 189.450 833.400 ;
        RECT 188.400 830.400 192.450 831.450 ;
        RECT 167.400 829.050 168.600 829.800 ;
        RECT 166.950 826.950 169.050 829.050 ;
        RECT 175.950 814.950 178.050 817.050 ;
        RECT 157.950 811.950 160.050 814.050 ;
        RECT 166.950 811.950 169.050 814.050 ;
        RECT 160.950 806.100 163.050 808.200 ;
        RECT 167.400 807.600 168.450 811.950 ;
        RECT 161.400 805.350 162.600 806.100 ;
        RECT 167.400 805.350 168.600 807.600 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 166.950 802.950 169.050 805.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 143.400 800.400 147.450 801.450 ;
        RECT 134.400 796.050 135.450 800.400 ;
        RECT 151.950 799.950 154.050 802.050 ;
        RECT 158.400 801.000 159.600 802.650 ;
        RECT 164.400 801.900 165.600 802.650 ;
        RECT 170.400 801.900 171.600 802.650 ;
        RECT 176.400 801.900 177.450 814.950 ;
        RECT 178.950 808.950 181.050 811.050 ;
        RECT 157.950 796.950 160.050 801.000 ;
        RECT 163.950 799.800 166.050 801.900 ;
        RECT 169.950 799.800 172.050 801.900 ;
        RECT 175.950 799.800 178.050 801.900 ;
        RECT 133.950 793.950 136.050 796.050 ;
        RECT 157.950 790.950 160.050 793.050 ;
        RECT 136.950 778.950 139.050 781.050 ;
        RECT 133.950 775.950 136.050 778.050 ;
        RECT 124.950 772.950 127.050 775.050 ;
        RECT 115.950 766.950 118.050 769.050 ;
        RECT 116.400 763.050 117.450 766.950 ;
        RECT 115.950 760.950 118.050 763.050 ;
        RECT 118.950 761.100 121.050 766.050 ;
        RECT 125.400 762.600 126.450 772.950 ;
        RECT 134.400 772.050 135.450 775.950 ;
        RECT 133.950 769.950 136.050 772.050 ;
        RECT 119.400 760.350 120.600 761.100 ;
        RECT 125.400 760.350 126.600 762.600 ;
        RECT 118.950 757.950 121.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 127.950 757.950 130.050 760.050 ;
        RECT 115.950 751.950 118.050 757.050 ;
        RECT 122.400 756.900 123.600 757.650 ;
        RECT 128.400 756.900 129.600 757.650 ;
        RECT 121.950 754.800 124.050 756.900 ;
        RECT 127.950 754.800 130.050 756.900 ;
        RECT 130.950 754.950 133.050 757.050 ;
        RECT 113.400 749.400 117.450 750.450 ;
        RECT 109.950 739.950 112.050 742.050 ;
        RECT 110.400 732.450 111.450 739.950 ;
        RECT 110.400 731.400 114.450 732.450 ;
        RECT 113.400 730.200 114.450 731.400 ;
        RECT 106.950 728.100 109.050 730.200 ;
        RECT 112.950 728.100 115.050 730.200 ;
        RECT 116.400 730.050 117.450 749.400 ;
        RECT 118.950 742.950 121.050 745.050 ;
        RECT 119.400 736.050 120.450 742.950 ;
        RECT 131.400 742.050 132.450 754.950 ;
        RECT 130.950 739.950 133.050 742.050 ;
        RECT 134.400 736.050 135.450 769.950 ;
        RECT 137.400 763.050 138.450 778.950 ;
        RECT 142.950 766.950 145.050 769.050 ;
        RECT 154.950 766.950 157.050 769.050 ;
        RECT 136.950 760.950 139.050 763.050 ;
        RECT 143.400 762.600 144.450 766.950 ;
        RECT 143.400 760.350 144.600 762.600 ;
        RECT 148.950 761.100 151.050 763.200 ;
        RECT 149.400 760.350 150.600 761.100 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 140.400 756.900 141.600 757.650 ;
        RECT 146.400 756.900 147.600 757.650 ;
        RECT 139.950 754.800 142.050 756.900 ;
        RECT 145.950 754.800 148.050 756.900 ;
        RECT 118.950 733.950 121.050 736.050 ;
        RECT 124.950 733.950 127.050 736.050 ;
        RECT 133.950 733.950 136.050 736.050 ;
        RECT 125.400 730.200 126.450 733.950 ;
        RECT 140.400 730.200 141.450 754.800 ;
        RECT 155.400 754.050 156.450 766.950 ;
        RECT 158.400 756.450 159.450 790.950 ;
        RECT 179.400 765.450 180.450 808.950 ;
        RECT 184.950 807.000 187.050 811.050 ;
        RECT 191.400 808.200 192.450 830.400 ;
        RECT 200.400 829.050 201.450 850.950 ;
        RECT 281.400 847.050 282.450 878.400 ;
        RECT 290.400 874.050 291.450 886.950 ;
        RECT 296.400 885.600 297.450 892.950 ;
        RECT 308.400 892.050 309.450 917.400 ;
        RECT 340.950 917.100 343.050 919.200 ;
        RECT 341.400 916.350 342.600 917.100 ;
        RECT 347.100 916.950 349.200 919.050 ;
        RECT 317.100 913.950 319.200 916.050 ;
        RECT 322.500 913.950 324.600 916.050 ;
        RECT 337.950 913.950 340.050 916.050 ;
        RECT 340.950 913.950 343.050 916.050 ;
        RECT 347.400 915.000 348.600 916.650 ;
        RECT 323.400 912.900 324.600 913.650 ;
        RECT 338.400 912.900 339.600 913.650 ;
        RECT 322.950 910.800 325.050 912.900 ;
        RECT 337.950 910.800 340.050 912.900 ;
        RECT 346.950 910.950 349.050 915.000 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 353.400 915.450 354.450 928.950 ;
        RECT 366.300 925.500 367.800 930.300 ;
        RECT 365.700 923.400 367.800 925.500 ;
        RECT 356.100 916.950 358.200 919.050 ;
        RECT 356.400 915.450 357.600 916.650 ;
        RECT 353.400 914.400 357.600 915.450 ;
        RECT 307.950 889.950 310.050 892.050 ;
        RECT 337.950 889.950 340.050 892.050 ;
        RECT 296.400 883.350 297.600 885.600 ;
        RECT 310.950 884.100 313.050 886.200 ;
        RECT 316.950 884.100 319.050 886.200 ;
        RECT 322.950 884.100 325.050 886.200 ;
        RECT 338.400 885.600 339.450 889.950 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 301.950 880.950 304.050 883.050 ;
        RECT 299.400 879.900 300.600 880.650 ;
        RECT 311.400 880.050 312.450 884.100 ;
        RECT 317.400 883.350 318.600 884.100 ;
        RECT 323.400 883.350 324.600 884.100 ;
        RECT 338.400 883.350 339.600 885.600 ;
        RECT 343.950 884.100 346.050 886.200 ;
        RECT 344.400 883.350 345.600 884.100 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 298.950 877.800 301.050 879.900 ;
        RECT 310.950 877.950 313.050 880.050 ;
        RECT 320.400 878.400 321.600 880.650 ;
        RECT 335.400 879.900 336.600 880.650 ;
        RECT 341.400 879.900 342.600 880.650 ;
        RECT 289.950 871.950 292.050 874.050 ;
        RECT 320.400 847.050 321.450 878.400 ;
        RECT 334.950 877.800 337.050 879.900 ;
        RECT 340.950 877.800 343.050 879.900 ;
        RECT 335.400 868.050 336.450 877.800 ;
        RECT 350.400 874.050 351.450 913.950 ;
        RECT 366.300 905.700 367.800 923.400 ;
        RECT 365.700 903.600 367.800 905.700 ;
        RECT 368.700 927.300 370.800 932.400 ;
        RECT 371.700 930.300 373.800 932.400 ;
        RECT 390.600 930.300 392.700 932.400 ;
        RECT 393.600 930.300 396.600 932.400 ;
        RECT 368.700 905.700 369.900 927.300 ;
        RECT 371.700 925.500 373.200 930.300 ;
        RECT 374.100 927.300 376.200 929.400 ;
        RECT 371.100 923.400 373.200 925.500 ;
        RECT 371.700 905.700 373.200 923.400 ;
        RECT 374.700 920.100 375.900 927.300 ;
        RECT 379.500 925.800 381.600 927.900 ;
        RECT 388.200 927.300 390.300 929.400 ;
        RECT 374.100 918.000 376.200 920.100 ;
        RECT 380.700 919.200 381.600 925.800 ;
        RECT 374.700 905.700 375.900 918.000 ;
        RECT 379.500 917.100 381.600 919.200 ;
        RECT 376.800 910.500 378.900 912.600 ;
        RECT 380.700 906.600 381.600 917.100 ;
        RECT 382.950 914.100 385.050 916.200 ;
        RECT 383.400 913.350 384.600 914.100 ;
        RECT 383.100 910.950 385.200 913.050 ;
        RECT 368.700 903.600 370.800 905.700 ;
        RECT 371.700 903.600 373.800 905.700 ;
        RECT 374.700 903.600 376.800 905.700 ;
        RECT 380.100 904.500 382.200 906.600 ;
        RECT 389.100 905.700 390.300 927.300 ;
        RECT 391.500 924.300 392.700 930.300 ;
        RECT 391.500 922.200 393.600 924.300 ;
        RECT 391.500 905.700 392.700 922.200 ;
        RECT 395.100 911.400 396.600 930.300 ;
        RECT 442.950 928.950 445.050 931.050 ;
        RECT 455.700 930.300 457.800 932.400 ;
        RECT 406.950 920.100 409.050 922.200 ;
        RECT 412.950 920.100 415.050 922.200 ;
        RECT 407.400 919.350 408.600 920.100 ;
        RECT 401.100 916.950 403.200 919.050 ;
        RECT 407.100 916.950 409.200 919.050 ;
        RECT 394.500 909.300 396.600 911.400 ;
        RECT 397.950 910.950 400.050 913.050 ;
        RECT 394.500 905.700 395.700 909.300 ;
        RECT 388.200 903.600 390.300 905.700 ;
        RECT 391.200 903.600 393.300 905.700 ;
        RECT 394.200 903.600 396.300 905.700 ;
        RECT 367.950 898.950 370.050 901.050 ;
        RECT 361.950 884.100 364.050 886.200 ;
        RECT 368.400 885.600 369.450 898.950 ;
        RECT 388.950 895.950 391.050 898.050 ;
        RECT 379.950 886.950 382.050 889.050 ;
        RECT 362.400 883.350 363.600 884.100 ;
        RECT 368.400 883.350 369.600 885.600 ;
        RECT 376.950 884.100 379.050 886.200 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 361.950 880.950 364.050 883.050 ;
        RECT 364.950 880.950 367.050 883.050 ;
        RECT 367.950 880.950 370.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 359.400 879.900 360.600 880.650 ;
        RECT 365.400 879.900 366.600 880.650 ;
        RECT 352.950 877.800 355.050 879.900 ;
        RECT 358.950 877.800 361.050 879.900 ;
        RECT 364.950 877.800 367.050 879.900 ;
        RECT 371.400 879.000 372.600 880.650 ;
        RECT 337.950 871.950 340.050 874.050 ;
        RECT 349.950 871.950 352.050 874.050 ;
        RECT 334.950 865.950 337.050 868.050 ;
        RECT 338.400 865.050 339.450 871.950 ;
        RECT 337.950 862.950 340.050 865.050 ;
        RECT 214.950 844.950 217.050 847.050 ;
        RECT 208.950 839.100 211.050 841.200 ;
        RECT 215.400 840.600 216.450 844.950 ;
        RECT 250.800 844.500 252.900 846.600 ;
        RECT 209.400 838.350 210.600 839.100 ;
        RECT 215.400 838.350 216.600 840.600 ;
        RECT 232.950 839.100 235.050 841.200 ;
        RECT 233.400 838.350 234.600 839.100 ;
        RECT 244.950 838.950 247.050 841.050 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 206.400 834.900 207.600 835.650 ;
        RECT 212.400 834.900 213.600 835.650 ;
        RECT 205.950 832.800 208.050 834.900 ;
        RECT 211.950 832.800 214.050 834.900 ;
        RECT 230.400 833.400 231.600 835.650 ;
        RECT 245.400 834.900 246.450 838.950 ;
        RECT 248.100 835.950 250.200 838.050 ;
        RECT 251.100 837.300 252.300 844.500 ;
        RECT 254.400 841.350 255.600 843.600 ;
        RECT 260.400 843.300 262.500 845.400 ;
        RECT 271.950 844.950 274.050 847.050 ;
        RECT 280.950 844.950 283.050 847.050 ;
        RECT 295.950 844.950 298.050 847.050 ;
        RECT 319.950 844.950 322.050 847.050 ;
        RECT 334.950 844.950 337.050 847.050 ;
        RECT 254.100 838.950 256.200 841.050 ;
        RECT 257.100 839.700 259.200 841.800 ;
        RECT 257.100 837.300 258.000 839.700 ;
        RECT 251.100 836.100 258.000 837.300 ;
        RECT 244.950 834.450 247.050 834.900 ;
        RECT 248.400 834.450 249.600 835.650 ;
        RECT 244.950 833.400 249.600 834.450 ;
        RECT 199.950 826.950 202.050 829.050 ;
        RECT 230.400 808.200 231.450 833.400 ;
        RECT 244.950 832.800 247.050 833.400 ;
        RECT 251.100 830.700 252.000 836.100 ;
        RECT 252.900 834.300 255.000 835.200 ;
        RECT 260.700 834.300 261.600 843.300 ;
        RECT 272.400 841.200 273.450 844.950 ;
        RECT 262.950 839.100 265.050 841.200 ;
        RECT 271.950 839.100 274.050 841.200 ;
        RECT 280.950 839.100 283.050 841.200 ;
        RECT 263.400 838.350 264.600 839.100 ;
        RECT 262.800 835.950 264.900 838.050 ;
        RECT 252.900 833.100 261.600 834.300 ;
        RECT 250.800 828.600 252.900 830.700 ;
        RECT 254.100 830.100 256.200 832.200 ;
        RECT 258.000 831.300 260.100 833.100 ;
        RECT 254.400 829.050 255.600 829.800 ;
        RECT 253.950 826.950 256.050 829.050 ;
        RECT 265.950 826.950 271.050 829.050 ;
        RECT 272.400 817.050 273.450 839.100 ;
        RECT 281.400 838.350 282.600 839.100 ;
        RECT 292.950 838.950 295.050 841.050 ;
        RECT 296.400 840.600 297.450 844.950 ;
        RECT 277.950 835.950 280.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 283.950 835.950 286.050 838.050 ;
        RECT 278.400 833.400 279.600 835.650 ;
        RECT 284.400 834.000 285.600 835.650 ;
        RECT 278.400 829.050 279.450 833.400 ;
        RECT 283.950 829.950 286.050 834.000 ;
        RECT 293.400 829.050 294.450 838.950 ;
        RECT 296.400 838.350 297.600 840.600 ;
        RECT 305.400 840.450 306.600 840.600 ;
        RECT 305.400 839.400 309.450 840.450 ;
        RECT 305.400 838.350 306.600 839.400 ;
        RECT 296.100 835.950 298.200 838.050 ;
        RECT 301.500 835.950 303.600 838.050 ;
        RECT 304.800 835.950 306.900 838.050 ;
        RECT 302.400 834.900 303.600 835.650 ;
        RECT 301.950 832.800 304.050 834.900 ;
        RECT 295.950 829.950 298.050 832.050 ;
        RECT 277.950 826.950 280.050 829.050 ;
        RECT 292.950 826.950 295.050 829.050 ;
        RECT 235.950 814.950 238.050 817.050 ;
        RECT 271.950 814.950 274.050 817.050 ;
        RECT 185.400 805.350 186.600 807.000 ;
        RECT 190.950 806.100 193.050 808.200 ;
        RECT 199.950 806.100 202.050 808.200 ;
        RECT 205.950 806.100 208.050 808.200 ;
        RECT 211.950 806.100 214.050 808.200 ;
        RECT 229.950 806.100 232.050 808.200 ;
        RECT 236.400 807.600 237.450 814.950 ;
        RECT 191.400 805.350 192.600 806.100 ;
        RECT 184.950 802.950 187.050 805.050 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 188.400 800.400 189.600 802.650 ;
        RECT 194.400 801.900 195.600 802.650 ;
        RECT 200.400 802.050 201.450 806.100 ;
        RECT 206.400 805.350 207.600 806.100 ;
        RECT 212.400 805.350 213.600 806.100 ;
        RECT 230.400 805.350 231.600 806.100 ;
        RECT 236.400 805.350 237.600 807.600 ;
        RECT 244.950 806.100 247.050 808.200 ;
        RECT 250.950 806.100 253.050 808.200 ;
        RECT 272.400 807.600 273.450 814.950 ;
        RECT 205.950 802.950 208.050 805.050 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 188.400 793.050 189.450 800.400 ;
        RECT 193.950 799.800 196.050 801.900 ;
        RECT 199.950 799.950 202.050 802.050 ;
        RECT 209.400 800.400 210.600 802.650 ;
        RECT 215.400 801.900 216.600 802.650 ;
        RECT 187.950 790.950 190.050 793.050 ;
        RECT 194.400 772.050 195.450 799.800 ;
        RECT 209.400 793.050 210.450 800.400 ;
        RECT 214.950 799.800 217.050 801.900 ;
        RECT 233.400 800.400 234.600 802.650 ;
        RECT 239.400 801.900 240.600 802.650 ;
        RECT 229.950 793.950 232.050 796.050 ;
        RECT 208.950 790.950 211.050 793.050 ;
        RECT 193.950 769.950 196.050 772.050 ;
        RECT 202.950 769.950 205.050 772.050 ;
        RECT 179.400 764.400 183.450 765.450 ;
        RECT 166.950 761.100 169.050 763.200 ;
        RECT 172.950 761.100 175.050 763.200 ;
        RECT 178.950 761.100 181.050 763.200 ;
        RECT 167.400 760.350 168.600 761.100 ;
        RECT 173.400 760.350 174.600 761.100 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 169.950 757.950 172.050 760.050 ;
        RECT 172.950 757.950 175.050 760.050 ;
        RECT 164.400 756.450 165.600 757.650 ;
        RECT 158.400 755.400 165.600 756.450 ;
        RECT 170.400 756.000 171.600 757.650 ;
        RECT 154.950 751.950 157.050 754.050 ;
        RECT 163.950 751.950 166.050 754.050 ;
        RECT 169.950 751.950 172.050 756.000 ;
        RECT 175.950 754.950 178.050 757.050 ;
        RECT 160.950 742.950 163.050 745.050 ;
        RECT 107.400 727.350 108.600 728.100 ;
        RECT 113.400 727.350 114.600 728.100 ;
        RECT 115.950 727.950 118.050 730.050 ;
        RECT 118.950 727.950 121.050 730.050 ;
        RECT 121.950 727.950 124.050 730.050 ;
        RECT 124.950 728.100 127.050 730.200 ;
        RECT 130.950 728.100 133.050 730.200 ;
        RECT 139.950 728.100 142.050 730.200 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 100.950 721.950 103.050 724.050 ;
        RECT 104.400 722.400 105.600 724.650 ;
        RECT 110.400 723.900 111.600 724.650 ;
        RECT 85.950 706.950 88.050 709.050 ;
        RECT 97.950 706.950 100.050 709.050 ;
        RECT 71.400 682.350 72.600 684.600 ;
        RECT 77.400 682.350 78.600 684.600 ;
        RECT 82.950 683.100 85.050 685.200 ;
        RECT 86.400 684.450 87.450 706.950 ;
        RECT 86.400 683.400 90.450 684.450 ;
        RECT 94.950 684.000 97.050 688.050 ;
        RECT 101.400 684.600 102.450 721.950 ;
        RECT 104.400 718.050 105.450 722.400 ;
        RECT 109.950 721.800 112.050 723.900 ;
        RECT 108.000 720.750 111.000 721.050 ;
        RECT 108.000 720.300 112.050 720.750 ;
        RECT 107.400 718.950 112.050 720.300 ;
        RECT 103.950 715.950 106.050 718.050 ;
        RECT 103.950 700.950 106.050 703.050 ;
        RECT 104.400 685.050 105.450 700.950 ;
        RECT 83.400 682.350 84.600 683.100 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 73.950 679.950 76.050 682.050 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 64.950 676.950 67.050 679.050 ;
        RECT 74.400 677.400 75.600 679.650 ;
        RECT 80.400 677.400 81.600 679.650 ;
        RECT 74.400 664.050 75.450 677.400 ;
        RECT 80.400 664.050 81.450 677.400 ;
        RECT 85.950 676.950 88.050 679.050 ;
        RECT 82.950 664.950 85.050 667.050 ;
        RECT 73.950 663.450 76.050 664.050 ;
        RECT 73.950 662.400 78.450 663.450 ;
        RECT 73.950 661.950 76.050 662.400 ;
        RECT 61.950 655.950 64.050 658.050 ;
        RECT 67.950 655.950 70.050 658.050 ;
        RECT 59.400 649.350 60.600 651.600 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 62.400 645.000 63.600 646.650 ;
        RECT 61.950 640.950 64.050 645.000 ;
        RECT 68.400 640.050 69.450 655.950 ;
        RECT 77.400 651.600 78.450 662.400 ;
        RECT 79.950 661.950 82.050 664.050 ;
        RECT 83.400 651.600 84.450 664.950 ;
        RECT 86.400 658.050 87.450 676.950 ;
        RECT 89.400 667.050 90.450 683.400 ;
        RECT 95.400 682.350 96.600 684.000 ;
        RECT 101.400 682.350 102.600 684.600 ;
        RECT 103.950 682.950 106.050 685.050 ;
        RECT 94.950 679.950 97.050 682.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 98.400 678.900 99.600 679.650 ;
        RECT 97.950 676.800 100.050 678.900 ;
        RECT 107.400 678.450 108.450 718.950 ;
        RECT 109.950 718.650 112.050 718.950 ;
        RECT 115.950 715.950 118.050 718.050 ;
        RECT 109.950 703.950 112.050 706.050 ;
        RECT 104.400 677.400 108.450 678.450 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 88.950 664.950 91.050 667.050 ;
        RECT 88.950 658.950 91.050 661.050 ;
        RECT 85.950 655.950 88.050 658.050 ;
        RECT 89.400 652.050 90.450 658.950 ;
        RECT 77.400 649.350 78.600 651.600 ;
        RECT 83.400 649.350 84.600 651.600 ;
        RECT 88.950 649.950 91.050 652.050 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 74.400 645.900 75.600 646.650 ;
        RECT 73.950 643.800 76.050 645.900 ;
        RECT 80.400 644.400 81.600 646.650 ;
        RECT 86.400 644.400 87.600 646.650 ;
        RECT 70.950 640.950 73.050 643.050 ;
        RECT 64.800 637.950 66.900 640.050 ;
        RECT 67.950 637.950 70.050 640.050 ;
        RECT 58.950 631.950 61.050 634.050 ;
        RECT 49.950 628.950 52.050 631.050 ;
        RECT 59.400 613.050 60.450 631.950 ;
        RECT 65.400 619.050 66.450 637.950 ;
        RECT 71.400 637.050 72.450 640.950 ;
        RECT 70.950 634.950 73.050 637.050 ;
        RECT 80.400 634.050 81.450 644.400 ;
        RECT 86.400 642.450 87.450 644.400 ;
        RECT 88.950 643.950 91.050 646.050 ;
        RECT 83.400 641.400 87.450 642.450 ;
        RECT 79.950 631.950 82.050 634.050 ;
        RECT 73.950 628.950 76.050 631.050 ;
        RECT 74.400 622.050 75.450 628.950 ;
        RECT 79.950 625.950 82.050 628.050 ;
        RECT 73.950 619.950 76.050 622.050 ;
        RECT 61.800 616.950 63.900 619.050 ;
        RECT 64.950 616.950 67.050 619.050 ;
        RECT 58.950 610.950 61.050 613.050 ;
        RECT 37.950 610.050 40.050 610.200 ;
        RECT 35.400 608.700 40.050 610.050 ;
        RECT 36.000 608.100 40.050 608.700 ;
        RECT 36.000 607.950 39.000 608.100 ;
        RECT 49.950 607.950 52.050 610.050 ;
        RECT 32.400 604.350 33.600 606.600 ;
        RECT 37.950 604.950 40.050 607.050 ;
        RECT 38.400 604.350 39.600 604.950 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 19.950 601.950 22.050 604.050 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 46.950 601.950 49.050 604.050 ;
        RECT 10.950 598.950 13.050 601.050 ;
        RECT 17.400 600.900 18.600 601.650 ;
        RECT 35.400 600.900 36.600 601.650 ;
        RECT 11.400 592.050 12.450 598.950 ;
        RECT 16.950 598.800 19.050 600.900 ;
        RECT 34.950 598.800 37.050 600.900 ;
        RECT 41.400 600.450 42.600 601.650 ;
        RECT 41.400 599.400 45.450 600.450 ;
        RECT 40.950 592.950 43.050 595.050 ;
        RECT 10.950 589.950 13.050 592.050 ;
        RECT 22.950 589.950 25.050 592.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 14.400 567.900 15.600 568.650 ;
        RECT 23.400 568.050 24.450 589.950 ;
        RECT 31.950 572.100 34.050 574.200 ;
        RECT 32.400 571.350 33.600 572.100 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 4.950 565.800 7.050 567.900 ;
        RECT 13.950 565.800 16.050 567.900 ;
        RECT 22.950 565.950 25.050 568.050 ;
        RECT 29.400 567.900 30.600 568.650 ;
        RECT 28.950 565.800 31.050 567.900 ;
        RECT 35.400 567.000 36.600 568.650 ;
        RECT 41.400 568.050 42.450 592.950 ;
        RECT 44.400 592.050 45.450 599.400 ;
        RECT 47.400 595.050 48.450 601.950 ;
        RECT 46.950 592.950 49.050 595.050 ;
        RECT 43.950 589.950 46.050 592.050 ;
        RECT 50.400 577.050 51.450 607.950 ;
        RECT 58.950 606.000 61.050 609.900 ;
        RECT 62.400 609.450 63.450 616.950 ;
        RECT 70.950 610.950 73.050 613.050 ;
        RECT 62.400 608.400 66.450 609.450 ;
        RECT 65.400 607.050 66.450 608.400 ;
        RECT 59.400 604.350 60.600 606.000 ;
        RECT 65.400 604.950 70.050 607.050 ;
        RECT 65.400 604.350 66.600 604.950 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 56.400 599.400 57.600 601.650 ;
        RECT 62.400 599.400 63.600 601.650 ;
        RECT 56.400 589.050 57.450 599.400 ;
        RECT 62.400 592.050 63.450 599.400 ;
        RECT 67.950 598.950 70.050 601.050 ;
        RECT 61.950 589.950 64.050 592.050 ;
        RECT 55.950 586.950 58.050 589.050 ;
        RECT 64.950 583.950 67.050 586.050 ;
        RECT 58.950 577.950 61.050 580.050 ;
        RECT 43.950 574.950 46.050 577.050 ;
        RECT 49.950 574.950 52.050 577.050 ;
        RECT 37.800 567.000 39.900 568.050 ;
        RECT 4.950 544.950 7.050 547.050 ;
        RECT 5.400 466.050 6.450 544.950 ;
        RECT 19.950 528.000 22.050 532.050 ;
        RECT 20.400 526.350 21.600 528.000 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 19.950 523.950 22.050 526.050 ;
        RECT 22.950 523.950 25.050 526.050 ;
        RECT 17.400 521.400 18.600 523.650 ;
        RECT 23.400 521.400 24.600 523.650 ;
        RECT 7.950 505.950 10.050 508.050 ;
        RECT 8.400 469.050 9.450 505.950 ;
        RECT 17.400 498.450 18.450 521.400 ;
        RECT 23.400 517.050 24.450 521.400 ;
        RECT 22.950 514.950 25.050 517.050 ;
        RECT 29.400 508.050 30.450 565.800 ;
        RECT 34.950 562.950 37.050 567.000 ;
        RECT 37.800 565.950 40.050 567.000 ;
        RECT 40.950 565.950 43.050 568.050 ;
        RECT 37.950 562.950 40.050 565.950 ;
        RECT 44.400 565.050 45.450 574.950 ;
        RECT 52.950 573.000 55.050 577.050 ;
        RECT 59.400 573.600 60.450 577.950 ;
        RECT 65.400 574.050 66.450 583.950 ;
        RECT 68.400 577.050 69.450 598.950 ;
        RECT 67.950 574.950 70.050 577.050 ;
        RECT 71.400 574.200 72.450 610.950 ;
        RECT 74.400 576.450 75.450 619.950 ;
        RECT 80.400 607.200 81.450 625.950 ;
        RECT 83.400 610.050 84.450 641.400 ;
        RECT 89.400 610.050 90.450 643.950 ;
        RECT 92.400 628.050 93.450 670.950 ;
        RECT 94.950 667.950 97.050 670.050 ;
        RECT 95.400 645.900 96.450 667.950 ;
        RECT 104.400 651.600 105.450 677.400 ;
        RECT 110.400 664.050 111.450 703.950 ;
        RECT 116.400 684.600 117.450 715.950 ;
        RECT 119.400 703.050 120.450 727.950 ;
        RECT 122.400 721.050 123.450 727.950 ;
        RECT 121.950 718.950 124.050 721.050 ;
        RECT 125.400 706.050 126.450 728.100 ;
        RECT 131.400 727.350 132.600 728.100 ;
        RECT 128.100 724.950 130.200 727.050 ;
        RECT 131.400 724.950 133.500 727.050 ;
        RECT 136.800 724.950 138.900 727.050 ;
        RECT 128.400 723.900 129.600 724.650 ;
        RECT 137.400 723.900 138.600 724.650 ;
        RECT 127.950 721.800 130.050 723.900 ;
        RECT 136.950 721.800 139.050 723.900 ;
        RECT 140.400 721.050 141.450 728.100 ;
        RECT 149.100 724.950 151.200 727.050 ;
        RECT 154.500 724.950 156.600 727.050 ;
        RECT 142.950 721.800 145.050 723.900 ;
        RECT 149.400 723.000 150.600 724.650 ;
        RECT 139.950 718.950 142.050 721.050 ;
        RECT 133.950 715.950 136.050 718.050 ;
        RECT 134.400 709.050 135.450 715.950 ;
        RECT 133.950 706.950 136.050 709.050 ;
        RECT 124.950 703.950 127.050 706.050 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 119.400 688.050 120.450 700.950 ;
        RECT 143.400 697.050 144.450 721.800 ;
        RECT 148.950 718.950 151.050 723.000 ;
        RECT 161.400 721.050 162.450 742.950 ;
        RECT 160.950 718.950 163.050 721.050 ;
        RECT 164.400 715.050 165.450 751.950 ;
        RECT 176.400 738.450 177.450 754.950 ;
        RECT 179.400 745.050 180.450 761.100 ;
        RECT 182.400 756.900 183.450 764.400 ;
        RECT 190.950 761.100 193.050 766.050 ;
        RECT 196.950 761.100 199.050 763.200 ;
        RECT 191.400 760.350 192.600 761.100 ;
        RECT 197.400 760.350 198.600 761.100 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 188.400 756.900 189.600 757.650 ;
        RECT 181.950 754.800 184.050 756.900 ;
        RECT 187.950 754.800 190.050 756.900 ;
        RECT 194.400 755.400 195.600 757.650 ;
        RECT 194.400 748.050 195.450 755.400 ;
        RECT 184.950 745.950 187.050 748.050 ;
        RECT 193.950 745.950 196.050 748.050 ;
        RECT 178.950 742.950 181.050 745.050 ;
        RECT 176.400 737.400 180.450 738.450 ;
        RECT 172.950 733.950 175.050 736.050 ;
        RECT 173.400 729.600 174.450 733.950 ;
        RECT 179.400 730.200 180.450 737.400 ;
        RECT 173.400 727.350 174.600 729.600 ;
        RECT 178.950 728.100 181.050 730.200 ;
        RECT 179.400 727.350 180.600 728.100 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 170.400 723.000 171.600 724.650 ;
        RECT 176.400 723.900 177.600 724.650 ;
        RECT 169.950 718.950 172.050 723.000 ;
        RECT 175.950 721.800 178.050 723.900 ;
        RECT 163.950 712.950 166.050 715.050 ;
        RECT 172.950 712.950 175.050 715.050 ;
        RECT 145.950 700.950 148.050 703.050 ;
        RECT 136.950 694.950 139.050 697.050 ;
        RECT 142.950 694.950 145.050 697.050 ;
        RECT 127.950 688.950 130.050 691.050 ;
        RECT 118.950 685.950 121.050 688.050 ;
        RECT 116.400 682.350 117.600 684.600 ;
        RECT 121.950 684.000 124.050 688.050 ;
        RECT 128.400 685.050 129.450 688.950 ;
        RECT 122.400 682.350 123.600 684.000 ;
        RECT 127.950 682.950 130.050 685.050 ;
        RECT 133.950 682.950 136.050 688.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 121.950 679.950 124.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 119.400 677.400 120.600 679.650 ;
        RECT 125.400 678.900 126.600 679.650 ;
        RECT 109.950 661.950 112.050 664.050 ;
        RECT 119.400 658.050 120.450 677.400 ;
        RECT 124.950 676.800 127.050 678.900 ;
        RECT 112.950 655.950 115.050 658.050 ;
        RECT 118.950 655.950 121.050 658.050 ;
        RECT 121.950 655.950 124.050 658.050 ;
        RECT 104.400 649.350 105.600 651.600 ;
        RECT 110.400 651.450 111.600 651.600 ;
        RECT 113.400 651.450 114.450 655.950 ;
        RECT 115.950 652.950 118.050 655.050 ;
        RECT 110.400 650.400 114.450 651.450 ;
        RECT 110.400 649.350 111.600 650.400 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 101.400 645.900 102.600 646.650 ;
        RECT 94.950 643.800 97.050 645.900 ;
        RECT 100.950 643.800 103.050 645.900 ;
        RECT 107.400 644.400 108.600 646.650 ;
        RECT 116.400 645.900 117.450 652.950 ;
        RECT 122.400 651.450 123.450 655.950 ;
        RECT 125.400 655.050 126.450 676.800 ;
        RECT 124.950 652.950 127.050 655.050 ;
        RECT 119.400 650.400 123.450 651.450 ;
        RECT 127.950 651.000 130.050 655.050 ;
        RECT 134.400 652.050 135.450 682.950 ;
        RECT 107.400 634.050 108.450 644.400 ;
        RECT 115.950 643.800 118.050 645.900 ;
        RECT 106.950 631.950 109.050 634.050 ;
        RECT 115.950 633.450 118.050 634.050 ;
        RECT 119.400 633.450 120.450 650.400 ;
        RECT 128.400 649.350 129.600 651.000 ;
        RECT 133.950 649.950 136.050 652.050 ;
        RECT 137.400 649.050 138.450 694.950 ;
        RECT 146.400 688.050 147.450 700.950 ;
        RECT 148.950 694.950 151.050 697.050 ;
        RECT 145.950 685.950 148.050 688.050 ;
        RECT 139.950 683.100 142.050 685.200 ;
        RECT 149.400 684.600 150.450 694.950 ;
        RECT 154.950 685.950 157.050 688.050 ;
        RECT 140.400 682.350 141.600 683.100 ;
        RECT 149.400 682.350 150.600 684.600 ;
        RECT 140.100 679.950 142.200 682.050 ;
        RECT 143.400 679.950 145.500 682.050 ;
        RECT 148.800 679.950 150.900 682.050 ;
        RECT 143.400 677.400 144.600 679.650 ;
        RECT 143.400 667.050 144.450 677.400 ;
        RECT 142.950 664.950 145.050 667.050 ;
        RECT 148.950 658.950 151.050 661.050 ;
        RECT 149.400 655.050 150.450 658.950 ;
        RECT 139.950 652.950 142.050 655.050 ;
        RECT 148.950 652.950 151.050 655.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 130.950 646.950 133.050 649.050 ;
        RECT 136.950 646.950 139.050 649.050 ;
        RECT 125.400 645.900 126.600 646.650 ;
        RECT 131.400 645.900 132.600 646.650 ;
        RECT 124.950 643.800 127.050 645.900 ;
        RECT 130.950 643.800 133.050 645.900 ;
        RECT 127.950 637.950 130.050 640.050 ;
        RECT 115.950 632.400 120.450 633.450 ;
        RECT 115.950 631.950 118.050 632.400 ;
        RECT 91.950 625.950 94.050 628.050 ;
        RECT 106.950 616.950 109.050 619.050 ;
        RECT 94.950 610.950 97.050 613.050 ;
        RECT 82.950 607.950 85.050 610.050 ;
        RECT 88.950 607.950 91.050 610.050 ;
        RECT 79.950 605.100 82.050 607.200 ;
        RECT 80.400 604.350 81.600 605.100 ;
        RECT 88.950 604.800 91.050 606.900 ;
        RECT 95.400 606.600 96.450 610.950 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 76.950 598.950 79.050 601.050 ;
        RECT 83.400 600.000 84.600 601.650 ;
        RECT 77.400 589.050 78.450 598.950 ;
        RECT 82.950 595.950 85.050 600.000 ;
        RECT 85.950 598.950 88.050 601.050 ;
        RECT 86.400 594.450 87.450 598.950 ;
        RECT 83.400 593.400 87.450 594.450 ;
        RECT 76.950 586.950 79.050 589.050 ;
        RECT 83.400 580.050 84.450 593.400 ;
        RECT 89.400 586.050 90.450 604.800 ;
        RECT 95.400 604.350 96.600 606.600 ;
        RECT 100.950 605.100 103.050 607.200 ;
        RECT 107.400 607.050 108.450 616.950 ;
        RECT 116.400 610.050 117.450 631.950 ;
        RECT 124.950 625.950 127.050 628.050 ;
        RECT 121.950 622.950 124.050 625.050 ;
        RECT 122.400 619.050 123.450 622.950 ;
        RECT 121.950 616.950 124.050 619.050 ;
        RECT 115.950 607.950 118.050 610.050 ;
        RECT 101.400 604.350 102.600 605.100 ;
        RECT 106.950 604.950 109.050 607.050 ;
        RECT 118.950 605.100 121.050 607.200 ;
        RECT 119.400 604.350 120.600 605.100 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 98.400 599.400 99.600 601.650 ;
        RECT 104.400 599.400 105.600 601.650 ;
        RECT 91.950 595.950 94.050 598.050 ;
        RECT 92.400 586.050 93.450 595.950 ;
        RECT 88.800 583.950 90.900 586.050 ;
        RECT 91.950 583.950 94.050 586.050 ;
        RECT 98.400 583.050 99.450 599.400 ;
        RECT 100.950 595.950 103.050 598.050 ;
        RECT 85.950 580.950 88.050 583.050 ;
        RECT 97.950 580.950 100.050 583.050 ;
        RECT 82.950 577.950 85.050 580.050 ;
        RECT 76.950 576.450 79.050 577.050 ;
        RECT 74.400 575.400 79.050 576.450 ;
        RECT 53.400 571.350 54.600 573.000 ;
        RECT 59.400 571.350 60.600 573.600 ;
        RECT 64.800 571.950 66.900 574.050 ;
        RECT 70.950 573.450 73.050 574.200 ;
        RECT 68.400 572.400 73.050 573.450 ;
        RECT 76.950 573.000 79.050 575.400 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 50.400 567.000 51.600 568.650 ;
        RECT 56.400 567.900 57.600 568.650 ;
        RECT 62.400 567.900 63.600 568.650 ;
        RECT 43.950 562.950 46.050 565.050 ;
        RECT 49.950 562.950 52.050 567.000 ;
        RECT 55.950 565.800 58.050 567.900 ;
        RECT 61.950 565.800 64.050 567.900 ;
        RECT 64.950 565.950 67.050 568.050 ;
        RECT 62.400 559.050 63.450 565.800 ;
        RECT 61.950 556.950 64.050 559.050 ;
        RECT 65.400 547.050 66.450 565.950 ;
        RECT 64.950 544.950 67.050 547.050 ;
        RECT 46.950 541.950 49.050 544.050 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 37.950 527.100 40.050 529.200 ;
        RECT 32.400 517.050 33.450 526.950 ;
        RECT 38.400 526.350 39.600 527.100 ;
        RECT 37.950 523.950 40.050 526.050 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 41.400 522.000 42.600 523.650 ;
        RECT 40.950 517.950 43.050 522.000 ;
        RECT 31.950 514.950 34.050 517.050 ;
        RECT 28.950 505.950 31.050 508.050 ;
        RECT 32.400 499.200 33.450 514.950 ;
        RECT 47.400 514.050 48.450 541.950 ;
        RECT 49.950 538.950 52.050 541.050 ;
        RECT 46.950 511.950 49.050 514.050 ;
        RECT 37.950 502.950 40.050 505.050 ;
        RECT 14.400 497.400 18.450 498.450 ;
        RECT 14.400 495.600 15.450 497.400 ;
        RECT 31.950 497.100 34.050 499.200 ;
        RECT 14.400 493.350 15.600 495.600 ;
        RECT 25.950 493.950 28.050 496.050 ;
        RECT 31.950 493.950 34.050 496.050 ;
        RECT 38.400 495.600 39.450 502.950 ;
        RECT 46.950 496.950 49.050 499.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 17.400 488.400 18.600 490.650 ;
        RECT 17.400 481.050 18.450 488.400 ;
        RECT 16.950 478.950 19.050 481.050 ;
        RECT 7.950 466.950 10.050 469.050 ;
        RECT 4.950 463.950 7.050 466.050 ;
        RECT 19.950 463.950 22.050 466.050 ;
        RECT 4.950 457.950 7.050 460.050 ;
        RECT 5.400 391.050 6.450 457.950 ;
        RECT 13.950 450.000 16.050 454.050 ;
        RECT 20.400 451.200 21.450 463.950 ;
        RECT 26.400 454.050 27.450 493.950 ;
        RECT 32.400 493.350 33.600 493.950 ;
        RECT 38.400 493.350 39.600 495.600 ;
        RECT 31.950 490.950 34.050 493.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 35.400 489.000 36.600 490.650 ;
        RECT 41.400 490.050 42.600 490.650 ;
        RECT 34.950 484.950 37.050 489.000 ;
        RECT 41.400 488.400 46.050 490.050 ;
        RECT 42.000 487.950 46.050 488.400 ;
        RECT 47.400 487.050 48.450 496.950 ;
        RECT 46.950 484.950 49.050 487.050 ;
        RECT 46.950 481.800 49.050 483.900 ;
        RECT 40.950 457.950 43.050 460.050 ;
        RECT 41.400 454.050 42.450 457.950 ;
        RECT 25.950 451.950 28.050 454.050 ;
        RECT 14.400 448.350 15.600 450.000 ;
        RECT 19.950 449.100 22.050 451.200 ;
        RECT 20.400 448.350 21.600 449.100 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 17.400 444.900 18.600 445.650 ;
        RECT 26.400 445.050 27.450 451.950 ;
        RECT 28.950 449.100 31.050 451.200 ;
        RECT 34.950 449.100 37.050 451.200 ;
        RECT 40.950 450.000 43.050 454.050 ;
        RECT 29.400 445.050 30.450 449.100 ;
        RECT 35.400 448.350 36.600 449.100 ;
        RECT 41.400 448.350 42.600 450.000 ;
        RECT 34.950 445.950 37.050 448.050 ;
        RECT 37.950 445.950 40.050 448.050 ;
        RECT 40.950 445.950 43.050 448.050 ;
        RECT 16.950 442.800 19.050 444.900 ;
        RECT 25.950 442.950 28.050 445.050 ;
        RECT 28.950 442.950 31.050 445.050 ;
        RECT 31.950 442.950 34.050 445.050 ;
        RECT 38.400 443.400 39.600 445.650 ;
        RECT 47.400 445.050 48.450 481.800 ;
        RECT 50.400 454.050 51.450 538.950 ;
        RECT 68.400 538.050 69.450 572.400 ;
        RECT 70.950 572.100 73.050 572.400 ;
        RECT 77.400 571.350 78.600 573.000 ;
        RECT 82.950 571.950 85.050 576.900 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 80.400 566.400 81.600 568.650 ;
        RECT 86.400 567.900 87.450 580.950 ;
        RECT 88.950 577.950 91.050 580.050 ;
        RECT 80.400 556.050 81.450 566.400 ;
        RECT 85.950 565.800 88.050 567.900 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 73.950 544.950 76.050 547.050 ;
        RECT 67.950 535.950 70.050 538.050 ;
        RECT 64.950 529.950 67.050 532.050 ;
        RECT 55.950 527.100 58.050 529.200 ;
        RECT 56.400 526.350 57.600 527.100 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 52.950 520.950 55.050 523.050 ;
        RECT 59.400 522.450 60.600 523.650 ;
        RECT 59.400 521.400 63.450 522.450 ;
        RECT 53.400 496.050 54.450 520.950 ;
        RECT 58.950 514.950 61.050 520.050 ;
        RECT 62.400 517.050 63.450 521.400 ;
        RECT 61.950 514.950 64.050 517.050 ;
        RECT 52.950 493.950 55.050 496.050 ;
        RECT 58.950 494.100 61.050 496.200 ;
        RECT 65.400 496.050 66.450 529.950 ;
        RECT 68.400 520.050 69.450 535.950 ;
        RECT 74.400 532.050 75.450 544.950 ;
        RECT 79.950 535.950 82.050 538.050 ;
        RECT 80.400 532.050 81.450 535.950 ;
        RECT 73.950 529.950 76.050 532.050 ;
        RECT 79.950 529.950 82.050 532.050 ;
        RECT 74.400 528.600 75.450 529.950 ;
        RECT 80.400 528.600 81.450 529.950 ;
        RECT 74.400 526.350 75.600 528.600 ;
        RECT 80.400 526.350 81.600 528.600 ;
        RECT 86.400 528.450 87.450 565.800 ;
        RECT 89.400 559.050 90.450 577.950 ;
        RECT 94.950 572.100 97.050 574.200 ;
        RECT 101.400 573.600 102.450 595.950 ;
        RECT 104.400 595.050 105.450 599.400 ;
        RECT 109.950 598.950 112.050 601.050 ;
        RECT 116.400 599.400 117.600 601.650 ;
        RECT 103.950 592.950 106.050 595.050 ;
        RECT 106.950 586.950 109.050 589.050 ;
        RECT 107.400 580.050 108.450 586.950 ;
        RECT 106.950 577.950 109.050 580.050 ;
        RECT 95.400 571.350 96.600 572.100 ;
        RECT 101.400 571.350 102.600 573.600 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 91.950 565.950 94.050 568.050 ;
        RECT 98.400 567.900 99.600 568.650 ;
        RECT 88.950 556.950 91.050 559.050 ;
        RECT 92.400 535.050 93.450 565.950 ;
        RECT 97.950 565.800 100.050 567.900 ;
        RECT 104.400 567.450 105.600 568.650 ;
        RECT 110.400 567.450 111.450 598.950 ;
        RECT 112.950 595.950 115.050 598.050 ;
        RECT 113.400 574.050 114.450 595.950 ;
        RECT 116.400 595.050 117.450 599.400 ;
        RECT 125.400 595.050 126.450 625.950 ;
        RECT 128.400 598.050 129.450 637.950 ;
        RECT 140.400 634.050 141.450 652.950 ;
        RECT 142.950 649.950 145.050 652.050 ;
        RECT 143.400 645.900 144.450 649.950 ;
        RECT 146.100 646.950 148.200 649.050 ;
        RECT 151.500 646.950 153.600 649.050 ;
        RECT 142.950 643.800 145.050 645.900 ;
        RECT 146.400 644.400 147.600 646.650 ;
        RECT 139.950 631.950 142.050 634.050 ;
        RECT 136.950 622.950 139.050 625.050 ;
        RECT 137.400 609.450 138.450 622.950 ;
        RECT 146.400 613.050 147.450 644.400 ;
        RECT 148.950 637.950 151.050 640.050 ;
        RECT 145.950 610.950 148.050 613.050 ;
        RECT 137.400 608.400 141.450 609.450 ;
        RECT 133.950 605.100 136.050 607.200 ;
        RECT 140.400 606.600 141.450 608.400 ;
        RECT 134.400 604.350 135.600 605.100 ;
        RECT 140.400 604.350 141.600 606.600 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 137.400 600.900 138.600 601.650 ;
        RECT 143.400 600.900 144.600 601.650 ;
        RECT 136.950 598.800 139.050 600.900 ;
        RECT 142.950 598.800 145.050 600.900 ;
        RECT 127.950 595.950 130.050 598.050 ;
        RECT 115.950 592.950 118.050 595.050 ;
        RECT 124.950 592.950 127.050 595.050 ;
        RECT 115.950 580.950 118.050 583.050 ;
        RECT 112.950 571.950 115.050 574.050 ;
        RECT 116.400 573.600 117.450 580.950 ;
        RECT 143.400 574.050 144.450 598.800 ;
        RECT 149.400 591.450 150.450 637.950 ;
        RECT 155.400 637.050 156.450 685.950 ;
        RECT 163.950 683.100 166.050 685.200 ;
        RECT 169.950 683.100 172.050 685.200 ;
        RECT 164.400 682.350 165.600 683.100 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 676.950 169.050 679.050 ;
        RECT 163.950 664.950 166.050 667.050 ;
        RECT 164.400 652.050 165.450 664.950 ;
        RECT 167.400 658.050 168.450 676.950 ;
        RECT 170.400 676.050 171.450 683.100 ;
        RECT 169.950 673.950 172.050 676.050 ;
        RECT 169.950 660.450 172.050 661.050 ;
        RECT 173.400 660.450 174.450 712.950 ;
        RECT 176.400 703.050 177.450 721.800 ;
        RECT 178.950 706.950 181.050 709.050 ;
        RECT 175.950 700.950 178.050 703.050 ;
        RECT 179.400 700.050 180.450 706.950 ;
        RECT 185.400 706.050 186.450 745.950 ;
        RECT 190.950 742.950 193.050 745.050 ;
        RECT 191.400 729.600 192.450 742.950 ;
        RECT 191.400 727.350 192.600 729.600 ;
        RECT 196.950 728.100 199.050 730.200 ;
        RECT 203.400 730.050 204.450 769.950 ;
        RECT 205.950 761.100 208.050 763.200 ;
        RECT 214.950 762.000 217.050 766.050 ;
        RECT 206.400 757.050 207.450 761.100 ;
        RECT 215.400 760.350 216.600 762.000 ;
        RECT 220.950 761.100 223.050 763.200 ;
        RECT 226.950 761.100 229.050 763.200 ;
        RECT 221.400 760.350 222.600 761.100 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 220.950 757.950 223.050 760.050 ;
        RECT 205.950 754.950 208.050 757.050 ;
        RECT 212.400 756.900 213.600 757.650 ;
        RECT 211.950 754.800 214.050 756.900 ;
        RECT 218.400 755.400 219.600 757.650 ;
        RECT 208.950 739.950 211.050 742.050 ;
        RECT 205.950 733.950 208.050 736.050 ;
        RECT 197.400 727.350 198.600 728.100 ;
        RECT 202.950 727.950 205.050 730.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 194.400 723.000 195.600 724.650 ;
        RECT 193.950 718.950 196.050 723.000 ;
        RECT 200.400 722.400 201.600 724.650 ;
        RECT 200.400 718.050 201.450 722.400 ;
        RECT 202.950 721.950 205.050 724.050 ;
        RECT 199.950 715.950 202.050 718.050 ;
        RECT 187.950 712.950 190.050 715.050 ;
        RECT 184.950 703.950 187.050 706.050 ;
        RECT 188.400 700.050 189.450 712.950 ;
        RECT 200.400 709.050 201.450 715.950 ;
        RECT 199.950 706.950 202.050 709.050 ;
        RECT 178.950 697.950 181.050 700.050 ;
        RECT 187.950 697.950 190.050 700.050 ;
        RECT 189.000 696.900 192.000 697.050 ;
        RECT 187.950 694.950 193.050 696.900 ;
        RECT 196.950 694.950 199.050 700.050 ;
        RECT 187.950 694.800 190.050 694.950 ;
        RECT 190.950 694.800 193.050 694.950 ;
        RECT 196.950 691.800 199.050 693.900 ;
        RECT 178.950 688.950 181.050 691.050 ;
        RECT 190.950 688.950 193.050 691.050 ;
        RECT 179.400 684.600 180.450 688.950 ;
        RECT 179.400 682.350 180.600 684.600 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 182.400 677.400 183.600 679.650 ;
        RECT 178.950 673.950 181.050 676.050 ;
        RECT 175.950 667.950 178.050 670.050 ;
        RECT 169.950 659.400 174.450 660.450 ;
        RECT 169.950 658.950 172.050 659.400 ;
        RECT 166.950 655.950 169.050 658.050 ;
        RECT 160.950 649.950 163.050 652.050 ;
        RECT 163.950 649.950 166.050 652.050 ;
        RECT 170.400 651.600 171.450 658.950 ;
        RECT 176.400 651.600 177.450 667.950 ;
        RECT 179.400 664.050 180.450 673.950 ;
        RECT 178.950 661.950 181.050 664.050 ;
        RECT 182.400 658.050 183.450 677.400 ;
        RECT 184.950 673.950 187.050 676.050 ;
        RECT 181.950 655.950 184.050 658.050 ;
        RECT 185.400 652.050 186.450 673.950 ;
        RECT 187.950 655.950 190.050 658.050 ;
        RECT 154.950 634.950 157.050 637.050 ;
        RECT 151.950 610.950 154.050 613.050 ;
        RECT 152.400 607.050 153.450 610.950 ;
        RECT 161.400 607.200 162.450 649.950 ;
        RECT 170.400 649.350 171.600 651.600 ;
        RECT 176.400 649.350 177.600 651.600 ;
        RECT 184.950 649.950 187.050 652.050 ;
        RECT 166.950 646.950 169.050 649.050 ;
        RECT 169.950 646.950 172.050 649.050 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 163.950 643.950 166.050 646.050 ;
        RECT 167.400 644.400 168.600 646.650 ;
        RECT 173.400 645.900 174.600 646.650 ;
        RECT 164.400 637.050 165.450 643.950 ;
        RECT 163.950 634.950 166.050 637.050 ;
        RECT 167.400 634.050 168.450 644.400 ;
        RECT 172.950 643.800 175.050 645.900 ;
        RECT 179.400 645.450 180.600 646.650 ;
        RECT 184.950 645.450 187.050 648.900 ;
        RECT 179.400 645.000 187.050 645.450 ;
        RECT 179.400 644.400 186.450 645.000 ;
        RECT 188.400 643.050 189.450 655.950 ;
        RECT 191.400 652.050 192.450 688.950 ;
        RECT 193.950 685.950 196.050 688.050 ;
        RECT 194.400 678.450 195.450 685.950 ;
        RECT 197.400 685.050 198.450 691.800 ;
        RECT 203.400 688.050 204.450 721.950 ;
        RECT 206.400 721.050 207.450 733.950 ;
        RECT 209.400 723.450 210.450 739.950 ;
        RECT 212.400 733.050 213.450 754.800 ;
        RECT 218.400 751.050 219.450 755.400 ;
        RECT 217.950 748.950 220.050 751.050 ;
        RECT 227.400 748.050 228.450 761.100 ;
        RECT 226.950 745.950 229.050 748.050 ;
        RECT 230.400 742.050 231.450 793.950 ;
        RECT 233.400 775.050 234.450 800.400 ;
        RECT 238.950 799.800 241.050 801.900 ;
        RECT 232.950 772.950 235.050 775.050 ;
        RECT 245.400 769.050 246.450 806.100 ;
        RECT 251.400 805.350 252.600 806.100 ;
        RECT 272.400 805.350 273.600 807.600 ;
        RECT 277.950 806.100 280.050 808.200 ;
        RECT 296.400 807.600 297.450 829.950 ;
        RECT 308.400 829.050 309.450 839.400 ;
        RECT 319.950 839.100 322.050 841.200 ;
        RECT 325.800 839.100 327.900 841.200 ;
        RECT 320.400 838.350 321.600 839.100 ;
        RECT 326.400 838.350 327.600 839.100 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 323.400 833.400 324.600 835.650 ;
        RECT 307.950 826.950 310.050 829.050 ;
        RECT 323.400 823.050 324.450 833.400 ;
        RECT 322.950 820.950 325.050 823.050 ;
        RECT 335.400 820.050 336.450 844.950 ;
        RECT 343.950 839.100 346.050 841.200 ;
        RECT 344.400 838.350 345.600 839.100 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 341.400 833.400 342.600 835.650 ;
        RECT 337.950 829.950 340.050 832.050 ;
        RECT 334.950 817.950 337.050 820.050 ;
        RECT 334.950 814.800 337.050 816.900 ;
        RECT 322.950 811.950 325.050 814.050 ;
        RECT 278.400 805.350 279.600 806.100 ;
        RECT 296.400 805.350 297.600 807.600 ;
        RECT 313.950 806.100 316.050 808.200 ;
        RECT 314.400 805.350 315.600 806.100 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 277.950 802.950 280.050 805.050 ;
        RECT 292.950 802.950 295.050 805.050 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 298.950 802.950 301.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 313.950 802.950 316.050 805.050 ;
        RECT 316.950 802.950 319.050 805.050 ;
        RECT 254.400 801.900 255.600 802.650 ;
        RECT 269.400 801.900 270.600 802.650 ;
        RECT 253.950 799.800 256.050 801.900 ;
        RECT 268.950 799.800 271.050 801.900 ;
        RECT 275.400 800.400 276.600 802.650 ;
        RECT 293.400 800.400 294.600 802.650 ;
        RECT 299.400 800.400 300.600 802.650 ;
        RECT 311.400 800.400 312.600 802.650 ;
        RECT 262.950 790.950 265.050 793.050 ;
        RECT 250.950 787.950 253.050 790.050 ;
        RECT 244.950 766.950 247.050 769.050 ;
        RECT 235.950 761.100 238.050 763.200 ;
        RECT 241.950 761.100 244.050 763.200 ;
        RECT 236.400 760.350 237.600 761.100 ;
        RECT 242.400 760.350 243.600 761.100 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 239.400 756.900 240.600 757.650 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 245.400 755.400 246.600 757.650 ;
        RECT 245.400 751.050 246.450 755.400 ;
        RECT 244.950 748.950 247.050 751.050 ;
        RECT 245.400 745.050 246.450 748.950 ;
        RECT 244.950 742.950 247.050 745.050 ;
        RECT 229.950 739.950 232.050 742.050 ;
        RECT 223.950 735.450 226.050 736.050 ;
        RECT 218.400 734.400 226.050 735.450 ;
        RECT 211.950 730.950 214.050 733.050 ;
        RECT 218.400 732.450 219.450 734.400 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 238.950 733.950 241.050 736.050 ;
        RECT 215.400 731.400 219.450 732.450 ;
        RECT 215.400 729.600 216.450 731.400 ;
        RECT 215.400 727.350 216.600 729.600 ;
        RECT 220.950 729.000 223.050 733.050 ;
        RECT 221.400 727.350 222.600 729.000 ;
        RECT 229.950 728.100 232.050 730.200 ;
        RECT 239.400 729.600 240.450 733.950 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 220.950 724.950 223.050 727.050 ;
        RECT 223.950 724.950 226.050 727.050 ;
        RECT 209.400 722.400 213.450 723.450 ;
        RECT 205.950 718.950 208.050 721.050 ;
        RECT 212.400 720.450 213.450 722.400 ;
        RECT 218.400 722.400 219.600 724.650 ;
        RECT 224.400 722.400 225.600 724.650 ;
        RECT 212.400 719.400 216.450 720.450 ;
        RECT 202.950 685.950 205.050 688.050 ;
        RECT 196.950 682.950 199.050 685.050 ;
        RECT 199.950 683.100 202.050 685.200 ;
        RECT 205.950 683.100 208.050 685.200 ;
        RECT 211.950 683.100 214.050 685.200 ;
        RECT 215.400 685.050 216.450 719.400 ;
        RECT 218.400 691.050 219.450 722.400 ;
        RECT 224.400 720.450 225.450 722.400 ;
        RECT 226.950 721.800 229.050 723.900 ;
        RECT 221.400 719.400 225.450 720.450 ;
        RECT 217.950 688.950 220.050 691.050 ;
        RECT 200.400 682.350 201.600 683.100 ;
        RECT 206.400 682.350 207.600 683.100 ;
        RECT 212.400 682.350 213.600 683.100 ;
        RECT 214.950 682.950 217.050 685.050 ;
        RECT 217.950 683.100 220.050 685.200 ;
        RECT 199.950 679.950 202.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 194.400 677.400 198.450 678.450 ;
        RECT 190.950 649.950 193.050 652.050 ;
        RECT 197.400 651.600 198.450 677.400 ;
        RECT 203.400 677.400 204.600 679.650 ;
        RECT 209.400 677.400 210.600 679.650 ;
        RECT 203.400 667.050 204.450 677.400 ;
        RECT 209.400 670.050 210.450 677.400 ;
        RECT 211.950 673.950 214.050 676.050 ;
        RECT 208.950 667.950 211.050 670.050 ;
        RECT 202.950 664.950 205.050 667.050 ;
        RECT 197.400 649.350 198.600 651.600 ;
        RECT 202.950 650.100 205.050 652.200 ;
        RECT 203.400 649.350 204.600 650.100 ;
        RECT 193.950 646.950 196.050 649.050 ;
        RECT 196.950 646.950 199.050 649.050 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 194.400 645.000 195.600 646.650 ;
        RECT 200.400 645.900 201.600 646.650 ;
        RECT 187.950 640.950 190.050 643.050 ;
        RECT 193.950 640.950 196.050 645.000 ;
        RECT 199.950 643.800 202.050 645.900 ;
        RECT 166.950 631.950 169.050 634.050 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 205.950 625.950 208.050 628.050 ;
        RECT 184.950 619.950 187.050 622.050 ;
        RECT 151.950 604.950 154.050 607.050 ;
        RECT 160.950 605.100 163.050 607.200 ;
        RECT 166.950 605.100 169.050 607.200 ;
        RECT 161.400 604.350 162.600 605.100 ;
        RECT 154.950 601.950 157.050 604.050 ;
        RECT 157.950 601.950 160.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 158.400 600.900 159.600 601.650 ;
        RECT 167.400 601.050 168.450 605.100 ;
        RECT 169.950 604.950 172.050 610.050 ;
        RECT 172.950 605.100 175.050 607.200 ;
        RECT 178.950 606.000 181.050 610.050 ;
        RECT 185.400 607.050 186.450 619.950 ;
        RECT 173.400 604.350 174.600 605.100 ;
        RECT 179.400 604.350 180.600 606.000 ;
        RECT 184.950 604.950 187.050 607.050 ;
        RECT 190.950 605.100 193.050 607.200 ;
        RECT 200.400 606.600 201.450 625.950 ;
        RECT 206.400 613.050 207.450 625.950 ;
        RECT 209.400 625.050 210.450 667.950 ;
        RECT 208.950 622.950 211.050 625.050 ;
        RECT 212.400 622.050 213.450 673.950 ;
        RECT 218.400 673.050 219.450 683.100 ;
        RECT 221.400 679.050 222.450 719.400 ;
        RECT 227.400 715.050 228.450 721.800 ;
        RECT 230.400 715.050 231.450 728.100 ;
        RECT 239.400 727.350 240.600 729.600 ;
        RECT 244.950 728.100 247.050 730.200 ;
        RECT 245.400 727.350 246.600 728.100 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 241.950 724.950 244.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 236.400 723.900 237.600 724.650 ;
        RECT 235.950 721.800 238.050 723.900 ;
        RECT 242.400 722.400 243.600 724.650 ;
        RECT 236.400 720.450 237.450 721.800 ;
        RECT 242.400 720.450 243.450 722.400 ;
        RECT 236.400 719.400 240.450 720.450 ;
        RECT 242.400 719.400 246.450 720.450 ;
        RECT 235.950 715.950 238.050 718.050 ;
        RECT 226.800 712.950 228.900 715.050 ;
        RECT 229.950 712.950 232.050 715.050 ;
        RECT 230.400 694.050 231.450 712.950 ;
        RECT 236.400 706.050 237.450 715.950 ;
        RECT 235.950 703.950 238.050 706.050 ;
        RECT 229.950 691.950 232.050 694.050 ;
        RECT 226.950 683.100 229.050 685.200 ;
        RECT 227.400 682.350 228.600 683.100 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 220.950 676.950 223.050 679.050 ;
        RECT 230.400 678.900 231.600 679.650 ;
        RECT 229.950 676.800 232.050 678.900 ;
        RECT 217.950 670.950 220.050 673.050 ;
        RECT 239.400 670.050 240.450 719.400 ;
        RECT 241.950 691.950 244.050 694.050 ;
        RECT 242.400 685.200 243.450 691.950 ;
        RECT 245.400 691.050 246.450 719.400 ;
        RECT 251.400 712.050 252.450 787.950 ;
        RECT 253.950 784.950 256.050 787.050 ;
        RECT 254.400 781.050 255.450 784.950 ;
        RECT 253.950 778.950 256.050 781.050 ;
        RECT 263.400 778.050 264.450 790.950 ;
        RECT 275.400 781.050 276.450 800.400 ;
        RECT 293.400 781.050 294.450 800.400 ;
        RECT 274.950 778.950 277.050 781.050 ;
        RECT 280.950 778.950 283.050 781.050 ;
        RECT 292.950 778.950 295.050 781.050 ;
        RECT 262.950 775.950 265.050 778.050 ;
        RECT 277.950 772.950 280.050 775.050 ;
        RECT 256.950 766.950 259.050 769.050 ;
        RECT 253.950 761.100 256.050 763.200 ;
        RECT 254.400 723.450 255.450 761.100 ;
        RECT 257.400 757.050 258.450 766.950 ;
        RECT 262.800 766.200 264.900 768.300 ;
        RECT 271.800 766.500 273.900 768.600 ;
        RECT 259.950 761.100 262.050 763.200 ;
        RECT 260.400 760.350 261.600 761.100 ;
        RECT 260.100 757.950 262.200 760.050 ;
        RECT 256.950 754.950 259.050 757.050 ;
        RECT 263.100 753.600 264.000 766.200 ;
        RECT 269.400 763.350 270.600 765.600 ;
        RECT 269.100 760.950 271.200 763.050 ;
        RECT 264.900 759.900 267.000 760.200 ;
        RECT 273.000 759.900 273.900 766.500 ;
        RECT 264.900 759.000 273.900 759.900 ;
        RECT 264.900 758.100 267.000 759.000 ;
        RECT 270.000 757.200 272.100 758.100 ;
        RECT 264.900 756.000 272.100 757.200 ;
        RECT 264.900 755.100 267.000 756.000 ;
        RECT 262.500 751.500 264.600 753.600 ;
        RECT 269.100 752.100 271.200 754.200 ;
        RECT 273.000 753.900 273.900 759.000 ;
        RECT 274.800 757.950 276.900 760.050 ;
        RECT 275.400 756.900 276.600 757.650 ;
        RECT 278.400 757.050 279.450 772.950 ;
        RECT 274.800 754.800 276.900 756.900 ;
        RECT 277.950 754.950 280.050 757.050 ;
        RECT 272.400 751.800 274.500 753.900 ;
        RECT 269.400 751.050 270.600 751.800 ;
        RECT 281.400 751.050 282.450 778.950 ;
        RECT 289.950 766.950 292.050 769.050 ;
        RECT 290.400 762.600 291.450 766.950 ;
        RECT 290.400 760.350 291.600 762.600 ;
        RECT 295.950 761.100 298.050 763.200 ;
        RECT 299.400 763.050 300.450 800.400 ;
        RECT 311.400 786.450 312.450 800.400 ;
        RECT 323.400 796.050 324.450 811.950 ;
        RECT 335.400 811.050 336.450 814.800 ;
        RECT 334.950 808.950 337.050 811.050 ;
        RECT 338.400 808.050 339.450 829.950 ;
        RECT 341.400 829.050 342.450 833.400 ;
        RECT 349.950 832.950 352.050 835.050 ;
        RECT 340.950 826.950 343.050 829.050 ;
        RECT 340.950 820.950 343.050 823.050 ;
        RECT 337.950 805.950 340.050 808.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 335.400 800.400 336.600 802.650 ;
        RECT 341.400 801.900 342.450 820.950 ;
        RECT 350.400 807.600 351.450 832.950 ;
        RECT 353.400 823.050 354.450 877.800 ;
        RECT 370.950 874.950 373.050 879.000 ;
        RECT 373.950 865.950 376.050 868.050 ;
        RECT 367.950 856.950 370.050 859.050 ;
        RECT 355.950 839.100 358.050 841.200 ;
        RECT 361.950 839.100 364.050 841.200 ;
        RECT 368.400 840.600 369.450 856.950 ;
        RECT 374.400 841.050 375.450 865.950 ;
        RECT 356.400 835.050 357.450 839.100 ;
        RECT 362.400 838.350 363.600 839.100 ;
        RECT 368.400 838.350 369.600 840.600 ;
        RECT 373.950 838.950 376.050 841.050 ;
        RECT 361.950 835.950 364.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 355.950 832.950 358.050 835.050 ;
        RECT 365.400 833.400 366.600 835.650 ;
        RECT 371.400 834.000 372.600 835.650 ;
        RECT 352.950 820.950 355.050 823.050 ;
        RECT 350.400 805.350 351.600 807.600 ;
        RECT 355.950 806.100 358.050 808.200 ;
        RECT 361.950 806.100 364.050 808.200 ;
        RECT 356.400 805.350 357.600 806.100 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 347.400 801.900 348.600 802.650 ;
        RECT 322.950 793.950 325.050 796.050 ;
        RECT 308.400 785.400 312.450 786.450 ;
        RECT 301.950 775.950 304.050 778.050 ;
        RECT 296.400 760.350 297.600 761.100 ;
        RECT 298.950 760.950 301.050 763.050 ;
        RECT 286.950 757.950 289.050 760.050 ;
        RECT 289.950 757.950 292.050 760.050 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 287.400 756.900 288.600 757.650 ;
        RECT 286.950 754.800 289.050 756.900 ;
        RECT 293.400 755.400 294.600 757.650 ;
        RECT 268.950 748.950 271.050 751.050 ;
        RECT 280.950 748.950 283.050 751.050 ;
        RECT 274.950 742.950 277.050 745.050 ;
        RECT 283.950 742.950 286.050 745.050 ;
        RECT 265.950 735.000 268.050 739.050 ;
        RECT 266.400 733.200 267.600 735.000 ;
        RECT 261.900 729.900 264.000 731.700 ;
        RECT 265.800 730.800 267.900 732.900 ;
        RECT 269.100 732.300 271.200 734.400 ;
        RECT 260.400 728.700 269.100 729.900 ;
        RECT 257.100 724.950 259.200 727.050 ;
        RECT 257.400 723.450 258.600 724.650 ;
        RECT 254.400 722.400 258.600 723.450 ;
        RECT 254.400 714.450 255.450 722.400 ;
        RECT 260.400 719.700 261.300 728.700 ;
        RECT 267.000 727.800 269.100 728.700 ;
        RECT 270.000 726.900 270.900 732.300 ;
        RECT 272.400 729.450 273.600 729.600 ;
        RECT 275.400 729.450 276.450 742.950 ;
        RECT 284.400 736.050 285.450 742.950 ;
        RECT 293.400 739.050 294.450 755.400 ;
        RECT 298.950 751.950 301.050 754.050 ;
        RECT 295.950 748.950 298.050 751.050 ;
        RECT 292.950 736.950 295.050 739.050 ;
        RECT 280.950 733.950 283.050 736.050 ;
        RECT 283.950 733.950 286.050 736.050 ;
        RECT 277.950 730.950 280.050 733.050 ;
        RECT 272.400 728.400 276.450 729.450 ;
        RECT 272.400 727.350 273.600 728.400 ;
        RECT 264.000 725.700 270.900 726.900 ;
        RECT 264.000 723.300 264.900 725.700 ;
        RECT 262.800 721.200 264.900 723.300 ;
        RECT 265.800 721.950 267.900 724.050 ;
        RECT 259.500 717.600 261.600 719.700 ;
        RECT 266.400 719.400 267.600 721.650 ;
        RECT 269.700 718.500 270.900 725.700 ;
        RECT 271.800 724.950 273.900 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 269.100 716.400 271.200 718.500 ;
        RECT 254.400 713.400 258.450 714.450 ;
        RECT 250.950 709.950 253.050 712.050 ;
        RECT 244.950 688.950 247.050 691.050 ;
        RECT 241.950 683.100 244.050 685.200 ;
        RECT 245.400 684.600 246.450 688.950 ;
        RECT 245.400 682.350 246.600 684.600 ;
        RECT 250.950 683.100 253.050 685.200 ;
        RECT 251.400 682.350 252.600 683.100 ;
        RECT 244.950 679.950 247.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 248.400 677.400 249.600 679.650 ;
        RECT 257.400 678.450 258.450 713.400 ;
        RECT 259.950 709.950 262.050 712.050 ;
        RECT 254.400 677.400 258.450 678.450 ;
        RECT 244.950 673.950 247.050 676.050 ;
        RECT 229.950 667.950 232.050 670.050 ;
        RECT 238.950 667.950 241.050 670.050 ;
        RECT 220.950 651.000 223.050 655.050 ;
        RECT 221.400 649.350 222.600 651.000 ;
        RECT 217.950 646.950 220.050 649.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 214.950 643.950 217.050 646.050 ;
        RECT 218.400 645.000 219.600 646.650 ;
        RECT 215.400 639.450 216.450 643.950 ;
        RECT 217.950 640.950 220.050 645.000 ;
        RECT 224.400 644.400 225.600 646.650 ;
        RECT 230.400 645.900 231.450 667.950 ;
        RECT 245.400 652.200 246.450 673.950 ;
        RECT 248.400 673.050 249.450 677.400 ;
        RECT 250.950 673.950 253.050 676.050 ;
        RECT 247.950 670.950 250.050 673.050 ;
        RECT 238.950 650.100 241.050 652.200 ;
        RECT 244.950 650.100 247.050 652.200 ;
        RECT 239.400 649.350 240.600 650.100 ;
        RECT 245.400 649.350 246.600 650.100 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 241.950 646.950 244.050 649.050 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 236.400 645.900 237.600 646.650 ;
        RECT 224.400 640.050 225.450 644.400 ;
        RECT 229.950 643.800 232.050 645.900 ;
        RECT 235.950 643.800 238.050 645.900 ;
        RECT 242.400 644.400 243.600 646.650 ;
        RECT 242.400 640.050 243.450 644.400 ;
        RECT 247.950 643.950 250.050 646.050 ;
        RECT 215.400 638.400 219.450 639.450 ;
        RECT 214.950 634.950 217.050 637.050 ;
        RECT 211.950 619.950 214.050 622.050 ;
        RECT 208.950 616.950 211.050 619.050 ;
        RECT 215.400 618.450 216.450 634.950 ;
        RECT 218.400 631.050 219.450 638.400 ;
        RECT 220.800 637.950 222.900 640.050 ;
        RECT 223.950 637.950 226.050 640.050 ;
        RECT 241.950 637.950 244.050 640.050 ;
        RECT 217.950 628.950 220.050 631.050 ;
        RECT 221.400 628.050 222.450 637.950 ;
        RECT 220.950 625.950 223.050 628.050 ;
        RECT 232.950 619.950 235.050 622.050 ;
        RECT 212.400 617.400 216.450 618.450 ;
        RECT 205.950 610.950 208.050 613.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 175.950 601.950 178.050 604.050 ;
        RECT 178.950 601.950 181.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 157.950 598.800 160.050 600.900 ;
        RECT 163.950 598.950 166.050 601.050 ;
        RECT 166.800 598.950 168.900 601.050 ;
        RECT 169.950 598.950 172.050 601.050 ;
        RECT 176.400 600.900 177.600 601.650 ;
        RECT 164.400 595.050 165.450 598.950 ;
        RECT 157.950 592.950 160.050 595.050 ;
        RECT 163.950 592.950 166.050 595.050 ;
        RECT 146.400 590.400 150.450 591.450 ;
        RECT 116.400 571.350 117.600 573.600 ;
        RECT 134.400 573.450 135.600 573.600 ;
        RECT 128.400 573.000 135.600 573.450 ;
        RECT 127.950 572.400 135.600 573.000 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 127.950 568.950 130.050 572.400 ;
        RECT 134.400 571.350 135.600 572.400 ;
        RECT 142.950 571.950 145.050 574.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 119.400 568.050 120.600 568.650 ;
        RECT 104.400 566.400 111.450 567.450 ;
        RECT 104.400 547.050 105.450 566.400 ;
        RECT 112.950 565.950 115.050 568.050 ;
        RECT 119.400 566.400 124.050 568.050 ;
        RECT 120.000 565.950 124.050 566.400 ;
        RECT 106.950 550.950 109.050 553.050 ;
        RECT 103.950 544.950 106.050 547.050 ;
        RECT 100.950 541.950 103.050 544.050 ;
        RECT 91.950 532.950 94.050 535.050 ;
        RECT 86.400 527.400 90.450 528.450 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 77.400 521.400 78.600 523.650 ;
        RECT 83.400 522.900 84.600 523.650 ;
        RECT 67.950 517.950 70.050 520.050 ;
        RECT 77.400 517.050 78.450 521.400 ;
        RECT 82.950 520.800 85.050 522.900 ;
        RECT 76.950 514.950 79.050 517.050 ;
        RECT 67.950 505.950 70.050 508.050 ;
        RECT 59.400 493.350 60.600 494.100 ;
        RECT 64.950 493.950 67.050 496.050 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 62.400 489.450 63.600 490.650 ;
        RECT 62.400 488.400 66.450 489.450 ;
        RECT 61.950 481.950 64.050 487.050 ;
        RECT 65.400 472.050 66.450 488.400 ;
        RECT 68.400 481.050 69.450 505.950 ;
        RECT 79.950 502.950 82.050 505.050 ;
        RECT 70.950 493.950 73.050 496.050 ;
        RECT 80.400 495.600 81.450 502.950 ;
        RECT 83.400 499.050 84.450 520.800 ;
        RECT 82.950 496.950 85.050 499.050 ;
        RECT 67.950 478.950 70.050 481.050 ;
        RECT 71.400 478.050 72.450 493.950 ;
        RECT 80.400 493.350 81.600 495.600 ;
        RECT 85.950 494.100 88.050 496.200 ;
        RECT 89.400 495.450 90.450 527.400 ;
        RECT 94.950 527.100 97.050 529.200 ;
        RECT 101.400 528.600 102.450 541.950 ;
        RECT 107.400 538.050 108.450 550.950 ;
        RECT 113.400 541.050 114.450 565.950 ;
        RECT 127.950 565.800 130.050 567.900 ;
        RECT 137.400 566.400 138.600 568.650 ;
        RECT 146.400 568.050 147.450 590.400 ;
        RECT 151.950 588.450 156.000 589.050 ;
        RECT 151.950 588.000 156.450 588.450 ;
        RECT 151.950 586.950 157.050 588.000 ;
        RECT 154.950 583.950 157.050 586.950 ;
        RECT 151.950 580.950 154.050 583.050 ;
        RECT 148.950 577.950 151.050 580.050 ;
        RECT 115.950 556.950 118.050 559.050 ;
        RECT 112.950 538.950 115.050 541.050 ;
        RECT 106.950 535.950 109.050 538.050 ;
        RECT 116.400 535.050 117.450 556.950 ;
        RECT 128.400 553.050 129.450 565.800 ;
        RECT 137.400 564.450 138.450 566.400 ;
        RECT 145.950 565.950 148.050 568.050 ;
        RECT 149.400 567.900 150.450 577.950 ;
        RECT 152.400 577.050 153.450 580.950 ;
        RECT 151.950 574.950 154.050 577.050 ;
        RECT 158.400 573.600 159.450 592.950 ;
        RECT 158.400 571.350 159.600 573.600 ;
        RECT 163.950 572.100 166.050 574.200 ;
        RECT 164.400 571.350 165.600 572.100 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 148.950 565.800 151.050 567.900 ;
        RECT 151.950 565.950 154.050 568.050 ;
        RECT 155.400 567.900 156.600 568.650 ;
        RECT 137.400 563.400 141.450 564.450 ;
        RECT 140.400 559.050 141.450 563.400 ;
        RECT 139.950 556.950 142.050 559.050 ;
        RECT 136.950 553.950 139.050 556.050 ;
        RECT 124.950 551.400 129.450 553.050 ;
        RECT 124.950 550.950 129.000 551.400 ;
        RECT 130.950 550.950 133.050 553.050 ;
        RECT 118.950 544.950 121.050 547.050 ;
        RECT 106.950 532.800 109.050 534.900 ;
        RECT 115.950 532.950 118.050 535.050 ;
        RECT 107.400 529.050 108.450 532.800 ;
        RECT 95.400 526.350 96.600 527.100 ;
        RECT 101.400 526.350 102.600 528.600 ;
        RECT 106.950 526.950 109.050 529.050 ;
        RECT 119.400 528.600 120.450 544.950 ;
        RECT 124.950 538.950 127.050 541.050 ;
        RECT 119.400 526.350 120.600 528.600 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 98.400 522.000 99.600 523.650 ;
        RECT 104.400 522.000 105.600 523.650 ;
        RECT 97.950 517.950 100.050 522.000 ;
        RECT 103.950 517.950 106.050 522.000 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 116.400 521.400 117.600 523.650 ;
        RECT 125.400 522.900 126.450 538.950 ;
        RECT 127.950 527.100 130.050 529.200 ;
        RECT 131.400 529.050 132.450 550.950 ;
        RECT 137.400 541.050 138.450 553.950 ;
        RECT 136.950 538.950 139.050 541.050 ;
        RECT 148.950 538.950 151.050 541.050 ;
        RECT 145.950 532.950 148.050 535.050 ;
        RECT 100.950 511.950 103.050 514.050 ;
        RECT 101.400 508.050 102.450 511.950 ;
        RECT 100.950 505.950 103.050 508.050 ;
        RECT 94.950 502.950 97.050 505.050 ;
        RECT 95.400 496.050 96.450 502.950 ;
        RECT 89.400 494.400 93.450 495.450 ;
        RECT 86.400 493.350 87.600 494.100 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 77.400 490.050 78.600 490.650 ;
        RECT 73.950 488.400 78.600 490.050 ;
        RECT 83.400 489.000 84.600 490.650 ;
        RECT 73.950 487.950 78.450 488.400 ;
        RECT 70.950 475.950 73.050 478.050 ;
        RECT 67.950 472.950 70.050 475.050 ;
        RECT 64.950 469.950 67.050 472.050 ;
        RECT 49.950 451.950 52.050 454.050 ;
        RECT 68.400 453.450 69.450 472.950 ;
        RECT 77.400 463.050 78.450 487.950 ;
        RECT 82.950 484.950 85.050 489.000 ;
        RECT 85.950 484.950 88.050 487.050 ;
        RECT 76.950 460.950 79.050 463.050 ;
        RECT 65.400 452.400 69.450 453.450 ;
        RECT 51.000 450.900 54.000 451.050 ;
        RECT 49.950 450.600 54.000 450.900 ;
        RECT 49.950 448.950 54.600 450.600 ;
        RECT 58.950 449.100 61.050 451.200 ;
        RECT 49.950 448.800 52.050 448.950 ;
        RECT 53.400 448.350 54.600 448.950 ;
        RECT 59.400 448.350 60.600 449.100 ;
        RECT 52.950 445.950 55.050 448.050 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 32.400 418.200 33.450 442.950 ;
        RECT 38.400 433.050 39.450 443.400 ;
        RECT 46.950 442.950 49.050 445.050 ;
        RECT 49.950 442.950 52.050 445.050 ;
        RECT 56.400 444.900 57.600 445.650 ;
        RECT 50.400 436.050 51.450 442.950 ;
        RECT 55.950 442.800 58.050 444.900 ;
        RECT 49.950 433.950 52.050 436.050 ;
        RECT 58.950 433.950 61.050 436.050 ;
        RECT 37.950 430.950 40.050 433.050 ;
        RECT 40.950 421.950 43.050 424.050 ;
        RECT 16.950 416.100 19.050 418.200 ;
        RECT 31.950 416.100 34.050 418.200 ;
        RECT 41.400 417.600 42.450 421.950 ;
        RECT 17.400 415.350 18.600 416.100 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 17.100 412.950 19.200 415.050 ;
        RECT 22.800 412.950 24.900 415.050 ;
        RECT 25.800 412.950 27.900 415.050 ;
        RECT 23.400 411.900 24.600 412.650 ;
        RECT 22.950 409.800 25.050 411.900 ;
        RECT 32.400 409.050 33.450 416.100 ;
        RECT 41.400 415.350 42.600 417.600 ;
        RECT 46.950 415.950 49.050 418.050 ;
        RECT 59.400 417.600 60.450 433.950 ;
        RECT 65.400 418.050 66.450 452.400 ;
        RECT 67.950 449.100 70.050 451.200 ;
        RECT 82.950 450.000 85.050 454.050 ;
        RECT 86.400 451.050 87.450 484.950 ;
        RECT 92.400 475.050 93.450 494.400 ;
        RECT 94.950 493.950 97.050 496.050 ;
        RECT 101.400 495.600 102.450 505.950 ;
        RECT 101.400 493.350 102.600 495.600 ;
        RECT 106.950 494.100 109.050 496.200 ;
        RECT 113.400 495.450 114.450 520.950 ;
        RECT 116.400 514.050 117.450 521.400 ;
        RECT 124.950 520.800 127.050 522.900 ;
        RECT 128.400 520.050 129.450 527.100 ;
        RECT 130.950 526.950 133.050 529.050 ;
        RECT 136.950 527.100 139.050 529.200 ;
        RECT 142.950 527.100 145.050 529.200 ;
        RECT 146.400 529.050 147.450 532.950 ;
        RECT 137.400 526.350 138.600 527.100 ;
        RECT 143.400 526.350 144.600 527.100 ;
        RECT 145.950 526.950 148.050 529.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 130.950 520.950 133.050 523.050 ;
        RECT 134.400 522.900 135.600 523.650 ;
        RECT 127.950 517.950 130.050 520.050 ;
        RECT 115.950 511.950 118.050 514.050 ;
        RECT 128.400 505.050 129.450 517.950 ;
        RECT 131.400 517.050 132.450 520.950 ;
        RECT 133.950 520.800 136.050 522.900 ;
        RECT 140.400 521.400 141.600 523.650 ;
        RECT 130.950 514.950 133.050 517.050 ;
        RECT 136.950 514.950 139.050 517.050 ;
        RECT 127.950 502.950 130.050 505.050 ;
        RECT 137.400 499.050 138.450 514.950 ;
        RECT 140.400 514.050 141.450 521.400 ;
        RECT 145.950 520.800 148.050 522.900 ;
        RECT 139.950 511.950 142.050 514.050 ;
        RECT 139.950 508.800 142.050 510.900 ;
        RECT 113.400 494.400 117.450 495.450 ;
        RECT 107.400 493.350 108.600 494.100 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 98.400 489.900 99.600 490.650 ;
        RECT 97.950 487.800 100.050 489.900 ;
        RECT 104.400 488.400 105.600 490.650 ;
        RECT 110.400 489.450 111.600 490.650 ;
        RECT 110.400 488.400 114.450 489.450 ;
        RECT 91.950 472.950 94.050 475.050 ;
        RECT 94.950 460.950 97.050 463.050 ;
        RECT 88.950 451.950 91.050 454.050 ;
        RECT 68.400 445.050 69.450 449.100 ;
        RECT 83.400 448.350 84.600 450.000 ;
        RECT 85.950 448.950 88.050 451.050 ;
        RECT 73.950 445.950 76.050 448.050 ;
        RECT 76.950 445.950 79.050 448.050 ;
        RECT 79.950 445.950 82.050 448.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 67.950 442.950 70.050 445.050 ;
        RECT 74.400 444.900 75.600 445.650 ;
        RECT 80.400 444.900 81.600 445.650 ;
        RECT 73.950 442.800 76.050 444.900 ;
        RECT 79.950 442.800 82.050 444.900 ;
        RECT 85.950 442.950 88.050 445.050 ;
        RECT 86.400 433.050 87.450 442.950 ;
        RECT 85.950 430.950 88.050 433.050 ;
        RECT 89.400 430.050 90.450 451.950 ;
        RECT 95.400 450.600 96.450 460.950 ;
        RECT 104.400 460.050 105.450 488.400 ;
        RECT 113.400 484.050 114.450 488.400 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 109.950 469.950 112.050 472.050 ;
        RECT 106.950 466.950 109.050 469.050 ;
        RECT 107.400 463.050 108.450 466.950 ;
        RECT 106.950 460.950 109.050 463.050 ;
        RECT 103.950 457.950 106.050 460.050 ;
        RECT 95.400 448.350 96.600 450.600 ;
        RECT 100.950 450.000 103.050 454.050 ;
        RECT 101.400 448.350 102.600 450.000 ;
        RECT 94.950 445.950 97.050 448.050 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 98.400 444.900 99.600 445.650 ;
        RECT 97.950 442.800 100.050 444.900 ;
        RECT 104.400 444.000 105.600 445.650 ;
        RECT 103.950 439.950 106.050 444.000 ;
        RECT 94.950 430.950 97.050 433.050 ;
        RECT 88.950 427.950 91.050 430.050 ;
        RECT 95.400 418.200 96.450 430.950 ;
        RECT 110.400 427.050 111.450 469.950 ;
        RECT 113.400 448.050 114.450 481.950 ;
        RECT 116.400 466.050 117.450 494.400 ;
        RECT 127.950 494.100 130.050 496.200 ;
        RECT 133.950 495.000 136.050 499.050 ;
        RECT 136.950 496.950 139.050 499.050 ;
        RECT 128.400 493.350 129.600 494.100 ;
        RECT 134.400 493.350 135.600 495.000 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 133.950 490.950 136.050 493.050 ;
        RECT 125.400 489.900 126.600 490.650 ;
        RECT 124.950 487.800 127.050 489.900 ;
        RECT 131.400 488.400 132.600 490.650 ;
        RECT 131.400 487.050 132.450 488.400 ;
        RECT 136.950 487.950 139.050 490.050 ;
        RECT 130.950 484.950 133.050 487.050 ;
        RECT 121.950 481.950 127.050 484.050 ;
        RECT 131.400 478.050 132.450 484.950 ;
        RECT 137.400 484.050 138.450 487.950 ;
        RECT 136.950 481.950 139.050 484.050 ;
        RECT 130.950 475.950 133.050 478.050 ;
        RECT 136.950 472.950 139.050 475.050 ;
        RECT 115.950 463.950 118.050 466.050 ;
        RECT 130.950 463.950 133.050 466.050 ;
        RECT 118.950 449.100 121.050 454.050 ;
        RECT 124.950 449.100 127.050 451.200 ;
        RECT 131.400 450.600 132.450 463.950 ;
        RECT 137.400 460.050 138.450 472.950 ;
        RECT 136.950 457.950 139.050 460.050 ;
        RECT 119.400 448.350 120.600 449.100 ;
        RECT 125.400 448.350 126.600 449.100 ;
        RECT 131.400 448.350 132.600 450.600 ;
        RECT 136.950 449.100 139.050 451.200 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 118.950 445.950 121.050 448.050 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 127.950 445.950 130.050 448.050 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 122.400 443.400 123.600 445.650 ;
        RECT 128.400 444.900 129.600 445.650 ;
        RECT 122.400 433.050 123.450 443.400 ;
        RECT 127.950 442.800 130.050 444.900 ;
        RECT 133.950 442.950 136.050 445.050 ;
        RECT 121.950 430.950 124.050 433.050 ;
        RECT 128.400 430.050 129.450 442.800 ;
        RECT 134.400 435.450 135.450 442.950 ;
        RECT 131.400 434.400 135.450 435.450 ;
        RECT 127.950 427.950 130.050 430.050 ;
        RECT 109.950 424.950 112.050 427.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 38.400 411.000 39.600 412.650 ;
        RECT 31.950 406.950 34.050 409.050 ;
        RECT 37.950 406.950 40.050 411.000 ;
        RECT 4.950 388.950 7.050 391.050 ;
        RECT 28.950 385.950 31.050 388.050 ;
        RECT 4.950 376.950 7.050 379.050 ;
        RECT 5.400 241.050 6.450 376.950 ;
        RECT 14.400 372.450 15.600 372.600 ;
        RECT 11.400 371.400 15.600 372.450 ;
        RECT 11.400 361.050 12.450 371.400 ;
        RECT 14.400 370.350 15.600 371.400 ;
        RECT 23.400 372.450 24.600 372.600 ;
        RECT 23.400 371.400 27.450 372.450 ;
        RECT 23.400 370.350 24.600 371.400 ;
        RECT 14.100 367.950 16.200 370.050 ;
        RECT 17.400 367.950 19.500 370.050 ;
        RECT 22.800 367.950 24.900 370.050 ;
        RECT 17.400 366.900 18.600 367.650 ;
        RECT 16.950 364.800 19.050 366.900 ;
        RECT 10.950 358.950 13.050 361.050 ;
        RECT 11.400 333.450 12.450 358.950 ;
        RECT 19.950 346.950 22.050 349.050 ;
        RECT 20.400 340.200 21.450 346.950 ;
        RECT 26.400 342.450 27.450 371.400 ;
        RECT 29.400 370.050 30.450 385.950 ;
        RECT 47.400 379.050 48.450 415.950 ;
        RECT 59.400 415.350 60.600 417.600 ;
        RECT 64.950 415.950 67.050 418.050 ;
        RECT 76.950 416.100 79.050 418.200 ;
        RECT 77.400 415.350 78.600 416.100 ;
        RECT 85.950 415.950 88.050 418.050 ;
        RECT 94.950 416.100 97.050 418.200 ;
        RECT 106.950 416.100 109.050 418.200 ;
        RECT 115.950 416.100 118.050 418.200 ;
        RECT 121.950 416.100 124.050 418.200 ;
        RECT 55.950 412.950 58.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 56.400 411.900 57.600 412.650 ;
        RECT 62.400 411.900 63.600 412.650 ;
        RECT 55.950 409.800 58.050 411.900 ;
        RECT 61.950 409.800 64.050 411.900 ;
        RECT 74.400 410.400 75.600 412.650 ;
        RECT 80.400 411.450 81.600 412.650 ;
        RECT 86.400 411.450 87.450 415.950 ;
        RECT 95.400 415.350 96.600 416.100 ;
        RECT 91.950 412.950 94.050 415.050 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 97.950 412.950 100.050 415.050 ;
        RECT 80.400 410.400 87.450 411.450 ;
        RECT 98.400 410.400 99.600 412.650 ;
        RECT 74.400 406.050 75.450 410.400 ;
        RECT 73.950 403.950 76.050 406.050 ;
        RECT 52.950 391.950 55.050 394.050 ;
        RECT 46.950 376.950 49.050 379.050 ;
        RECT 37.950 371.100 40.050 373.200 ;
        RECT 44.400 372.450 45.600 372.600 ;
        RECT 47.400 372.450 48.450 376.950 ;
        RECT 53.400 373.200 54.450 391.950 ;
        RECT 61.950 385.950 64.050 388.050 ;
        RECT 44.400 371.400 48.450 372.450 ;
        RECT 38.400 370.350 39.600 371.100 ;
        RECT 44.400 370.350 45.600 371.400 ;
        RECT 52.950 371.100 55.050 373.200 ;
        RECT 62.400 372.600 63.450 385.950 ;
        RECT 28.950 367.950 31.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 43.950 367.950 46.050 370.050 ;
        RECT 41.400 365.400 42.600 367.650 ;
        RECT 41.400 355.050 42.450 365.400 ;
        RECT 40.950 352.950 43.050 355.050 ;
        RECT 41.400 346.050 42.450 352.950 ;
        RECT 40.950 343.950 43.050 346.050 ;
        RECT 46.950 343.950 49.050 346.050 ;
        RECT 26.400 341.400 30.450 342.450 ;
        RECT 19.950 338.100 22.050 340.200 ;
        RECT 25.950 338.100 28.050 340.200 ;
        RECT 20.400 337.350 21.600 338.100 ;
        RECT 14.100 334.950 16.200 337.050 ;
        RECT 19.500 334.950 21.600 337.050 ;
        RECT 22.800 334.950 24.900 337.050 ;
        RECT 14.400 333.450 15.600 334.650 ;
        RECT 11.400 332.400 15.600 333.450 ;
        RECT 23.400 333.000 24.600 334.650 ;
        RECT 14.400 301.050 15.450 332.400 ;
        RECT 22.950 328.950 25.050 333.000 ;
        RECT 13.950 298.950 16.050 301.050 ;
        RECT 16.950 293.100 19.050 295.200 ;
        RECT 17.400 292.350 18.600 293.100 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 14.400 287.400 15.600 289.650 ;
        RECT 20.400 288.000 21.600 289.650 ;
        RECT 14.400 283.050 15.450 287.400 ;
        RECT 19.950 283.950 22.050 288.000 ;
        RECT 22.950 286.950 25.050 289.050 ;
        RECT 13.950 280.950 16.050 283.050 ;
        RECT 23.400 280.050 24.450 286.950 ;
        RECT 26.400 286.050 27.450 338.100 ;
        RECT 29.400 333.900 30.450 341.400 ;
        RECT 40.950 338.100 43.050 340.200 ;
        RECT 47.400 339.600 48.450 343.950 ;
        RECT 41.400 337.350 42.600 338.100 ;
        RECT 47.400 337.350 48.600 339.600 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 38.400 333.900 39.600 334.650 ;
        RECT 44.400 333.900 45.600 334.650 ;
        RECT 28.950 331.800 31.050 333.900 ;
        RECT 37.950 331.800 40.050 333.900 ;
        RECT 43.950 331.800 46.050 333.900 ;
        RECT 37.950 328.650 40.050 330.750 ;
        RECT 28.950 298.950 31.050 301.050 ;
        RECT 25.950 283.950 28.050 286.050 ;
        RECT 29.400 283.050 30.450 298.950 ;
        RECT 38.400 298.050 39.450 328.650 ;
        RECT 44.400 319.050 45.450 331.800 ;
        RECT 43.950 316.950 46.050 319.050 ;
        RECT 53.400 307.050 54.450 371.100 ;
        RECT 62.400 370.350 63.600 372.600 ;
        RECT 67.950 371.100 70.050 373.200 ;
        RECT 68.400 370.350 69.600 371.100 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 67.950 367.950 70.050 370.050 ;
        RECT 59.400 365.400 60.600 367.650 ;
        RECT 65.400 366.000 66.600 367.650 ;
        RECT 59.400 361.050 60.450 365.400 ;
        RECT 64.950 361.950 67.050 366.000 ;
        RECT 70.950 364.950 73.050 367.050 ;
        RECT 58.950 358.950 61.050 361.050 ;
        RECT 55.950 343.950 58.050 346.050 ;
        RECT 67.950 343.950 70.050 346.050 ;
        RECT 56.400 340.050 57.450 343.950 ;
        RECT 55.800 337.950 57.900 340.050 ;
        RECT 58.950 338.100 61.050 340.200 ;
        RECT 59.400 337.350 60.600 338.100 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 62.400 333.900 63.600 334.650 ;
        RECT 61.950 331.800 64.050 333.900 ;
        RECT 52.950 304.950 55.050 307.050 ;
        RECT 68.400 298.050 69.450 343.950 ;
        RECT 71.400 334.050 72.450 364.950 ;
        RECT 74.400 340.050 75.450 403.950 ;
        RECT 98.400 394.050 99.450 410.400 ;
        RECT 107.400 400.050 108.450 416.100 ;
        RECT 116.400 415.350 117.600 416.100 ;
        RECT 122.400 415.350 123.600 416.100 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 118.950 412.950 121.050 415.050 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 113.400 410.400 114.600 412.650 ;
        RECT 119.400 410.400 120.600 412.650 ;
        RECT 106.950 397.950 109.050 400.050 ;
        RECT 113.400 396.450 114.450 410.400 ;
        RECT 115.950 397.950 118.050 400.050 ;
        RECT 107.400 395.400 114.450 396.450 ;
        RECT 97.950 391.950 100.050 394.050 ;
        RECT 97.950 376.950 100.050 379.050 ;
        RECT 80.400 372.450 81.600 372.600 ;
        RECT 77.400 371.400 81.600 372.450 ;
        RECT 77.400 364.050 78.450 371.400 ;
        RECT 80.400 370.350 81.600 371.400 ;
        RECT 88.950 371.100 91.050 373.200 ;
        RECT 89.400 370.350 90.600 371.100 ;
        RECT 80.100 367.950 82.200 370.050 ;
        RECT 83.400 367.950 85.500 370.050 ;
        RECT 88.800 367.950 90.900 370.050 ;
        RECT 83.400 365.400 84.600 367.650 ;
        RECT 76.950 361.950 79.050 364.050 ;
        RECT 77.400 343.050 78.450 361.950 ;
        RECT 83.400 355.050 84.450 365.400 ;
        RECT 82.950 352.950 85.050 355.050 ;
        RECT 79.950 346.950 82.050 349.050 ;
        RECT 76.950 340.950 79.050 343.050 ;
        RECT 73.950 337.950 76.050 340.050 ;
        RECT 80.400 339.600 81.450 346.950 ;
        RECT 88.950 340.950 91.050 343.050 ;
        RECT 80.400 337.350 81.600 339.600 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 70.950 331.950 73.050 334.050 ;
        RECT 77.400 333.900 78.600 334.650 ;
        RECT 76.950 331.800 79.050 333.900 ;
        RECT 83.400 332.400 84.600 334.650 ;
        RECT 89.400 333.900 90.450 340.950 ;
        RECT 98.400 339.600 99.450 376.950 ;
        RECT 107.400 373.200 108.450 395.400 ;
        RECT 112.950 391.950 115.050 394.050 ;
        RECT 106.950 371.100 109.050 373.200 ;
        RECT 113.400 372.600 114.450 391.950 ;
        RECT 116.400 373.050 117.450 397.950 ;
        RECT 119.400 394.050 120.450 410.400 ;
        RECT 131.400 408.450 132.450 434.400 ;
        RECT 137.400 426.450 138.450 449.100 ;
        RECT 140.400 442.050 141.450 508.800 ;
        RECT 146.400 508.050 147.450 520.800 ;
        RECT 149.400 514.050 150.450 538.950 ;
        RECT 148.950 511.950 151.050 514.050 ;
        RECT 152.400 511.050 153.450 565.950 ;
        RECT 154.950 565.800 157.050 567.900 ;
        RECT 161.400 566.400 162.600 568.650 ;
        RECT 161.400 559.050 162.450 566.400 ;
        RECT 166.950 565.950 169.050 568.050 ;
        RECT 160.950 556.950 163.050 559.050 ;
        RECT 160.950 535.950 163.050 538.050 ;
        RECT 154.950 532.950 157.050 535.050 ;
        RECT 155.400 529.050 156.450 532.950 ;
        RECT 154.950 526.950 157.050 529.050 ;
        RECT 161.400 528.600 162.450 535.950 ;
        RECT 167.400 529.050 168.450 565.950 ;
        RECT 170.400 553.050 171.450 598.950 ;
        RECT 175.950 598.800 178.050 600.900 ;
        RECT 182.400 599.400 183.600 601.650 ;
        RECT 191.400 601.050 192.450 605.100 ;
        RECT 200.400 604.350 201.600 606.600 ;
        RECT 205.950 605.100 208.050 609.900 ;
        RECT 209.400 607.050 210.450 616.950 ;
        RECT 206.400 604.350 207.600 605.100 ;
        RECT 208.950 604.950 211.050 607.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 182.400 595.050 183.450 599.400 ;
        RECT 184.950 598.950 187.050 601.050 ;
        RECT 190.950 598.950 193.050 601.050 ;
        RECT 197.400 600.000 198.600 601.650 ;
        RECT 203.400 600.900 204.600 601.650 ;
        RECT 181.950 592.950 184.050 595.050 ;
        RECT 181.950 586.950 184.050 589.050 ;
        RECT 172.950 577.950 175.050 580.050 ;
        RECT 169.950 550.950 172.050 553.050 ;
        RECT 169.950 529.950 172.050 532.050 ;
        RECT 161.400 526.350 162.600 528.600 ;
        RECT 166.950 526.950 169.050 529.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 154.950 520.950 157.050 523.050 ;
        RECT 158.400 522.900 159.600 523.650 ;
        RECT 151.950 508.950 154.050 511.050 ;
        RECT 145.950 505.950 148.050 508.050 ;
        RECT 142.950 496.950 145.050 499.050 ;
        RECT 143.400 451.050 144.450 496.950 ;
        RECT 146.400 496.050 147.450 505.950 ;
        RECT 145.800 493.950 147.900 496.050 ;
        RECT 148.950 494.100 151.050 496.200 ;
        RECT 155.400 496.050 156.450 520.950 ;
        RECT 157.950 520.800 160.050 522.900 ;
        RECT 164.400 521.400 165.600 523.650 ;
        RECT 159.000 519.750 162.000 520.050 ;
        RECT 157.950 519.300 162.000 519.750 ;
        RECT 157.950 519.000 162.450 519.300 ;
        RECT 157.950 517.950 163.050 519.000 ;
        RECT 157.950 517.650 160.050 517.950 ;
        RECT 160.950 514.950 163.050 517.950 ;
        RECT 157.950 511.950 160.050 514.050 ;
        RECT 149.400 493.350 150.600 494.100 ;
        RECT 154.950 493.950 157.050 496.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 487.950 157.050 490.050 ;
        RECT 145.950 484.950 148.050 487.050 ;
        RECT 146.400 478.050 147.450 484.950 ;
        RECT 145.950 475.950 148.050 478.050 ;
        RECT 155.400 466.050 156.450 487.950 ;
        RECT 154.950 463.950 157.050 466.050 ;
        RECT 142.950 448.950 145.050 451.050 ;
        RECT 145.950 449.100 148.050 451.200 ;
        RECT 152.400 450.450 153.600 450.600 ;
        RECT 155.400 450.450 156.450 463.950 ;
        RECT 152.400 449.400 156.450 450.450 ;
        RECT 146.400 448.350 147.600 449.100 ;
        RECT 152.400 448.350 153.600 449.400 ;
        RECT 158.400 448.050 159.450 511.950 ;
        RECT 164.400 505.050 165.450 521.400 ;
        RECT 166.950 520.950 169.050 523.050 ;
        RECT 163.950 502.950 166.050 505.050 ;
        RECT 163.950 498.450 166.050 499.050 ;
        RECT 167.400 498.450 168.450 520.950 ;
        RECT 170.400 505.050 171.450 529.950 ;
        RECT 173.400 529.050 174.450 577.950 ;
        RECT 182.400 577.050 183.450 586.950 ;
        RECT 181.950 574.950 184.050 577.050 ;
        RECT 185.400 576.450 186.450 598.950 ;
        RECT 196.950 595.950 199.050 600.000 ;
        RECT 202.950 598.800 205.050 600.900 ;
        RECT 212.400 600.450 213.450 617.400 ;
        RECT 217.950 610.950 223.050 613.050 ;
        RECT 226.950 610.950 229.050 613.050 ;
        RECT 214.950 605.100 217.050 607.200 ;
        RECT 220.950 605.100 223.050 607.200 ;
        RECT 227.400 606.600 228.450 610.950 ;
        RECT 233.400 607.050 234.450 619.950 ;
        RECT 235.950 607.950 238.050 610.050 ;
        RECT 215.400 601.050 216.450 605.100 ;
        RECT 221.400 604.350 222.600 605.100 ;
        RECT 227.400 604.350 228.600 606.600 ;
        RECT 232.950 604.950 235.050 607.050 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 226.950 601.950 229.050 604.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 209.400 599.400 213.450 600.450 ;
        RECT 193.950 592.950 196.050 595.050 ;
        RECT 185.400 575.400 189.450 576.450 ;
        RECT 182.400 573.600 183.450 574.950 ;
        RECT 188.400 573.600 189.450 575.400 ;
        RECT 194.400 574.050 195.450 592.950 ;
        RECT 197.400 577.050 198.450 595.950 ;
        RECT 209.400 595.050 210.450 599.400 ;
        RECT 214.950 598.950 217.050 601.050 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 224.400 599.400 225.600 601.650 ;
        RECT 230.400 600.900 231.600 601.650 ;
        RECT 218.400 595.050 219.450 598.950 ;
        RECT 199.950 592.950 202.050 595.050 ;
        RECT 208.950 592.950 211.050 595.050 ;
        RECT 217.950 592.950 220.050 595.050 ;
        RECT 196.950 574.950 199.050 577.050 ;
        RECT 182.400 571.350 183.600 573.600 ;
        RECT 188.400 571.350 189.600 573.600 ;
        RECT 193.950 571.950 196.050 574.050 ;
        RECT 196.950 571.800 199.050 573.900 ;
        RECT 178.950 568.950 181.050 571.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 184.950 568.950 187.050 571.050 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 179.400 566.400 180.600 568.650 ;
        RECT 185.400 566.400 186.600 568.650 ;
        RECT 191.400 567.900 192.600 568.650 ;
        RECT 197.400 567.900 198.450 571.800 ;
        RECT 200.400 568.050 201.450 592.950 ;
        RECT 211.950 586.950 214.050 589.050 ;
        RECT 212.400 583.050 213.450 586.950 ;
        RECT 211.950 580.950 214.050 583.050 ;
        RECT 205.950 572.100 208.050 574.200 ;
        RECT 212.400 573.600 213.450 580.950 ;
        RECT 224.400 574.050 225.450 599.400 ;
        RECT 229.950 598.800 232.050 600.900 ;
        RECT 232.950 598.950 235.050 601.050 ;
        RECT 236.400 600.900 237.450 607.950 ;
        RECT 241.950 606.000 244.050 610.050 ;
        RECT 248.400 606.600 249.450 643.950 ;
        RECT 251.400 610.050 252.450 673.950 ;
        RECT 254.400 646.050 255.450 677.400 ;
        RECT 260.400 676.050 261.450 709.950 ;
        RECT 262.950 697.950 265.050 700.050 ;
        RECT 263.400 685.050 264.450 697.950 ;
        RECT 265.950 688.950 268.050 691.050 ;
        RECT 262.950 682.950 265.050 685.050 ;
        RECT 266.400 684.600 267.450 688.950 ;
        RECT 275.400 688.200 276.450 724.950 ;
        RECT 278.400 705.450 279.450 730.950 ;
        RECT 281.400 730.050 282.450 733.950 ;
        RECT 280.950 727.950 283.050 730.050 ;
        RECT 283.950 729.000 286.050 732.900 ;
        RECT 289.950 729.000 292.050 733.050 ;
        RECT 293.400 730.050 294.450 736.950 ;
        RECT 284.400 727.350 285.600 729.000 ;
        RECT 290.400 727.350 291.600 729.000 ;
        RECT 292.950 727.950 295.050 730.050 ;
        RECT 283.950 724.950 286.050 727.050 ;
        RECT 286.950 724.950 289.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 287.400 722.400 288.600 724.650 ;
        RECT 283.950 718.950 286.050 721.050 ;
        RECT 278.400 704.400 282.450 705.450 ;
        RECT 277.950 700.950 280.050 703.050 ;
        RECT 274.950 686.100 277.050 688.200 ;
        RECT 259.950 673.950 262.050 676.050 ;
        RECT 256.950 670.950 259.050 673.050 ;
        RECT 257.400 664.050 258.450 670.950 ;
        RECT 256.950 661.950 259.050 664.050 ;
        RECT 259.950 658.950 262.050 661.050 ;
        RECT 260.400 651.600 261.450 658.950 ;
        RECT 263.400 658.050 264.450 682.950 ;
        RECT 266.400 682.350 267.600 684.600 ;
        RECT 274.950 682.950 277.050 685.050 ;
        RECT 275.400 682.350 276.600 682.950 ;
        RECT 266.100 679.950 268.200 682.050 ;
        RECT 269.400 679.950 271.500 682.050 ;
        RECT 274.800 679.950 276.900 682.050 ;
        RECT 269.400 678.900 270.600 679.650 ;
        RECT 278.400 679.050 279.450 700.950 ;
        RECT 281.400 685.050 282.450 704.400 ;
        RECT 280.950 682.950 283.050 685.050 ;
        RECT 280.950 679.800 283.050 681.900 ;
        RECT 268.950 676.800 271.050 678.900 ;
        RECT 277.950 676.950 280.050 679.050 ;
        RECT 269.400 667.050 270.450 676.800 ;
        RECT 281.400 676.050 282.450 679.800 ;
        RECT 271.950 673.950 274.050 676.050 ;
        RECT 276.000 675.900 279.000 676.050 ;
        RECT 276.000 675.450 280.050 675.900 ;
        RECT 275.400 673.950 280.050 675.450 ;
        RECT 280.950 673.950 283.050 676.050 ;
        RECT 268.950 664.950 271.050 667.050 ;
        RECT 262.950 655.950 265.050 658.050 ;
        RECT 268.950 655.950 271.050 658.050 ;
        RECT 260.400 649.350 261.600 651.600 ;
        RECT 257.100 646.950 259.200 649.050 ;
        RECT 260.400 646.950 262.500 649.050 ;
        RECT 265.800 646.950 267.900 649.050 ;
        RECT 253.950 643.950 256.050 646.050 ;
        RECT 257.400 644.400 258.600 646.650 ;
        RECT 266.400 645.450 267.600 646.650 ;
        RECT 269.400 645.450 270.450 655.950 ;
        RECT 266.400 644.400 270.450 645.450 ;
        RECT 257.400 640.050 258.450 644.400 ;
        RECT 262.950 640.950 265.050 643.050 ;
        RECT 256.950 637.950 259.050 640.050 ;
        RECT 259.950 610.950 262.050 613.050 ;
        RECT 250.950 607.950 253.050 610.050 ;
        RECT 260.400 607.200 261.450 610.950 ;
        RECT 242.400 604.350 243.600 606.000 ;
        RECT 248.400 604.350 249.600 606.600 ;
        RECT 253.950 605.100 256.050 607.200 ;
        RECT 259.950 605.100 262.050 607.200 ;
        RECT 254.400 604.350 255.600 605.100 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 226.950 580.950 229.050 583.050 ;
        RECT 206.400 571.350 207.600 572.100 ;
        RECT 212.400 571.350 213.600 573.600 ;
        RECT 223.950 571.950 226.050 574.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 179.400 559.050 180.450 566.400 ;
        RECT 185.400 564.300 186.450 566.400 ;
        RECT 190.950 565.800 193.050 567.900 ;
        RECT 196.800 565.800 198.900 567.900 ;
        RECT 199.950 565.950 202.050 568.050 ;
        RECT 202.950 565.950 205.050 568.050 ;
        RECT 209.400 567.900 210.600 568.650 ;
        RECT 190.950 564.300 193.050 564.750 ;
        RECT 185.400 563.250 193.050 564.300 ;
        RECT 190.950 562.650 193.050 563.250 ;
        RECT 193.950 562.950 196.050 565.050 ;
        RECT 178.950 556.950 181.050 559.050 ;
        RECT 187.800 556.950 189.900 559.050 ;
        RECT 190.950 556.950 193.050 559.050 ;
        RECT 179.400 544.050 180.450 556.950 ;
        RECT 178.950 541.950 181.050 544.050 ;
        RECT 184.950 538.950 187.050 541.050 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 178.950 528.000 181.050 532.050 ;
        RECT 185.400 528.600 186.450 538.950 ;
        RECT 188.400 529.050 189.450 556.950 ;
        RECT 179.400 526.350 180.600 528.000 ;
        RECT 185.400 526.350 186.600 528.600 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 176.400 521.400 177.600 523.650 ;
        RECT 182.400 522.900 183.600 523.650 ;
        RECT 191.400 523.050 192.450 556.950 ;
        RECT 194.400 556.050 195.450 562.950 ;
        RECT 193.950 553.950 196.050 556.050 ;
        RECT 203.400 544.050 204.450 565.950 ;
        RECT 208.950 565.800 211.050 567.900 ;
        RECT 215.400 566.400 216.600 568.650 ;
        RECT 227.400 568.050 228.450 580.950 ;
        RECT 233.400 580.050 234.450 598.950 ;
        RECT 235.950 598.800 238.050 600.900 ;
        RECT 245.400 599.400 246.600 601.650 ;
        RECT 251.400 600.000 252.600 601.650 ;
        RECT 245.400 595.050 246.450 599.400 ;
        RECT 250.950 595.950 253.050 600.000 ;
        RECT 253.950 595.950 256.050 598.050 ;
        RECT 244.950 592.950 247.050 595.050 ;
        RECT 250.950 589.950 253.050 592.050 ;
        RECT 235.950 583.950 238.050 586.050 ;
        RECT 236.400 580.050 237.450 583.950 ;
        RECT 232.800 577.950 234.900 580.050 ;
        RECT 235.950 577.950 238.050 580.050 ;
        RECT 238.950 579.000 241.050 583.050 ;
        RECT 239.400 577.200 240.600 579.000 ;
        RECT 234.900 573.900 237.000 575.700 ;
        RECT 238.800 574.800 240.900 576.900 ;
        RECT 242.100 576.300 244.200 578.400 ;
        RECT 233.400 572.700 242.100 573.900 ;
        RECT 230.100 568.950 232.200 571.050 ;
        RECT 209.400 564.450 210.450 565.800 ;
        RECT 215.400 564.450 216.450 566.400 ;
        RECT 220.950 565.800 223.050 567.900 ;
        RECT 226.950 565.950 229.050 568.050 ;
        RECT 230.400 567.900 231.600 568.650 ;
        RECT 229.950 565.800 232.050 567.900 ;
        RECT 206.400 563.400 210.450 564.450 ;
        RECT 212.400 563.400 216.450 564.450 ;
        RECT 202.950 541.950 205.050 544.050 ;
        RECT 196.950 538.950 199.050 541.050 ;
        RECT 197.400 528.600 198.450 538.950 ;
        RECT 202.950 535.950 205.050 538.050 ;
        RECT 203.400 528.600 204.450 535.950 ;
        RECT 206.400 535.050 207.450 563.400 ;
        RECT 212.400 553.050 213.450 563.400 ;
        RECT 221.400 559.050 222.450 565.800 ;
        RECT 233.400 563.700 234.300 572.700 ;
        RECT 240.000 571.800 242.100 572.700 ;
        RECT 243.000 570.900 243.900 576.300 ;
        RECT 245.400 573.450 246.600 573.600 ;
        RECT 245.400 572.400 249.450 573.450 ;
        RECT 245.400 571.350 246.600 572.400 ;
        RECT 237.000 569.700 243.900 570.900 ;
        RECT 237.000 567.300 237.900 569.700 ;
        RECT 235.800 565.200 237.900 567.300 ;
        RECT 238.800 565.950 240.900 568.050 ;
        RECT 232.500 561.600 234.600 563.700 ;
        RECT 239.400 563.400 240.600 565.650 ;
        RECT 242.700 562.500 243.900 569.700 ;
        RECT 244.800 568.950 246.900 571.050 ;
        RECT 242.100 560.400 244.200 562.500 ;
        RECT 220.950 556.950 223.050 559.050 ;
        RECT 226.950 556.950 232.050 559.050 ;
        RECT 223.950 553.800 226.050 555.900 ;
        RECT 211.950 550.950 214.050 553.050 ;
        RECT 208.950 544.950 211.050 547.050 ;
        RECT 205.950 532.950 208.050 535.050 ;
        RECT 209.400 529.050 210.450 544.950 ;
        RECT 224.400 532.050 225.450 553.800 ;
        RECT 232.950 550.950 235.050 553.050 ;
        RECT 211.950 529.950 214.050 532.050 ;
        RECT 197.400 526.350 198.600 528.600 ;
        RECT 203.400 526.350 204.600 528.600 ;
        RECT 208.950 526.950 211.050 529.050 ;
        RECT 196.950 523.950 199.050 526.050 ;
        RECT 199.950 523.950 202.050 526.050 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 176.400 508.050 177.450 521.400 ;
        RECT 181.950 520.800 184.050 522.900 ;
        RECT 187.950 520.950 190.050 523.050 ;
        RECT 190.950 520.950 193.050 523.050 ;
        RECT 200.400 521.400 201.600 523.650 ;
        RECT 206.400 522.900 207.600 523.650 ;
        RECT 178.950 517.950 181.050 520.050 ;
        RECT 175.950 505.950 178.050 508.050 ;
        RECT 169.950 502.950 172.050 505.050 ;
        RECT 163.950 497.400 168.450 498.450 ;
        RECT 163.950 496.950 166.050 497.400 ;
        RECT 164.400 495.600 165.450 496.950 ;
        RECT 164.400 493.350 165.600 495.600 ;
        RECT 169.950 494.100 172.050 496.200 ;
        RECT 170.400 493.350 171.600 494.100 ;
        RECT 175.950 493.950 178.050 499.050 ;
        RECT 163.950 490.950 166.050 493.050 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 160.950 487.950 163.050 490.050 ;
        RECT 167.400 488.400 168.600 490.650 ;
        RECT 173.400 488.400 174.600 490.650 ;
        RECT 179.400 490.050 180.450 517.950 ;
        RECT 184.950 514.950 187.050 517.050 ;
        RECT 185.400 510.450 186.450 514.950 ;
        RECT 188.400 514.050 189.450 520.950 ;
        RECT 200.400 517.050 201.450 521.400 ;
        RECT 205.950 520.800 208.050 522.900 ;
        RECT 212.400 517.050 213.450 529.950 ;
        RECT 217.950 528.000 220.050 532.050 ;
        RECT 223.950 529.950 226.050 532.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 225.000 528.600 229.050 529.050 ;
        RECT 218.400 526.350 219.600 528.000 ;
        RECT 224.400 526.950 229.050 528.600 ;
        RECT 224.400 526.350 225.600 526.950 ;
        RECT 217.950 523.950 220.050 526.050 ;
        RECT 220.950 523.950 223.050 526.050 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 221.400 522.900 222.600 523.650 ;
        RECT 220.950 520.800 223.050 522.900 ;
        RECT 226.950 520.950 229.050 523.050 ;
        RECT 199.950 514.950 202.050 517.050 ;
        RECT 211.950 514.950 214.050 517.050 ;
        RECT 187.950 511.950 190.050 514.050 ;
        RECT 190.950 510.450 193.050 511.050 ;
        RECT 185.400 509.400 193.050 510.450 ;
        RECT 190.950 508.950 193.050 509.400 ;
        RECT 211.950 510.450 216.000 511.050 ;
        RECT 211.950 508.950 216.450 510.450 ;
        RECT 181.950 502.950 184.050 505.050 ;
        RECT 211.950 502.950 214.050 505.050 ;
        RECT 182.400 499.050 183.450 502.950 ;
        RECT 190.950 499.950 193.050 502.050 ;
        RECT 202.950 499.950 205.050 502.050 ;
        RECT 181.950 496.950 184.050 499.050 ;
        RECT 145.950 445.950 148.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 149.400 444.900 150.600 445.650 ;
        RECT 148.950 442.800 151.050 444.900 ;
        RECT 139.950 439.950 142.050 442.050 ;
        RECT 145.950 439.950 148.050 442.050 ;
        RECT 134.400 425.400 138.450 426.450 ;
        RECT 134.400 424.050 135.450 425.400 ;
        RECT 133.950 421.950 136.050 424.050 ;
        RECT 134.400 411.450 135.450 421.950 ;
        RECT 142.950 417.000 145.050 421.050 ;
        RECT 143.400 415.350 144.600 417.000 ;
        RECT 137.100 412.950 139.200 415.050 ;
        RECT 142.500 412.950 144.600 415.050 ;
        RECT 137.400 411.450 138.600 412.650 ;
        RECT 134.400 410.400 138.600 411.450 ;
        RECT 146.400 409.050 147.450 439.950 ;
        RECT 161.400 433.050 162.450 487.950 ;
        RECT 167.400 457.050 168.450 488.400 ;
        RECT 173.400 478.050 174.450 488.400 ;
        RECT 178.800 487.950 180.900 490.050 ;
        RECT 182.400 489.900 183.450 496.950 ;
        RECT 191.400 495.600 192.450 499.950 ;
        RECT 191.400 493.350 192.600 495.600 ;
        RECT 196.950 494.100 199.050 496.200 ;
        RECT 197.400 493.350 198.600 494.100 ;
        RECT 187.950 490.950 190.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 188.400 489.900 189.600 490.650 ;
        RECT 181.950 487.800 184.050 489.900 ;
        RECT 187.950 487.800 190.050 489.900 ;
        RECT 194.400 489.000 195.600 490.650 ;
        RECT 193.950 484.950 196.050 489.000 ;
        RECT 175.950 481.950 178.050 484.050 ;
        RECT 172.950 475.950 175.050 478.050 ;
        RECT 176.400 475.050 177.450 481.950 ;
        RECT 175.950 472.950 178.050 475.050 ;
        RECT 187.950 472.950 190.050 475.050 ;
        RECT 178.950 466.950 181.050 469.050 ;
        RECT 166.950 454.950 169.050 457.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 170.400 444.900 171.600 445.650 ;
        RECT 169.950 442.800 172.050 444.900 ;
        RECT 179.400 439.050 180.450 466.950 ;
        RECT 188.400 450.600 189.450 472.950 ;
        RECT 203.400 469.050 204.450 499.950 ;
        RECT 212.400 495.600 213.450 502.950 ;
        RECT 215.400 502.050 216.450 508.950 ;
        RECT 214.950 499.950 217.050 502.050 ;
        RECT 212.400 493.350 213.600 495.600 ;
        RECT 217.950 494.100 220.050 496.200 ;
        RECT 218.400 493.350 219.600 494.100 ;
        RECT 211.950 490.950 214.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 215.400 488.400 216.600 490.650 ;
        RECT 221.400 489.900 222.600 490.650 ;
        RECT 227.400 490.050 228.450 520.950 ;
        RECT 230.400 499.050 231.450 529.950 ;
        RECT 233.400 523.050 234.450 550.950 ;
        RECT 248.400 547.050 249.450 572.400 ;
        RECT 251.400 568.050 252.450 589.950 ;
        RECT 250.950 565.950 253.050 568.050 ;
        RECT 247.950 544.950 250.050 547.050 ;
        RECT 235.950 541.950 238.050 544.050 ;
        RECT 236.400 529.050 237.450 541.950 ;
        RECT 235.950 526.950 238.050 529.050 ;
        RECT 241.950 527.100 244.050 529.200 ;
        RECT 249.000 528.600 253.050 529.050 ;
        RECT 242.400 526.350 243.600 527.100 ;
        RECT 248.400 526.950 253.050 528.600 ;
        RECT 248.400 526.350 249.600 526.950 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 244.950 523.950 247.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 239.400 522.900 240.600 523.650 ;
        RECT 238.950 520.800 241.050 522.900 ;
        RECT 245.400 521.400 246.600 523.650 ;
        RECT 232.950 514.950 235.050 517.050 ;
        RECT 229.950 496.950 232.050 499.050 ;
        RECT 215.400 481.050 216.450 488.400 ;
        RECT 220.950 487.800 223.050 489.900 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 214.950 478.950 217.050 481.050 ;
        RECT 233.400 478.050 234.450 514.950 ;
        RECT 245.400 505.050 246.450 521.400 ;
        RECT 250.950 520.950 253.050 523.050 ;
        RECT 251.400 514.050 252.450 520.950 ;
        RECT 250.950 511.950 253.050 514.050 ;
        RECT 244.950 502.950 247.050 505.050 ;
        RECT 250.950 502.950 253.050 505.050 ;
        RECT 235.950 494.100 238.050 496.200 ;
        RECT 244.950 494.100 247.050 496.200 ;
        RECT 236.400 493.350 237.600 494.100 ;
        RECT 245.400 493.350 246.600 494.100 ;
        RECT 251.400 493.050 252.450 502.950 ;
        RECT 236.100 490.950 238.200 493.050 ;
        RECT 239.100 490.950 241.200 493.050 ;
        RECT 244.800 490.950 246.900 493.050 ;
        RECT 247.800 490.950 249.900 493.050 ;
        RECT 250.950 490.950 253.050 493.050 ;
        RECT 239.400 489.900 240.600 490.650 ;
        RECT 238.950 487.800 241.050 489.900 ;
        RECT 248.400 489.450 249.600 490.650 ;
        RECT 248.400 488.400 252.450 489.450 ;
        RECT 247.950 481.950 250.050 484.050 ;
        RECT 232.950 475.950 235.050 478.050 ;
        RECT 205.950 469.950 208.050 472.050 ;
        RECT 226.950 469.950 229.050 472.050 ;
        RECT 241.950 469.950 244.050 472.050 ;
        RECT 196.950 466.950 199.050 469.050 ;
        RECT 202.950 466.950 205.050 469.050 ;
        RECT 197.400 457.050 198.450 466.950 ;
        RECT 206.400 460.050 207.450 469.950 ;
        RECT 227.400 466.050 228.450 469.950 ;
        RECT 238.950 466.950 241.050 469.050 ;
        RECT 223.800 463.950 225.900 466.050 ;
        RECT 226.950 463.950 229.050 466.050 ;
        RECT 205.800 457.950 207.900 460.050 ;
        RECT 208.950 457.950 211.050 460.050 ;
        RECT 196.950 454.950 199.050 457.050 ;
        RECT 188.400 448.350 189.600 450.600 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 197.400 444.900 198.450 454.950 ;
        RECT 202.950 449.100 205.050 451.200 ;
        RECT 209.400 450.600 210.450 457.950 ;
        RECT 224.400 451.200 225.450 463.950 ;
        RECT 203.400 448.350 204.600 449.100 ;
        RECT 209.400 448.350 210.600 450.600 ;
        RECT 214.950 449.100 217.050 451.200 ;
        RECT 220.800 449.100 222.900 451.200 ;
        RECT 223.950 449.100 226.050 451.200 ;
        RECT 229.950 449.100 232.050 451.200 ;
        RECT 235.950 449.100 238.050 451.200 ;
        RECT 239.400 451.050 240.450 466.950 ;
        RECT 242.400 466.050 243.450 469.950 ;
        RECT 241.950 463.950 244.050 466.050 ;
        RECT 215.400 448.350 216.600 449.100 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 205.950 445.950 208.050 448.050 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 211.950 445.950 214.050 448.050 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 206.400 444.900 207.600 445.650 ;
        RECT 196.950 442.800 199.050 444.900 ;
        RECT 205.950 442.800 208.050 444.900 ;
        RECT 212.400 443.400 213.600 445.650 ;
        RECT 221.400 445.050 222.450 449.100 ;
        RECT 230.400 448.350 231.600 449.100 ;
        RECT 236.400 448.350 237.600 449.100 ;
        RECT 238.950 448.950 241.050 451.050 ;
        RECT 241.950 449.100 244.050 451.200 ;
        RECT 248.400 451.050 249.450 481.950 ;
        RECT 251.400 466.050 252.450 488.400 ;
        RECT 254.400 484.050 255.450 595.950 ;
        RECT 260.400 592.050 261.450 605.100 ;
        RECT 263.400 598.050 264.450 640.950 ;
        RECT 266.400 637.050 267.450 644.400 ;
        RECT 265.950 634.950 268.050 637.050 ;
        RECT 272.400 628.050 273.450 673.950 ;
        RECT 271.950 625.950 274.050 628.050 ;
        RECT 275.400 622.050 276.450 673.950 ;
        RECT 277.950 673.800 280.050 673.950 ;
        RECT 280.950 667.950 283.050 670.050 ;
        RECT 281.400 651.600 282.450 667.950 ;
        RECT 284.400 654.450 285.450 718.950 ;
        RECT 287.400 712.050 288.450 722.400 ;
        RECT 292.950 721.950 295.050 724.050 ;
        RECT 286.950 709.950 289.050 712.050 ;
        RECT 289.950 700.950 292.050 703.050 ;
        RECT 286.950 682.950 289.050 685.050 ;
        RECT 290.400 684.600 291.450 700.950 ;
        RECT 293.400 691.050 294.450 721.950 ;
        RECT 296.400 718.050 297.450 748.950 ;
        RECT 299.400 733.050 300.450 751.950 ;
        RECT 302.400 736.050 303.450 775.950 ;
        RECT 304.800 761.100 306.900 763.200 ;
        RECT 308.400 763.050 309.450 785.400 ;
        RECT 335.400 766.050 336.450 800.400 ;
        RECT 340.950 799.800 343.050 801.900 ;
        RECT 346.950 799.800 349.050 801.900 ;
        RECT 353.400 800.400 354.600 802.650 ;
        RECT 353.400 790.050 354.450 800.400 ;
        RECT 352.950 787.950 355.050 790.050 ;
        RECT 343.950 769.950 346.050 772.050 ;
        RECT 355.950 769.950 358.050 772.050 ;
        RECT 305.400 757.050 306.450 761.100 ;
        RECT 307.950 760.950 310.050 763.050 ;
        RECT 313.950 762.000 316.050 766.050 ;
        RECT 334.950 763.950 337.050 766.050 ;
        RECT 314.400 760.350 315.600 762.000 ;
        RECT 319.950 761.100 322.050 763.200 ;
        RECT 325.950 761.100 328.050 763.200 ;
        RECT 337.950 761.100 340.050 763.200 ;
        RECT 320.400 760.350 321.600 761.100 ;
        RECT 310.950 757.950 313.050 760.050 ;
        RECT 313.950 757.950 316.050 760.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 304.950 754.950 307.050 757.050 ;
        RECT 307.950 754.950 310.050 757.050 ;
        RECT 311.400 756.900 312.600 757.650 ;
        RECT 308.400 739.050 309.450 754.950 ;
        RECT 310.950 754.800 313.050 756.900 ;
        RECT 317.400 755.400 318.600 757.650 ;
        RECT 326.400 757.050 327.450 761.100 ;
        RECT 338.400 760.350 339.600 761.100 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 317.400 745.050 318.450 755.400 ;
        RECT 325.950 754.950 328.050 757.050 ;
        RECT 335.400 756.900 336.600 757.650 ;
        RECT 334.950 754.800 337.050 756.900 ;
        RECT 322.950 748.950 325.050 751.050 ;
        RECT 323.400 745.050 324.450 748.950 ;
        RECT 316.950 742.950 319.050 745.050 ;
        RECT 322.950 742.950 325.050 745.050 ;
        RECT 319.950 739.950 322.050 742.050 ;
        RECT 307.950 736.950 310.050 739.050 ;
        RECT 316.950 736.950 319.050 739.050 ;
        RECT 301.950 733.950 304.050 736.050 ;
        RECT 298.950 730.950 301.050 733.050 ;
        RECT 304.950 732.450 309.000 733.050 ;
        RECT 304.950 730.950 309.450 732.450 ;
        RECT 295.950 715.950 298.050 718.050 ;
        RECT 292.950 688.950 295.050 691.050 ;
        RECT 287.400 658.050 288.450 682.950 ;
        RECT 290.400 682.350 291.600 684.600 ;
        RECT 290.100 679.950 292.200 682.050 ;
        RECT 295.500 679.950 297.600 682.050 ;
        RECT 296.400 677.400 297.600 679.650 ;
        RECT 296.400 667.050 297.450 677.400 ;
        RECT 299.400 670.050 300.450 730.950 ;
        RECT 308.400 729.600 309.450 730.950 ;
        RECT 308.400 727.350 309.600 729.600 ;
        RECT 313.950 727.950 316.050 733.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 301.950 721.950 304.050 724.050 ;
        RECT 305.400 722.400 306.600 724.650 ;
        RECT 311.400 722.400 312.600 724.650 ;
        RECT 298.950 667.950 301.050 670.050 ;
        RECT 295.950 664.950 298.050 667.050 ;
        RECT 286.950 655.950 289.050 658.050 ;
        RECT 284.400 653.400 288.450 654.450 ;
        RECT 287.400 652.200 288.450 653.400 ;
        RECT 281.400 649.350 282.600 651.600 ;
        RECT 286.950 650.100 289.050 652.200 ;
        RECT 287.400 649.350 288.600 650.100 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 284.400 645.000 285.600 646.650 ;
        RECT 277.950 640.950 280.050 643.050 ;
        RECT 283.950 640.950 286.050 645.000 ;
        RECT 290.400 644.400 291.600 646.650 ;
        RECT 274.950 619.950 277.050 622.050 ;
        RECT 268.950 605.100 271.050 607.200 ;
        RECT 269.400 604.350 270.600 605.100 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 272.400 601.050 273.600 601.650 ;
        RECT 262.950 595.950 265.050 598.050 ;
        RECT 265.950 595.950 268.050 601.050 ;
        RECT 272.400 598.950 277.050 601.050 ;
        RECT 259.950 589.950 262.050 592.050 ;
        RECT 259.950 583.950 262.050 586.050 ;
        RECT 260.400 573.600 261.450 583.950 ;
        RECT 266.400 573.600 267.450 595.950 ;
        RECT 272.400 574.050 273.450 598.950 ;
        RECT 274.950 595.800 277.050 597.900 ;
        RECT 275.400 582.450 276.450 595.800 ;
        RECT 278.400 586.050 279.450 640.950 ;
        RECT 286.950 637.950 289.050 640.050 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 281.400 628.050 282.450 631.950 ;
        RECT 280.950 625.950 283.050 628.050 ;
        RECT 280.950 619.950 283.050 622.050 ;
        RECT 281.400 601.050 282.450 619.950 ;
        RECT 287.400 609.450 288.450 637.950 ;
        RECT 290.400 637.050 291.450 644.400 ;
        RECT 292.950 643.950 295.050 646.050 ;
        RECT 289.950 634.950 292.050 637.050 ;
        RECT 284.400 609.000 288.450 609.450 ;
        RECT 283.950 608.400 288.450 609.000 ;
        RECT 283.950 604.950 286.050 608.400 ;
        RECT 289.950 605.100 292.050 607.200 ;
        RECT 293.400 607.050 294.450 643.950 ;
        RECT 296.400 619.050 297.450 664.950 ;
        RECT 298.950 655.950 301.050 658.050 ;
        RECT 295.950 616.950 298.050 619.050 ;
        RECT 290.400 604.350 291.600 605.100 ;
        RECT 292.950 604.950 295.050 607.050 ;
        RECT 299.400 606.450 300.450 655.950 ;
        RECT 302.400 655.050 303.450 721.950 ;
        RECT 305.400 703.050 306.450 722.400 ;
        RECT 311.400 718.050 312.450 722.400 ;
        RECT 310.950 715.950 313.050 718.050 ;
        RECT 304.950 700.950 307.050 703.050 ;
        RECT 307.950 688.950 310.050 691.050 ;
        RECT 304.950 682.950 307.050 688.050 ;
        RECT 308.400 684.600 309.450 688.950 ;
        RECT 311.400 687.450 312.450 715.950 ;
        RECT 313.950 712.950 316.050 715.050 ;
        RECT 314.400 703.050 315.450 712.950 ;
        RECT 317.400 712.050 318.450 736.950 ;
        RECT 320.400 733.050 321.450 739.950 ;
        RECT 328.950 733.950 331.050 736.050 ;
        RECT 319.950 730.950 322.050 733.050 ;
        RECT 319.950 727.800 322.050 729.900 ;
        RECT 329.400 729.600 330.450 733.950 ;
        RECT 335.400 730.050 336.450 754.800 ;
        RECT 344.400 739.050 345.450 769.950 ;
        RECT 356.400 762.600 357.450 769.950 ;
        RECT 356.400 760.350 357.600 762.600 ;
        RECT 350.400 757.950 352.500 760.050 ;
        RECT 355.800 757.950 357.900 760.050 ;
        RECT 350.400 756.900 351.600 757.650 ;
        RECT 349.950 754.800 352.050 756.900 ;
        RECT 358.950 754.800 361.050 756.900 ;
        RECT 346.950 745.950 349.050 748.050 ;
        RECT 337.950 736.950 340.050 739.050 ;
        RECT 343.950 736.950 346.050 739.050 ;
        RECT 320.400 724.050 321.450 727.800 ;
        RECT 329.400 727.350 330.600 729.600 ;
        RECT 334.950 727.950 337.050 730.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 331.950 724.950 334.050 727.050 ;
        RECT 319.950 721.950 322.050 724.050 ;
        RECT 326.400 723.900 327.600 724.650 ;
        RECT 332.400 723.900 333.600 724.650 ;
        RECT 325.950 721.800 328.050 723.900 ;
        RECT 331.950 721.800 334.050 723.900 ;
        RECT 338.400 718.050 339.450 736.950 ;
        RECT 340.950 733.950 343.050 736.050 ;
        RECT 341.400 730.050 342.450 733.950 ;
        RECT 340.950 727.950 343.050 730.050 ;
        RECT 347.400 729.600 348.450 745.950 ;
        RECT 352.950 736.950 355.050 739.050 ;
        RECT 353.400 733.050 354.450 736.950 ;
        RECT 352.950 730.950 355.050 733.050 ;
        RECT 353.400 729.600 354.450 730.950 ;
        RECT 347.400 727.350 348.600 729.600 ;
        RECT 353.400 727.350 354.600 729.600 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 346.950 724.950 349.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 340.950 721.950 343.050 724.050 ;
        RECT 344.400 723.900 345.600 724.650 ;
        RECT 325.950 715.950 331.050 718.050 ;
        RECT 337.950 715.950 340.050 718.050 ;
        RECT 328.950 712.800 331.050 714.900 ;
        RECT 341.400 714.450 342.450 721.950 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 350.400 722.400 351.600 724.650 ;
        RECT 350.400 715.050 351.450 722.400 ;
        RECT 338.400 713.400 342.450 714.450 ;
        RECT 316.950 709.950 319.050 712.050 ;
        RECT 313.950 700.950 316.050 703.050 ;
        RECT 311.400 686.400 315.450 687.450 ;
        RECT 314.400 684.600 315.450 686.400 ;
        RECT 308.400 682.350 309.600 684.600 ;
        RECT 314.400 682.350 315.600 684.600 ;
        RECT 323.100 682.950 325.200 685.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 323.400 680.400 324.600 682.650 ;
        RECT 329.400 682.050 330.450 712.800 ;
        RECT 332.100 682.950 334.200 685.050 ;
        RECT 311.400 678.900 312.600 679.650 ;
        RECT 317.400 678.900 318.600 679.650 ;
        RECT 304.950 673.950 307.050 678.900 ;
        RECT 310.950 676.800 313.050 678.900 ;
        RECT 316.950 676.800 319.050 678.900 ;
        RECT 317.400 673.050 318.450 676.800 ;
        RECT 313.950 671.400 318.450 673.050 ;
        RECT 313.950 670.950 318.000 671.400 ;
        RECT 319.950 667.950 322.050 670.050 ;
        RECT 320.400 655.050 321.450 667.950 ;
        RECT 323.400 667.050 324.450 680.400 ;
        RECT 328.950 679.950 331.050 682.050 ;
        RECT 332.400 680.400 333.600 682.650 ;
        RECT 322.950 664.950 325.050 667.050 ;
        RECT 332.400 664.050 333.450 680.400 ;
        RECT 338.400 667.050 339.450 713.400 ;
        RECT 349.950 712.950 352.050 715.050 ;
        RECT 341.700 696.300 343.800 698.400 ;
        RECT 342.300 691.500 343.800 696.300 ;
        RECT 341.700 689.400 343.800 691.500 ;
        RECT 342.300 671.700 343.800 689.400 ;
        RECT 341.700 669.600 343.800 671.700 ;
        RECT 344.700 693.300 346.800 698.400 ;
        RECT 347.700 696.300 349.800 698.400 ;
        RECT 359.400 697.050 360.450 754.800 ;
        RECT 362.400 739.050 363.450 806.100 ;
        RECT 365.400 801.450 366.450 833.400 ;
        RECT 370.950 829.950 373.050 834.000 ;
        RECT 377.400 832.050 378.450 884.100 ;
        RECT 380.400 880.050 381.450 886.950 ;
        RECT 389.400 885.600 390.450 895.950 ;
        RECT 389.400 883.350 390.600 885.600 ;
        RECT 385.950 880.950 388.050 883.050 ;
        RECT 388.950 880.950 391.050 883.050 ;
        RECT 379.950 877.950 382.050 880.050 ;
        RECT 386.400 879.000 387.600 880.650 ;
        RECT 385.950 874.950 388.050 879.000 ;
        RECT 398.400 877.050 399.450 910.950 ;
        RECT 406.950 901.950 409.050 904.050 ;
        RECT 407.400 885.600 408.450 901.950 ;
        RECT 413.400 901.050 414.450 920.100 ;
        RECT 437.100 916.950 439.200 919.050 ;
        RECT 425.400 913.950 427.500 916.050 ;
        RECT 430.800 913.950 432.900 916.050 ;
        RECT 437.400 914.400 438.600 916.650 ;
        RECT 443.400 915.450 444.450 928.950 ;
        RECT 456.300 925.500 457.800 930.300 ;
        RECT 455.700 923.400 457.800 925.500 ;
        RECT 446.100 916.950 448.200 919.050 ;
        RECT 446.400 915.450 447.600 916.650 ;
        RECT 443.400 914.400 447.600 915.450 ;
        RECT 425.400 911.400 426.600 913.650 ;
        RECT 412.950 898.950 415.050 901.050 ;
        RECT 425.400 898.050 426.450 911.400 ;
        RECT 427.950 901.950 430.050 904.050 ;
        RECT 424.950 895.950 427.050 898.050 ;
        RECT 407.400 883.350 408.600 885.600 ;
        RECT 412.950 884.100 415.050 886.200 ;
        RECT 421.950 884.100 424.050 886.200 ;
        RECT 428.400 886.050 429.450 901.950 ;
        RECT 437.400 898.050 438.450 914.400 ;
        RECT 436.950 895.950 439.050 898.050 ;
        RECT 413.400 883.350 414.600 884.100 ;
        RECT 403.950 880.950 406.050 883.050 ;
        RECT 406.950 880.950 409.050 883.050 ;
        RECT 409.950 880.950 412.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 404.400 878.400 405.600 880.650 ;
        RECT 410.400 879.000 411.600 880.650 ;
        RECT 397.950 874.950 400.050 877.050 ;
        RECT 404.400 874.050 405.450 878.400 ;
        RECT 409.950 874.950 412.050 879.000 ;
        RECT 416.400 878.400 417.600 880.650 ;
        RECT 422.400 879.450 423.450 884.100 ;
        RECT 427.950 883.950 430.050 886.050 ;
        RECT 419.400 878.400 423.450 879.450 ;
        RECT 403.950 871.950 406.050 874.050 ;
        RECT 409.950 868.950 412.050 871.050 ;
        RECT 410.400 865.050 411.450 868.950 ;
        RECT 409.950 862.950 412.050 865.050 ;
        RECT 394.950 847.950 397.050 850.050 ;
        RECT 406.950 847.950 409.050 850.050 ;
        RECT 385.950 839.100 388.050 841.200 ;
        RECT 386.400 838.350 387.600 839.100 ;
        RECT 395.400 838.050 396.450 847.950 ;
        RECT 397.950 841.950 400.050 844.050 ;
        RECT 382.950 835.950 385.050 838.050 ;
        RECT 385.950 835.950 388.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 394.950 835.950 397.050 838.050 ;
        RECT 383.400 834.900 384.600 835.650 ;
        RECT 382.950 832.800 385.050 834.900 ;
        RECT 389.400 833.400 390.600 835.650 ;
        RECT 389.400 832.050 390.450 833.400 ;
        RECT 398.400 832.050 399.450 841.950 ;
        RECT 407.400 840.600 408.450 847.950 ;
        RECT 407.400 838.350 408.600 840.600 ;
        RECT 403.950 835.950 406.050 838.050 ;
        RECT 406.950 835.950 409.050 838.050 ;
        RECT 409.950 835.950 412.050 838.050 ;
        RECT 404.400 833.400 405.600 835.650 ;
        RECT 410.400 834.900 411.600 835.650 ;
        RECT 376.950 829.950 379.050 832.050 ;
        RECT 388.950 831.450 391.050 832.050 ;
        RECT 386.400 830.400 391.050 831.450 ;
        RECT 373.950 817.950 376.050 820.050 ;
        RECT 379.950 817.950 382.050 820.050 ;
        RECT 374.400 807.600 375.450 817.950 ;
        RECT 380.400 807.600 381.450 817.950 ;
        RECT 374.400 805.350 375.600 807.600 ;
        RECT 380.400 805.350 381.600 807.600 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 365.400 800.400 369.450 801.450 ;
        RECT 368.400 796.050 369.450 800.400 ;
        RECT 371.400 800.400 372.600 802.650 ;
        RECT 377.400 800.400 378.600 802.650 ;
        RECT 367.950 793.950 370.050 796.050 ;
        RECT 371.400 769.050 372.450 800.400 ;
        RECT 377.400 787.050 378.450 800.400 ;
        RECT 382.950 799.950 385.050 802.050 ;
        RECT 379.950 796.950 382.050 799.050 ;
        RECT 376.950 784.950 379.050 787.050 ;
        RECT 370.950 766.950 373.050 769.050 ;
        RECT 370.950 761.100 373.050 763.200 ;
        RECT 371.400 760.350 372.600 761.100 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 374.400 756.900 375.600 757.650 ;
        RECT 373.950 754.800 376.050 756.900 ;
        RECT 380.400 754.050 381.450 796.950 ;
        RECT 383.400 763.050 384.450 799.950 ;
        RECT 386.400 766.050 387.450 830.400 ;
        RECT 388.950 829.950 391.050 830.400 ;
        RECT 397.950 829.950 400.050 832.050 ;
        RECT 397.950 826.800 400.050 828.900 ;
        RECT 398.400 814.050 399.450 826.800 ;
        RECT 397.950 811.950 400.050 814.050 ;
        RECT 394.950 807.000 397.050 811.050 ;
        RECT 404.400 808.050 405.450 833.400 ;
        RECT 409.950 832.800 412.050 834.900 ;
        RECT 416.400 832.050 417.450 878.400 ;
        RECT 419.400 834.450 420.450 878.400 ;
        RECT 428.400 859.050 429.450 883.950 ;
        RECT 433.800 880.950 435.900 883.050 ;
        RECT 439.800 880.950 441.900 883.050 ;
        RECT 434.400 879.000 435.600 880.650 ;
        RECT 433.950 874.950 436.050 879.000 ;
        RECT 433.950 862.950 436.050 865.050 ;
        RECT 430.950 859.950 433.050 862.050 ;
        RECT 427.950 856.950 430.050 859.050 ;
        RECT 421.950 840.600 426.000 841.050 ;
        RECT 431.400 840.600 432.450 859.950 ;
        RECT 434.400 844.050 435.450 862.950 ;
        RECT 439.950 850.950 442.050 853.050 ;
        RECT 433.950 841.950 436.050 844.050 ;
        RECT 421.950 838.950 426.600 840.600 ;
        RECT 425.400 838.350 426.600 838.950 ;
        RECT 431.400 838.350 432.600 840.600 ;
        RECT 436.950 839.100 439.050 841.200 ;
        RECT 440.400 841.050 441.450 850.950 ;
        RECT 446.400 847.050 447.450 914.400 ;
        RECT 448.950 914.100 451.050 916.200 ;
        RECT 449.400 892.050 450.450 914.100 ;
        RECT 456.300 905.700 457.800 923.400 ;
        RECT 455.700 903.600 457.800 905.700 ;
        RECT 458.700 927.300 460.800 932.400 ;
        RECT 461.700 930.300 463.800 932.400 ;
        RECT 480.600 930.300 482.700 932.400 ;
        RECT 483.600 930.300 486.600 932.400 ;
        RECT 458.700 905.700 459.900 927.300 ;
        RECT 461.700 925.500 463.200 930.300 ;
        RECT 464.100 927.300 466.200 929.400 ;
        RECT 461.100 923.400 463.200 925.500 ;
        RECT 461.700 905.700 463.200 923.400 ;
        RECT 464.700 920.100 465.900 927.300 ;
        RECT 469.500 925.800 471.600 927.900 ;
        RECT 478.200 927.300 480.300 929.400 ;
        RECT 464.100 918.000 466.200 920.100 ;
        RECT 470.700 919.200 471.600 925.800 ;
        RECT 464.700 905.700 465.900 918.000 ;
        RECT 469.500 917.100 471.600 919.200 ;
        RECT 466.800 910.500 468.900 912.600 ;
        RECT 470.700 906.600 471.600 917.100 ;
        RECT 472.950 914.100 475.050 916.200 ;
        RECT 473.400 913.350 474.600 914.100 ;
        RECT 473.100 910.950 475.200 913.050 ;
        RECT 458.700 903.600 460.800 905.700 ;
        RECT 461.700 903.600 463.800 905.700 ;
        RECT 464.700 903.600 466.800 905.700 ;
        RECT 470.100 904.500 472.200 906.600 ;
        RECT 479.100 905.700 480.300 927.300 ;
        RECT 481.500 924.300 482.700 930.300 ;
        RECT 481.500 922.200 483.600 924.300 ;
        RECT 481.500 905.700 482.700 922.200 ;
        RECT 485.100 911.400 486.600 930.300 ;
        RECT 518.400 930.300 521.400 932.400 ;
        RECT 522.300 930.300 524.400 932.400 ;
        RECT 541.200 930.300 543.300 932.400 ;
        RECT 496.950 920.100 499.050 922.200 ;
        RECT 505.950 920.100 508.050 922.200 ;
        RECT 497.400 919.350 498.600 920.100 ;
        RECT 506.400 919.350 507.600 920.100 ;
        RECT 491.100 916.950 493.200 919.050 ;
        RECT 497.100 916.950 499.200 919.050 ;
        RECT 505.800 916.950 507.900 919.050 ;
        RECT 511.800 916.950 513.900 919.050 ;
        RECT 493.950 913.950 496.050 916.050 ;
        RECT 484.500 909.300 486.600 911.400 ;
        RECT 490.950 910.950 493.050 913.050 ;
        RECT 484.500 905.700 485.700 909.300 ;
        RECT 478.200 903.600 480.300 905.700 ;
        RECT 481.200 903.600 483.300 905.700 ;
        RECT 484.200 903.600 486.300 905.700 ;
        RECT 454.950 898.950 457.050 901.050 ;
        RECT 448.950 889.950 451.050 892.050 ;
        RECT 455.400 879.450 456.450 898.950 ;
        RECT 491.400 898.050 492.450 910.950 ;
        RECT 494.400 901.050 495.450 913.950 ;
        RECT 518.400 911.400 519.900 930.300 ;
        RECT 522.300 924.300 523.500 930.300 ;
        RECT 521.400 922.200 523.500 924.300 ;
        RECT 518.400 909.300 520.500 911.400 ;
        RECT 519.300 905.700 520.500 909.300 ;
        RECT 522.300 905.700 523.500 922.200 ;
        RECT 524.700 927.300 526.800 929.400 ;
        RECT 524.700 905.700 525.900 927.300 ;
        RECT 533.400 925.800 535.500 927.900 ;
        RECT 538.800 927.300 540.900 929.400 ;
        RECT 533.400 919.200 534.300 925.800 ;
        RECT 539.100 920.100 540.300 927.300 ;
        RECT 541.800 925.500 543.300 930.300 ;
        RECT 544.200 927.300 546.300 932.400 ;
        RECT 541.800 923.400 543.900 925.500 ;
        RECT 533.400 917.100 535.500 919.200 ;
        RECT 538.800 918.000 540.900 920.100 ;
        RECT 529.950 914.100 532.050 916.200 ;
        RECT 530.400 913.350 531.600 914.100 ;
        RECT 529.800 910.950 531.900 913.050 ;
        RECT 533.400 906.600 534.300 917.100 ;
        RECT 536.100 910.500 538.200 912.600 ;
        RECT 511.950 901.950 514.050 904.050 ;
        RECT 518.700 903.600 520.800 905.700 ;
        RECT 521.700 903.600 523.800 905.700 ;
        RECT 524.700 903.600 526.800 905.700 ;
        RECT 532.800 904.500 534.900 906.600 ;
        RECT 539.100 905.700 540.300 918.000 ;
        RECT 541.800 905.700 543.300 923.400 ;
        RECT 545.100 905.700 546.300 927.300 ;
        RECT 538.200 903.600 540.300 905.700 ;
        RECT 541.200 903.600 543.300 905.700 ;
        RECT 544.200 903.600 546.300 905.700 ;
        RECT 547.200 930.300 549.300 932.400 ;
        RECT 608.400 930.300 611.400 932.400 ;
        RECT 612.300 930.300 614.400 932.400 ;
        RECT 631.200 930.300 633.300 932.400 ;
        RECT 547.200 925.500 548.700 930.300 ;
        RECT 547.200 923.400 549.300 925.500 ;
        RECT 547.200 905.700 548.700 923.400 ;
        RECT 580.950 919.950 583.050 922.050 ;
        RECT 595.950 920.100 598.050 922.200 ;
        RECT 556.800 916.950 558.900 919.050 ;
        RECT 565.800 916.950 567.900 919.050 ;
        RECT 557.400 915.000 558.600 916.650 ;
        RECT 556.950 910.950 559.050 915.000 ;
        RECT 566.400 914.400 567.600 916.650 ;
        RECT 566.400 910.050 567.450 914.400 ;
        RECT 574.950 914.100 577.050 916.200 ;
        RECT 565.950 907.950 568.050 910.050 ;
        RECT 547.200 903.600 549.300 905.700 ;
        RECT 566.400 904.050 567.450 907.950 ;
        RECT 565.950 901.950 568.050 904.050 ;
        RECT 493.950 898.950 496.050 901.050 ;
        RECT 481.950 895.950 484.050 898.050 ;
        RECT 490.950 895.950 493.050 898.050 ;
        RECT 463.950 891.450 466.050 892.050 ;
        RECT 463.950 890.400 468.450 891.450 ;
        RECT 463.950 889.950 466.050 890.400 ;
        RECT 464.400 885.600 465.450 889.950 ;
        RECT 464.400 883.350 465.600 885.600 ;
        RECT 458.100 880.950 460.200 883.050 ;
        RECT 463.500 880.950 465.600 883.050 ;
        RECT 458.400 879.450 459.600 880.650 ;
        RECT 455.400 878.400 459.600 879.450 ;
        RECT 467.400 877.050 468.450 890.400 ;
        RECT 469.950 884.100 472.050 886.200 ;
        RECT 475.950 884.100 478.050 886.200 ;
        RECT 482.400 885.600 483.450 895.950 ;
        RECT 499.950 894.450 502.050 895.050 ;
        RECT 494.400 893.400 502.050 894.450 ;
        RECT 466.950 874.950 469.050 877.050 ;
        RECT 470.400 874.050 471.450 884.100 ;
        RECT 476.400 883.350 477.600 884.100 ;
        RECT 482.400 883.350 483.600 885.600 ;
        RECT 475.950 880.950 478.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 481.950 880.950 484.050 883.050 ;
        RECT 484.950 880.950 487.050 883.050 ;
        RECT 479.400 878.400 480.600 880.650 ;
        RECT 485.400 879.900 486.600 880.650 ;
        RECT 494.400 879.900 495.450 893.400 ;
        RECT 499.950 892.950 502.050 893.400 ;
        RECT 496.950 889.950 499.050 892.050 ;
        RECT 497.400 886.200 498.450 889.950 ;
        RECT 496.950 884.100 499.050 886.200 ;
        RECT 505.950 884.100 508.050 886.200 ;
        RECT 512.400 886.050 513.450 901.950 ;
        RECT 517.950 892.950 520.050 895.050 ;
        RECT 497.400 883.350 498.600 884.100 ;
        RECT 497.400 880.950 499.500 883.050 ;
        RECT 502.800 880.950 504.900 883.050 ;
        RECT 469.950 871.950 472.050 874.050 ;
        RECT 460.950 868.950 463.050 871.050 ;
        RECT 445.950 844.950 448.050 847.050 ;
        RECT 437.400 838.350 438.600 839.100 ;
        RECT 439.950 838.950 442.050 841.050 ;
        RECT 445.950 838.950 448.050 841.050 ;
        RECT 454.950 839.100 457.050 841.200 ;
        RECT 424.950 835.950 427.050 838.050 ;
        RECT 427.950 835.950 430.050 838.050 ;
        RECT 430.950 835.950 433.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 428.400 834.900 429.600 835.650 ;
        RECT 434.400 834.900 435.600 835.650 ;
        RECT 419.400 833.400 423.450 834.450 ;
        RECT 409.950 826.950 412.050 831.750 ;
        RECT 415.950 829.950 418.050 832.050 ;
        RECT 406.950 814.950 409.050 817.050 ;
        RECT 395.400 805.350 396.600 807.000 ;
        RECT 403.950 805.950 406.050 808.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 398.400 800.400 399.600 802.650 ;
        RECT 398.400 766.050 399.450 800.400 ;
        RECT 407.400 799.050 408.450 814.950 ;
        RECT 415.950 806.100 418.050 808.200 ;
        RECT 422.400 807.600 423.450 833.400 ;
        RECT 427.950 832.800 430.050 834.900 ;
        RECT 433.950 832.800 436.050 834.900 ;
        RECT 439.950 832.950 442.050 835.050 ;
        RECT 446.400 834.900 447.450 838.950 ;
        RECT 455.400 838.350 456.600 839.100 ;
        RECT 451.950 835.950 454.050 838.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 452.400 834.900 453.600 835.650 ;
        RECT 427.950 829.650 430.050 831.750 ;
        RECT 416.400 805.350 417.600 806.100 ;
        RECT 422.400 805.350 423.600 807.600 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 413.400 800.400 414.600 802.650 ;
        RECT 419.400 800.400 420.600 802.650 ;
        RECT 406.950 796.950 409.050 799.050 ;
        RECT 413.400 781.050 414.450 800.400 ;
        RECT 419.400 798.450 420.450 800.400 ;
        RECT 419.400 797.400 423.450 798.450 ;
        RECT 418.950 787.950 421.050 790.050 ;
        RECT 412.950 778.950 415.050 781.050 ;
        RECT 403.950 769.950 406.050 772.050 ;
        RECT 385.950 763.950 388.050 766.050 ;
        RECT 397.950 763.950 400.050 766.050 ;
        RECT 382.950 760.950 385.050 763.050 ;
        RECT 388.950 761.100 391.050 763.200 ;
        RECT 389.400 760.350 390.600 761.100 ;
        RECT 397.950 760.800 400.050 762.900 ;
        RECT 404.400 762.600 405.450 769.950 ;
        RECT 419.400 766.050 420.450 787.950 ;
        RECT 422.400 787.050 423.450 797.400 ;
        RECT 421.950 784.950 424.050 787.050 ;
        RECT 422.400 772.050 423.450 784.950 ;
        RECT 428.400 778.050 429.450 829.650 ;
        RECT 440.400 811.050 441.450 832.950 ;
        RECT 445.950 832.800 448.050 834.900 ;
        RECT 451.950 832.800 454.050 834.900 ;
        RECT 457.950 826.950 460.050 829.050 ;
        RECT 454.950 823.950 457.050 826.050 ;
        RECT 445.950 820.950 448.050 823.050 ;
        RECT 451.950 820.950 454.050 823.050 ;
        RECT 446.400 814.050 447.450 820.950 ;
        RECT 445.950 811.950 448.050 814.050 ;
        RECT 439.950 808.950 442.050 811.050 ;
        RECT 430.950 805.950 433.050 808.050 ;
        RECT 431.400 796.050 432.450 805.950 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 445.950 803.100 448.050 805.200 ;
        RECT 437.400 800.400 438.600 802.650 ;
        RECT 446.400 802.350 447.600 803.100 ;
        RECT 430.950 793.950 433.050 796.050 ;
        RECT 437.400 790.050 438.450 800.400 ;
        RECT 446.100 799.950 448.200 802.050 ;
        RECT 439.950 796.950 442.050 799.050 ;
        RECT 436.950 787.950 439.050 790.050 ;
        RECT 440.400 787.050 441.450 796.950 ;
        RECT 442.950 787.950 445.050 790.050 ;
        RECT 439.950 784.950 442.050 787.050 ;
        RECT 427.950 775.950 430.050 778.050 ;
        RECT 430.950 772.950 433.050 775.050 ;
        RECT 421.950 769.950 424.050 772.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 386.400 757.050 387.600 757.650 ;
        RECT 382.950 755.400 387.600 757.050 ;
        RECT 392.400 757.050 393.600 757.650 ;
        RECT 392.400 755.400 397.050 757.050 ;
        RECT 382.950 754.950 387.450 755.400 ;
        RECT 393.000 754.950 397.050 755.400 ;
        RECT 379.950 751.950 382.050 754.050 ;
        RECT 367.950 739.950 370.050 742.050 ;
        RECT 361.950 736.950 364.050 739.050 ;
        RECT 368.400 732.450 369.450 739.950 ;
        RECT 373.950 736.950 376.050 739.050 ;
        RECT 374.400 733.050 375.450 736.950 ;
        RECT 365.400 731.400 369.450 732.450 ;
        RECT 365.400 729.600 366.450 731.400 ;
        RECT 373.950 730.950 376.050 733.050 ;
        RECT 365.400 727.350 366.600 729.600 ;
        RECT 370.950 728.100 373.050 730.200 ;
        RECT 386.400 730.050 387.450 754.950 ;
        RECT 394.950 751.800 397.050 753.900 ;
        RECT 388.950 736.950 391.050 739.050 ;
        RECT 371.400 727.350 372.600 728.100 ;
        RECT 382.800 727.950 384.900 730.050 ;
        RECT 385.950 727.950 388.050 730.050 ;
        RECT 389.400 729.600 390.450 736.950 ;
        RECT 395.400 729.600 396.450 751.800 ;
        RECT 398.400 732.450 399.450 760.800 ;
        RECT 404.400 760.350 405.600 762.600 ;
        RECT 409.950 762.000 412.050 766.050 ;
        RECT 415.950 763.950 418.050 766.050 ;
        RECT 418.950 763.950 421.050 766.050 ;
        RECT 410.400 760.350 411.600 762.000 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 407.400 756.900 408.600 757.650 ;
        RECT 406.950 754.800 409.050 756.900 ;
        RECT 416.400 748.050 417.450 763.950 ;
        RECT 419.400 757.050 420.450 763.950 ;
        RECT 424.950 761.100 427.050 763.200 ;
        RECT 431.400 762.600 432.450 772.950 ;
        RECT 425.400 760.350 426.600 761.100 ;
        RECT 431.400 760.350 432.600 762.600 ;
        RECT 439.950 761.100 442.050 763.200 ;
        RECT 443.400 763.050 444.450 787.950 ;
        RECT 452.400 784.050 453.450 820.950 ;
        RECT 455.400 804.600 456.450 823.950 ;
        RECT 458.400 820.050 459.450 826.950 ;
        RECT 461.400 823.050 462.450 868.950 ;
        RECT 469.950 865.950 472.050 868.050 ;
        RECT 463.950 862.950 466.050 865.050 ;
        RECT 464.400 856.050 465.450 862.950 ;
        RECT 463.950 853.950 466.050 856.050 ;
        RECT 464.400 834.900 465.450 853.950 ;
        RECT 470.400 840.600 471.450 865.950 ;
        RECT 479.400 862.050 480.450 878.400 ;
        RECT 484.950 877.800 487.050 879.900 ;
        RECT 493.950 877.800 496.050 879.900 ;
        RECT 503.400 879.000 504.600 880.650 ;
        RECT 502.950 874.950 505.050 879.000 ;
        RECT 496.950 871.950 499.050 874.050 ;
        RECT 478.950 859.950 481.050 862.050 ;
        RECT 487.950 844.950 490.050 847.050 ;
        RECT 470.400 838.350 471.600 840.600 ;
        RECT 478.950 839.100 481.050 841.200 ;
        RECT 488.400 840.450 489.450 844.950 ;
        RECT 491.400 840.450 492.600 840.600 ;
        RECT 488.400 839.400 492.600 840.450 ;
        RECT 469.950 835.950 472.050 838.050 ;
        RECT 472.950 835.950 475.050 838.050 ;
        RECT 473.400 834.900 474.600 835.650 ;
        RECT 479.400 835.050 480.450 839.100 ;
        RECT 463.950 832.800 466.050 834.900 ;
        RECT 472.950 832.800 475.050 834.900 ;
        RECT 478.950 832.950 481.050 835.050 ;
        RECT 475.950 829.950 478.050 832.050 ;
        RECT 460.950 820.950 463.050 823.050 ;
        RECT 476.400 820.050 477.450 829.950 ;
        RECT 488.400 826.050 489.450 839.400 ;
        RECT 491.400 838.350 492.600 839.400 ;
        RECT 491.100 835.950 493.200 838.050 ;
        RECT 490.950 829.950 493.050 832.050 ;
        RECT 487.950 823.950 490.050 826.050 ;
        RECT 488.400 820.050 489.450 823.950 ;
        RECT 491.400 823.050 492.450 829.950 ;
        RECT 490.950 820.950 493.050 823.050 ;
        RECT 457.950 817.950 460.050 820.050 ;
        RECT 462.000 819.450 466.050 820.050 ;
        RECT 461.400 817.950 466.050 819.450 ;
        RECT 475.950 817.950 478.050 820.050 ;
        RECT 487.950 817.950 490.050 820.050 ;
        RECT 461.400 811.050 462.450 817.950 ;
        RECT 464.700 813.300 466.800 815.400 ;
        RECT 460.950 808.950 463.050 811.050 ;
        RECT 455.400 802.350 456.600 804.600 ;
        RECT 460.950 803.100 463.050 805.200 ;
        RECT 455.100 799.950 457.200 802.050 ;
        RECT 457.950 790.950 460.050 793.050 ;
        RECT 451.950 781.950 454.050 784.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 427.950 757.950 430.050 760.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 433.950 757.950 436.050 760.050 ;
        RECT 418.950 754.950 421.050 757.050 ;
        RECT 428.400 756.000 429.600 757.650 ;
        RECT 434.400 757.050 435.600 757.650 ;
        RECT 427.950 751.950 430.050 756.000 ;
        RECT 434.400 755.400 439.050 757.050 ;
        RECT 435.000 754.950 439.050 755.400 ;
        RECT 406.950 745.950 409.050 748.050 ;
        RECT 415.950 745.950 418.050 748.050 ;
        RECT 430.950 745.950 433.050 748.050 ;
        RECT 403.950 736.950 406.050 739.050 ;
        RECT 398.400 732.000 402.450 732.450 ;
        RECT 398.400 731.400 403.050 732.000 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 724.950 373.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 374.400 723.900 375.600 724.650 ;
        RECT 373.950 721.800 376.050 723.900 ;
        RECT 383.400 721.050 384.450 727.950 ;
        RECT 389.400 727.350 390.600 729.600 ;
        RECT 395.400 727.350 396.600 729.600 ;
        RECT 400.950 727.950 403.050 731.400 ;
        RECT 388.950 724.950 391.050 727.050 ;
        RECT 391.950 724.950 394.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 392.400 723.000 393.600 724.650 ;
        RECT 398.400 723.900 399.600 724.650 ;
        RECT 391.950 721.050 394.050 723.000 ;
        RECT 397.950 721.800 400.050 723.900 ;
        RECT 382.950 718.950 385.050 721.050 ;
        RECT 391.800 720.000 394.050 721.050 ;
        RECT 391.800 718.950 393.900 720.000 ;
        RECT 394.950 718.950 397.050 721.050 ;
        RECT 391.950 712.950 394.050 715.050 ;
        RECT 344.700 671.700 345.900 693.300 ;
        RECT 347.700 691.500 349.200 696.300 ;
        RECT 350.100 693.300 352.200 695.400 ;
        RECT 358.950 694.950 361.050 697.050 ;
        RECT 366.600 696.300 368.700 698.400 ;
        RECT 369.600 696.300 372.600 698.400 ;
        RECT 347.100 689.400 349.200 691.500 ;
        RECT 347.700 671.700 349.200 689.400 ;
        RECT 350.700 686.100 351.900 693.300 ;
        RECT 355.500 691.800 357.600 693.900 ;
        RECT 364.200 693.300 366.300 695.400 ;
        RECT 350.100 684.000 352.200 686.100 ;
        RECT 356.700 685.200 357.600 691.800 ;
        RECT 350.700 671.700 351.900 684.000 ;
        RECT 355.500 683.100 357.600 685.200 ;
        RECT 352.800 676.500 354.900 678.600 ;
        RECT 356.700 672.600 357.600 683.100 ;
        RECT 358.950 681.000 361.050 685.050 ;
        RECT 359.400 679.350 360.600 681.000 ;
        RECT 359.100 676.950 361.200 679.050 ;
        RECT 344.700 669.600 346.800 671.700 ;
        RECT 347.700 669.600 349.800 671.700 ;
        RECT 350.700 669.600 352.800 671.700 ;
        RECT 356.100 670.500 358.200 672.600 ;
        RECT 365.100 671.700 366.300 693.300 ;
        RECT 367.500 690.300 368.700 696.300 ;
        RECT 367.500 688.200 369.600 690.300 ;
        RECT 367.500 671.700 368.700 688.200 ;
        RECT 371.100 677.400 372.600 696.300 ;
        RECT 373.950 694.950 376.050 697.050 ;
        RECT 370.500 675.300 372.600 677.400 ;
        RECT 370.500 671.700 371.700 675.300 ;
        RECT 364.200 669.600 366.300 671.700 ;
        RECT 367.200 669.600 369.300 671.700 ;
        RECT 370.200 669.600 372.300 671.700 ;
        RECT 337.950 664.950 340.050 667.050 ;
        RECT 343.950 664.950 346.050 667.050 ;
        RECT 370.950 664.950 373.050 667.050 ;
        RECT 331.950 661.950 334.050 664.050 ;
        RECT 344.400 657.450 345.450 664.950 ;
        RECT 364.950 661.950 367.050 664.050 ;
        RECT 301.950 652.950 304.050 655.050 ;
        RECT 313.950 652.950 316.050 655.050 ;
        RECT 319.950 652.950 322.050 655.050 ;
        RECT 340.800 654.300 342.900 656.400 ;
        RECT 344.400 655.200 345.600 657.450 ;
        RECT 304.950 650.100 307.050 652.200 ;
        RECT 305.400 649.350 306.600 650.100 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 307.950 646.950 310.050 649.050 ;
        RECT 308.400 645.900 309.600 646.650 ;
        RECT 301.950 643.800 304.050 645.900 ;
        RECT 307.800 643.800 309.900 645.900 ;
        RECT 310.950 643.950 313.050 646.050 ;
        RECT 296.400 605.400 300.450 606.450 ;
        RECT 302.400 606.600 303.450 643.800 ;
        RECT 311.400 637.050 312.450 643.950 ;
        RECT 310.950 634.950 313.050 637.050 ;
        RECT 314.400 625.050 315.450 652.950 ;
        RECT 322.950 650.100 325.050 652.200 ;
        RECT 338.400 651.450 339.600 651.600 ;
        RECT 335.400 650.400 339.600 651.450 ;
        RECT 323.400 649.350 324.600 650.100 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 325.950 646.950 328.050 649.050 ;
        RECT 320.400 644.400 321.600 646.650 ;
        RECT 326.400 644.400 327.600 646.650 ;
        RECT 320.400 640.050 321.450 644.400 ;
        RECT 319.950 637.950 322.050 640.050 ;
        RECT 307.950 622.950 310.050 625.050 ;
        RECT 313.950 622.950 316.050 625.050 ;
        RECT 308.400 606.600 309.450 622.950 ;
        RECT 313.950 616.950 316.050 619.050 ;
        RECT 286.950 601.950 289.050 604.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 280.950 598.950 283.050 601.050 ;
        RECT 292.950 598.950 295.050 601.050 ;
        RECT 286.950 595.950 289.050 598.050 ;
        RECT 277.950 583.950 280.050 586.050 ;
        RECT 275.400 581.400 279.450 582.450 ;
        RECT 274.950 577.950 277.050 580.050 ;
        RECT 260.400 571.350 261.600 573.600 ;
        RECT 266.400 571.350 267.600 573.600 ;
        RECT 271.950 571.950 274.050 574.050 ;
        RECT 275.400 571.050 276.450 577.950 ;
        RECT 259.950 568.950 262.050 571.050 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 256.950 565.950 259.050 568.050 ;
        RECT 263.400 566.400 264.600 568.650 ;
        RECT 269.400 566.400 270.600 568.650 ;
        RECT 257.400 529.050 258.450 565.950 ;
        RECT 263.400 556.050 264.450 566.400 ;
        RECT 262.950 553.950 265.050 556.050 ;
        RECT 269.400 541.050 270.450 566.400 ;
        RECT 274.950 565.800 277.050 567.900 ;
        RECT 268.950 538.950 271.050 541.050 ;
        RECT 256.950 526.950 259.050 529.050 ;
        RECT 262.950 527.100 265.050 529.200 ;
        RECT 269.400 529.050 270.450 538.950 ;
        RECT 271.950 529.950 274.050 532.050 ;
        RECT 263.400 526.350 264.600 527.100 ;
        RECT 268.950 526.950 271.050 529.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 260.400 523.050 261.600 523.650 ;
        RECT 256.950 521.400 261.600 523.050 ;
        RECT 266.400 521.400 267.600 523.650 ;
        RECT 256.950 520.950 261.450 521.400 ;
        RECT 256.950 514.950 259.050 517.050 ;
        RECT 257.400 496.050 258.450 514.950 ;
        RECT 260.400 505.050 261.450 520.950 ;
        RECT 262.950 517.950 265.050 520.050 ;
        RECT 263.400 511.050 264.450 517.950 ;
        RECT 262.950 508.950 265.050 511.050 ;
        RECT 259.950 502.950 262.050 505.050 ;
        RECT 262.950 498.450 265.050 499.050 ;
        RECT 266.400 498.450 267.450 521.400 ;
        RECT 268.950 517.950 271.050 523.050 ;
        RECT 272.400 510.450 273.450 529.950 ;
        RECT 262.950 497.400 267.450 498.450 ;
        RECT 269.400 509.400 273.450 510.450 ;
        RECT 256.950 493.950 259.050 496.050 ;
        RECT 262.950 495.000 265.050 497.400 ;
        RECT 263.400 493.350 264.600 495.000 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 256.950 484.950 259.050 490.050 ;
        RECT 260.400 489.900 261.600 490.650 ;
        RECT 259.950 487.800 262.050 489.900 ;
        RECT 253.950 481.950 256.050 484.050 ;
        RECT 250.950 463.950 253.050 466.050 ;
        RECT 250.950 457.950 253.050 460.050 ;
        RECT 251.400 454.050 252.450 457.950 ;
        RECT 250.950 451.950 253.050 454.050 ;
        RECT 226.950 445.950 229.050 448.050 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 232.950 445.950 235.050 448.050 ;
        RECT 235.950 445.950 238.050 448.050 ;
        RECT 212.400 439.050 213.450 443.400 ;
        RECT 220.950 442.950 223.050 445.050 ;
        RECT 227.400 444.900 228.600 445.650 ;
        RECT 233.400 444.900 234.600 445.650 ;
        RECT 226.950 442.800 229.050 444.900 ;
        RECT 232.950 442.800 235.050 444.900 ;
        RECT 214.950 439.950 217.050 442.050 ;
        RECT 238.950 439.950 241.050 444.900 ;
        RECT 178.950 436.950 181.050 439.050 ;
        RECT 211.950 436.950 214.050 439.050 ;
        RECT 160.950 430.950 163.050 433.050 ;
        RECT 181.950 430.950 184.050 433.050 ;
        RECT 193.950 430.950 196.050 433.050 ;
        RECT 157.950 423.450 160.050 424.050 ;
        RECT 152.400 422.400 160.050 423.450 ;
        RECT 152.400 418.050 153.450 422.400 ;
        RECT 157.950 421.950 160.050 422.400 ;
        RECT 175.950 421.950 178.050 424.050 ;
        RECT 151.950 415.950 154.050 418.050 ;
        RECT 154.950 417.000 157.050 421.050 ;
        RECT 163.950 418.950 166.050 421.050 ;
        RECT 155.400 415.350 156.600 417.000 ;
        RECT 155.400 412.950 157.500 415.050 ;
        RECT 160.800 412.950 162.900 415.050 ;
        RECT 161.400 410.400 162.600 412.650 ;
        RECT 131.400 407.400 135.450 408.450 ;
        RECT 127.950 400.950 130.050 403.050 ;
        RECT 118.950 391.950 121.050 394.050 ;
        RECT 107.400 370.350 108.600 371.100 ;
        RECT 113.400 370.350 114.600 372.600 ;
        RECT 115.950 370.950 118.050 373.050 ;
        RECT 128.400 372.600 129.450 400.950 ;
        RECT 128.400 370.350 129.600 372.600 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 106.950 367.950 109.050 370.050 ;
        RECT 109.950 367.950 112.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 104.400 365.400 105.600 367.650 ;
        RECT 110.400 366.900 111.600 367.650 ;
        RECT 125.400 366.900 126.600 367.650 ;
        RECT 104.400 361.050 105.450 365.400 ;
        RECT 109.950 364.800 112.050 366.900 ;
        RECT 115.950 364.800 118.050 366.900 ;
        RECT 124.950 364.800 127.050 366.900 ;
        RECT 134.400 366.450 135.450 407.400 ;
        RECT 145.950 406.950 148.050 409.050 ;
        RECT 154.950 406.950 157.050 409.050 ;
        RECT 139.950 371.100 142.050 373.200 ;
        RECT 145.950 372.000 148.050 376.050 ;
        RECT 151.950 373.950 154.050 376.050 ;
        RECT 140.400 370.350 141.600 371.100 ;
        RECT 146.400 370.350 147.600 372.000 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 143.400 366.900 144.600 367.650 ;
        RECT 131.400 365.400 135.450 366.450 ;
        RECT 103.950 358.950 106.050 361.050 ;
        RECT 103.950 346.950 106.050 349.050 ;
        RECT 98.400 337.350 99.600 339.600 ;
        RECT 94.950 334.950 97.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 77.400 304.050 78.450 331.800 ;
        RECT 83.400 310.050 84.450 332.400 ;
        RECT 88.950 331.800 91.050 333.900 ;
        RECT 95.400 332.400 96.600 334.650 ;
        RECT 95.400 328.050 96.450 332.400 ;
        RECT 94.950 325.950 97.050 328.050 ;
        RECT 82.950 307.950 85.050 310.050 ;
        RECT 76.950 301.950 79.050 304.050 ;
        RECT 104.400 301.050 105.450 346.950 ;
        RECT 116.400 339.600 117.450 364.800 ;
        RECT 125.400 361.050 126.450 364.800 ;
        RECT 124.950 358.950 127.050 361.050 ;
        RECT 116.400 337.350 117.600 339.600 ;
        RECT 121.950 338.100 124.050 340.200 ;
        RECT 127.950 338.100 130.050 340.200 ;
        RECT 122.400 337.350 123.600 338.100 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 115.950 334.950 118.050 337.050 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 121.950 334.950 124.050 337.050 ;
        RECT 113.400 333.900 114.600 334.650 ;
        RECT 112.950 331.800 115.050 333.900 ;
        RECT 119.400 332.400 120.600 334.650 ;
        RECT 119.400 328.050 120.450 332.400 ;
        RECT 128.400 331.050 129.450 338.100 ;
        RECT 131.400 333.450 132.450 365.400 ;
        RECT 142.950 364.800 145.050 366.900 ;
        RECT 152.400 361.050 153.450 373.950 ;
        RECT 155.400 367.050 156.450 406.950 ;
        RECT 161.400 406.050 162.450 410.400 ;
        RECT 160.950 403.950 163.050 406.050 ;
        RECT 164.400 400.050 165.450 418.950 ;
        RECT 176.400 417.600 177.450 421.950 ;
        RECT 182.400 417.600 183.450 430.950 ;
        RECT 176.400 415.350 177.600 417.600 ;
        RECT 182.400 415.350 183.600 417.600 ;
        RECT 175.950 412.950 178.050 415.050 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 179.400 410.400 180.600 412.650 ;
        RECT 179.400 403.050 180.450 410.400 ;
        RECT 187.950 409.950 190.050 412.050 ;
        RECT 178.950 400.950 181.050 403.050 ;
        RECT 163.950 397.950 166.050 400.050 ;
        RECT 160.950 371.100 163.050 373.200 ;
        RECT 167.400 372.450 168.600 372.600 ;
        RECT 167.400 371.400 174.450 372.450 ;
        RECT 161.400 370.350 162.600 371.100 ;
        RECT 167.400 370.350 168.600 371.400 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 154.950 364.950 157.050 367.050 ;
        RECT 164.400 366.900 165.600 367.650 ;
        RECT 163.950 364.800 166.050 366.900 ;
        RECT 139.950 358.950 142.050 361.050 ;
        RECT 151.950 358.950 154.050 361.050 ;
        RECT 140.400 339.600 141.450 358.950 ;
        RECT 148.950 346.950 151.050 349.050 ;
        RECT 140.400 337.350 141.600 339.600 ;
        RECT 136.950 334.950 139.050 337.050 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 131.400 332.400 135.450 333.450 ;
        RECT 127.950 328.950 130.050 331.050 ;
        RECT 118.950 325.950 121.050 328.050 ;
        RECT 124.950 316.950 127.050 319.050 ;
        RECT 115.950 301.950 118.050 304.050 ;
        RECT 103.950 298.950 106.050 301.050 ;
        RECT 112.950 298.950 115.050 301.050 ;
        RECT 37.950 295.950 40.050 298.050 ;
        RECT 67.950 295.950 70.050 298.050 ;
        RECT 73.950 295.950 76.050 298.050 ;
        RECT 38.400 294.600 39.450 295.950 ;
        RECT 38.400 292.350 39.600 294.600 ;
        RECT 43.950 293.100 46.050 295.200 ;
        RECT 49.950 293.100 52.050 295.200 ;
        RECT 55.950 293.100 58.050 295.200 ;
        RECT 61.950 293.100 64.050 295.200 ;
        RECT 70.950 293.100 73.050 295.200 ;
        RECT 44.400 292.350 45.600 293.100 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 31.950 286.950 34.050 289.050 ;
        RECT 35.400 287.400 36.600 289.650 ;
        RECT 41.400 287.400 42.600 289.650 ;
        RECT 28.950 280.950 31.050 283.050 ;
        RECT 22.950 277.950 25.050 280.050 ;
        RECT 23.400 265.050 24.450 277.950 ;
        RECT 28.950 277.800 31.050 279.900 ;
        RECT 29.400 265.050 30.450 277.800 ;
        RECT 22.950 262.950 25.050 265.050 ;
        RECT 28.950 262.950 31.050 265.050 ;
        RECT 7.950 260.100 10.050 262.200 ;
        RECT 16.950 260.100 19.050 262.200 ;
        RECT 24.000 261.600 28.050 262.050 ;
        RECT 8.400 250.050 9.450 260.100 ;
        RECT 17.400 259.350 18.600 260.100 ;
        RECT 23.400 259.950 28.050 261.600 ;
        RECT 28.950 261.450 31.050 261.900 ;
        RECT 32.400 261.450 33.450 286.950 ;
        RECT 35.400 280.050 36.450 287.400 ;
        RECT 41.400 280.050 42.450 287.400 ;
        RECT 50.400 280.050 51.450 293.100 ;
        RECT 56.400 292.350 57.600 293.100 ;
        RECT 62.400 292.350 63.600 293.100 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 59.400 288.900 60.600 289.650 ;
        RECT 58.950 286.800 61.050 288.900 ;
        RECT 65.400 287.400 66.600 289.650 ;
        RECT 71.400 288.450 72.450 293.100 ;
        RECT 74.400 288.900 75.450 295.950 ;
        RECT 79.950 293.100 82.050 295.200 ;
        RECT 85.950 294.000 88.050 298.050 ;
        RECT 104.400 297.450 105.450 298.950 ;
        RECT 101.400 296.400 105.450 297.450 ;
        RECT 80.400 292.350 81.600 293.100 ;
        RECT 86.400 292.350 87.600 294.000 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 94.950 289.950 97.050 295.200 ;
        RECT 101.400 294.600 102.450 296.400 ;
        RECT 101.400 292.350 102.600 294.600 ;
        RECT 106.950 293.100 109.050 295.200 ;
        RECT 107.400 292.350 108.600 293.100 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 68.400 287.400 72.450 288.450 ;
        RECT 55.950 283.950 58.050 286.050 ;
        RECT 34.950 277.950 37.050 280.050 ;
        RECT 40.950 277.950 43.050 280.050 ;
        RECT 49.950 277.950 52.050 280.050 ;
        RECT 49.950 265.950 52.050 268.050 ;
        RECT 28.950 260.400 33.450 261.450 ;
        RECT 23.400 259.350 24.600 259.950 ;
        RECT 28.950 259.800 31.050 260.400 ;
        RECT 34.950 260.100 37.050 262.200 ;
        RECT 40.950 260.100 43.050 262.200 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 14.400 255.450 15.600 256.650 ;
        RECT 20.400 255.900 21.600 256.650 ;
        RECT 11.400 254.400 15.600 255.450 ;
        RECT 7.950 247.950 10.050 250.050 ;
        RECT 11.400 247.050 12.450 254.400 ;
        RECT 19.950 253.800 22.050 255.900 ;
        RECT 25.950 253.950 28.050 256.050 ;
        RECT 10.950 244.950 13.050 247.050 ;
        RECT 4.950 238.950 7.050 241.050 ;
        RECT 11.400 216.600 12.450 244.950 ;
        RECT 11.400 214.350 12.600 216.600 ;
        RECT 26.400 216.450 27.450 253.950 ;
        RECT 29.400 244.050 30.450 259.800 ;
        RECT 35.400 259.350 36.600 260.100 ;
        RECT 41.400 259.350 42.600 260.100 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 38.400 255.900 39.600 256.650 ;
        RECT 44.400 255.900 45.600 256.650 ;
        RECT 50.400 255.900 51.450 265.950 ;
        RECT 56.400 265.050 57.450 283.950 ;
        RECT 65.400 274.050 66.450 287.400 ;
        RECT 64.950 271.950 67.050 274.050 ;
        RECT 55.950 262.950 58.050 265.050 ;
        RECT 52.950 259.950 55.050 262.050 ;
        RECT 61.950 260.100 64.050 262.200 ;
        RECT 68.400 261.600 69.450 287.400 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 83.400 287.400 84.600 289.650 ;
        RECT 89.400 287.400 90.600 289.650 ;
        RECT 76.950 283.950 79.050 286.050 ;
        RECT 73.950 265.950 76.050 268.050 ;
        RECT 37.950 253.800 40.050 255.900 ;
        RECT 43.950 253.800 46.050 255.900 ;
        RECT 49.950 253.800 52.050 255.900 ;
        RECT 28.950 241.950 31.050 244.050 ;
        RECT 40.950 241.950 43.050 244.050 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 28.950 229.950 31.050 232.050 ;
        RECT 23.400 215.400 27.450 216.450 ;
        RECT 29.400 216.600 30.450 229.950 ;
        RECT 35.400 217.200 36.450 235.950 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 14.400 210.900 15.600 211.650 ;
        RECT 13.950 208.800 16.050 210.900 ;
        RECT 23.400 187.050 24.450 215.400 ;
        RECT 29.400 214.350 30.600 216.600 ;
        RECT 34.950 215.100 37.050 217.200 ;
        RECT 35.400 214.350 36.600 215.100 ;
        RECT 28.950 211.950 31.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 32.400 210.900 33.600 211.650 ;
        RECT 41.400 211.050 42.450 241.950 ;
        RECT 49.950 223.950 52.050 226.050 ;
        RECT 50.400 216.600 51.450 223.950 ;
        RECT 53.400 223.050 54.450 259.950 ;
        RECT 62.400 259.350 63.600 260.100 ;
        RECT 68.400 259.350 69.600 261.600 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 55.950 253.950 58.050 256.050 ;
        RECT 59.400 255.000 60.600 256.650 ;
        RECT 65.400 255.900 66.600 256.650 ;
        RECT 74.400 256.050 75.450 265.950 ;
        RECT 56.400 247.050 57.450 253.950 ;
        RECT 58.950 247.950 61.050 255.000 ;
        RECT 64.950 253.800 67.050 255.900 ;
        RECT 73.950 253.950 76.050 256.050 ;
        RECT 64.950 247.950 67.050 252.750 ;
        RECT 55.950 244.950 58.050 247.050 ;
        RECT 64.950 241.950 67.050 244.050 ;
        RECT 52.950 220.950 55.050 223.050 ;
        RECT 61.950 220.950 64.050 223.050 ;
        RECT 50.400 214.350 51.600 216.600 ;
        RECT 55.950 215.100 58.050 217.200 ;
        RECT 56.400 214.350 57.600 215.100 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 31.950 208.800 34.050 210.900 ;
        RECT 40.950 208.950 43.050 211.050 ;
        RECT 53.400 209.400 54.600 211.650 ;
        RECT 53.400 207.450 54.450 209.400 ;
        RECT 50.400 206.400 54.450 207.450 ;
        RECT 22.950 184.950 25.050 187.050 ;
        RECT 28.950 184.950 31.050 187.050 ;
        RECT 31.950 184.950 34.050 187.050 ;
        RECT 4.950 182.100 7.050 184.200 ;
        RECT 16.950 182.100 19.050 184.200 ;
        RECT 24.000 183.600 28.050 184.050 ;
        RECT 5.400 100.050 6.450 182.100 ;
        RECT 17.400 181.350 18.600 182.100 ;
        RECT 23.400 181.950 28.050 183.600 ;
        RECT 23.400 181.350 24.600 181.950 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 14.400 176.400 15.600 178.650 ;
        RECT 20.400 176.400 21.600 178.650 ;
        RECT 14.400 169.050 15.450 176.400 ;
        RECT 13.950 166.950 16.050 169.050 ;
        RECT 20.400 163.050 21.450 176.400 ;
        RECT 29.400 175.050 30.450 184.950 ;
        RECT 28.950 172.950 31.050 175.050 ;
        RECT 19.950 160.950 22.050 163.050 ;
        RECT 28.950 139.950 31.050 142.050 ;
        RECT 7.950 137.100 10.050 139.200 ;
        RECT 13.950 137.100 16.050 139.200 ;
        RECT 19.950 137.100 22.050 139.200 ;
        RECT 8.400 124.050 9.450 137.100 ;
        RECT 14.400 136.350 15.600 137.100 ;
        RECT 20.400 136.350 21.600 137.100 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 17.400 132.900 18.600 133.650 ;
        RECT 23.400 133.050 24.600 133.650 ;
        RECT 16.950 130.800 19.050 132.900 ;
        RECT 23.400 131.400 28.050 133.050 ;
        RECT 24.000 130.950 28.050 131.400 ;
        RECT 7.950 121.950 10.050 124.050 ;
        RECT 17.400 108.450 18.450 130.800 ;
        RECT 29.400 124.050 30.450 139.950 ;
        RECT 32.400 139.200 33.450 184.950 ;
        RECT 40.950 183.000 43.050 187.050 ;
        RECT 41.400 181.350 42.600 183.000 ;
        RECT 46.950 182.100 49.050 184.200 ;
        RECT 50.400 184.050 51.450 206.400 ;
        RECT 62.400 187.050 63.450 220.950 ;
        RECT 65.400 217.050 66.450 241.950 ;
        RECT 70.950 238.950 73.050 241.050 ;
        RECT 64.950 214.950 67.050 217.050 ;
        RECT 71.400 216.600 72.450 238.950 ;
        RECT 77.400 226.050 78.450 283.950 ;
        RECT 83.400 280.050 84.450 287.400 ;
        RECT 89.400 280.050 90.450 287.400 ;
        RECT 91.950 286.950 94.050 289.050 ;
        RECT 82.950 277.950 85.050 280.050 ;
        RECT 88.950 277.950 91.050 280.050 ;
        RECT 92.400 268.050 93.450 286.950 ;
        RECT 94.950 286.800 97.050 288.900 ;
        RECT 104.400 287.400 105.600 289.650 ;
        RECT 91.950 265.950 94.050 268.050 ;
        RECT 85.950 261.000 88.050 265.050 ;
        RECT 86.400 259.350 87.600 261.000 ;
        RECT 80.100 256.950 82.200 259.050 ;
        RECT 85.500 256.950 87.600 259.050 ;
        RECT 88.800 256.950 90.900 259.050 ;
        RECT 80.400 255.900 81.600 256.650 ;
        RECT 89.400 255.900 90.600 256.650 ;
        RECT 79.950 253.800 82.050 255.900 ;
        RECT 88.950 253.800 91.050 255.900 ;
        RECT 88.950 235.950 91.050 238.050 ;
        RECT 76.950 223.950 79.050 226.050 ;
        RECT 89.400 223.050 90.450 235.950 ;
        RECT 88.950 220.950 91.050 223.050 ;
        RECT 92.400 219.450 93.450 265.950 ;
        RECT 95.400 232.050 96.450 286.800 ;
        RECT 97.950 283.950 100.050 286.050 ;
        RECT 98.400 277.050 99.450 283.950 ;
        RECT 104.400 283.050 105.450 287.400 ;
        RECT 113.400 283.050 114.450 298.950 ;
        RECT 116.400 295.050 117.450 301.950 ;
        RECT 115.950 292.950 118.050 295.050 ;
        RECT 118.950 293.100 121.050 295.200 ;
        RECT 125.400 294.600 126.450 316.950 ;
        RECT 134.400 310.050 135.450 332.400 ;
        RECT 137.400 332.400 138.600 334.650 ;
        RECT 143.400 332.400 144.600 334.650 ;
        RECT 149.400 333.900 150.450 346.950 ;
        RECT 173.400 343.050 174.450 371.400 ;
        RECT 179.400 349.050 180.450 400.950 ;
        RECT 188.400 388.050 189.450 409.950 ;
        RECT 187.950 385.950 190.050 388.050 ;
        RECT 181.950 371.100 184.050 373.200 ;
        RECT 182.400 370.350 183.600 371.100 ;
        RECT 182.100 367.950 184.200 370.050 ;
        RECT 187.500 367.950 189.600 370.050 ;
        RECT 188.400 365.400 189.600 367.650 ;
        RECT 188.400 349.050 189.450 365.400 ;
        RECT 194.400 352.050 195.450 430.950 ;
        RECT 211.950 424.950 214.050 427.050 ;
        RECT 199.950 416.100 202.050 418.200 ;
        RECT 205.950 417.000 208.050 421.050 ;
        RECT 212.400 418.200 213.450 424.950 ;
        RECT 200.400 415.350 201.600 416.100 ;
        RECT 206.400 415.350 207.600 417.000 ;
        RECT 211.950 416.100 214.050 418.200 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 203.400 410.400 204.600 412.650 ;
        RECT 212.400 412.050 213.450 416.100 ;
        RECT 203.400 394.050 204.450 410.400 ;
        RECT 208.800 409.950 210.900 412.050 ;
        RECT 211.950 409.950 214.050 412.050 ;
        RECT 209.400 406.050 210.450 409.950 ;
        RECT 208.950 403.950 211.050 406.050 ;
        RECT 205.950 397.950 208.050 400.050 ;
        RECT 202.950 391.950 205.050 394.050 ;
        RECT 206.400 391.050 207.450 397.950 ;
        RECT 199.950 388.950 202.050 391.050 ;
        RECT 205.950 388.950 208.050 391.050 ;
        RECT 200.400 382.050 201.450 388.950 ;
        RECT 202.950 382.950 205.050 385.050 ;
        RECT 199.950 379.950 202.050 382.050 ;
        RECT 196.950 376.950 199.050 379.050 ;
        RECT 193.950 349.950 196.050 352.050 ;
        RECT 178.950 346.950 181.050 349.050 ;
        RECT 187.950 346.950 190.050 349.050 ;
        RECT 151.950 338.100 154.050 340.200 ;
        RECT 160.950 338.100 163.050 340.200 ;
        RECT 166.950 339.000 169.050 343.050 ;
        RECT 172.950 340.950 175.050 343.050 ;
        RECT 190.950 342.450 193.050 343.050 ;
        RECT 179.400 341.400 193.050 342.450 ;
        RECT 179.400 340.200 180.450 341.400 ;
        RECT 190.950 340.950 193.050 341.400 ;
        RECT 193.950 340.950 196.050 343.050 ;
        RECT 137.400 325.050 138.450 332.400 ;
        RECT 143.400 328.050 144.450 332.400 ;
        RECT 148.950 331.800 151.050 333.900 ;
        RECT 152.400 333.450 153.450 338.100 ;
        RECT 161.400 337.350 162.600 338.100 ;
        RECT 167.400 337.350 168.600 339.000 ;
        RECT 172.950 337.800 175.050 339.900 ;
        RECT 178.950 338.100 181.050 340.200 ;
        RECT 184.950 338.100 187.050 340.200 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 158.400 333.900 159.600 334.650 ;
        RECT 152.400 332.400 156.450 333.450 ;
        RECT 145.950 328.950 148.050 331.050 ;
        RECT 142.950 325.950 145.050 328.050 ;
        RECT 136.950 322.950 139.050 325.050 ;
        RECT 146.400 319.050 147.450 328.950 ;
        RECT 151.950 325.950 154.050 328.050 ;
        RECT 145.950 316.950 148.050 319.050 ;
        RECT 136.950 313.950 139.050 316.050 ;
        RECT 133.950 307.950 136.050 310.050 ;
        RECT 130.950 301.950 133.050 304.050 ;
        RECT 131.400 294.600 132.450 301.950 ;
        RECT 134.400 295.050 135.450 307.950 ;
        RECT 119.400 292.350 120.600 293.100 ;
        RECT 125.400 292.350 126.600 294.600 ;
        RECT 131.400 292.350 132.600 294.600 ;
        RECT 133.950 292.950 136.050 295.050 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 115.950 286.950 118.050 289.050 ;
        RECT 122.400 288.900 123.600 289.650 ;
        RECT 103.950 280.950 106.050 283.050 ;
        RECT 112.950 280.950 115.050 283.050 ;
        RECT 97.950 274.950 100.050 277.050 ;
        RECT 104.400 265.050 105.450 280.950 ;
        RECT 113.400 277.050 114.450 280.950 ;
        RECT 112.950 274.950 115.050 277.050 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 97.950 262.950 100.050 265.050 ;
        RECT 103.950 262.950 106.050 265.050 ;
        RECT 98.400 255.900 99.450 262.950 ;
        RECT 107.400 261.600 108.450 268.950 ;
        RECT 116.400 262.200 117.450 286.950 ;
        RECT 121.950 286.800 124.050 288.900 ;
        RECT 128.400 287.400 129.600 289.650 ;
        RECT 137.400 289.050 138.450 313.950 ;
        RECT 146.400 294.600 147.450 316.950 ;
        RECT 148.950 304.950 151.050 307.050 ;
        RECT 149.400 295.050 150.450 304.950 ;
        RECT 146.400 292.350 147.600 294.600 ;
        RECT 148.950 292.950 151.050 295.050 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 128.400 283.050 129.450 287.400 ;
        RECT 133.950 286.950 136.050 289.050 ;
        RECT 136.950 286.950 139.050 289.050 ;
        RECT 143.400 288.900 144.600 289.650 ;
        RECT 127.950 280.950 130.050 283.050 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 107.400 259.350 108.600 261.600 ;
        RECT 112.800 260.100 114.900 262.200 ;
        RECT 115.950 260.100 118.050 262.200 ;
        RECT 113.400 259.350 114.600 260.100 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 104.400 255.900 105.600 256.650 ;
        RECT 97.950 253.800 100.050 255.900 ;
        RECT 103.950 253.800 106.050 255.900 ;
        RECT 110.400 254.400 111.600 256.650 ;
        RECT 110.400 238.050 111.450 254.400 ;
        RECT 119.400 250.050 120.450 268.950 ;
        RECT 121.950 259.950 124.050 262.050 ;
        RECT 130.800 260.100 132.900 262.200 ;
        RECT 134.400 262.050 135.450 286.950 ;
        RECT 142.950 286.800 145.050 288.900 ;
        RECT 152.400 286.050 153.450 325.950 ;
        RECT 155.400 325.050 156.450 332.400 ;
        RECT 157.950 331.800 160.050 333.900 ;
        RECT 164.400 332.400 165.600 334.650 ;
        RECT 164.400 328.050 165.450 332.400 ;
        RECT 173.400 330.450 174.450 337.800 ;
        RECT 179.400 337.350 180.600 338.100 ;
        RECT 185.400 337.350 186.600 338.100 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 170.400 329.400 174.450 330.450 ;
        RECT 182.400 332.400 183.600 334.650 ;
        RECT 188.400 333.900 189.600 334.650 ;
        RECT 194.400 333.900 195.450 340.950 ;
        RECT 163.950 325.950 166.050 328.050 ;
        RECT 154.950 322.950 157.050 325.050 ;
        RECT 155.400 289.050 156.450 322.950 ;
        RECT 163.950 293.100 166.050 295.200 ;
        RECT 164.400 292.350 165.600 293.100 ;
        RECT 160.950 289.950 163.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 154.950 286.950 157.050 289.050 ;
        RECT 161.400 287.400 162.600 289.650 ;
        RECT 151.950 283.950 154.050 286.050 ;
        RECT 139.950 280.950 142.050 283.050 ;
        RECT 136.950 262.950 139.050 265.050 ;
        RECT 118.950 247.950 121.050 250.050 ;
        RECT 109.950 235.950 112.050 238.050 ;
        RECT 94.950 229.950 97.050 232.050 ;
        RECT 100.950 229.950 103.050 232.050 ;
        RECT 89.400 218.400 93.450 219.450 ;
        RECT 71.400 214.350 72.600 216.600 ;
        RECT 76.950 215.100 79.050 217.200 ;
        RECT 82.950 215.100 85.050 217.200 ;
        RECT 89.400 216.600 90.450 218.400 ;
        RECT 77.400 214.350 78.600 215.100 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 68.400 210.900 69.600 211.650 ;
        RECT 67.950 208.800 70.050 210.900 ;
        RECT 74.400 209.400 75.600 211.650 ;
        RECT 83.400 211.050 84.450 215.100 ;
        RECT 89.400 214.350 90.600 216.600 ;
        RECT 94.950 215.100 97.050 217.200 ;
        RECT 95.400 214.350 96.600 215.100 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 67.950 187.950 70.050 190.050 ;
        RECT 61.950 184.950 64.050 187.050 ;
        RECT 47.400 181.350 48.600 182.100 ;
        RECT 49.950 181.950 52.050 184.050 ;
        RECT 52.950 182.100 55.050 184.200 ;
        RECT 62.400 183.600 63.450 184.950 ;
        RECT 68.400 183.600 69.450 187.950 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 38.400 177.900 39.600 178.650 ;
        RECT 44.400 177.900 45.600 178.650 ;
        RECT 53.400 178.050 54.450 182.100 ;
        RECT 62.400 181.350 63.600 183.600 ;
        RECT 68.400 181.350 69.600 183.600 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 67.950 178.950 70.050 181.050 ;
        RECT 37.950 175.800 40.050 177.900 ;
        RECT 43.950 175.800 46.050 177.900 ;
        RECT 49.950 175.950 52.050 178.050 ;
        RECT 52.950 175.950 55.050 178.050 ;
        RECT 59.400 176.400 60.600 178.650 ;
        RECT 65.400 176.400 66.600 178.650 ;
        RECT 38.400 157.050 39.450 175.800 ;
        RECT 40.950 172.950 43.050 175.050 ;
        RECT 41.400 160.050 42.450 172.950 ;
        RECT 40.950 157.950 43.050 160.050 ;
        RECT 37.950 154.950 40.050 157.050 ;
        RECT 34.950 145.950 37.050 148.050 ;
        RECT 31.950 137.100 34.050 139.200 ;
        RECT 35.400 139.050 36.450 145.950 ;
        RECT 34.950 136.950 37.050 139.050 ;
        RECT 37.950 137.100 40.050 139.200 ;
        RECT 43.950 138.000 46.050 142.050 ;
        RECT 50.400 139.050 51.450 175.950 ;
        RECT 52.950 166.950 55.050 169.050 ;
        RECT 38.400 136.350 39.600 137.100 ;
        RECT 44.400 136.350 45.600 138.000 ;
        RECT 49.950 136.950 52.050 139.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 43.950 133.950 46.050 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 41.400 132.900 42.600 133.650 ;
        RECT 40.950 130.800 43.050 132.900 ;
        RECT 47.400 132.450 48.600 133.650 ;
        RECT 53.400 133.050 54.450 166.950 ;
        RECT 55.950 160.950 58.050 163.050 ;
        RECT 47.400 131.400 51.450 132.450 ;
        RECT 46.950 127.950 49.050 130.050 ;
        RECT 28.950 121.950 31.050 124.050 ;
        RECT 37.950 108.450 40.050 112.050 ;
        RECT 14.400 107.400 18.450 108.450 ;
        RECT 35.400 108.000 40.050 108.450 ;
        RECT 35.400 107.400 39.450 108.000 ;
        RECT 14.400 105.600 15.450 107.400 ;
        RECT 14.400 103.350 15.600 105.600 ;
        RECT 19.950 104.100 22.050 106.200 ;
        RECT 20.400 103.350 21.600 104.100 ;
        RECT 25.950 103.950 28.050 106.050 ;
        RECT 35.400 105.600 36.450 107.400 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 4.950 97.950 7.050 100.050 ;
        RECT 11.400 99.900 12.600 100.650 ;
        RECT 10.950 97.800 13.050 99.900 ;
        RECT 17.400 98.400 18.600 100.650 ;
        RECT 11.400 60.450 12.450 97.800 ;
        RECT 17.400 85.050 18.450 98.400 ;
        RECT 26.400 97.050 27.450 103.950 ;
        RECT 35.400 103.350 36.600 105.600 ;
        RECT 40.950 104.100 43.050 106.200 ;
        RECT 41.400 103.350 42.600 104.100 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 32.400 99.900 33.600 100.650 ;
        RECT 31.950 97.800 34.050 99.900 ;
        RECT 38.400 99.000 39.600 100.650 ;
        RECT 47.400 99.900 48.450 127.950 ;
        RECT 50.400 115.050 51.450 131.400 ;
        RECT 52.950 130.950 55.050 133.050 ;
        RECT 49.950 112.950 52.050 115.050 ;
        RECT 56.400 109.050 57.450 160.950 ;
        RECT 59.400 160.050 60.450 176.400 ;
        RECT 58.950 157.950 61.050 160.050 ;
        RECT 59.400 139.050 60.450 157.950 ;
        RECT 65.400 157.050 66.450 176.400 ;
        RECT 74.400 169.050 75.450 209.400 ;
        RECT 82.950 208.950 85.050 211.050 ;
        RECT 92.400 210.900 93.600 211.650 ;
        RECT 91.950 208.800 94.050 210.900 ;
        RECT 88.950 199.950 91.050 202.050 ;
        RECT 76.950 182.100 79.050 184.200 ;
        RECT 82.950 182.100 85.050 184.200 ;
        RECT 89.400 183.600 90.450 199.950 ;
        RECT 92.400 187.050 93.450 208.800 ;
        RECT 101.400 208.050 102.450 229.950 ;
        RECT 109.950 220.950 112.050 223.050 ;
        RECT 110.400 216.600 111.450 220.950 ;
        RECT 122.400 220.050 123.450 259.950 ;
        RECT 131.400 259.350 132.600 260.100 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 128.400 256.050 129.600 256.650 ;
        RECT 124.950 254.400 129.600 256.050 ;
        RECT 124.950 253.950 129.000 254.400 ;
        RECT 133.950 253.950 136.050 256.050 ;
        RECT 125.400 244.050 126.450 253.950 ;
        RECT 124.950 241.950 127.050 244.050 ;
        RECT 134.400 220.050 135.450 253.950 ;
        RECT 110.400 214.350 111.600 216.600 ;
        RECT 115.950 215.100 118.050 220.050 ;
        RECT 121.950 217.950 124.050 220.050 ;
        RECT 133.950 217.950 136.050 220.050 ;
        RECT 137.400 217.200 138.450 262.950 ;
        RECT 140.400 238.050 141.450 280.950 ;
        RECT 161.400 280.050 162.450 287.400 ;
        RECT 166.950 283.950 169.050 286.050 ;
        RECT 160.950 277.950 163.050 280.050 ;
        RECT 145.950 271.950 148.050 274.050 ;
        RECT 146.400 261.600 147.450 271.950 ;
        RECT 154.950 268.950 157.050 271.050 ;
        RECT 146.400 259.350 147.600 261.600 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 149.400 255.900 150.600 256.650 ;
        RECT 148.950 253.800 151.050 255.900 ;
        RECT 155.400 250.050 156.450 268.950 ;
        RECT 161.400 261.600 162.450 277.950 ;
        RECT 167.400 261.600 168.450 283.950 ;
        RECT 170.400 271.050 171.450 329.400 ;
        RECT 182.400 325.050 183.450 332.400 ;
        RECT 187.950 331.800 190.050 333.900 ;
        RECT 193.950 331.800 196.050 333.900 ;
        RECT 181.950 322.950 184.050 325.050 ;
        RECT 193.950 322.950 196.050 325.050 ;
        RECT 172.950 301.950 175.050 304.050 ;
        RECT 169.950 268.950 172.050 271.050 ;
        RECT 161.400 259.350 162.600 261.600 ;
        RECT 167.400 259.350 168.600 261.600 ;
        RECT 173.400 261.450 174.450 301.950 ;
        RECT 181.950 293.100 184.050 295.200 ;
        RECT 187.950 293.100 190.050 295.200 ;
        RECT 182.400 292.350 183.600 293.100 ;
        RECT 188.400 292.350 189.600 293.100 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 179.400 288.900 180.600 289.650 ;
        RECT 178.950 286.800 181.050 288.900 ;
        RECT 185.400 287.400 186.600 289.650 ;
        RECT 194.400 289.050 195.450 322.950 ;
        RECT 185.400 274.050 186.450 287.400 ;
        RECT 190.950 286.950 193.050 289.050 ;
        RECT 193.950 286.950 196.050 289.050 ;
        RECT 187.950 277.950 190.050 280.050 ;
        RECT 178.950 271.950 181.050 274.050 ;
        RECT 184.950 271.950 187.050 274.050 ;
        RECT 179.400 262.050 180.450 271.950 ;
        RECT 188.400 265.050 189.450 277.950 ;
        RECT 191.400 271.050 192.450 286.950 ;
        RECT 193.950 283.800 196.050 285.900 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 184.800 264.000 186.900 265.050 ;
        RECT 184.800 262.950 187.050 264.000 ;
        RECT 187.950 262.950 190.050 265.050 ;
        RECT 173.400 260.400 177.450 261.450 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 164.400 255.900 165.600 256.650 ;
        RECT 163.950 253.800 166.050 255.900 ;
        RECT 170.400 254.400 171.600 256.650 ;
        RECT 170.400 250.050 171.450 254.400 ;
        RECT 148.950 247.950 151.050 250.050 ;
        RECT 154.950 247.950 157.050 250.050 ;
        RECT 169.950 247.950 172.050 250.050 ;
        RECT 139.950 235.950 142.050 238.050 ;
        RECT 124.950 215.100 127.050 217.200 ;
        RECT 130.950 215.100 133.050 217.200 ;
        RECT 136.950 215.100 139.050 217.200 ;
        RECT 116.400 214.350 117.600 215.100 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 113.400 209.400 114.600 211.650 ;
        RECT 100.950 205.950 103.050 208.050 ;
        RECT 113.400 199.050 114.450 209.400 ;
        RECT 125.400 202.050 126.450 215.100 ;
        RECT 131.400 214.350 132.600 215.100 ;
        RECT 137.400 214.350 138.600 215.100 ;
        RECT 145.950 214.950 148.050 217.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 134.400 209.400 135.600 211.650 ;
        RECT 140.400 210.900 141.600 211.650 ;
        RECT 124.950 199.950 127.050 202.050 ;
        RECT 112.950 196.950 115.050 199.050 ;
        RECT 121.950 196.950 124.050 199.050 ;
        RECT 103.950 190.950 106.050 193.050 ;
        RECT 97.950 187.950 100.050 190.050 ;
        RECT 91.950 184.950 94.050 187.050 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 64.950 154.950 67.050 157.050 ;
        RECT 77.400 148.050 78.450 182.100 ;
        RECT 83.400 181.350 84.600 182.100 ;
        RECT 89.400 181.350 90.600 183.600 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 88.950 178.950 91.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 86.400 177.900 87.600 178.650 ;
        RECT 92.400 178.050 93.600 178.650 ;
        RECT 85.950 175.800 88.050 177.900 ;
        RECT 92.400 176.400 97.050 178.050 ;
        RECT 93.000 175.950 97.050 176.400 ;
        RECT 86.400 169.050 87.450 175.800 ;
        RECT 98.400 175.050 99.450 187.950 ;
        RECT 104.400 184.200 105.450 190.950 ;
        RECT 109.950 187.950 112.050 190.050 ;
        RECT 118.950 187.950 121.050 190.050 ;
        RECT 103.950 182.100 106.050 184.200 ;
        RECT 110.400 183.600 111.450 187.950 ;
        RECT 104.400 181.350 105.600 182.100 ;
        RECT 110.400 181.350 111.600 183.600 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 109.950 178.950 112.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 107.400 176.400 108.600 178.650 ;
        RECT 113.400 176.400 114.600 178.650 ;
        RECT 91.950 172.950 94.050 175.050 ;
        RECT 97.950 172.950 100.050 175.050 ;
        RECT 85.950 166.950 88.050 169.050 ;
        RECT 79.950 160.950 82.050 163.050 ;
        RECT 76.950 145.950 79.050 148.050 ;
        RECT 80.400 142.050 81.450 160.950 ;
        RECT 92.400 151.050 93.450 172.950 ;
        RECT 107.400 169.050 108.450 176.400 ;
        RECT 113.400 175.050 114.450 176.400 ;
        RECT 112.950 172.950 115.050 175.050 ;
        RECT 106.950 166.950 109.050 169.050 ;
        RECT 91.950 148.950 94.050 151.050 ;
        RECT 97.950 148.950 100.050 151.050 ;
        RECT 58.950 136.950 61.050 139.050 ;
        RECT 64.950 138.000 67.050 142.050 ;
        RECT 65.400 136.350 66.600 138.000 ;
        RECT 70.950 137.100 73.050 139.200 ;
        RECT 79.950 138.450 82.050 142.050 ;
        RECT 92.400 138.600 93.450 148.950 ;
        RECT 94.950 139.950 97.050 142.050 ;
        RECT 83.400 138.450 84.600 138.600 ;
        RECT 79.950 138.000 84.600 138.450 ;
        RECT 80.400 137.400 84.600 138.000 ;
        RECT 71.400 136.350 72.600 137.100 ;
        RECT 83.400 136.350 84.600 137.400 ;
        RECT 92.400 136.350 93.600 138.600 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 67.950 133.950 70.050 136.050 ;
        RECT 70.950 133.950 73.050 136.050 ;
        RECT 83.100 133.950 85.200 136.050 ;
        RECT 88.500 133.950 90.600 136.050 ;
        RECT 91.800 133.950 93.900 136.050 ;
        RECT 58.950 130.950 61.050 133.050 ;
        RECT 62.400 131.400 63.600 133.650 ;
        RECT 68.400 132.900 69.600 133.650 ;
        RECT 49.950 106.950 52.050 109.050 ;
        RECT 55.950 106.950 58.050 109.050 ;
        RECT 25.950 94.950 28.050 97.050 ;
        RECT 37.950 91.950 40.050 99.000 ;
        RECT 46.950 97.800 49.050 99.900 ;
        RECT 16.950 82.950 19.050 85.050 ;
        RECT 17.400 64.050 18.450 82.950 ;
        RECT 40.950 70.950 43.050 73.050 ;
        RECT 16.950 61.950 19.050 64.050 ;
        RECT 14.400 60.450 15.600 60.600 ;
        RECT 11.400 59.400 15.600 60.450 ;
        RECT 14.400 58.350 15.600 59.400 ;
        RECT 22.950 59.100 25.050 61.200 ;
        RECT 34.950 60.000 37.050 64.050 ;
        RECT 41.400 60.600 42.450 70.950 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 17.400 54.000 18.600 55.650 ;
        RECT 16.950 49.950 19.050 54.000 ;
        RECT 23.400 40.050 24.450 59.100 ;
        RECT 35.400 58.350 36.600 60.000 ;
        RECT 41.400 58.350 42.600 60.600 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 32.400 54.000 33.600 55.650 ;
        RECT 31.950 49.950 34.050 54.000 ;
        RECT 38.400 53.400 39.600 55.650 ;
        RECT 38.400 49.050 39.450 53.400 ;
        RECT 43.950 52.950 46.050 55.050 ;
        RECT 37.950 46.950 40.050 49.050 ;
        RECT 22.950 37.950 25.050 40.050 ;
        RECT 16.950 26.100 19.050 28.200 ;
        RECT 23.400 27.600 24.450 37.950 ;
        RECT 17.400 25.350 18.600 26.100 ;
        RECT 23.400 25.350 24.600 27.600 ;
        RECT 28.950 26.100 31.050 28.200 ;
        RECT 37.950 26.100 40.050 31.050 ;
        RECT 44.400 27.600 45.450 52.950 ;
        RECT 47.400 52.050 48.450 97.800 ;
        RECT 50.400 73.050 51.450 106.950 ;
        RECT 59.400 105.600 60.450 130.950 ;
        RECT 62.400 124.050 63.450 131.400 ;
        RECT 67.950 130.800 70.050 132.900 ;
        RECT 89.400 131.400 90.600 133.650 ;
        RECT 61.950 121.950 64.050 124.050 ;
        RECT 68.400 112.050 69.450 130.800 ;
        RECT 89.400 124.050 90.450 131.400 ;
        RECT 88.950 121.950 91.050 124.050 ;
        RECT 89.400 112.050 90.450 121.950 ;
        RECT 67.950 109.950 70.050 112.050 ;
        RECT 79.950 109.950 82.050 112.050 ;
        RECT 88.950 109.950 91.050 112.050 ;
        RECT 59.400 103.350 60.600 105.600 ;
        RECT 64.950 104.100 67.050 106.200 ;
        RECT 70.950 104.100 73.050 106.200 ;
        RECT 80.400 105.600 81.450 109.950 ;
        RECT 65.400 103.350 66.600 104.100 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 56.400 99.900 57.600 100.650 ;
        RECT 55.950 97.800 58.050 99.900 ;
        RECT 62.400 98.400 63.600 100.650 ;
        RECT 62.400 85.050 63.450 98.400 ;
        RECT 71.400 94.050 72.450 104.100 ;
        RECT 80.400 103.350 81.600 105.600 ;
        RECT 88.950 103.950 91.050 106.050 ;
        RECT 77.100 100.950 79.200 103.050 ;
        RECT 80.400 100.950 82.500 103.050 ;
        RECT 85.800 100.950 87.900 103.050 ;
        RECT 77.400 98.400 78.600 100.650 ;
        RECT 86.400 99.450 87.600 100.650 ;
        RECT 89.400 99.450 90.450 103.950 ;
        RECT 86.400 98.400 90.450 99.450 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 67.950 85.950 70.050 88.050 ;
        RECT 61.950 82.950 64.050 85.050 ;
        RECT 49.950 70.950 52.050 73.050 ;
        RECT 58.950 64.950 61.050 67.050 ;
        RECT 59.400 61.200 60.450 64.950 ;
        RECT 52.950 59.100 55.050 61.200 ;
        RECT 58.950 59.100 61.050 61.200 ;
        RECT 53.400 58.350 54.600 59.100 ;
        RECT 59.400 58.350 60.600 59.100 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 56.400 53.400 57.600 55.650 ;
        RECT 62.400 54.900 63.600 55.650 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 49.950 46.950 52.050 49.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 22.950 22.950 25.050 25.050 ;
        RECT 14.400 21.000 15.600 22.650 ;
        RECT 13.950 16.950 16.050 21.000 ;
        RECT 20.400 20.400 21.600 22.650 ;
        RECT 29.400 22.050 30.450 26.100 ;
        RECT 38.400 25.350 39.600 26.100 ;
        RECT 44.400 25.350 45.600 27.600 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 40.950 22.950 43.050 25.050 ;
        RECT 43.950 22.950 46.050 25.050 ;
        RECT 20.400 18.450 21.450 20.400 ;
        RECT 20.400 17.400 24.450 18.450 ;
        RECT 23.400 15.450 24.450 17.400 ;
        RECT 25.950 16.950 28.050 22.050 ;
        RECT 28.950 19.950 31.050 22.050 ;
        RECT 35.400 21.900 36.600 22.650 ;
        RECT 41.400 21.900 42.600 22.650 ;
        RECT 50.400 22.050 51.450 46.950 ;
        RECT 56.400 46.050 57.450 53.400 ;
        RECT 61.950 52.800 64.050 54.900 ;
        RECT 64.950 46.950 67.050 49.050 ;
        RECT 55.950 43.950 58.050 46.050 ;
        RECT 58.950 40.950 61.050 43.050 ;
        RECT 52.950 25.950 55.050 28.050 ;
        RECT 59.400 27.600 60.450 40.950 ;
        RECT 65.400 28.200 66.450 46.950 ;
        RECT 68.400 43.050 69.450 85.950 ;
        RECT 77.400 85.050 78.450 98.400 ;
        RECT 91.950 97.950 94.050 100.050 ;
        RECT 88.950 88.950 91.050 91.050 ;
        RECT 76.950 82.950 79.050 85.050 ;
        RECT 76.950 73.950 79.050 76.050 ;
        RECT 70.950 70.950 73.050 73.050 ;
        RECT 71.400 46.050 72.450 70.950 ;
        RECT 77.400 61.200 78.450 73.950 ;
        RECT 89.400 72.450 90.450 88.950 ;
        RECT 92.400 82.050 93.450 97.950 ;
        RECT 91.950 79.950 94.050 82.050 ;
        RECT 89.400 71.400 93.450 72.450 ;
        RECT 76.950 59.100 79.050 61.200 ;
        RECT 82.950 59.100 85.050 61.200 ;
        RECT 77.400 58.350 78.600 59.100 ;
        RECT 83.400 58.350 84.600 59.100 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 73.950 52.950 76.050 55.050 ;
        RECT 80.400 53.400 81.600 55.650 ;
        RECT 86.400 54.900 87.600 55.650 ;
        RECT 92.400 55.050 93.450 71.400 ;
        RECT 95.400 61.200 96.450 139.950 ;
        RECT 98.400 106.050 99.450 148.950 ;
        RECT 106.950 145.950 109.050 148.050 ;
        RECT 107.400 138.600 108.450 145.950 ;
        RECT 113.400 145.050 114.450 172.950 ;
        RECT 119.400 154.050 120.450 187.950 ;
        RECT 122.400 163.050 123.450 196.950 ;
        RECT 134.400 187.050 135.450 209.400 ;
        RECT 139.950 208.800 142.050 210.900 ;
        RECT 142.950 199.950 145.050 202.050 ;
        RECT 136.950 196.950 139.050 199.050 ;
        RECT 133.950 184.950 136.050 187.050 ;
        RECT 130.950 182.100 133.050 184.200 ;
        RECT 137.400 183.600 138.450 196.950 ;
        RECT 131.400 181.350 132.600 182.100 ;
        RECT 137.400 181.350 138.600 183.600 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 128.400 177.900 129.600 178.650 ;
        RECT 134.400 177.900 135.600 178.650 ;
        RECT 143.400 177.900 144.450 199.950 ;
        RECT 146.400 184.200 147.450 214.950 ;
        RECT 149.400 211.050 150.450 247.950 ;
        RECT 172.950 241.950 175.050 244.050 ;
        RECT 160.950 229.950 163.050 232.050 ;
        RECT 154.950 216.000 157.050 220.050 ;
        RECT 161.400 216.600 162.450 229.950 ;
        RECT 166.950 220.950 169.050 223.050 ;
        RECT 155.400 214.350 156.600 216.000 ;
        RECT 161.400 214.350 162.600 216.600 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 160.950 211.950 163.050 214.050 ;
        RECT 148.950 208.950 151.050 211.050 ;
        RECT 158.400 209.400 159.600 211.650 ;
        RECT 151.950 190.950 154.050 193.050 ;
        RECT 145.950 182.100 148.050 184.200 ;
        RECT 152.400 183.600 153.450 190.950 ;
        RECT 158.400 187.050 159.450 209.400 ;
        RECT 167.400 207.450 168.450 220.950 ;
        RECT 173.400 216.600 174.450 241.950 ;
        RECT 176.400 241.050 177.450 260.400 ;
        RECT 178.950 259.950 181.050 262.050 ;
        RECT 184.950 261.000 187.050 262.950 ;
        RECT 185.400 259.350 186.600 261.000 ;
        RECT 190.950 260.100 193.050 262.200 ;
        RECT 194.400 262.050 195.450 283.800 ;
        RECT 191.400 259.350 192.600 260.100 ;
        RECT 193.950 259.950 196.050 262.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 182.400 255.900 183.600 256.650 ;
        RECT 188.400 255.900 189.600 256.650 ;
        RECT 181.950 253.800 184.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 193.950 253.950 196.050 256.050 ;
        RECT 190.950 250.950 193.050 253.050 ;
        RECT 184.950 247.950 187.050 250.050 ;
        RECT 175.950 238.950 178.050 241.050 ;
        RECT 181.950 238.950 184.050 241.050 ;
        RECT 173.400 214.350 174.600 216.600 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 176.400 209.400 177.600 211.650 ;
        RECT 169.950 207.450 172.050 208.050 ;
        RECT 167.400 206.400 172.050 207.450 ;
        RECT 169.950 205.950 172.050 206.400 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 160.950 187.950 163.050 190.050 ;
        RECT 157.950 184.950 160.050 187.050 ;
        RECT 152.400 181.350 153.600 183.600 ;
        RECT 158.400 183.450 159.600 183.600 ;
        RECT 161.400 183.450 162.450 187.950 ;
        RECT 163.950 184.950 166.050 187.050 ;
        RECT 158.400 182.400 162.450 183.450 ;
        RECT 158.400 181.350 159.600 182.400 ;
        RECT 148.950 178.950 151.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 127.950 175.800 130.050 177.900 ;
        RECT 133.950 175.800 136.050 177.900 ;
        RECT 142.950 175.800 145.050 177.900 ;
        RECT 149.400 177.000 150.600 178.650 ;
        RECT 128.400 172.050 129.450 175.800 ;
        RECT 148.950 172.950 151.050 177.000 ;
        RECT 155.400 176.400 156.600 178.650 ;
        RECT 155.400 172.050 156.450 176.400 ;
        RECT 157.950 172.950 160.050 175.050 ;
        RECT 127.950 169.950 130.050 172.050 ;
        RECT 139.950 169.950 142.050 172.050 ;
        RECT 154.950 169.950 157.050 172.050 ;
        RECT 121.950 160.950 124.050 163.050 ;
        RECT 118.950 151.950 121.050 154.050 ;
        RECT 124.950 145.950 127.050 148.050 ;
        RECT 112.950 142.950 115.050 145.050 ;
        RECT 118.950 142.950 121.050 145.050 ;
        RECT 107.400 136.350 108.600 138.600 ;
        RECT 112.950 137.100 115.050 139.200 ;
        RECT 113.400 136.350 114.600 137.100 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 104.400 131.400 105.600 133.650 ;
        RECT 110.400 132.900 111.600 133.650 ;
        RECT 104.400 118.050 105.450 131.400 ;
        RECT 109.950 130.800 112.050 132.900 ;
        RECT 106.950 121.950 109.050 124.050 ;
        RECT 103.950 115.950 106.050 118.050 ;
        RECT 97.950 105.450 100.050 106.050 ;
        RECT 107.400 105.600 108.450 121.950 ;
        RECT 110.400 115.050 111.450 130.800 ;
        RECT 109.950 112.950 112.050 115.050 ;
        RECT 101.400 105.450 102.600 105.600 ;
        RECT 97.950 104.400 102.600 105.450 ;
        RECT 97.950 103.950 100.050 104.400 ;
        RECT 101.400 103.350 102.600 104.400 ;
        RECT 107.400 103.350 108.600 105.600 ;
        RECT 112.950 103.950 115.050 106.050 ;
        RECT 115.950 104.100 118.050 106.200 ;
        RECT 119.400 106.050 120.450 142.950 ;
        RECT 125.400 139.200 126.450 145.950 ;
        RECT 130.950 142.950 133.050 145.050 ;
        RECT 124.950 137.100 127.050 139.200 ;
        RECT 131.400 138.600 132.450 142.950 ;
        RECT 125.400 136.350 126.600 137.100 ;
        RECT 131.400 136.350 132.600 138.600 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 128.400 132.900 129.600 133.650 ;
        RECT 134.400 132.900 135.600 133.650 ;
        RECT 140.400 133.050 141.450 169.950 ;
        RECT 142.950 160.950 145.050 163.050 ;
        RECT 127.950 130.800 130.050 132.900 ;
        RECT 133.950 130.800 136.050 132.900 ;
        RECT 139.950 130.950 142.050 133.050 ;
        RECT 134.400 108.450 135.450 130.800 ;
        RECT 139.950 112.950 142.050 115.050 ;
        RECT 131.400 107.400 135.450 108.450 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 106.950 100.950 109.050 103.050 ;
        RECT 104.400 98.400 105.600 100.650 ;
        RECT 104.400 94.050 105.450 98.400 ;
        RECT 113.400 97.050 114.450 103.950 ;
        RECT 112.950 94.950 115.050 97.050 ;
        RECT 103.950 91.950 106.050 94.050 ;
        RECT 116.400 91.050 117.450 104.100 ;
        RECT 118.950 103.950 121.050 106.050 ;
        RECT 124.950 104.100 127.050 106.200 ;
        RECT 131.400 105.600 132.450 107.400 ;
        RECT 125.400 103.350 126.600 104.100 ;
        RECT 131.400 103.350 132.600 105.600 ;
        RECT 121.950 100.950 124.050 103.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 127.950 100.950 130.050 103.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 122.400 99.900 123.600 100.650 ;
        RECT 121.950 97.800 124.050 99.900 ;
        RECT 128.400 98.400 129.600 100.650 ;
        RECT 134.400 99.000 135.600 100.650 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 122.400 85.050 123.450 97.800 ;
        RECT 128.400 97.050 129.450 98.400 ;
        RECT 128.400 95.400 133.050 97.050 ;
        RECT 129.000 94.950 133.050 95.400 ;
        RECT 133.950 94.950 136.050 99.000 ;
        RECT 136.950 97.950 139.050 100.050 ;
        RECT 115.950 82.950 118.050 85.050 ;
        RECT 121.950 82.950 124.050 85.050 ;
        RECT 130.950 82.950 133.050 85.050 ;
        RECT 103.950 64.950 106.050 67.050 ;
        RECT 94.950 59.100 97.050 61.200 ;
        RECT 104.400 60.600 105.450 64.950 ;
        RECT 74.400 49.050 75.450 52.950 ;
        RECT 80.400 51.450 81.450 53.400 ;
        RECT 85.950 52.800 88.050 54.900 ;
        RECT 91.950 52.950 94.050 55.050 ;
        RECT 77.400 50.400 81.450 51.450 ;
        RECT 73.950 46.950 76.050 49.050 ;
        RECT 70.950 43.950 73.050 46.050 ;
        RECT 67.950 40.950 70.050 43.050 ;
        RECT 77.400 40.050 78.450 50.400 ;
        RECT 76.950 37.950 79.050 40.050 ;
        RECT 73.950 28.950 76.050 31.050 ;
        RECT 34.950 19.800 37.050 21.900 ;
        RECT 28.950 15.450 31.050 18.900 ;
        RECT 35.400 16.050 36.450 19.800 ;
        RECT 40.950 16.950 43.050 21.900 ;
        RECT 49.950 19.950 52.050 22.050 ;
        RECT 23.400 15.000 31.050 15.450 ;
        RECT 23.400 14.400 30.450 15.000 ;
        RECT 34.950 13.950 37.050 16.050 ;
        RECT 53.400 13.050 54.450 25.950 ;
        RECT 59.400 25.350 60.600 27.600 ;
        RECT 64.950 26.100 67.050 28.200 ;
        RECT 65.400 25.350 66.600 26.100 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 62.400 21.000 63.600 22.650 ;
        RECT 68.400 21.900 69.600 22.650 ;
        RECT 61.950 16.950 64.050 21.000 ;
        RECT 67.950 19.800 70.050 21.900 ;
        RECT 74.400 19.050 75.450 28.950 ;
        RECT 77.400 22.050 78.450 37.950 ;
        RECT 91.950 34.950 94.050 37.050 ;
        RECT 85.950 26.100 88.050 31.050 ;
        RECT 92.400 27.600 93.450 34.950 ;
        RECT 95.400 28.200 96.450 59.100 ;
        RECT 104.400 58.350 105.600 60.600 ;
        RECT 109.950 59.100 112.050 61.200 ;
        RECT 110.400 58.350 111.600 59.100 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 101.400 53.400 102.600 55.650 ;
        RECT 107.400 54.900 108.600 55.650 ;
        RECT 116.400 55.050 117.450 82.950 ;
        RECT 131.400 76.050 132.450 82.950 ;
        RECT 130.950 73.950 133.050 76.050 ;
        RECT 127.950 70.950 130.050 73.050 ;
        RECT 128.400 67.050 129.450 70.950 ;
        RECT 124.800 64.950 126.900 67.050 ;
        RECT 127.950 64.950 130.050 67.050 ;
        RECT 125.400 60.600 126.450 64.950 ;
        RECT 131.400 60.600 132.450 73.950 ;
        RECT 125.400 58.350 126.600 60.600 ;
        RECT 131.400 58.350 132.600 60.600 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 101.400 46.050 102.450 53.400 ;
        RECT 106.950 52.800 109.050 54.900 ;
        RECT 115.950 52.950 118.050 55.050 ;
        RECT 122.400 53.400 123.600 55.650 ;
        RECT 128.400 54.900 129.600 55.650 ;
        RECT 118.950 49.950 121.050 52.050 ;
        RECT 100.950 45.450 103.050 46.050 ;
        RECT 98.400 44.400 103.050 45.450 ;
        RECT 86.400 25.350 87.600 26.100 ;
        RECT 92.400 25.350 93.600 27.600 ;
        RECT 94.950 26.100 97.050 28.200 ;
        RECT 98.400 25.050 99.450 44.400 ;
        RECT 100.950 43.950 103.050 44.400 ;
        RECT 106.950 26.100 109.050 28.200 ;
        RECT 112.950 27.000 115.050 31.050 ;
        RECT 107.400 25.350 108.600 26.100 ;
        RECT 113.400 25.350 114.600 27.000 ;
        RECT 119.400 25.050 120.450 49.950 ;
        RECT 122.400 46.050 123.450 53.400 ;
        RECT 127.950 52.800 130.050 54.900 ;
        RECT 121.950 43.950 124.050 46.050 ;
        RECT 137.400 40.050 138.450 97.950 ;
        RECT 140.400 97.050 141.450 112.950 ;
        RECT 143.400 106.050 144.450 160.950 ;
        RECT 151.950 157.950 154.050 160.050 ;
        RECT 152.400 142.050 153.450 157.950 ;
        RECT 145.950 138.000 148.050 142.050 ;
        RECT 151.950 139.950 154.050 142.050 ;
        RECT 146.400 136.350 147.600 138.000 ;
        RECT 154.950 137.100 157.050 139.200 ;
        RECT 155.400 136.350 156.600 137.100 ;
        RECT 146.100 133.950 148.200 136.050 ;
        RECT 149.400 133.950 151.500 136.050 ;
        RECT 154.800 133.950 156.900 136.050 ;
        RECT 149.400 132.900 150.600 133.650 ;
        RECT 158.400 133.050 159.450 172.950 ;
        RECT 148.950 130.800 151.050 132.900 ;
        RECT 157.950 130.950 160.050 133.050 ;
        RECT 164.400 124.050 165.450 184.950 ;
        RECT 167.400 139.200 168.450 199.950 ;
        RECT 170.400 184.050 171.450 205.950 ;
        RECT 176.400 199.050 177.450 209.400 ;
        RECT 175.950 196.950 178.050 199.050 ;
        RECT 175.950 187.950 178.050 190.050 ;
        RECT 176.400 184.200 177.450 187.950 ;
        RECT 169.950 181.950 172.050 184.050 ;
        RECT 175.950 182.100 178.050 184.200 ;
        RECT 182.400 184.050 183.450 238.950 ;
        RECT 176.400 181.350 177.600 182.100 ;
        RECT 181.950 181.950 184.050 184.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 173.400 177.000 174.600 178.650 ;
        RECT 172.950 172.950 175.050 177.000 ;
        RECT 179.400 176.400 180.600 178.650 ;
        RECT 179.400 174.450 180.450 176.400 ;
        RECT 181.950 175.950 184.050 178.050 ;
        RECT 176.400 173.400 180.450 174.450 ;
        RECT 176.400 171.450 177.450 173.400 ;
        RECT 173.400 170.400 177.450 171.450 ;
        RECT 173.400 142.050 174.450 170.400 ;
        RECT 175.950 157.950 178.050 160.050 ;
        RECT 172.950 139.950 175.050 142.050 ;
        RECT 166.950 138.450 169.050 139.200 ;
        RECT 176.400 138.600 177.450 157.950 ;
        RECT 170.400 138.450 171.600 138.600 ;
        RECT 166.950 137.400 171.600 138.450 ;
        RECT 166.950 137.100 169.050 137.400 ;
        RECT 170.400 136.350 171.600 137.400 ;
        RECT 176.400 136.350 177.600 138.600 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 173.400 131.400 174.600 133.650 ;
        RECT 182.400 133.050 183.450 175.950 ;
        RECT 185.400 172.050 186.450 247.950 ;
        RECT 191.400 232.050 192.450 250.950 ;
        RECT 194.400 250.050 195.450 253.950 ;
        RECT 193.950 247.950 196.050 250.050 ;
        RECT 197.400 247.050 198.450 376.950 ;
        RECT 203.400 373.200 204.450 382.950 ;
        RECT 202.950 371.100 205.050 373.200 ;
        RECT 208.950 371.100 211.050 373.200 ;
        RECT 203.400 370.350 204.600 371.100 ;
        RECT 209.400 370.350 210.600 371.100 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 205.950 367.950 208.050 370.050 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 206.400 365.400 207.600 367.650 ;
        RECT 206.400 355.050 207.450 365.400 ;
        RECT 215.400 361.050 216.450 439.950 ;
        RECT 226.950 436.950 229.050 439.050 ;
        RECT 242.400 438.450 243.450 449.100 ;
        RECT 247.950 448.950 250.050 451.050 ;
        RECT 253.950 450.000 256.050 454.050 ;
        RECT 254.400 448.350 255.600 450.000 ;
        RECT 259.950 449.100 262.050 451.200 ;
        RECT 265.950 449.100 268.050 451.200 ;
        RECT 260.400 448.350 261.600 449.100 ;
        RECT 250.950 445.950 253.050 448.050 ;
        RECT 253.950 445.950 256.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 247.950 442.950 250.050 445.050 ;
        RECT 251.400 444.900 252.600 445.650 ;
        RECT 257.400 444.900 258.600 445.650 ;
        RECT 248.400 439.050 249.450 442.950 ;
        RECT 250.950 442.800 253.050 444.900 ;
        RECT 256.950 442.800 259.050 444.900 ;
        RECT 266.400 442.050 267.450 449.100 ;
        RECT 265.950 439.950 268.050 442.050 ;
        RECT 239.400 437.400 243.450 438.450 ;
        RECT 217.950 433.950 220.050 436.050 ;
        RECT 218.400 421.050 219.450 433.950 ;
        RECT 217.950 418.950 220.050 421.050 ;
        RECT 220.950 416.100 223.050 418.200 ;
        RECT 227.400 417.600 228.450 436.950 ;
        RECT 229.950 430.950 232.050 433.050 ;
        RECT 230.400 427.050 231.450 430.950 ;
        RECT 229.950 424.950 232.050 427.050 ;
        RECT 239.400 418.050 240.450 437.400 ;
        RECT 247.950 436.950 250.050 439.050 ;
        RECT 256.950 436.950 259.050 439.050 ;
        RECT 221.400 415.350 222.600 416.100 ;
        RECT 227.400 415.350 228.600 417.600 ;
        RECT 238.950 415.950 241.050 418.050 ;
        RECT 247.950 417.000 250.050 421.050 ;
        RECT 253.950 418.950 256.050 421.050 ;
        RECT 248.400 415.350 249.600 417.000 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 244.950 412.950 247.050 415.050 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 217.950 409.950 220.050 412.050 ;
        RECT 224.400 411.900 225.600 412.650 ;
        RECT 218.400 364.050 219.450 409.950 ;
        RECT 223.950 409.800 226.050 411.900 ;
        RECT 230.400 410.400 231.600 412.650 ;
        RECT 245.400 411.900 246.600 412.650 ;
        RECT 254.400 412.050 255.450 418.950 ;
        RECT 230.400 408.450 231.450 410.400 ;
        RECT 244.950 409.800 247.050 411.900 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 227.400 407.400 231.450 408.450 ;
        RECT 223.950 382.950 226.050 385.050 ;
        RECT 224.400 372.600 225.450 382.950 ;
        RECT 227.400 382.050 228.450 407.400 ;
        RECT 257.400 391.050 258.450 436.950 ;
        RECT 269.400 433.050 270.450 509.400 ;
        RECT 275.400 508.050 276.450 565.800 ;
        RECT 278.400 550.050 279.450 581.400 ;
        RECT 287.400 573.600 288.450 595.950 ;
        RECT 293.400 579.450 294.450 598.950 ;
        RECT 296.400 583.050 297.450 605.400 ;
        RECT 302.400 604.350 303.600 606.600 ;
        RECT 308.400 604.350 309.600 606.600 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 307.950 601.950 310.050 604.050 ;
        RECT 298.950 595.950 301.050 601.050 ;
        RECT 305.400 599.400 306.600 601.650 ;
        RECT 295.950 580.950 298.050 583.050 ;
        RECT 305.400 580.050 306.450 599.400 ;
        RECT 314.400 589.050 315.450 616.950 ;
        RECT 322.950 613.950 325.050 616.050 ;
        RECT 316.950 607.950 319.050 610.050 ;
        RECT 317.400 600.450 318.450 607.950 ;
        RECT 323.400 606.600 324.450 613.950 ;
        RECT 326.400 613.050 327.450 644.400 ;
        RECT 328.950 643.950 331.050 646.050 ;
        RECT 329.400 637.050 330.450 643.950 ;
        RECT 335.400 640.050 336.450 650.400 ;
        RECT 338.400 649.350 339.600 650.400 ;
        RECT 338.100 646.950 340.200 649.050 ;
        RECT 341.100 648.900 342.000 654.300 ;
        RECT 344.100 652.800 346.200 654.900 ;
        RECT 348.000 651.900 350.100 653.700 ;
        RECT 342.900 650.700 351.600 651.900 ;
        RECT 342.900 649.800 345.000 650.700 ;
        RECT 341.100 647.700 348.000 648.900 ;
        RECT 341.100 640.500 342.300 647.700 ;
        RECT 344.100 643.950 346.200 646.050 ;
        RECT 347.100 645.300 348.000 647.700 ;
        RECT 344.400 641.400 345.600 643.650 ;
        RECT 347.100 643.200 349.200 645.300 ;
        RECT 350.700 641.700 351.600 650.700 ;
        RECT 352.800 646.950 354.900 649.050 ;
        RECT 358.950 647.100 361.050 649.200 ;
        RECT 365.400 648.450 366.450 661.950 ;
        RECT 371.400 649.050 372.450 664.950 ;
        RECT 368.400 648.450 369.600 648.600 ;
        RECT 365.400 647.400 369.600 648.450 ;
        RECT 353.400 645.450 354.600 646.650 ;
        RECT 359.400 646.350 360.600 647.100 ;
        RECT 353.400 644.400 357.450 645.450 ;
        RECT 334.950 637.950 337.050 640.050 ;
        RECT 340.800 638.400 342.900 640.500 ;
        RECT 350.400 639.600 352.500 641.700 ;
        RECT 328.950 634.950 331.050 637.050 ;
        RECT 356.400 636.450 357.450 644.400 ;
        RECT 359.100 643.950 361.200 646.050 ;
        RECT 353.400 635.400 357.450 636.450 ;
        RECT 329.400 628.050 330.450 634.950 ;
        RECT 328.950 625.950 331.050 628.050 ;
        RECT 325.950 610.950 328.050 613.050 ;
        RECT 329.400 606.600 330.450 625.950 ;
        RECT 337.950 616.950 340.050 619.050 ;
        RECT 334.950 613.950 337.050 616.050 ;
        RECT 323.400 604.350 324.600 606.600 ;
        RECT 329.400 604.350 330.600 606.600 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 326.400 600.900 327.600 601.650 ;
        RECT 317.400 599.400 321.450 600.450 ;
        RECT 313.950 586.950 316.050 589.050 ;
        RECT 293.400 578.400 297.450 579.450 ;
        RECT 287.400 571.350 288.600 573.600 ;
        RECT 283.950 568.950 286.050 571.050 ;
        RECT 286.950 568.950 289.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 280.950 565.950 283.050 568.050 ;
        RECT 284.400 567.900 285.600 568.650 ;
        RECT 277.950 547.950 280.050 550.050 ;
        RECT 281.400 547.050 282.450 565.950 ;
        RECT 283.950 565.800 286.050 567.900 ;
        RECT 290.400 566.400 291.600 568.650 ;
        RECT 286.950 556.950 289.050 559.050 ;
        RECT 287.400 553.050 288.450 556.950 ;
        RECT 290.400 556.050 291.450 566.400 ;
        RECT 296.400 559.050 297.450 578.400 ;
        RECT 304.950 577.950 307.050 580.050 ;
        RECT 310.950 577.950 313.050 580.050 ;
        RECT 311.400 574.050 312.450 577.950 ;
        RECT 320.400 574.050 321.450 599.400 ;
        RECT 325.950 598.800 328.050 600.900 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 328.950 595.950 331.050 598.050 ;
        RECT 331.950 595.950 334.050 598.050 ;
        RECT 323.400 592.050 324.450 595.950 ;
        RECT 322.950 589.950 325.050 592.050 ;
        RECT 310.950 571.950 313.050 574.050 ;
        RECT 319.950 571.950 322.050 574.050 ;
        RECT 329.400 573.600 330.450 595.950 ;
        RECT 329.400 571.350 330.600 573.600 ;
        RECT 304.950 568.950 307.050 571.050 ;
        RECT 307.950 568.950 310.050 571.050 ;
        RECT 313.950 569.100 316.050 571.200 ;
        RECT 308.400 566.400 309.600 568.650 ;
        RECT 295.950 556.950 298.050 559.050 ;
        RECT 289.950 553.950 292.050 556.050 ;
        RECT 308.400 553.050 309.450 566.400 ;
        RECT 310.950 565.950 313.050 568.050 ;
        RECT 286.950 550.950 289.050 553.050 ;
        RECT 292.950 550.950 295.050 553.050 ;
        RECT 307.950 550.950 310.050 553.050 ;
        RECT 280.950 544.950 283.050 547.050 ;
        RECT 293.400 544.050 294.450 550.950 ;
        RECT 295.950 547.950 298.050 550.050 ;
        RECT 292.950 541.950 295.050 544.050 ;
        RECT 289.950 538.950 292.050 541.050 ;
        RECT 283.950 527.100 286.050 532.050 ;
        RECT 290.400 528.600 291.450 538.950 ;
        RECT 284.400 526.350 285.600 527.100 ;
        RECT 290.400 526.350 291.600 528.600 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 277.950 520.950 280.050 523.050 ;
        RECT 281.400 522.900 282.600 523.650 ;
        RECT 278.400 517.050 279.450 520.950 ;
        RECT 280.950 520.800 283.050 522.900 ;
        RECT 287.400 521.400 288.600 523.650 ;
        RECT 283.950 517.950 286.050 520.050 ;
        RECT 277.950 514.950 280.050 517.050 ;
        RECT 274.950 505.950 277.050 508.050 ;
        RECT 277.950 502.950 280.050 505.050 ;
        RECT 271.950 496.950 274.050 499.050 ;
        RECT 272.400 489.900 273.450 496.950 ;
        RECT 278.400 496.200 279.450 502.950 ;
        RECT 277.950 494.100 280.050 496.200 ;
        RECT 284.400 495.600 285.450 517.950 ;
        RECT 287.400 514.050 288.450 521.400 ;
        RECT 296.400 514.050 297.450 547.950 ;
        RECT 301.950 527.100 304.050 529.200 ;
        RECT 307.950 527.100 310.050 529.200 ;
        RECT 311.400 529.050 312.450 565.950 ;
        RECT 302.400 526.350 303.600 527.100 ;
        RECT 308.400 526.350 309.600 527.100 ;
        RECT 310.950 526.950 313.050 529.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 304.950 523.950 307.050 526.050 ;
        RECT 307.950 523.950 310.050 526.050 ;
        RECT 305.400 521.400 306.600 523.650 ;
        RECT 314.400 523.050 315.450 569.100 ;
        RECT 323.100 568.950 325.200 571.050 ;
        RECT 328.500 568.950 330.600 571.050 ;
        RECT 316.950 562.950 319.050 568.050 ;
        RECT 323.400 567.900 324.600 568.650 ;
        RECT 322.950 565.800 325.050 567.900 ;
        RECT 322.950 562.650 325.050 564.750 ;
        RECT 316.950 556.950 319.050 559.050 ;
        RECT 286.950 511.950 289.050 514.050 ;
        RECT 295.950 511.950 298.050 514.050 ;
        RECT 298.950 508.950 301.050 511.050 ;
        RECT 299.400 502.050 300.450 508.950 ;
        RECT 305.400 508.050 306.450 521.400 ;
        RECT 310.950 520.950 313.050 523.050 ;
        RECT 313.950 520.950 316.050 523.050 ;
        RECT 304.950 505.950 307.050 508.050 ;
        RECT 304.950 502.800 307.050 504.900 ;
        RECT 289.950 499.950 295.050 502.050 ;
        RECT 295.950 499.950 298.050 502.050 ;
        RECT 298.950 499.950 301.050 502.050 ;
        RECT 278.400 493.350 279.600 494.100 ;
        RECT 284.400 493.350 285.600 495.600 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 281.400 489.900 282.600 490.650 ;
        RECT 271.950 487.800 274.050 489.900 ;
        RECT 280.950 487.800 283.050 489.900 ;
        RECT 287.400 489.000 288.600 490.650 ;
        RECT 286.950 484.950 289.050 489.000 ;
        RECT 289.950 487.950 292.050 490.050 ;
        RECT 286.950 481.800 289.050 483.900 ;
        RECT 280.950 475.950 283.050 478.050 ;
        RECT 271.950 463.950 274.050 466.050 ;
        RECT 272.400 451.050 273.450 463.950 ;
        RECT 281.400 454.050 282.450 475.950 ;
        RECT 271.950 448.950 274.050 451.050 ;
        RECT 280.950 450.000 283.050 454.050 ;
        RECT 281.400 448.350 282.600 450.000 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 278.400 444.000 279.600 445.650 ;
        RECT 277.950 439.950 280.050 444.000 ;
        RECT 283.950 442.950 286.050 445.050 ;
        RECT 284.400 436.050 285.450 442.950 ;
        RECT 287.400 439.050 288.450 481.800 ;
        RECT 290.400 466.050 291.450 487.950 ;
        RECT 293.400 484.050 294.450 490.950 ;
        RECT 296.400 489.900 297.450 499.950 ;
        RECT 305.400 495.600 306.450 502.800 ;
        RECT 311.400 502.050 312.450 520.950 ;
        RECT 317.400 505.050 318.450 556.950 ;
        RECT 323.400 529.200 324.450 562.650 ;
        RECT 332.400 538.050 333.450 595.950 ;
        RECT 335.400 580.050 336.450 613.950 ;
        RECT 338.400 607.050 339.450 616.950 ;
        RECT 346.950 613.950 349.050 616.050 ;
        RECT 347.400 607.200 348.450 613.950 ;
        RECT 353.400 613.050 354.450 635.400 ;
        RECT 358.950 634.950 361.050 637.050 ;
        RECT 355.950 628.950 358.050 631.050 ;
        RECT 352.950 610.950 355.050 613.050 ;
        RECT 337.950 604.950 340.050 607.050 ;
        RECT 340.950 605.100 343.050 607.200 ;
        RECT 346.950 605.100 349.050 607.200 ;
        RECT 341.400 604.350 342.600 605.100 ;
        RECT 347.400 604.350 348.600 605.100 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 344.400 599.400 345.600 601.650 ;
        RECT 350.400 599.400 351.600 601.650 ;
        RECT 344.400 595.050 345.450 599.400 ;
        RECT 346.950 595.950 349.050 598.050 ;
        RECT 343.950 592.950 346.050 595.050 ;
        RECT 334.950 577.950 337.050 580.050 ;
        RECT 340.950 577.950 343.050 580.050 ;
        RECT 334.950 569.100 337.050 571.200 ;
        RECT 335.400 568.350 336.600 569.100 ;
        RECT 341.400 568.050 342.450 577.950 ;
        RECT 344.400 570.450 345.600 570.600 ;
        RECT 347.400 570.450 348.450 595.950 ;
        RECT 350.400 592.050 351.450 599.400 ;
        RECT 356.400 598.050 357.450 628.950 ;
        RECT 359.400 613.050 360.450 634.950 ;
        RECT 365.400 631.050 366.450 647.400 ;
        RECT 368.400 646.350 369.600 647.400 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 368.100 643.950 370.200 646.050 ;
        RECT 370.950 640.950 373.050 643.050 ;
        RECT 364.950 628.950 367.050 631.050 ;
        RECT 358.950 610.950 361.050 613.050 ;
        RECT 371.400 610.050 372.450 640.950 ;
        RECT 374.400 619.050 375.450 694.950 ;
        RECT 382.950 691.950 385.050 694.050 ;
        RECT 383.400 687.600 384.450 691.950 ;
        RECT 383.400 685.350 384.600 687.600 ;
        RECT 377.100 682.950 379.200 685.050 ;
        RECT 383.100 682.950 385.200 685.050 ;
        RECT 392.400 664.050 393.450 712.950 ;
        RECT 395.400 670.050 396.450 718.950 ;
        RECT 404.400 718.050 405.450 736.950 ;
        RECT 407.400 718.050 408.450 745.950 ;
        RECT 415.950 728.100 418.050 730.200 ;
        RECT 421.950 729.000 424.050 733.050 ;
        RECT 416.400 727.350 417.600 728.100 ;
        RECT 422.400 727.350 423.600 729.000 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 415.950 724.950 418.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 413.400 724.050 414.600 724.650 ;
        RECT 409.950 722.400 414.600 724.050 ;
        RECT 419.400 723.000 420.600 724.650 ;
        RECT 409.950 721.950 414.000 722.400 ;
        RECT 418.950 721.050 421.050 723.000 ;
        RECT 431.400 721.050 432.450 745.950 ;
        RECT 433.950 736.950 436.050 739.050 ;
        RECT 418.800 720.000 421.050 721.050 ;
        RECT 418.800 718.950 420.900 720.000 ;
        RECT 421.950 718.950 424.050 721.050 ;
        RECT 430.950 718.950 433.050 721.050 ;
        RECT 403.800 715.950 405.900 718.050 ;
        RECT 406.950 715.950 409.050 718.050 ;
        RECT 400.950 712.950 403.050 715.050 ;
        RECT 408.000 714.900 412.050 715.050 ;
        RECT 406.950 712.950 412.050 714.900 ;
        RECT 401.400 709.050 402.450 712.950 ;
        RECT 406.950 712.800 409.050 712.950 ;
        RECT 400.950 706.950 403.050 709.050 ;
        RECT 418.950 706.950 421.050 709.050 ;
        RECT 403.950 703.950 406.050 706.050 ;
        RECT 400.950 700.950 403.050 703.050 ;
        RECT 401.400 691.050 402.450 700.950 ;
        RECT 400.950 688.950 403.050 691.050 ;
        RECT 404.400 684.600 405.450 703.950 ;
        RECT 419.400 697.050 420.450 706.950 ;
        RECT 418.950 694.950 421.050 697.050 ;
        RECT 409.950 688.950 412.050 694.050 ;
        RECT 418.950 691.800 421.050 693.900 ;
        RECT 404.400 682.350 405.600 684.600 ;
        RECT 409.950 683.100 412.050 685.200 ;
        RECT 410.400 682.350 411.600 683.100 ;
        RECT 415.950 682.950 418.050 685.050 ;
        RECT 419.400 684.450 420.450 691.800 ;
        RECT 422.400 688.050 423.450 718.950 ;
        RECT 424.950 706.950 427.050 712.050 ;
        RECT 430.950 709.950 433.050 712.050 ;
        RECT 424.950 703.800 427.050 705.900 ;
        RECT 425.400 694.050 426.450 703.800 ;
        RECT 424.950 691.950 427.050 694.050 ;
        RECT 427.950 690.450 430.050 691.050 ;
        RECT 431.400 690.450 432.450 709.950 ;
        RECT 434.400 709.050 435.450 736.950 ;
        RECT 440.400 733.050 441.450 761.100 ;
        RECT 442.950 760.950 445.050 763.050 ;
        RECT 445.950 761.100 448.050 763.200 ;
        RECT 452.400 762.600 453.450 781.950 ;
        RECT 458.400 766.200 459.450 790.950 ;
        RECT 461.400 781.050 462.450 803.100 ;
        RECT 465.300 795.600 466.800 813.300 ;
        RECT 464.700 793.500 466.800 795.600 ;
        RECT 465.300 788.700 466.800 793.500 ;
        RECT 464.700 786.600 466.800 788.700 ;
        RECT 467.700 813.300 469.800 815.400 ;
        RECT 470.700 813.300 472.800 815.400 ;
        RECT 473.700 813.300 475.800 815.400 ;
        RECT 467.700 791.700 468.900 813.300 ;
        RECT 470.700 795.600 472.200 813.300 ;
        RECT 473.700 801.000 474.900 813.300 ;
        RECT 479.100 812.400 481.200 814.500 ;
        RECT 487.200 813.300 489.300 815.400 ;
        RECT 490.200 813.300 492.300 815.400 ;
        RECT 493.200 813.300 495.300 815.400 ;
        RECT 475.800 806.400 477.900 808.500 ;
        RECT 479.700 801.900 480.600 812.400 ;
        RECT 482.100 805.950 484.200 808.050 ;
        RECT 482.400 804.900 483.600 805.650 ;
        RECT 481.950 802.800 484.050 804.900 ;
        RECT 473.100 798.900 475.200 801.000 ;
        RECT 478.500 799.800 480.600 801.900 ;
        RECT 470.100 793.500 472.200 795.600 ;
        RECT 467.700 786.600 469.800 791.700 ;
        RECT 470.700 788.700 472.200 793.500 ;
        RECT 473.700 791.700 474.900 798.900 ;
        RECT 479.700 793.200 480.600 799.800 ;
        RECT 481.950 796.950 484.050 799.050 ;
        RECT 473.100 789.600 475.200 791.700 ;
        RECT 478.500 791.100 480.600 793.200 ;
        RECT 470.700 786.600 472.800 788.700 ;
        RECT 460.950 778.950 463.050 781.050 ;
        RECT 470.400 774.300 473.400 776.400 ;
        RECT 474.300 774.300 476.400 776.400 ;
        RECT 457.950 764.100 460.050 766.200 ;
        RECT 458.400 763.350 459.600 764.100 ;
        RECT 466.950 763.950 469.050 766.050 ;
        RECT 446.400 760.350 447.600 761.100 ;
        RECT 452.400 760.350 453.600 762.600 ;
        RECT 457.800 760.950 459.900 763.050 ;
        RECT 463.800 760.950 465.900 763.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 442.950 754.950 445.050 757.050 ;
        RECT 449.400 755.400 450.600 757.650 ;
        RECT 443.400 751.050 444.450 754.950 ;
        RECT 442.950 748.950 445.050 751.050 ;
        RECT 445.950 742.950 448.050 745.050 ;
        RECT 439.950 730.950 442.050 733.050 ;
        RECT 436.950 728.100 439.050 730.200 ;
        RECT 437.400 727.350 438.600 728.100 ;
        RECT 437.400 724.950 439.500 727.050 ;
        RECT 442.800 724.950 444.900 727.050 ;
        RECT 443.400 722.400 444.600 724.650 ;
        RECT 443.400 709.050 444.450 722.400 ;
        RECT 433.950 706.950 436.050 709.050 ;
        RECT 442.950 706.950 445.050 709.050 ;
        RECT 427.950 689.400 432.450 690.450 ;
        RECT 427.950 688.950 430.050 689.400 ;
        RECT 421.950 685.950 424.050 688.050 ;
        RECT 428.400 684.600 429.450 688.950 ;
        RECT 434.400 687.600 435.450 706.950 ;
        RECT 442.950 703.800 445.050 705.900 ;
        RECT 434.400 685.350 435.600 687.600 ;
        RECT 422.400 684.450 423.600 684.600 ;
        RECT 419.400 683.400 423.600 684.450 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 401.400 678.900 402.600 679.650 ;
        RECT 400.950 676.800 403.050 678.900 ;
        RECT 407.400 677.400 408.600 679.650 ;
        RECT 407.400 673.050 408.450 677.400 ;
        RECT 416.400 673.050 417.450 682.950 ;
        RECT 422.400 682.350 423.600 683.400 ;
        RECT 428.400 682.350 429.600 684.600 ;
        RECT 433.800 682.950 435.900 685.050 ;
        RECT 439.800 682.950 441.900 685.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 418.950 676.950 421.050 679.050 ;
        RECT 425.400 678.900 426.600 679.650 ;
        RECT 406.950 670.950 409.050 673.050 ;
        RECT 415.950 670.950 418.050 673.050 ;
        RECT 394.950 667.950 397.050 670.050 ;
        RECT 419.400 664.050 420.450 676.950 ;
        RECT 424.950 676.800 427.050 678.900 ;
        RECT 424.950 667.950 427.050 670.050 ;
        RECT 430.950 667.950 433.050 670.050 ;
        RECT 391.950 661.950 394.050 664.050 ;
        RECT 418.950 661.950 421.050 664.050 ;
        RECT 377.700 657.300 379.800 659.400 ;
        RECT 378.300 639.600 379.800 657.300 ;
        RECT 377.700 637.500 379.800 639.600 ;
        RECT 378.300 632.700 379.800 637.500 ;
        RECT 377.700 630.600 379.800 632.700 ;
        RECT 380.700 657.300 382.800 659.400 ;
        RECT 383.700 657.300 385.800 659.400 ;
        RECT 386.700 657.300 388.800 659.400 ;
        RECT 380.700 635.700 381.900 657.300 ;
        RECT 383.700 639.600 385.200 657.300 ;
        RECT 386.700 645.000 387.900 657.300 ;
        RECT 392.100 656.400 394.200 658.500 ;
        RECT 400.200 657.300 402.300 659.400 ;
        RECT 403.200 657.300 405.300 659.400 ;
        RECT 406.200 657.300 408.300 659.400 ;
        RECT 409.950 658.950 412.050 661.050 ;
        RECT 388.800 650.400 390.900 652.500 ;
        RECT 392.700 645.900 393.600 656.400 ;
        RECT 395.100 649.950 397.200 652.050 ;
        RECT 386.100 642.900 388.200 645.000 ;
        RECT 391.500 643.800 393.600 645.900 ;
        RECT 383.100 637.500 385.200 639.600 ;
        RECT 380.700 630.600 382.800 635.700 ;
        RECT 383.700 632.700 385.200 637.500 ;
        RECT 386.700 635.700 387.900 642.900 ;
        RECT 392.700 637.200 393.600 643.800 ;
        RECT 386.100 633.600 388.200 635.700 ;
        RECT 391.500 635.100 393.600 637.200 ;
        RECT 395.400 647.400 396.600 649.650 ;
        RECT 383.700 630.600 385.800 632.700 ;
        RECT 373.950 616.950 376.050 619.050 ;
        RECT 367.800 609.000 369.900 610.050 ;
        RECT 367.800 607.950 370.050 609.000 ;
        RECT 370.950 607.950 373.050 610.050 ;
        RECT 361.950 605.100 364.050 607.200 ;
        RECT 367.950 605.100 370.050 607.950 ;
        RECT 382.950 605.100 385.050 607.200 ;
        RECT 388.950 606.000 391.050 610.050 ;
        RECT 395.400 606.450 396.450 647.400 ;
        RECT 401.100 635.700 402.300 657.300 ;
        RECT 400.200 633.600 402.300 635.700 ;
        RECT 403.500 640.800 404.700 657.300 ;
        RECT 406.500 653.700 407.700 657.300 ;
        RECT 406.500 651.600 408.600 653.700 ;
        RECT 403.500 638.700 405.600 640.800 ;
        RECT 403.500 632.700 404.700 638.700 ;
        RECT 407.100 632.700 408.600 651.600 ;
        RECT 402.600 630.600 404.700 632.700 ;
        RECT 405.600 630.600 408.600 632.700 ;
        RECT 410.400 625.050 411.450 658.950 ;
        RECT 413.100 643.950 415.200 646.050 ;
        RECT 419.100 643.950 421.200 646.050 ;
        RECT 419.400 642.900 420.600 643.650 ;
        RECT 418.950 640.800 421.050 642.900 ;
        RECT 421.950 631.950 424.050 634.050 ;
        RECT 400.950 622.950 403.050 625.050 ;
        RECT 409.950 622.950 412.050 625.050 ;
        RECT 418.950 622.950 421.050 625.050 ;
        RECT 362.400 604.350 363.600 605.100 ;
        RECT 368.400 604.350 369.600 605.100 ;
        RECT 383.400 604.350 384.600 605.100 ;
        RECT 389.400 604.350 390.600 606.000 ;
        RECT 395.400 605.400 399.450 606.450 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 382.950 601.950 385.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 365.400 599.400 366.600 601.650 ;
        RECT 386.400 599.400 387.600 601.650 ;
        RECT 392.400 600.900 393.600 601.650 ;
        RECT 355.950 595.950 358.050 598.050 ;
        RECT 349.950 589.950 352.050 592.050 ;
        RECT 349.950 586.800 352.050 588.900 ;
        RECT 344.400 569.400 348.450 570.450 ;
        RECT 344.400 568.350 345.600 569.400 ;
        RECT 335.100 565.950 337.200 568.050 ;
        RECT 340.950 565.950 343.050 568.050 ;
        RECT 344.100 565.950 346.200 568.050 ;
        RECT 337.950 559.950 340.050 562.050 ;
        RECT 331.950 535.950 334.050 538.050 ;
        RECT 338.400 532.050 339.450 559.950 ;
        RECT 337.950 529.950 340.050 532.050 ;
        RECT 322.950 527.100 325.050 529.200 ;
        RECT 323.400 526.350 324.600 527.100 ;
        RECT 331.950 526.950 334.050 529.050 ;
        RECT 335.100 526.950 337.200 529.050 ;
        RECT 323.100 523.950 325.200 526.050 ;
        RECT 328.500 523.950 330.600 526.050 ;
        RECT 329.400 522.900 330.600 523.650 ;
        RECT 328.950 520.800 331.050 522.900 ;
        RECT 332.400 522.450 333.450 526.950 ;
        RECT 335.400 525.900 336.600 526.650 ;
        RECT 334.800 523.800 336.900 525.900 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 332.400 521.400 336.450 522.450 ;
        RECT 329.400 519.450 330.450 520.800 ;
        RECT 329.400 518.400 333.450 519.450 ;
        RECT 316.950 502.950 319.050 505.050 ;
        RECT 310.950 499.950 313.050 502.050 ;
        RECT 327.000 498.450 331.050 499.050 ;
        RECT 326.400 496.950 331.050 498.450 ;
        RECT 305.400 493.350 306.600 495.600 ;
        RECT 310.950 494.100 313.050 496.200 ;
        RECT 316.950 494.100 319.050 496.200 ;
        RECT 326.400 495.600 327.450 496.950 ;
        RECT 332.400 496.050 333.450 518.400 ;
        RECT 311.400 493.350 312.600 494.100 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 304.950 490.950 307.050 493.050 ;
        RECT 307.950 490.950 310.050 493.050 ;
        RECT 310.950 490.950 313.050 493.050 ;
        RECT 302.400 489.900 303.600 490.650 ;
        RECT 295.950 487.800 298.050 489.900 ;
        RECT 301.950 487.800 304.050 489.900 ;
        RECT 308.400 488.400 309.600 490.650 ;
        RECT 308.400 486.450 309.450 488.400 ;
        RECT 305.400 485.400 309.450 486.450 ;
        RECT 292.950 481.950 295.050 484.050 ;
        RECT 295.950 469.950 298.050 472.050 ;
        RECT 296.400 466.050 297.450 469.950 ;
        RECT 289.950 463.950 292.050 466.050 ;
        RECT 295.950 463.950 298.050 466.050 ;
        RECT 289.950 451.950 292.050 454.050 ;
        RECT 286.950 436.950 289.050 439.050 ;
        RECT 283.950 433.950 286.050 436.050 ;
        RECT 268.950 430.950 271.050 433.050 ;
        RECT 274.950 418.950 277.050 421.050 ;
        RECT 265.950 416.100 268.050 418.200 ;
        RECT 271.950 416.100 274.050 418.200 ;
        RECT 266.400 415.350 267.600 416.100 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 263.400 411.900 264.600 412.650 ;
        RECT 272.400 412.050 273.450 416.100 ;
        RECT 262.950 409.800 265.050 411.900 ;
        RECT 271.950 409.950 274.050 412.050 ;
        RECT 275.400 406.050 276.450 418.950 ;
        RECT 284.400 417.600 285.450 433.950 ;
        RECT 290.400 427.050 291.450 451.950 ;
        RECT 305.400 450.600 306.450 485.400 ;
        RECT 317.400 456.450 318.450 494.100 ;
        RECT 326.400 493.350 327.600 495.600 ;
        RECT 331.950 493.950 334.050 496.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 323.400 489.900 324.600 490.650 ;
        RECT 322.950 487.800 325.050 489.900 ;
        RECT 329.400 488.400 330.600 490.650 ;
        RECT 329.400 484.050 330.450 488.400 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 329.400 469.050 330.450 481.950 ;
        RECT 328.950 466.950 331.050 469.050 ;
        RECT 314.400 455.400 318.450 456.450 ;
        RECT 296.400 450.450 297.600 450.600 ;
        RECT 293.400 449.400 297.600 450.450 ;
        RECT 293.400 442.050 294.450 449.400 ;
        RECT 296.400 448.350 297.600 449.400 ;
        RECT 305.400 448.350 306.600 450.600 ;
        RECT 296.100 445.950 298.200 448.050 ;
        RECT 301.500 445.950 303.600 448.050 ;
        RECT 304.800 445.950 306.900 448.050 ;
        RECT 302.400 444.900 303.600 445.650 ;
        RECT 314.400 445.050 315.450 455.400 ;
        RECT 322.950 449.100 325.050 451.200 ;
        RECT 323.400 448.350 324.600 449.100 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 301.950 442.800 304.050 444.900 ;
        RECT 313.950 442.950 316.050 445.050 ;
        RECT 320.400 444.000 321.600 445.650 ;
        RECT 326.400 444.900 327.600 445.650 ;
        RECT 292.950 439.950 295.050 442.050 ;
        RECT 301.950 439.650 304.050 441.750 ;
        RECT 319.950 439.950 322.050 444.000 ;
        RECT 325.950 442.800 328.050 444.900 ;
        RECT 292.950 430.950 295.050 433.050 ;
        RECT 289.950 424.950 292.050 427.050 ;
        RECT 284.400 415.350 285.600 417.600 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 281.400 411.900 282.600 412.650 ;
        RECT 280.950 409.800 283.050 411.900 ;
        RECT 287.400 411.450 288.600 412.650 ;
        RECT 287.400 410.400 291.450 411.450 ;
        RECT 274.950 403.950 277.050 406.050 ;
        RECT 268.950 397.950 271.050 400.050 ;
        RECT 256.950 388.950 259.050 391.050 ;
        RECT 226.950 379.950 229.050 382.050 ;
        RECT 247.950 379.950 250.050 382.050 ;
        RECT 259.950 379.950 262.050 382.050 ;
        RECT 229.950 376.950 232.050 379.050 ;
        RECT 230.400 372.600 231.450 376.950 ;
        RECT 248.400 376.050 249.450 379.950 ;
        RECT 224.400 370.350 225.600 372.600 ;
        RECT 230.400 370.350 231.600 372.600 ;
        RECT 235.950 372.000 238.050 376.050 ;
        RECT 241.950 373.950 244.050 376.050 ;
        RECT 247.950 373.950 250.050 376.050 ;
        RECT 236.400 370.350 237.600 372.000 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 226.950 367.950 229.050 370.050 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 227.400 366.000 228.600 367.650 ;
        RECT 233.400 366.900 234.600 367.650 ;
        RECT 217.950 361.950 220.050 364.050 ;
        RECT 223.950 361.950 226.050 364.050 ;
        RECT 226.950 361.950 229.050 366.000 ;
        RECT 232.950 364.800 235.050 366.900 ;
        RECT 214.950 358.950 217.050 361.050 ;
        RECT 205.950 352.950 208.050 355.050 ;
        RECT 211.950 349.950 214.050 352.050 ;
        RECT 202.950 339.000 205.050 343.050 ;
        RECT 212.400 339.600 213.450 349.950 ;
        RECT 214.950 346.950 217.050 349.050 ;
        RECT 215.400 343.050 216.450 346.950 ;
        RECT 214.950 340.950 217.050 343.050 ;
        RECT 220.950 340.950 223.050 343.050 ;
        RECT 203.400 337.350 204.600 339.000 ;
        RECT 212.400 337.350 213.600 339.600 ;
        RECT 202.800 334.950 204.900 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 217.500 334.950 219.600 337.050 ;
        RECT 205.950 331.950 208.050 334.050 ;
        RECT 209.400 333.000 210.600 334.650 ;
        RECT 218.400 333.450 219.600 334.650 ;
        RECT 221.400 333.450 222.450 340.950 ;
        RECT 206.400 328.050 207.450 331.950 ;
        RECT 208.950 328.950 211.050 333.000 ;
        RECT 218.400 332.400 222.450 333.450 ;
        RECT 214.950 328.950 217.050 331.050 ;
        RECT 205.950 325.950 208.050 328.050 ;
        RECT 211.950 316.950 214.050 319.050 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 206.400 298.050 207.450 307.950 ;
        RECT 205.950 294.000 208.050 298.050 ;
        RECT 206.400 292.350 207.600 294.000 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 199.950 286.950 202.050 289.050 ;
        RECT 203.400 287.400 204.600 289.650 ;
        RECT 196.950 244.950 199.050 247.050 ;
        RECT 200.400 244.050 201.450 286.950 ;
        RECT 203.400 283.050 204.450 287.400 ;
        RECT 202.950 280.950 205.050 283.050 ;
        RECT 212.400 277.050 213.450 316.950 ;
        RECT 215.400 288.450 216.450 328.950 ;
        RECT 224.400 316.050 225.450 361.950 ;
        RECT 232.950 361.650 235.050 363.750 ;
        RECT 226.950 349.950 229.050 352.050 ;
        RECT 227.400 325.050 228.450 349.950 ;
        RECT 229.950 343.950 232.050 346.050 ;
        RECT 226.950 322.950 229.050 325.050 ;
        RECT 223.950 313.950 226.050 316.050 ;
        RECT 230.400 307.050 231.450 343.950 ;
        RECT 233.400 340.050 234.450 361.650 ;
        RECT 238.950 358.950 241.050 361.050 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 239.400 339.600 240.450 358.950 ;
        RECT 242.400 346.050 243.450 373.950 ;
        RECT 260.400 372.600 261.450 379.950 ;
        RECT 251.400 372.450 252.600 372.600 ;
        RECT 248.400 371.400 252.600 372.450 ;
        RECT 244.950 355.950 247.050 358.050 ;
        RECT 245.400 349.050 246.450 355.950 ;
        RECT 244.950 346.950 247.050 349.050 ;
        RECT 241.950 343.950 244.050 346.050 ;
        RECT 239.400 337.350 240.600 339.600 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 232.950 331.950 235.050 334.050 ;
        RECT 236.400 332.400 237.600 334.650 ;
        RECT 242.400 333.900 243.600 334.650 ;
        RECT 233.400 322.050 234.450 331.950 ;
        RECT 236.400 328.050 237.450 332.400 ;
        RECT 241.950 331.800 244.050 333.900 ;
        RECT 235.950 325.950 238.050 328.050 ;
        RECT 232.950 319.950 235.050 322.050 ;
        RECT 248.400 313.050 249.450 371.400 ;
        RECT 251.400 370.350 252.600 371.400 ;
        RECT 260.400 370.350 261.600 372.600 ;
        RECT 265.950 370.950 268.050 373.050 ;
        RECT 251.100 367.950 253.200 370.050 ;
        RECT 254.400 367.950 256.500 370.050 ;
        RECT 259.800 367.950 261.900 370.050 ;
        RECT 254.400 366.900 255.600 367.650 ;
        RECT 253.950 364.800 256.050 366.900 ;
        RECT 266.400 360.450 267.450 370.950 ;
        RECT 269.400 366.900 270.450 397.950 ;
        RECT 281.400 385.050 282.450 409.800 ;
        RECT 286.950 406.950 289.050 409.050 ;
        RECT 280.950 382.950 283.050 385.050 ;
        RECT 271.950 371.100 274.050 373.200 ;
        RECT 272.400 370.350 273.600 371.100 ;
        RECT 272.100 367.950 274.200 370.050 ;
        RECT 277.500 367.950 279.600 370.050 ;
        RECT 283.950 367.950 286.050 370.050 ;
        RECT 268.950 364.800 271.050 366.900 ;
        RECT 278.400 366.450 279.600 367.650 ;
        RECT 278.400 365.400 282.450 366.450 ;
        RECT 263.400 359.400 267.450 360.450 ;
        RECT 250.950 346.950 253.050 349.050 ;
        RECT 241.950 310.950 244.050 313.050 ;
        RECT 247.950 310.950 250.050 313.050 ;
        RECT 229.950 304.950 232.050 307.050 ;
        RECT 223.950 294.450 226.050 295.200 ;
        RECT 223.950 293.400 228.450 294.450 ;
        RECT 223.950 293.100 226.050 293.400 ;
        RECT 224.400 292.350 225.600 293.100 ;
        RECT 218.400 289.950 220.500 292.050 ;
        RECT 223.800 289.950 225.900 292.050 ;
        RECT 218.400 288.450 219.600 289.650 ;
        RECT 215.400 287.400 219.600 288.450 ;
        RECT 217.950 283.950 220.050 286.050 ;
        RECT 211.950 274.950 214.050 277.050 ;
        RECT 205.950 268.950 208.050 271.050 ;
        RECT 206.400 261.600 207.450 268.950 ;
        RECT 206.400 259.350 207.600 261.600 ;
        RECT 214.950 260.100 217.050 262.200 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 209.400 255.900 210.600 256.650 ;
        RECT 208.950 253.800 211.050 255.900 ;
        RECT 208.950 244.950 211.050 247.050 ;
        RECT 199.950 241.950 202.050 244.050 ;
        RECT 205.950 241.950 208.050 244.050 ;
        RECT 193.950 232.950 196.050 235.050 ;
        RECT 190.950 229.950 193.050 232.050 ;
        RECT 194.400 222.450 195.450 232.950 ;
        RECT 196.950 229.950 199.050 232.050 ;
        RECT 191.400 221.400 195.450 222.450 ;
        RECT 191.400 216.600 192.450 221.400 ;
        RECT 197.400 216.600 198.450 229.950 ;
        RECT 191.400 214.350 192.600 216.600 ;
        RECT 197.400 214.350 198.600 216.600 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 199.950 211.950 202.050 214.050 ;
        RECT 194.400 210.900 195.600 211.650 ;
        RECT 193.950 208.800 196.050 210.900 ;
        RECT 200.400 209.400 201.600 211.650 ;
        RECT 193.950 202.950 196.050 205.050 ;
        RECT 187.950 182.100 190.050 184.200 ;
        RECT 194.400 183.600 195.450 202.950 ;
        RECT 200.400 202.050 201.450 209.400 ;
        RECT 199.950 199.950 202.050 202.050 ;
        RECT 184.950 169.950 187.050 172.050 ;
        RECT 188.400 169.050 189.450 182.100 ;
        RECT 194.400 181.350 195.600 183.600 ;
        RECT 199.950 182.100 202.050 184.200 ;
        RECT 206.400 184.050 207.450 241.950 ;
        RECT 200.400 181.350 201.600 182.100 ;
        RECT 205.950 181.950 208.050 184.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 197.400 176.400 198.600 178.650 ;
        RECT 203.400 177.000 204.600 178.650 ;
        RECT 209.400 177.450 210.450 244.950 ;
        RECT 215.400 235.050 216.450 260.100 ;
        RECT 218.400 241.050 219.450 283.950 ;
        RECT 220.950 277.950 223.050 280.050 ;
        RECT 221.400 262.050 222.450 277.950 ;
        RECT 227.400 268.050 228.450 293.400 ;
        RECT 230.400 280.050 231.450 304.950 ;
        RECT 235.950 293.100 238.050 295.200 ;
        RECT 242.400 294.600 243.450 310.950 ;
        RECT 236.400 292.350 237.600 293.100 ;
        RECT 242.400 292.350 243.600 294.600 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 238.950 289.950 241.050 292.050 ;
        RECT 241.950 289.950 244.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 239.400 288.900 240.600 289.650 ;
        RECT 238.950 286.800 241.050 288.900 ;
        RECT 245.400 288.000 246.600 289.650 ;
        RECT 244.950 283.950 247.050 288.000 ;
        RECT 229.950 277.950 232.050 280.050 ;
        RECT 235.950 274.950 238.050 277.050 ;
        RECT 241.950 274.950 244.050 277.050 ;
        RECT 226.950 265.950 229.050 268.050 ;
        RECT 220.950 259.950 223.050 262.050 ;
        RECT 226.950 260.100 229.050 262.200 ;
        RECT 227.400 259.350 228.600 260.100 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 224.400 256.050 225.600 256.650 ;
        RECT 220.950 254.400 225.600 256.050 ;
        RECT 230.400 254.400 231.600 256.650 ;
        RECT 220.950 253.950 225.000 254.400 ;
        RECT 230.400 241.050 231.450 254.400 ;
        RECT 232.950 241.950 235.050 244.050 ;
        RECT 217.950 238.950 220.050 241.050 ;
        RECT 229.950 238.950 232.050 241.050 ;
        RECT 214.950 232.950 217.050 235.050 ;
        RECT 226.950 232.950 229.050 235.050 ;
        RECT 214.950 226.950 217.050 229.050 ;
        RECT 211.950 223.950 214.050 226.050 ;
        RECT 212.400 217.050 213.450 223.950 ;
        RECT 211.950 214.950 214.050 217.050 ;
        RECT 215.400 216.600 216.450 226.950 ;
        RECT 215.400 214.350 216.600 216.600 ;
        RECT 220.950 215.100 223.050 217.200 ;
        RECT 227.400 217.050 228.450 232.950 ;
        RECT 229.950 217.950 232.050 220.050 ;
        RECT 221.400 214.350 222.600 215.100 ;
        RECT 226.950 214.950 229.050 217.050 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 211.950 208.950 214.050 211.050 ;
        RECT 218.400 210.900 219.600 211.650 ;
        RECT 212.400 202.050 213.450 208.950 ;
        RECT 217.950 208.800 220.050 210.900 ;
        RECT 224.400 210.450 225.600 211.650 ;
        RECT 226.950 210.450 229.050 211.050 ;
        RECT 224.400 209.400 229.050 210.450 ;
        RECT 226.950 208.950 229.050 209.400 ;
        RECT 223.950 205.950 226.050 208.050 ;
        RECT 211.950 199.950 214.050 202.050 ;
        RECT 220.950 199.950 223.050 202.050 ;
        RECT 211.950 181.950 214.050 184.050 ;
        RECT 221.400 183.600 222.450 199.950 ;
        RECT 224.400 193.050 225.450 205.950 ;
        RECT 223.950 190.950 226.050 193.050 ;
        RECT 224.400 187.050 225.450 190.950 ;
        RECT 223.950 184.950 226.050 187.050 ;
        RECT 227.400 183.600 228.450 208.950 ;
        RECT 230.400 205.050 231.450 217.950 ;
        RECT 233.400 217.050 234.450 241.950 ;
        RECT 236.400 220.050 237.450 274.950 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 239.400 262.050 240.450 268.950 ;
        RECT 238.950 259.950 241.050 262.050 ;
        RECT 242.400 261.600 243.450 274.950 ;
        RECT 242.400 259.350 243.600 261.600 ;
        RECT 247.950 261.000 250.050 265.050 ;
        RECT 251.400 264.450 252.450 346.950 ;
        RECT 256.950 339.000 259.050 343.050 ;
        RECT 263.400 340.050 264.450 359.400 ;
        RECT 265.950 352.950 268.050 355.050 ;
        RECT 257.400 337.350 258.600 339.000 ;
        RECT 262.950 337.950 265.050 340.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 260.400 333.900 261.600 334.650 ;
        RECT 259.800 331.800 261.900 333.900 ;
        RECT 262.950 331.950 265.050 334.050 ;
        RECT 253.950 319.950 256.050 322.050 ;
        RECT 254.400 295.050 255.450 319.950 ;
        RECT 263.400 295.050 264.450 331.950 ;
        RECT 266.400 325.050 267.450 352.950 ;
        RECT 281.400 352.050 282.450 365.400 ;
        RECT 280.950 349.950 283.050 352.050 ;
        RECT 277.950 346.950 280.050 349.050 ;
        RECT 268.950 343.950 271.050 346.050 ;
        RECT 265.950 322.950 268.050 325.050 ;
        RECT 253.950 292.950 256.050 295.050 ;
        RECT 260.400 294.450 261.600 294.600 ;
        RECT 262.950 294.450 265.050 295.050 ;
        RECT 260.400 293.400 265.050 294.450 ;
        RECT 260.400 292.350 261.600 293.400 ;
        RECT 262.950 292.950 265.050 293.400 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 257.400 287.400 258.600 289.650 ;
        RECT 257.400 283.050 258.450 287.400 ;
        RECT 262.950 286.950 265.050 289.050 ;
        RECT 256.950 280.950 259.050 283.050 ;
        RECT 251.400 263.400 255.450 264.450 ;
        RECT 248.400 259.350 249.600 261.000 ;
        RECT 241.950 256.950 244.050 259.050 ;
        RECT 244.950 256.950 247.050 259.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 245.400 255.900 246.600 256.650 ;
        RECT 244.950 253.800 247.050 255.900 ;
        RECT 247.950 250.950 250.050 253.050 ;
        RECT 244.950 247.950 247.050 250.050 ;
        RECT 235.950 217.950 238.050 220.050 ;
        RECT 232.950 214.950 235.050 217.050 ;
        RECT 238.950 215.100 241.050 217.200 ;
        RECT 239.400 214.350 240.600 215.100 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 236.400 210.900 237.600 211.650 ;
        RECT 235.950 208.800 238.050 210.900 ;
        RECT 245.400 210.450 246.450 247.950 ;
        RECT 248.400 223.050 249.450 250.950 ;
        RECT 254.400 250.050 255.450 263.400 ;
        RECT 256.950 262.950 259.050 265.050 ;
        RECT 263.400 264.450 264.450 286.950 ;
        RECT 269.400 274.050 270.450 343.950 ;
        RECT 278.400 340.200 279.450 346.950 ;
        RECT 284.400 346.050 285.450 367.950 ;
        RECT 287.400 358.050 288.450 406.950 ;
        RECT 290.400 405.450 291.450 410.400 ;
        RECT 293.400 409.050 294.450 430.950 ;
        RECT 295.950 427.950 298.050 430.050 ;
        RECT 296.400 418.050 297.450 427.950 ;
        RECT 302.400 424.050 303.450 439.650 ;
        RECT 335.400 436.050 336.450 521.400 ;
        RECT 338.400 511.050 339.450 523.950 ;
        RECT 337.950 508.950 340.050 511.050 ;
        RECT 337.950 496.950 340.050 499.050 ;
        RECT 338.400 489.900 339.450 496.950 ;
        RECT 341.400 496.050 342.450 565.950 ;
        RECT 350.400 564.450 351.450 586.800 ;
        RECT 365.400 586.050 366.450 599.400 ;
        RECT 364.950 583.950 367.050 586.050 ;
        RECT 353.700 579.300 355.800 581.400 ;
        RECT 347.400 563.400 351.450 564.450 ;
        RECT 347.400 532.050 348.450 563.400 ;
        RECT 354.300 561.600 355.800 579.300 ;
        RECT 353.700 559.500 355.800 561.600 ;
        RECT 354.300 554.700 355.800 559.500 ;
        RECT 353.700 552.600 355.800 554.700 ;
        RECT 356.700 579.300 358.800 581.400 ;
        RECT 359.700 579.300 361.800 581.400 ;
        RECT 362.700 579.300 364.800 581.400 ;
        RECT 356.700 557.700 357.900 579.300 ;
        RECT 359.700 561.600 361.200 579.300 ;
        RECT 362.700 567.000 363.900 579.300 ;
        RECT 368.100 578.400 370.200 580.500 ;
        RECT 376.200 579.300 378.300 581.400 ;
        RECT 379.200 579.300 381.300 581.400 ;
        RECT 382.200 579.300 384.300 581.400 ;
        RECT 364.800 572.400 366.900 574.500 ;
        RECT 368.700 567.900 369.600 578.400 ;
        RECT 371.100 571.950 373.200 574.050 ;
        RECT 371.400 570.900 372.600 571.650 ;
        RECT 370.950 568.800 373.050 570.900 ;
        RECT 362.100 564.900 364.200 567.000 ;
        RECT 367.500 565.800 369.600 567.900 ;
        RECT 359.100 559.500 361.200 561.600 ;
        RECT 356.700 552.600 358.800 557.700 ;
        RECT 359.700 554.700 361.200 559.500 ;
        RECT 362.700 557.700 363.900 564.900 ;
        RECT 368.700 559.200 369.600 565.800 ;
        RECT 362.100 555.600 364.200 557.700 ;
        RECT 367.500 557.100 369.600 559.200 ;
        RECT 377.100 557.700 378.300 579.300 ;
        RECT 376.200 555.600 378.300 557.700 ;
        RECT 379.500 562.800 380.700 579.300 ;
        RECT 382.500 575.700 383.700 579.300 ;
        RECT 382.500 573.600 384.600 575.700 ;
        RECT 379.500 560.700 381.600 562.800 ;
        RECT 379.500 554.700 380.700 560.700 ;
        RECT 383.100 554.700 384.600 573.600 ;
        RECT 359.700 552.600 361.800 554.700 ;
        RECT 378.600 552.600 380.700 554.700 ;
        RECT 381.600 552.600 384.600 554.700 ;
        RECT 386.400 547.050 387.450 599.400 ;
        RECT 391.950 598.800 394.050 600.900 ;
        RECT 398.400 595.050 399.450 605.400 ;
        RECT 401.400 601.050 402.450 622.950 ;
        RECT 415.950 619.800 418.050 621.900 ;
        RECT 403.950 604.950 406.050 607.050 ;
        RECT 412.950 606.000 415.050 610.050 ;
        RECT 400.950 598.950 403.050 601.050 ;
        RECT 397.950 592.950 400.050 595.050 ;
        RECT 400.950 583.950 403.050 586.050 ;
        RECT 391.950 574.950 394.050 577.050 ;
        RECT 392.400 571.050 393.450 574.950 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 401.400 568.050 402.450 583.950 ;
        RECT 389.100 565.950 391.200 568.050 ;
        RECT 395.100 565.950 397.200 568.050 ;
        RECT 400.950 565.950 403.050 568.050 ;
        RECT 395.400 565.050 396.600 565.650 ;
        RECT 395.400 562.950 400.050 565.050 ;
        RECT 385.950 544.950 388.050 547.050 ;
        RECT 353.700 540.300 355.800 542.400 ;
        RECT 349.950 535.950 352.050 538.050 ;
        RECT 346.950 529.950 349.050 532.050 ;
        RECT 344.100 526.950 346.200 529.050 ;
        RECT 344.400 525.450 345.600 526.650 ;
        RECT 350.400 525.450 351.450 535.950 ;
        RECT 354.300 535.500 355.800 540.300 ;
        RECT 353.700 533.400 355.800 535.500 ;
        RECT 344.400 524.400 351.450 525.450 ;
        RECT 346.950 520.950 349.050 523.050 ;
        RECT 343.950 517.950 346.050 520.050 ;
        RECT 344.400 499.050 345.450 517.950 ;
        RECT 343.950 496.950 346.050 499.050 ;
        RECT 340.950 493.950 343.050 496.050 ;
        RECT 347.400 495.600 348.450 520.950 ;
        RECT 354.300 515.700 355.800 533.400 ;
        RECT 353.700 513.600 355.800 515.700 ;
        RECT 356.700 537.300 358.800 542.400 ;
        RECT 359.700 540.300 361.800 542.400 ;
        RECT 378.600 540.300 380.700 542.400 ;
        RECT 381.600 540.300 384.600 542.400 ;
        RECT 385.950 541.800 388.050 543.900 ;
        RECT 356.700 515.700 357.900 537.300 ;
        RECT 359.700 535.500 361.200 540.300 ;
        RECT 362.100 537.300 364.200 539.400 ;
        RECT 359.100 533.400 361.200 535.500 ;
        RECT 359.700 515.700 361.200 533.400 ;
        RECT 362.700 530.100 363.900 537.300 ;
        RECT 367.500 535.800 369.600 537.900 ;
        RECT 376.200 537.300 378.300 539.400 ;
        RECT 362.100 528.000 364.200 530.100 ;
        RECT 368.700 529.200 369.600 535.800 ;
        RECT 362.700 515.700 363.900 528.000 ;
        RECT 367.500 527.100 369.600 529.200 ;
        RECT 364.800 520.500 366.900 522.600 ;
        RECT 368.700 516.600 369.600 527.100 ;
        RECT 370.950 524.100 373.050 526.200 ;
        RECT 371.400 523.350 372.600 524.100 ;
        RECT 371.100 520.950 373.200 523.050 ;
        RECT 356.700 513.600 358.800 515.700 ;
        RECT 359.700 513.600 361.800 515.700 ;
        RECT 362.700 513.600 364.800 515.700 ;
        RECT 368.100 514.500 370.200 516.600 ;
        RECT 377.100 515.700 378.300 537.300 ;
        RECT 379.500 534.300 380.700 540.300 ;
        RECT 379.500 532.200 381.600 534.300 ;
        RECT 379.500 515.700 380.700 532.200 ;
        RECT 383.100 521.400 384.600 540.300 ;
        RECT 386.400 523.050 387.450 541.800 ;
        RECT 395.400 531.600 396.450 562.950 ;
        RECT 400.950 562.800 403.050 564.900 ;
        RECT 401.400 555.450 402.450 562.800 ;
        RECT 398.400 555.000 402.450 555.450 ;
        RECT 397.950 554.400 402.450 555.000 ;
        RECT 397.950 550.950 400.050 554.400 ;
        RECT 404.400 553.050 405.450 604.950 ;
        RECT 413.400 604.350 414.600 606.000 ;
        RECT 407.400 601.950 409.500 604.050 ;
        RECT 412.500 601.950 414.600 604.050 ;
        RECT 407.400 600.900 408.600 601.650 ;
        RECT 416.400 601.050 417.450 619.800 ;
        RECT 406.950 598.800 409.050 600.900 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 419.400 589.050 420.450 622.950 ;
        RECT 422.400 601.050 423.450 631.950 ;
        RECT 425.400 616.050 426.450 667.950 ;
        RECT 427.950 661.950 430.050 664.050 ;
        RECT 428.400 622.050 429.450 661.950 ;
        RECT 427.950 619.950 430.050 622.050 ;
        RECT 424.950 613.950 427.050 616.050 ;
        RECT 431.400 610.200 432.450 667.950 ;
        RECT 437.400 655.050 438.450 679.950 ;
        RECT 439.950 655.950 442.050 658.050 ;
        RECT 436.950 652.950 439.050 655.050 ;
        RECT 440.400 651.600 441.450 655.950 ;
        RECT 443.400 654.450 444.450 703.800 ;
        RECT 446.400 703.050 447.450 742.950 ;
        RECT 449.400 723.900 450.450 755.400 ;
        RECT 460.950 745.950 463.050 748.050 ;
        RECT 461.400 729.600 462.450 745.950 ;
        RECT 467.400 742.050 468.450 763.950 ;
        RECT 470.400 755.400 471.900 774.300 ;
        RECT 474.300 768.300 475.500 774.300 ;
        RECT 473.400 766.200 475.500 768.300 ;
        RECT 470.400 753.300 472.500 755.400 ;
        RECT 471.300 749.700 472.500 753.300 ;
        RECT 474.300 749.700 475.500 766.200 ;
        RECT 476.700 771.300 478.800 773.400 ;
        RECT 482.400 772.050 483.450 796.950 ;
        RECT 488.100 791.700 489.300 813.300 ;
        RECT 487.200 789.600 489.300 791.700 ;
        RECT 490.500 796.800 491.700 813.300 ;
        RECT 493.500 809.700 494.700 813.300 ;
        RECT 493.500 807.600 495.600 809.700 ;
        RECT 490.500 794.700 492.600 796.800 ;
        RECT 490.500 788.700 491.700 794.700 ;
        RECT 494.100 788.700 495.600 807.600 ;
        RECT 497.400 799.050 498.450 871.950 ;
        RECT 502.950 811.950 505.050 814.050 ;
        RECT 503.400 805.050 504.450 811.950 ;
        RECT 506.400 811.050 507.450 884.100 ;
        RECT 511.950 883.950 514.050 886.050 ;
        RECT 518.400 885.600 519.450 892.950 ;
        RECT 518.400 883.350 519.600 885.600 ;
        RECT 523.950 884.100 526.050 886.200 ;
        RECT 535.950 884.100 538.050 889.050 ;
        RECT 541.950 884.100 544.050 886.200 ;
        RECT 547.950 884.100 550.050 886.200 ;
        RECT 556.950 885.000 559.050 889.050 ;
        RECT 575.400 885.600 576.450 914.100 ;
        RECT 581.400 892.050 582.450 919.950 ;
        RECT 596.400 919.350 597.600 920.100 ;
        RECT 595.800 916.950 597.900 919.050 ;
        RECT 601.800 916.950 603.900 919.050 ;
        RECT 584.400 913.950 586.500 916.050 ;
        RECT 589.800 913.950 591.900 916.050 ;
        RECT 584.400 912.000 585.600 913.650 ;
        RECT 583.950 907.950 586.050 912.000 ;
        RECT 608.400 911.400 609.900 930.300 ;
        RECT 612.300 924.300 613.500 930.300 ;
        RECT 611.400 922.200 613.500 924.300 ;
        RECT 608.400 909.300 610.500 911.400 ;
        RECT 609.300 905.700 610.500 909.300 ;
        RECT 612.300 905.700 613.500 922.200 ;
        RECT 614.700 927.300 616.800 929.400 ;
        RECT 614.700 905.700 615.900 927.300 ;
        RECT 623.400 925.800 625.500 927.900 ;
        RECT 628.800 927.300 630.900 929.400 ;
        RECT 623.400 919.200 624.300 925.800 ;
        RECT 629.100 920.100 630.300 927.300 ;
        RECT 631.800 925.500 633.300 930.300 ;
        RECT 634.200 927.300 636.300 932.400 ;
        RECT 631.800 923.400 633.900 925.500 ;
        RECT 623.400 917.100 625.500 919.200 ;
        RECT 628.800 918.000 630.900 920.100 ;
        RECT 619.950 914.100 622.050 916.200 ;
        RECT 620.400 913.350 621.600 914.100 ;
        RECT 619.800 910.950 621.900 913.050 ;
        RECT 623.400 906.600 624.300 917.100 ;
        RECT 626.100 910.500 628.200 912.600 ;
        RECT 608.700 903.600 610.800 905.700 ;
        RECT 611.700 903.600 613.800 905.700 ;
        RECT 614.700 903.600 616.800 905.700 ;
        RECT 622.800 904.500 624.900 906.600 ;
        RECT 629.100 905.700 630.300 918.000 ;
        RECT 631.800 905.700 633.300 923.400 ;
        RECT 635.100 905.700 636.300 927.300 ;
        RECT 628.200 903.600 630.300 905.700 ;
        RECT 631.200 903.600 633.300 905.700 ;
        RECT 634.200 903.600 636.300 905.700 ;
        RECT 637.200 930.300 639.300 932.400 ;
        RECT 737.700 930.300 739.800 932.400 ;
        RECT 637.200 925.500 638.700 930.300 ;
        RECT 658.950 925.950 661.050 928.050 ;
        RECT 637.200 923.400 639.300 925.500 ;
        RECT 637.200 905.700 638.700 923.400 ;
        RECT 646.800 916.950 648.900 919.050 ;
        RECT 655.800 916.950 657.900 919.050 ;
        RECT 647.400 915.450 648.600 916.650 ;
        RECT 644.400 914.400 648.600 915.450 ;
        RECT 656.400 914.400 657.600 916.650 ;
        RECT 644.400 913.050 645.450 914.400 ;
        RECT 643.950 910.950 646.050 913.050 ;
        RECT 637.200 903.600 639.300 905.700 ;
        RECT 598.950 898.950 601.050 901.050 ;
        RECT 580.950 889.950 583.050 892.050 ;
        RECT 589.950 889.950 592.050 892.050 ;
        RECT 524.400 883.350 525.600 884.100 ;
        RECT 536.400 883.350 537.600 884.100 ;
        RECT 542.400 883.350 543.600 884.100 ;
        RECT 514.950 880.950 517.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 515.400 879.900 516.600 880.650 ;
        RECT 521.400 879.900 522.600 880.650 ;
        RECT 514.950 877.800 517.050 879.900 ;
        RECT 520.950 877.800 523.050 879.900 ;
        RECT 539.400 878.400 540.600 880.650 ;
        RECT 548.400 880.050 549.450 884.100 ;
        RECT 557.400 883.350 558.600 885.000 ;
        RECT 575.400 883.350 576.600 885.600 ;
        RECT 580.950 884.100 583.050 886.200 ;
        RECT 581.400 883.350 582.600 884.100 ;
        RECT 586.950 883.950 589.050 886.050 ;
        RECT 553.950 880.950 556.050 883.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 571.950 880.950 574.050 883.050 ;
        RECT 574.950 880.950 577.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 539.400 871.050 540.450 878.400 ;
        RECT 547.950 877.950 550.050 880.050 ;
        RECT 554.400 878.400 555.600 880.650 ;
        RECT 572.400 878.400 573.600 880.650 ;
        RECT 578.400 878.400 579.600 880.650 ;
        RECT 587.400 879.900 588.450 883.950 ;
        RECT 548.400 874.050 549.450 877.950 ;
        RECT 547.950 871.950 550.050 874.050 ;
        RECT 538.950 868.950 541.050 871.050 ;
        RECT 547.950 859.950 550.050 862.050 ;
        RECT 548.400 841.200 549.450 859.950 ;
        RECT 554.400 856.050 555.450 878.400 ;
        RECT 553.950 853.950 556.050 856.050 ;
        RECT 554.400 844.050 555.450 853.950 ;
        RECT 553.950 841.950 556.050 844.050 ;
        RECT 529.950 839.100 532.050 841.200 ;
        RECT 530.400 838.350 531.600 839.100 ;
        RECT 535.800 838.950 537.900 841.050 ;
        RECT 538.950 838.950 541.050 841.050 ;
        RECT 547.950 839.100 550.050 841.200 ;
        RECT 562.950 840.000 565.050 844.050 ;
        RECT 509.100 835.950 511.200 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 527.400 834.900 528.600 835.650 ;
        RECT 526.950 832.800 529.050 834.900 ;
        RECT 508.950 826.950 511.050 829.050 ;
        RECT 505.950 808.950 508.050 811.050 ;
        RECT 509.400 805.050 510.450 826.950 ;
        RECT 536.400 823.050 537.450 838.950 ;
        RECT 529.950 820.950 532.050 823.050 ;
        RECT 535.950 820.950 538.050 823.050 ;
        RECT 514.950 811.950 517.050 814.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 500.100 799.950 502.200 802.050 ;
        RECT 506.100 799.950 508.200 802.050 ;
        RECT 496.950 796.950 499.050 799.050 ;
        RECT 506.400 798.900 507.600 799.650 ;
        RECT 505.950 796.800 508.050 798.900 ;
        RECT 511.950 796.950 514.050 802.050 ;
        RECT 506.400 793.050 507.450 796.800 ;
        RECT 505.950 790.950 508.050 793.050 ;
        RECT 489.600 786.600 491.700 788.700 ;
        RECT 492.600 786.600 495.600 788.700 ;
        RECT 515.400 781.050 516.450 811.950 ;
        RECT 517.950 805.950 520.050 808.050 ;
        RECT 520.950 807.600 525.000 808.050 ;
        RECT 530.400 807.600 531.450 820.950 ;
        RECT 535.950 817.800 538.050 819.900 ;
        RECT 536.400 808.050 537.450 817.800 ;
        RECT 520.950 805.950 525.600 807.600 ;
        RECT 518.400 798.900 519.450 805.950 ;
        RECT 524.400 805.350 525.600 805.950 ;
        RECT 530.400 805.350 531.600 807.600 ;
        RECT 535.950 805.950 538.050 808.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 529.950 802.950 532.050 805.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 520.950 799.950 523.050 802.050 ;
        RECT 527.400 801.900 528.600 802.650 ;
        RECT 517.950 796.800 520.050 798.900 ;
        RECT 521.400 790.050 522.450 799.950 ;
        RECT 526.950 799.800 529.050 801.900 ;
        RECT 533.400 800.400 534.600 802.650 ;
        RECT 539.400 802.050 540.450 838.950 ;
        RECT 548.400 838.350 549.600 839.100 ;
        RECT 563.400 838.350 564.600 840.000 ;
        RECT 568.950 839.100 571.050 841.200 ;
        RECT 572.400 841.050 573.450 878.400 ;
        RECT 578.400 871.050 579.450 878.400 ;
        RECT 586.950 877.800 589.050 879.900 ;
        RECT 577.950 868.950 580.050 871.050 ;
        RECT 578.400 847.050 579.450 868.950 ;
        RECT 590.400 850.050 591.450 889.950 ;
        RECT 599.400 885.600 600.450 898.950 ;
        RECT 616.950 895.950 619.050 898.050 ;
        RECT 607.950 886.950 610.050 889.050 ;
        RECT 599.400 883.350 600.600 885.600 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 598.950 880.950 601.050 883.050 ;
        RECT 596.400 879.900 597.600 880.650 ;
        RECT 608.400 879.900 609.450 886.950 ;
        RECT 617.400 885.600 618.450 895.950 ;
        RECT 617.400 883.350 618.600 885.600 ;
        RECT 622.950 884.100 625.050 886.200 ;
        RECT 623.400 883.350 624.600 884.100 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 628.950 881.100 631.050 883.200 ;
        RECT 638.400 882.450 639.600 882.600 ;
        RECT 635.400 881.400 639.600 882.450 ;
        RECT 595.950 877.800 598.050 879.900 ;
        RECT 607.950 877.800 610.050 879.900 ;
        RECT 614.400 878.400 615.600 880.650 ;
        RECT 620.400 879.900 621.600 880.650 ;
        RECT 629.400 880.350 630.600 881.100 ;
        RECT 614.400 874.050 615.450 878.400 ;
        RECT 619.950 877.800 622.050 879.900 ;
        RECT 629.100 877.950 631.200 880.050 ;
        RECT 601.950 871.950 604.050 874.050 ;
        RECT 613.950 871.950 616.050 874.050 ;
        RECT 589.950 847.950 592.050 850.050 ;
        RECT 577.950 844.950 580.050 847.050 ;
        RECT 578.400 843.450 579.450 844.950 ;
        RECT 575.400 842.400 579.450 843.450 ;
        RECT 569.400 838.350 570.600 839.100 ;
        RECT 571.950 838.950 574.050 841.050 ;
        RECT 542.400 835.950 544.500 838.050 ;
        RECT 547.800 835.950 549.900 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 542.400 834.900 543.600 835.650 ;
        RECT 566.400 834.900 567.600 835.650 ;
        RECT 541.950 832.800 544.050 834.900 ;
        RECT 565.950 832.800 568.050 834.900 ;
        RECT 571.950 832.950 574.050 835.050 ;
        RECT 566.400 831.450 567.450 832.800 ;
        RECT 566.400 830.400 570.450 831.450 ;
        RECT 565.950 823.950 568.050 826.050 ;
        RECT 556.950 814.950 559.050 817.050 ;
        RECT 547.950 811.950 550.050 814.050 ;
        RECT 548.400 807.600 549.450 811.950 ;
        RECT 548.400 805.350 549.600 807.600 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 550.950 802.950 553.050 805.050 ;
        RECT 523.800 793.950 525.900 796.050 ;
        RECT 526.950 793.950 529.050 798.750 ;
        RECT 520.950 787.950 523.050 790.050 ;
        RECT 484.950 778.950 487.050 781.050 ;
        RECT 514.950 778.950 517.050 781.050 ;
        RECT 485.400 775.050 486.450 778.950 ;
        RECT 484.950 772.950 487.050 775.050 ;
        RECT 493.200 774.300 495.300 776.400 ;
        RECT 476.700 749.700 477.900 771.300 ;
        RECT 481.950 769.950 484.050 772.050 ;
        RECT 482.400 766.050 483.450 769.950 ;
        RECT 485.400 769.800 487.500 771.900 ;
        RECT 490.800 771.300 492.900 773.400 ;
        RECT 481.950 763.950 484.050 766.050 ;
        RECT 485.400 763.200 486.300 769.800 ;
        RECT 491.100 764.100 492.300 771.300 ;
        RECT 493.800 769.500 495.300 774.300 ;
        RECT 496.200 771.300 498.300 776.400 ;
        RECT 493.800 767.400 495.900 769.500 ;
        RECT 485.400 761.100 487.500 763.200 ;
        RECT 490.800 762.000 492.900 764.100 ;
        RECT 481.950 758.100 484.050 760.200 ;
        RECT 482.400 757.350 483.600 758.100 ;
        RECT 481.800 754.950 483.900 757.050 ;
        RECT 485.400 750.600 486.300 761.100 ;
        RECT 488.100 754.500 490.200 756.600 ;
        RECT 470.700 747.600 472.800 749.700 ;
        RECT 473.700 747.600 475.800 749.700 ;
        RECT 476.700 747.600 478.800 749.700 ;
        RECT 484.800 748.500 486.900 750.600 ;
        RECT 491.100 749.700 492.300 762.000 ;
        RECT 493.800 749.700 495.300 767.400 ;
        RECT 497.100 749.700 498.300 771.300 ;
        RECT 490.200 747.600 492.300 749.700 ;
        RECT 493.200 747.600 495.300 749.700 ;
        RECT 496.200 747.600 498.300 749.700 ;
        RECT 499.200 774.300 501.300 776.400 ;
        RECT 499.200 769.500 500.700 774.300 ;
        RECT 520.950 772.950 523.050 775.050 ;
        RECT 499.200 767.400 501.300 769.500 ;
        RECT 499.200 749.700 500.700 767.400 ;
        RECT 511.950 766.950 514.050 769.050 ;
        RECT 502.950 760.950 505.050 763.050 ;
        RECT 508.800 760.950 510.900 763.050 ;
        RECT 499.200 747.600 501.300 749.700 ;
        RECT 503.400 745.050 504.450 760.950 ;
        RECT 509.400 759.450 510.600 760.650 ;
        RECT 512.400 759.450 513.450 766.950 ;
        RECT 517.800 760.950 519.900 763.050 ;
        RECT 509.400 758.400 513.450 759.450 ;
        RECT 518.400 758.400 519.600 760.650 ;
        RECT 518.400 754.050 519.450 758.400 ;
        RECT 511.950 751.950 514.050 754.050 ;
        RECT 517.950 751.950 520.050 754.050 ;
        RECT 481.950 742.950 484.050 745.050 ;
        RECT 502.950 742.950 505.050 745.050 ;
        RECT 466.950 739.950 469.050 742.050 ;
        RECT 466.950 736.800 469.050 738.900 ;
        RECT 467.400 733.050 468.450 736.800 ;
        RECT 461.400 727.350 462.600 729.600 ;
        RECT 466.950 729.000 469.050 733.050 ;
        RECT 482.400 730.200 483.450 742.950 ;
        RECT 502.950 739.800 505.050 741.900 ;
        RECT 467.400 727.350 468.600 729.000 ;
        RECT 481.950 728.100 484.050 730.200 ;
        RECT 503.400 729.600 504.450 739.800 ;
        RECT 482.400 727.350 483.600 728.100 ;
        RECT 503.400 727.350 504.600 729.600 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 460.950 724.950 463.050 727.050 ;
        RECT 463.950 724.950 466.050 727.050 ;
        RECT 466.950 724.950 469.050 727.050 ;
        RECT 482.400 724.950 484.500 727.050 ;
        RECT 487.800 724.950 489.900 727.050 ;
        RECT 499.950 724.950 502.050 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 458.400 723.900 459.600 724.650 ;
        RECT 448.950 721.800 451.050 723.900 ;
        RECT 457.950 721.800 460.050 723.900 ;
        RECT 464.400 723.000 465.600 724.650 ;
        RECT 488.400 723.900 489.600 724.650 ;
        RECT 500.400 723.900 501.600 724.650 ;
        RECT 506.400 723.900 507.600 724.650 ;
        RECT 463.950 718.950 466.050 723.000 ;
        RECT 487.950 721.800 490.050 723.900 ;
        RECT 499.950 721.800 502.050 723.900 ;
        RECT 505.950 721.800 508.050 723.900 ;
        RECT 512.400 723.450 513.450 751.950 ;
        RECT 514.950 745.950 517.050 748.050 ;
        RECT 515.400 723.900 516.450 745.950 ;
        RECT 521.400 745.050 522.450 772.950 ;
        RECT 520.950 742.950 523.050 745.050 ;
        RECT 524.400 729.600 525.450 793.950 ;
        RECT 529.950 787.950 532.050 790.050 ;
        RECT 530.400 775.050 531.450 787.950 ;
        RECT 533.400 781.050 534.450 800.400 ;
        RECT 538.950 799.950 541.050 802.050 ;
        RECT 545.400 801.450 546.600 802.650 ;
        RECT 551.400 801.900 552.600 802.650 ;
        RECT 557.400 801.900 558.450 814.950 ;
        RECT 566.400 807.600 567.450 823.950 ;
        RECT 569.400 810.450 570.450 830.400 ;
        RECT 572.400 826.050 573.450 832.950 ;
        RECT 571.950 823.950 574.050 826.050 ;
        RECT 569.400 810.000 573.450 810.450 ;
        RECT 569.400 809.400 574.050 810.000 ;
        RECT 566.400 805.350 567.600 807.600 ;
        RECT 571.950 805.950 574.050 809.400 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 568.950 802.950 571.050 805.050 ;
        RECT 563.400 801.900 564.600 802.650 ;
        RECT 569.400 801.900 570.600 802.650 ;
        RECT 575.400 802.050 576.450 842.400 ;
        RECT 583.950 839.100 586.050 841.200 ;
        RECT 602.400 840.600 603.450 871.950 ;
        RECT 613.950 853.950 616.050 856.050 ;
        RECT 614.400 841.050 615.450 853.950 ;
        RECT 635.400 850.050 636.450 881.400 ;
        RECT 638.400 880.350 639.600 881.400 ;
        RECT 638.100 877.950 640.200 880.050 ;
        RECT 644.400 862.050 645.450 910.950 ;
        RECT 656.400 910.050 657.450 914.400 ;
        RECT 659.400 913.050 660.450 925.950 ;
        RECT 738.300 925.500 739.800 930.300 ;
        RECT 737.700 923.400 739.800 925.500 ;
        RECT 673.950 917.100 676.050 919.200 ;
        RECT 674.400 916.350 675.600 917.100 ;
        RECT 694.950 916.950 697.050 919.050 ;
        RECT 719.100 916.950 721.200 919.050 ;
        RECT 728.100 916.950 730.200 919.050 ;
        RECT 670.950 913.950 673.050 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 686.100 913.950 688.200 916.050 ;
        RECT 691.500 913.950 693.600 916.050 ;
        RECT 658.950 910.950 661.050 913.050 ;
        RECT 671.400 912.900 672.600 913.650 ;
        RECT 670.950 910.800 673.050 912.900 ;
        RECT 692.400 911.400 693.600 913.650 ;
        RECT 655.950 907.950 658.050 910.050 ;
        RECT 656.400 901.050 657.450 907.950 ;
        RECT 655.950 898.950 658.050 901.050 ;
        RECT 647.700 891.300 649.800 893.400 ;
        RECT 648.300 873.600 649.800 891.300 ;
        RECT 647.700 871.500 649.800 873.600 ;
        RECT 648.300 866.700 649.800 871.500 ;
        RECT 647.700 864.600 649.800 866.700 ;
        RECT 650.700 891.300 652.800 893.400 ;
        RECT 653.700 891.300 655.800 893.400 ;
        RECT 656.700 891.300 658.800 893.400 ;
        RECT 650.700 869.700 651.900 891.300 ;
        RECT 653.700 873.600 655.200 891.300 ;
        RECT 656.700 879.000 657.900 891.300 ;
        RECT 662.100 890.400 664.200 892.500 ;
        RECT 670.200 891.300 672.300 893.400 ;
        RECT 673.200 891.300 675.300 893.400 ;
        RECT 676.200 891.300 678.300 893.400 ;
        RECT 658.800 884.400 660.900 886.500 ;
        RECT 662.700 879.900 663.600 890.400 ;
        RECT 665.100 883.950 667.200 886.050 ;
        RECT 665.400 882.900 666.600 883.650 ;
        RECT 664.950 880.800 667.050 882.900 ;
        RECT 656.100 876.900 658.200 879.000 ;
        RECT 661.500 877.800 663.600 879.900 ;
        RECT 653.100 871.500 655.200 873.600 ;
        RECT 650.700 864.600 652.800 869.700 ;
        RECT 653.700 866.700 655.200 871.500 ;
        RECT 656.700 869.700 657.900 876.900 ;
        RECT 662.700 871.200 663.600 877.800 ;
        RECT 656.100 867.600 658.200 869.700 ;
        RECT 661.500 869.100 663.600 871.200 ;
        RECT 671.100 869.700 672.300 891.300 ;
        RECT 670.200 867.600 672.300 869.700 ;
        RECT 673.500 874.800 674.700 891.300 ;
        RECT 676.500 887.700 677.700 891.300 ;
        RECT 685.950 889.950 688.050 892.050 ;
        RECT 676.500 885.600 678.600 887.700 ;
        RECT 673.500 872.700 675.600 874.800 ;
        RECT 673.500 866.700 674.700 872.700 ;
        RECT 677.100 866.700 678.600 885.600 ;
        RECT 686.400 883.050 687.450 889.950 ;
        RECT 692.400 883.050 693.450 911.400 ;
        RECT 683.400 882.450 684.600 882.600 ;
        RECT 680.400 881.400 684.600 882.450 ;
        RECT 680.400 877.050 681.450 881.400 ;
        RECT 683.400 880.350 684.600 881.400 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 691.950 880.950 694.050 883.050 ;
        RECT 683.100 877.950 685.200 880.050 ;
        RECT 689.100 877.950 691.200 880.050 ;
        RECT 679.950 874.950 682.050 877.050 ;
        RECT 685.950 874.950 688.050 877.050 ;
        RECT 682.950 868.950 685.050 871.050 ;
        RECT 653.700 864.600 655.800 866.700 ;
        RECT 672.600 864.600 674.700 866.700 ;
        RECT 675.600 864.600 678.600 866.700 ;
        RECT 637.950 859.950 640.050 862.050 ;
        RECT 643.950 859.950 646.050 862.050 ;
        RECT 673.950 859.950 676.050 862.050 ;
        RECT 638.400 853.050 639.450 859.950 ;
        RECT 637.950 850.950 640.050 853.050 ;
        RECT 641.400 852.300 644.400 854.400 ;
        RECT 645.300 852.300 647.400 854.400 ;
        RECT 664.200 852.300 666.300 854.400 ;
        RECT 628.950 847.950 631.050 850.050 ;
        RECT 634.950 847.950 637.050 850.050 ;
        RECT 629.400 843.600 630.450 847.950 ;
        RECT 629.400 841.350 630.600 843.600 ;
        RECT 584.400 838.350 585.600 839.100 ;
        RECT 602.400 838.350 603.600 840.600 ;
        RECT 610.950 838.950 613.050 841.050 ;
        RECT 613.950 838.950 616.050 841.050 ;
        RECT 619.950 839.100 622.050 841.200 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 581.400 833.400 582.600 835.650 ;
        RECT 587.400 834.000 588.600 835.650 ;
        RECT 605.400 834.000 606.600 835.650 ;
        RECT 577.950 805.950 580.050 808.050 ;
        RECT 578.400 802.050 579.450 805.950 ;
        RECT 542.400 800.400 546.600 801.450 ;
        RECT 538.950 796.800 541.050 798.900 ;
        RECT 535.950 793.950 538.050 796.050 ;
        RECT 532.950 778.950 535.050 781.050 ;
        RECT 536.400 775.050 537.450 793.950 ;
        RECT 529.950 772.950 532.050 775.050 ;
        RECT 535.950 772.950 538.050 775.050 ;
        RECT 539.400 769.050 540.450 796.800 ;
        RECT 542.400 790.050 543.450 800.400 ;
        RECT 550.950 799.800 553.050 801.900 ;
        RECT 556.950 799.800 559.050 801.900 ;
        RECT 562.950 799.800 565.050 801.900 ;
        RECT 568.950 799.800 571.050 801.900 ;
        RECT 574.800 799.950 576.900 802.050 ;
        RECT 577.950 799.950 580.050 802.050 ;
        RECT 577.950 796.800 580.050 798.900 ;
        RECT 547.950 793.950 550.050 796.050 ;
        RECT 541.950 787.950 544.050 790.050 ;
        RECT 541.950 784.800 544.050 786.900 ;
        RECT 532.950 766.950 535.050 769.050 ;
        RECT 538.950 766.950 541.050 769.050 ;
        RECT 527.100 760.950 529.200 763.050 ;
        RECT 527.400 758.400 528.600 760.650 ;
        RECT 527.400 733.050 528.450 758.400 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 533.400 759.450 534.450 766.950 ;
        RECT 536.100 760.950 538.200 763.050 ;
        RECT 536.400 759.450 537.600 760.650 ;
        RECT 533.400 758.400 537.600 759.450 ;
        RECT 530.400 738.450 531.450 757.950 ;
        RECT 538.950 754.950 541.050 757.050 ;
        RECT 535.950 751.950 538.050 754.050 ;
        RECT 530.400 737.400 534.450 738.450 ;
        RECT 529.950 733.950 532.050 736.050 ;
        RECT 526.950 730.950 529.050 733.050 ;
        RECT 530.400 729.600 531.450 733.950 ;
        RECT 533.400 730.050 534.450 737.400 ;
        RECT 536.400 733.050 537.450 751.950 ;
        RECT 539.400 748.050 540.450 754.950 ;
        RECT 538.950 745.950 541.050 748.050 ;
        RECT 538.950 739.950 541.050 742.050 ;
        RECT 535.950 730.950 538.050 733.050 ;
        RECT 524.400 727.350 525.600 729.600 ;
        RECT 530.400 727.350 531.600 729.600 ;
        RECT 532.800 727.950 534.900 730.050 ;
        RECT 535.950 727.800 538.050 729.900 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 523.950 724.950 526.050 727.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 521.400 723.900 522.600 724.650 ;
        RECT 527.400 723.900 528.600 724.650 ;
        RECT 509.400 722.400 513.450 723.450 ;
        RECT 484.950 718.950 487.050 721.050 ;
        RECT 457.950 706.950 460.050 709.050 ;
        RECT 478.950 706.950 481.050 709.050 ;
        RECT 445.950 700.950 448.050 703.050 ;
        RECT 446.400 696.300 449.400 698.400 ;
        RECT 450.300 696.300 452.400 698.400 ;
        RECT 446.400 677.400 447.900 696.300 ;
        RECT 450.300 690.300 451.500 696.300 ;
        RECT 449.400 688.200 451.500 690.300 ;
        RECT 446.400 675.300 448.500 677.400 ;
        RECT 447.300 671.700 448.500 675.300 ;
        RECT 450.300 671.700 451.500 688.200 ;
        RECT 452.700 693.300 454.800 695.400 ;
        RECT 452.700 671.700 453.900 693.300 ;
        RECT 454.950 685.950 457.050 688.050 ;
        RECT 455.400 681.450 456.450 685.950 ;
        RECT 458.400 685.050 459.450 706.950 ;
        RECT 469.200 696.300 471.300 698.400 ;
        RECT 461.400 691.800 463.500 693.900 ;
        RECT 466.800 693.300 468.900 695.400 ;
        RECT 461.400 685.200 462.300 691.800 ;
        RECT 467.100 686.100 468.300 693.300 ;
        RECT 469.800 691.500 471.300 696.300 ;
        RECT 472.200 693.300 474.300 698.400 ;
        RECT 469.800 689.400 471.900 691.500 ;
        RECT 457.950 682.950 460.050 685.050 ;
        RECT 461.400 683.100 463.500 685.200 ;
        RECT 466.800 684.000 468.900 686.100 ;
        RECT 458.400 681.450 459.600 681.600 ;
        RECT 455.400 680.400 459.600 681.450 ;
        RECT 458.400 679.350 459.600 680.400 ;
        RECT 457.800 676.950 459.900 679.050 ;
        RECT 461.400 672.600 462.300 683.100 ;
        RECT 464.100 676.500 466.200 678.600 ;
        RECT 446.700 669.600 448.800 671.700 ;
        RECT 449.700 669.600 451.800 671.700 ;
        RECT 452.700 669.600 454.800 671.700 ;
        RECT 460.800 670.500 462.900 672.600 ;
        RECT 467.100 671.700 468.300 684.000 ;
        RECT 469.800 671.700 471.300 689.400 ;
        RECT 473.100 671.700 474.300 693.300 ;
        RECT 466.200 669.600 468.300 671.700 ;
        RECT 469.200 669.600 471.300 671.700 ;
        RECT 472.200 669.600 474.300 671.700 ;
        RECT 475.200 696.300 477.300 698.400 ;
        RECT 475.200 691.500 476.700 696.300 ;
        RECT 475.200 689.400 477.300 691.500 ;
        RECT 475.200 671.700 476.700 689.400 ;
        RECT 475.200 669.600 477.300 671.700 ;
        RECT 463.950 664.950 466.050 667.050 ;
        RECT 448.950 655.950 451.050 658.050 ;
        RECT 443.400 654.000 447.450 654.450 ;
        RECT 443.400 653.400 448.050 654.000 ;
        RECT 440.400 649.350 441.600 651.600 ;
        RECT 445.950 649.950 448.050 653.400 ;
        RECT 436.950 646.950 439.050 649.050 ;
        RECT 439.950 646.950 442.050 649.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 437.400 644.400 438.600 646.650 ;
        RECT 443.400 645.900 444.600 646.650 ;
        RECT 437.400 637.050 438.450 644.400 ;
        RECT 442.950 643.800 445.050 645.900 ;
        RECT 439.950 640.950 442.050 643.050 ;
        RECT 436.950 634.950 439.050 637.050 ;
        RECT 437.400 628.050 438.450 634.950 ;
        RECT 436.950 625.950 439.050 628.050 ;
        RECT 436.950 619.950 439.050 622.050 ;
        RECT 433.950 616.950 436.050 619.050 ;
        RECT 430.950 608.100 433.050 610.200 ;
        RECT 434.400 610.050 435.450 616.950 ;
        RECT 433.950 607.950 436.050 610.050 ;
        RECT 430.950 604.950 433.050 607.050 ;
        RECT 437.400 606.600 438.450 619.950 ;
        RECT 440.400 607.050 441.450 640.950 ;
        RECT 449.400 622.050 450.450 655.950 ;
        RECT 451.950 652.950 454.050 655.050 ;
        RECT 448.950 619.950 451.050 622.050 ;
        RECT 452.400 619.050 453.450 652.950 ;
        RECT 460.950 651.000 463.050 655.050 ;
        RECT 461.400 649.350 462.600 651.000 ;
        RECT 464.400 649.050 465.450 664.950 ;
        RECT 472.950 658.950 475.050 661.050 ;
        RECT 455.100 646.950 457.200 649.050 ;
        RECT 460.500 646.950 462.600 649.050 ;
        RECT 463.950 646.950 466.050 649.050 ;
        RECT 455.400 645.000 456.600 646.650 ;
        RECT 454.950 640.800 457.050 645.000 ;
        RECT 457.950 634.950 460.050 637.050 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 455.400 622.050 456.450 628.950 ;
        RECT 454.950 619.950 457.050 622.050 ;
        RECT 451.950 616.950 454.050 619.050 ;
        RECT 448.950 610.950 451.050 613.050 ;
        RECT 431.400 604.350 432.600 604.950 ;
        RECT 437.400 604.350 438.600 606.600 ;
        RECT 439.950 604.950 442.050 607.050 ;
        RECT 443.100 604.950 445.200 607.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 443.400 602.400 444.600 604.650 ;
        RECT 421.950 598.950 424.050 601.050 ;
        RECT 424.950 598.950 427.050 601.050 ;
        RECT 428.400 599.400 429.600 601.650 ;
        RECT 434.400 599.400 435.600 601.650 ;
        RECT 418.950 586.950 421.050 589.050 ;
        RECT 406.950 577.950 409.050 580.050 ;
        RECT 421.950 577.950 424.050 580.050 ;
        RECT 407.400 568.050 408.450 577.950 ;
        RECT 415.950 573.000 418.050 577.050 ;
        RECT 422.400 573.600 423.450 577.950 ;
        RECT 425.400 574.050 426.450 598.950 ;
        RECT 428.400 595.050 429.450 599.400 ;
        RECT 427.950 592.950 430.050 595.050 ;
        RECT 434.400 592.050 435.450 599.400 ;
        RECT 433.950 589.950 436.050 592.050 ;
        RECT 427.950 586.950 430.050 589.050 ;
        RECT 416.400 571.350 417.600 573.000 ;
        RECT 422.400 571.350 423.600 573.600 ;
        RECT 424.950 571.950 427.050 574.050 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 418.950 568.950 421.050 571.050 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 406.950 565.950 409.050 568.050 ;
        RECT 413.400 567.900 414.600 568.650 ;
        RECT 412.950 565.800 415.050 567.900 ;
        RECT 419.400 567.000 420.600 568.650 ;
        RECT 406.950 562.800 409.050 564.900 ;
        RECT 418.950 562.950 421.050 567.000 ;
        RECT 428.400 565.050 429.450 586.950 ;
        RECT 443.400 586.050 444.450 602.400 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 442.950 583.950 445.050 586.050 ;
        RECT 433.950 577.950 436.050 580.050 ;
        RECT 434.400 573.600 435.450 577.950 ;
        RECT 434.400 571.350 435.600 573.600 ;
        RECT 439.950 573.000 442.050 577.050 ;
        RECT 446.400 574.050 447.450 601.950 ;
        RECT 440.400 571.350 441.600 573.000 ;
        RECT 445.950 571.950 448.050 574.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 439.950 568.950 442.050 571.050 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 430.950 565.950 433.050 568.050 ;
        RECT 437.400 566.400 438.600 568.650 ;
        RECT 443.400 566.400 444.600 568.650 ;
        RECT 427.950 562.950 430.050 565.050 ;
        RECT 407.400 559.050 408.450 562.800 ;
        RECT 406.950 556.950 409.050 559.050 ;
        RECT 424.950 556.950 427.050 559.050 ;
        RECT 415.950 553.950 418.050 556.050 ;
        RECT 404.400 552.450 409.050 553.050 ;
        RECT 401.400 551.400 409.050 552.450 ;
        RECT 401.400 549.450 402.450 551.400 ;
        RECT 405.000 550.950 409.050 551.400 ;
        RECT 398.400 548.400 402.450 549.450 ;
        RECT 398.400 532.050 399.450 548.400 ;
        RECT 403.950 547.950 406.050 550.050 ;
        RECT 400.950 541.950 403.050 547.050 ;
        RECT 400.950 532.950 403.050 535.050 ;
        RECT 395.400 529.350 396.600 531.600 ;
        RECT 397.950 529.950 400.050 532.050 ;
        RECT 389.100 526.950 391.200 529.050 ;
        RECT 395.100 526.950 397.200 529.050 ;
        RECT 401.400 526.050 402.450 532.950 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 382.500 519.300 384.600 521.400 ;
        RECT 385.950 520.950 388.050 523.050 ;
        RECT 382.500 515.700 383.700 519.300 ;
        RECT 376.200 513.600 378.300 515.700 ;
        RECT 379.200 513.600 381.300 515.700 ;
        RECT 382.200 513.600 384.300 515.700 ;
        RECT 385.950 511.950 388.050 514.050 ;
        RECT 373.950 508.950 376.050 511.050 ;
        RECT 354.000 495.600 358.050 496.050 ;
        RECT 347.400 493.350 348.600 495.600 ;
        RECT 353.400 495.450 358.050 495.600 ;
        RECT 353.400 494.400 360.450 495.450 ;
        RECT 353.400 493.950 358.050 494.400 ;
        RECT 353.400 493.350 354.600 493.950 ;
        RECT 343.950 490.950 346.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 349.950 490.950 352.050 493.050 ;
        RECT 352.950 490.950 355.050 493.050 ;
        RECT 344.400 489.900 345.600 490.650 ;
        RECT 350.400 489.900 351.600 490.650 ;
        RECT 337.950 487.800 340.050 489.900 ;
        RECT 343.950 487.800 346.050 489.900 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 343.950 481.950 346.050 484.050 ;
        RECT 340.950 478.950 343.050 481.050 ;
        RECT 310.950 433.950 313.050 436.050 ;
        RECT 334.950 433.950 337.050 436.050 ;
        RECT 301.950 421.950 304.050 424.050 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 302.400 417.600 303.450 421.950 ;
        RECT 302.400 415.350 303.600 417.600 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 299.400 411.900 300.600 412.650 ;
        RECT 305.400 411.900 306.600 412.650 ;
        RECT 311.400 411.900 312.450 433.950 ;
        RECT 316.950 417.000 319.050 421.050 ;
        RECT 325.950 418.950 328.050 421.050 ;
        RECT 317.400 415.350 318.600 417.000 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 298.950 409.800 301.050 411.900 ;
        RECT 304.950 409.800 307.050 411.900 ;
        RECT 310.950 409.800 313.050 411.900 ;
        RECT 320.400 410.400 321.600 412.650 ;
        RECT 292.950 406.950 295.050 409.050 ;
        RECT 290.400 404.400 294.450 405.450 ;
        RECT 289.950 388.950 292.050 391.050 ;
        RECT 290.400 361.050 291.450 388.950 ;
        RECT 293.400 388.050 294.450 404.400 ;
        RECT 298.950 400.950 301.050 403.050 ;
        RECT 292.950 385.950 295.050 388.050 ;
        RECT 293.400 376.050 294.450 385.950 ;
        RECT 292.950 373.950 295.050 376.050 ;
        RECT 299.400 375.450 300.450 400.950 ;
        RECT 305.400 382.050 306.450 409.800 ;
        RECT 320.400 406.050 321.450 410.400 ;
        RECT 319.950 403.950 322.050 406.050 ;
        RECT 307.950 394.950 310.050 397.050 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 299.400 374.400 303.450 375.450 ;
        RECT 298.950 371.100 301.050 373.200 ;
        RECT 299.400 370.350 300.600 371.100 ;
        RECT 293.400 367.950 295.500 370.050 ;
        RECT 298.800 367.950 300.900 370.050 ;
        RECT 293.400 366.900 294.600 367.650 ;
        RECT 302.400 366.900 303.450 374.400 ;
        RECT 292.950 364.800 295.050 366.900 ;
        RECT 301.950 364.800 304.050 366.900 ;
        RECT 289.950 358.950 292.050 361.050 ;
        RECT 286.950 355.950 289.050 358.050 ;
        RECT 293.400 352.050 294.450 364.800 ;
        RECT 301.950 357.450 304.050 361.050 ;
        RECT 301.950 357.000 306.450 357.450 ;
        RECT 302.400 356.400 306.450 357.000 ;
        RECT 292.950 349.950 295.050 352.050 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 283.950 343.950 286.050 346.050 ;
        RECT 277.950 338.100 280.050 340.200 ;
        RECT 284.400 339.600 285.450 343.950 ;
        RECT 299.400 343.050 300.450 349.950 ;
        RECT 305.400 343.050 306.450 356.400 ;
        RECT 289.950 340.950 292.050 343.050 ;
        RECT 298.950 340.950 301.050 343.050 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 278.400 337.350 279.600 338.100 ;
        RECT 284.400 337.350 285.600 339.600 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 277.950 334.950 280.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 275.400 332.400 276.600 334.650 ;
        RECT 281.400 333.900 282.600 334.650 ;
        RECT 290.400 333.900 291.450 340.950 ;
        RECT 301.950 338.100 304.050 340.200 ;
        RECT 308.400 339.600 309.450 394.950 ;
        RECT 316.950 391.950 319.050 394.050 ;
        RECT 317.400 372.600 318.450 391.950 ;
        RECT 317.400 370.350 318.600 372.600 ;
        RECT 326.400 370.050 327.450 418.950 ;
        RECT 328.950 416.100 331.050 418.200 ;
        RECT 334.950 416.100 337.050 418.200 ;
        RECT 341.400 417.600 342.450 478.950 ;
        RECT 344.400 450.600 345.450 481.950 ;
        RECT 344.400 448.350 345.600 450.600 ;
        RECT 344.100 445.950 346.200 448.050 ;
        RECT 349.500 445.950 351.600 448.050 ;
        RECT 350.400 443.400 351.600 445.650 ;
        RECT 356.400 445.050 357.450 487.950 ;
        RECT 359.400 475.050 360.450 494.400 ;
        RECT 367.950 494.100 370.050 496.200 ;
        RECT 374.400 495.600 375.450 508.950 ;
        RECT 382.950 505.950 385.050 508.050 ;
        RECT 368.400 493.350 369.600 494.100 ;
        RECT 374.400 493.350 375.600 495.600 ;
        RECT 367.950 490.950 370.050 493.050 ;
        RECT 370.950 490.950 373.050 493.050 ;
        RECT 373.950 490.950 376.050 493.050 ;
        RECT 376.950 490.950 379.050 493.050 ;
        RECT 371.400 489.000 372.600 490.650 ;
        RECT 377.400 489.900 378.600 490.650 ;
        RECT 370.950 484.950 373.050 489.000 ;
        RECT 376.950 487.800 379.050 489.900 ;
        RECT 376.950 484.650 379.050 486.750 ;
        RECT 358.950 472.950 361.050 475.050 ;
        RECT 364.950 469.950 367.050 472.050 ;
        RECT 365.400 466.050 366.450 469.950 ;
        RECT 364.950 463.950 367.050 466.050 ;
        RECT 373.950 463.950 376.050 466.050 ;
        RECT 367.950 460.950 370.050 463.050 ;
        RECT 358.950 454.950 361.050 457.050 ;
        RECT 350.400 433.050 351.450 443.400 ;
        RECT 355.950 442.950 358.050 445.050 ;
        RECT 359.400 441.450 360.450 454.950 ;
        RECT 368.400 450.600 369.450 460.950 ;
        RECT 368.400 448.350 369.600 450.600 ;
        RECT 362.400 445.950 364.500 448.050 ;
        RECT 367.800 445.950 369.900 448.050 ;
        RECT 362.400 444.900 363.600 445.650 ;
        RECT 361.950 442.800 364.050 444.900 ;
        RECT 359.400 440.400 363.450 441.450 ;
        RECT 349.950 430.950 352.050 433.050 ;
        RECT 329.400 373.050 330.450 416.100 ;
        RECT 335.400 415.350 336.600 416.100 ;
        RECT 341.400 415.350 342.600 417.600 ;
        RECT 349.950 416.100 352.050 418.200 ;
        RECT 355.950 416.100 358.050 418.200 ;
        RECT 362.400 417.600 363.450 440.400 ;
        RECT 367.950 424.950 370.050 427.050 ;
        RECT 368.400 418.050 369.450 424.950 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 338.400 410.400 339.600 412.650 ;
        RECT 334.950 403.950 337.050 406.050 ;
        RECT 328.950 370.950 331.050 373.050 ;
        RECT 335.400 372.600 336.450 403.950 ;
        RECT 338.400 394.050 339.450 410.400 ;
        RECT 346.950 403.950 349.050 406.050 ;
        RECT 337.950 391.950 340.050 394.050 ;
        RECT 342.000 372.600 346.050 373.050 ;
        RECT 335.400 370.350 336.600 372.600 ;
        RECT 341.400 370.950 346.050 372.600 ;
        RECT 341.400 370.350 342.600 370.950 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 337.950 367.950 340.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 314.400 366.900 315.600 367.650 ;
        RECT 313.950 364.800 316.050 366.900 ;
        RECT 320.400 366.000 321.600 367.650 ;
        RECT 332.400 367.050 333.600 367.650 ;
        RECT 319.950 361.950 322.050 366.000 ;
        RECT 328.950 365.400 333.600 367.050 ;
        RECT 338.400 366.000 339.600 367.650 ;
        RECT 328.950 364.950 333.000 365.400 ;
        RECT 325.950 361.950 328.050 364.050 ;
        RECT 334.950 361.950 337.050 364.050 ;
        RECT 337.950 361.950 340.050 366.000 ;
        RECT 313.950 349.950 316.050 352.050 ;
        RECT 302.400 337.350 303.600 338.100 ;
        RECT 308.400 337.350 309.600 339.600 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 304.950 334.950 307.050 337.050 ;
        RECT 307.950 334.950 310.050 337.050 ;
        RECT 275.400 328.050 276.450 332.400 ;
        RECT 280.950 331.800 283.050 333.900 ;
        RECT 289.950 331.800 292.050 333.900 ;
        RECT 299.400 333.000 300.600 334.650 ;
        RECT 305.400 333.900 306.600 334.650 ;
        RECT 314.400 333.900 315.450 349.950 ;
        RECT 316.950 337.950 319.050 340.050 ;
        RECT 326.400 339.600 327.450 361.950 ;
        RECT 295.950 328.950 298.050 331.050 ;
        RECT 298.950 328.950 301.050 333.000 ;
        RECT 304.950 331.800 307.050 333.900 ;
        RECT 313.950 331.800 316.050 333.900 ;
        RECT 317.400 333.450 318.450 337.950 ;
        RECT 326.400 337.350 327.600 339.600 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 328.950 334.950 331.050 337.050 ;
        RECT 323.400 333.450 324.600 334.650 ;
        RECT 317.400 332.400 324.600 333.450 ;
        RECT 329.400 333.000 330.600 334.650 ;
        RECT 301.950 328.950 304.050 331.050 ;
        RECT 307.950 328.950 310.050 331.050 ;
        RECT 274.950 325.950 277.050 328.050 ;
        RECT 296.400 319.050 297.450 328.950 ;
        RECT 298.950 322.800 301.050 324.900 ;
        RECT 277.950 316.950 280.050 319.050 ;
        RECT 295.950 316.950 298.050 319.050 ;
        RECT 278.400 295.050 279.450 316.950 ;
        RECT 280.950 313.950 283.050 316.050 ;
        RECT 277.950 292.950 280.050 295.050 ;
        RECT 281.400 294.600 282.450 313.950 ;
        RECT 289.950 307.950 292.050 310.050 ;
        RECT 290.400 294.600 291.450 307.950 ;
        RECT 295.950 301.950 298.050 304.050 ;
        RECT 292.950 298.950 295.050 301.050 ;
        RECT 281.400 292.350 282.600 294.600 ;
        RECT 290.400 292.350 291.600 294.600 ;
        RECT 274.800 289.950 276.900 292.050 ;
        RECT 280.950 289.950 283.050 292.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 289.500 289.950 291.600 292.050 ;
        RECT 275.400 288.450 276.600 289.650 ;
        RECT 277.950 288.450 280.050 289.050 ;
        RECT 284.400 288.900 285.600 289.650 ;
        RECT 275.400 287.400 280.050 288.450 ;
        RECT 277.950 286.950 280.050 287.400 ;
        RECT 278.400 277.050 279.450 286.950 ;
        RECT 283.950 286.800 286.050 288.900 ;
        RECT 283.950 280.950 286.050 283.050 ;
        RECT 271.950 274.950 274.050 277.050 ;
        RECT 277.950 274.950 280.050 277.050 ;
        RECT 268.950 271.950 271.050 274.050 ;
        RECT 272.400 271.050 273.450 274.950 ;
        RECT 271.950 268.950 274.050 271.050 ;
        RECT 260.400 264.000 264.450 264.450 ;
        RECT 259.950 263.400 264.450 264.000 ;
        RECT 257.400 250.050 258.450 262.950 ;
        RECT 259.950 259.950 262.050 263.400 ;
        RECT 265.950 260.100 268.050 262.200 ;
        RECT 274.950 260.100 277.050 262.200 ;
        RECT 266.400 259.350 267.600 260.100 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 265.950 256.950 268.050 259.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 259.950 253.950 262.050 256.050 ;
        RECT 263.400 255.900 264.600 256.650 ;
        RECT 253.800 247.950 255.900 250.050 ;
        RECT 256.950 247.950 259.050 250.050 ;
        RECT 257.400 244.050 258.450 247.950 ;
        RECT 256.950 241.950 259.050 244.050 ;
        RECT 260.400 235.050 261.450 253.950 ;
        RECT 262.950 253.800 265.050 255.900 ;
        RECT 269.400 254.400 270.600 256.650 ;
        RECT 269.400 247.050 270.450 254.400 ;
        RECT 271.950 247.950 274.050 250.050 ;
        RECT 268.950 244.950 271.050 247.050 ;
        RECT 262.950 241.950 265.050 244.050 ;
        RECT 259.950 232.950 262.050 235.050 ;
        RECT 250.950 223.950 253.050 226.050 ;
        RECT 256.950 223.950 259.050 226.050 ;
        RECT 247.950 220.950 250.050 223.050 ;
        RECT 251.400 216.600 252.450 223.950 ;
        RECT 257.400 216.600 258.450 223.950 ;
        RECT 263.400 217.050 264.450 241.950 ;
        RECT 269.400 229.050 270.450 244.950 ;
        RECT 268.950 226.950 271.050 229.050 ;
        RECT 265.950 220.950 268.050 226.050 ;
        RECT 269.400 222.450 270.450 226.950 ;
        RECT 272.400 226.050 273.450 247.950 ;
        RECT 271.950 223.950 274.050 226.050 ;
        RECT 269.400 221.400 273.450 222.450 ;
        RECT 265.950 217.800 268.050 219.900 ;
        RECT 251.400 214.350 252.600 216.600 ;
        RECT 257.400 214.350 258.600 216.600 ;
        RECT 262.950 214.950 265.050 217.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 256.950 211.950 259.050 214.050 ;
        RECT 259.950 211.950 262.050 214.050 ;
        RECT 254.400 210.900 255.600 211.650 ;
        RECT 245.400 209.400 249.450 210.450 ;
        RECT 229.950 202.950 232.050 205.050 ;
        RECT 229.950 196.950 232.050 199.050 ;
        RECT 230.400 184.050 231.450 196.950 ;
        RECT 232.950 193.950 235.050 196.050 ;
        RECT 193.950 172.950 196.050 175.050 ;
        RECT 187.950 166.950 190.050 169.050 ;
        RECT 194.400 157.050 195.450 172.950 ;
        RECT 197.400 172.050 198.450 176.400 ;
        RECT 199.800 172.950 201.900 175.050 ;
        RECT 202.950 172.950 205.050 177.000 ;
        RECT 206.400 176.400 210.450 177.450 ;
        RECT 196.950 169.950 199.050 172.050 ;
        RECT 200.400 163.050 201.450 172.950 ;
        RECT 199.950 160.950 202.050 163.050 ;
        RECT 193.950 154.950 196.050 157.050 ;
        RECT 199.950 154.950 202.050 157.050 ;
        RECT 184.950 151.950 187.050 154.050 ;
        RECT 163.950 121.950 166.050 124.050 ;
        RECT 154.950 118.950 157.050 121.050 ;
        RECT 142.950 103.950 145.050 106.050 ;
        RECT 148.950 104.100 151.050 106.200 ;
        RECT 155.400 105.600 156.450 118.950 ;
        RECT 160.950 115.950 163.050 118.050 ;
        RECT 149.400 103.350 150.600 104.100 ;
        RECT 155.400 103.350 156.600 105.600 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 154.950 100.950 157.050 103.050 ;
        RECT 146.400 98.400 147.600 100.650 ;
        RECT 152.400 99.900 153.600 100.650 ;
        RECT 161.400 99.900 162.450 115.950 ;
        RECT 173.400 112.050 174.450 131.400 ;
        RECT 181.950 130.950 184.050 133.050 ;
        RECT 185.400 129.450 186.450 151.950 ;
        RECT 187.950 145.950 190.050 148.050 ;
        RECT 196.950 145.950 199.050 148.050 ;
        RECT 188.400 138.600 189.450 145.950 ;
        RECT 197.400 138.600 198.450 145.950 ;
        RECT 188.400 136.350 189.600 138.600 ;
        RECT 197.400 136.350 198.600 138.600 ;
        RECT 188.100 133.950 190.200 136.050 ;
        RECT 191.400 133.950 193.500 136.050 ;
        RECT 196.800 133.950 198.900 136.050 ;
        RECT 191.400 132.900 192.600 133.650 ;
        RECT 190.950 130.800 193.050 132.900 ;
        RECT 200.400 130.050 201.450 154.950 ;
        RECT 202.950 148.950 205.050 151.050 ;
        RECT 203.400 142.050 204.450 148.950 ;
        RECT 202.950 139.950 205.050 142.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 185.400 128.400 189.450 129.450 ;
        RECT 163.950 109.950 166.050 112.050 ;
        RECT 172.950 109.950 175.050 112.050 ;
        RECT 178.950 109.950 181.050 112.050 ;
        RECT 139.950 94.950 142.050 97.050 ;
        RECT 146.400 91.050 147.450 98.400 ;
        RECT 151.950 97.800 154.050 99.900 ;
        RECT 160.950 97.800 163.050 99.900 ;
        RECT 145.950 88.950 148.050 91.050 ;
        RECT 164.400 85.050 165.450 109.950 ;
        RECT 172.950 104.100 175.050 106.200 ;
        RECT 179.400 105.600 180.450 109.950 ;
        RECT 173.400 103.350 174.600 104.100 ;
        RECT 179.400 103.350 180.600 105.600 ;
        RECT 184.950 104.100 187.050 106.200 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 175.950 100.950 178.050 103.050 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 170.400 98.400 171.600 100.650 ;
        RECT 176.400 99.900 177.600 100.650 ;
        RECT 170.400 88.050 171.450 98.400 ;
        RECT 175.950 97.800 178.050 99.900 ;
        RECT 185.400 94.050 186.450 104.100 ;
        RECT 188.400 99.450 189.450 128.400 ;
        RECT 199.950 127.950 202.050 130.050 ;
        RECT 199.950 121.950 202.050 124.050 ;
        RECT 200.400 115.050 201.450 121.950 ;
        RECT 203.400 121.050 204.450 133.950 ;
        RECT 202.950 118.950 205.050 121.050 ;
        RECT 202.950 115.800 205.050 117.900 ;
        RECT 206.400 117.450 207.450 176.400 ;
        RECT 208.950 145.950 211.050 148.050 ;
        RECT 209.400 138.450 210.450 145.950 ;
        RECT 212.400 142.050 213.450 181.950 ;
        RECT 221.400 181.350 222.600 183.600 ;
        RECT 227.400 181.350 228.600 183.600 ;
        RECT 229.950 181.950 232.050 184.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 218.400 176.400 219.600 178.650 ;
        RECT 224.400 177.900 225.600 178.650 ;
        RECT 218.400 169.050 219.450 176.400 ;
        RECT 223.950 175.800 226.050 177.900 ;
        RECT 233.400 175.050 234.450 193.950 ;
        RECT 241.950 183.000 244.050 187.050 ;
        RECT 248.400 183.600 249.450 209.400 ;
        RECT 253.950 208.800 256.050 210.900 ;
        RECT 260.400 209.400 261.600 211.650 ;
        RECT 256.950 205.950 259.050 208.050 ;
        RECT 253.950 184.950 256.050 187.050 ;
        RECT 242.400 181.350 243.600 183.000 ;
        RECT 248.400 181.350 249.600 183.600 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 244.950 178.950 247.050 181.050 ;
        RECT 247.950 178.950 250.050 181.050 ;
        RECT 239.400 177.900 240.600 178.650 ;
        RECT 238.950 175.800 241.050 177.900 ;
        RECT 245.400 176.400 246.600 178.650 ;
        RECT 232.950 172.950 235.050 175.050 ;
        RECT 217.950 166.950 220.050 169.050 ;
        RECT 223.950 166.950 226.050 169.050 ;
        RECT 220.950 163.050 223.050 166.050 ;
        RECT 217.950 162.000 223.050 163.050 ;
        RECT 217.950 161.400 222.450 162.000 ;
        RECT 217.950 160.950 222.000 161.400 ;
        RECT 224.400 151.050 225.450 166.950 ;
        RECT 232.950 160.950 235.050 163.050 ;
        RECT 223.950 148.950 226.050 151.050 ;
        RECT 229.950 142.950 232.050 145.050 ;
        RECT 211.950 139.950 214.050 142.050 ;
        RECT 212.400 138.450 213.600 138.600 ;
        RECT 209.400 137.400 213.600 138.450 ;
        RECT 212.400 136.350 213.600 137.400 ;
        RECT 217.950 137.100 220.050 139.200 ;
        RECT 218.400 136.350 219.600 137.100 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 215.400 131.400 216.600 133.650 ;
        RECT 221.400 132.900 222.600 133.650 ;
        RECT 211.950 127.950 214.050 130.050 ;
        RECT 208.950 118.950 211.050 124.050 ;
        RECT 206.400 116.400 210.450 117.450 ;
        RECT 199.950 112.950 202.050 115.050 ;
        RECT 196.950 104.100 199.050 106.200 ;
        RECT 203.400 105.600 204.450 115.800 ;
        RECT 197.400 103.350 198.600 104.100 ;
        RECT 203.400 103.350 204.600 105.600 ;
        RECT 209.400 103.050 210.450 116.400 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 190.950 99.450 193.050 100.050 ;
        RECT 188.400 98.400 193.050 99.450 ;
        RECT 190.950 94.950 193.050 98.400 ;
        RECT 194.400 98.400 195.600 100.650 ;
        RECT 200.400 99.000 201.600 100.650 ;
        RECT 194.400 94.050 195.450 98.400 ;
        RECT 196.950 94.950 199.050 97.050 ;
        RECT 199.950 94.950 202.050 99.000 ;
        RECT 175.950 91.950 178.050 94.050 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 193.950 91.950 196.050 94.050 ;
        RECT 169.950 85.950 172.050 88.050 ;
        RECT 163.950 82.950 166.050 85.050 ;
        RECT 145.950 76.950 148.050 79.050 ;
        RECT 169.950 76.950 172.050 79.050 ;
        RECT 139.950 70.950 142.050 73.050 ;
        RECT 140.400 61.050 141.450 70.950 ;
        RECT 139.950 58.950 142.050 61.050 ;
        RECT 146.400 60.600 147.450 76.950 ;
        RECT 154.950 64.950 157.050 70.050 ;
        RECT 160.950 67.950 166.050 70.050 ;
        RECT 146.400 58.350 147.600 60.600 ;
        RECT 151.950 60.000 154.050 64.050 ;
        RECT 160.950 61.950 163.050 66.900 ;
        RECT 152.400 58.350 153.600 60.000 ;
        RECT 160.950 58.800 163.050 60.900 ;
        RECT 170.400 60.600 171.450 76.950 ;
        RECT 176.400 73.050 177.450 91.950 ;
        RECT 197.400 88.050 198.450 94.950 ;
        RECT 202.950 88.950 205.050 91.050 ;
        RECT 196.950 85.950 199.050 88.050 ;
        RECT 178.950 73.950 181.050 76.050 ;
        RECT 175.950 70.950 178.050 73.050 ;
        RECT 179.400 67.050 180.450 73.950 ;
        RECT 178.950 64.950 181.050 67.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 143.400 53.400 144.600 55.650 ;
        RECT 149.400 54.900 150.600 55.650 ;
        RECT 161.400 54.900 162.450 58.800 ;
        RECT 170.400 58.350 171.600 60.600 ;
        RECT 175.950 59.100 178.050 61.200 ;
        RECT 179.400 61.050 180.450 64.950 ;
        RECT 176.400 58.350 177.600 59.100 ;
        RECT 178.950 58.950 181.050 61.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 181.950 57.450 184.050 61.050 ;
        RECT 190.950 59.100 193.050 61.200 ;
        RECT 196.950 59.100 199.050 61.200 ;
        RECT 203.400 61.050 204.450 88.950 ;
        RECT 209.400 69.450 210.450 100.950 ;
        RECT 212.400 100.050 213.450 127.950 ;
        RECT 215.400 112.050 216.450 131.400 ;
        RECT 220.950 130.800 223.050 132.900 ;
        RECT 223.950 124.950 226.050 127.050 ;
        RECT 214.950 109.950 217.050 112.050 ;
        RECT 217.950 105.000 220.050 109.050 ;
        RECT 224.400 105.600 225.450 124.950 ;
        RECT 227.400 115.050 228.450 133.950 ;
        RECT 230.400 124.050 231.450 142.950 ;
        RECT 233.400 139.050 234.450 160.950 ;
        RECT 245.400 151.050 246.450 176.400 ;
        RECT 247.950 172.950 250.050 175.050 ;
        RECT 244.950 148.950 247.050 151.050 ;
        RECT 244.950 144.450 247.050 145.050 ;
        RECT 248.400 144.450 249.450 172.950 ;
        RECT 254.400 163.050 255.450 184.950 ;
        RECT 257.400 184.050 258.450 205.950 ;
        RECT 260.400 187.050 261.450 209.400 ;
        RECT 266.400 205.050 267.450 217.800 ;
        RECT 268.950 214.950 271.050 220.050 ;
        RECT 272.400 216.600 273.450 221.400 ;
        RECT 275.400 220.050 276.450 260.100 ;
        RECT 278.400 244.050 279.450 274.950 ;
        RECT 280.950 268.950 283.050 271.050 ;
        RECT 281.400 250.050 282.450 268.950 ;
        RECT 284.400 268.050 285.450 280.950 ;
        RECT 293.400 280.050 294.450 298.950 ;
        RECT 296.400 283.050 297.450 301.950 ;
        RECT 295.950 280.950 298.050 283.050 ;
        RECT 292.950 277.950 295.050 280.050 ;
        RECT 299.400 271.050 300.450 322.800 ;
        RECT 302.400 319.050 303.450 328.950 ;
        RECT 301.950 316.950 304.050 319.050 ;
        RECT 301.950 295.950 304.050 298.050 ;
        RECT 302.400 288.900 303.450 295.950 ;
        RECT 308.400 295.200 309.450 328.950 ;
        RECT 310.950 297.450 315.000 298.050 ;
        RECT 310.950 295.950 315.450 297.450 ;
        RECT 307.950 293.100 310.050 295.200 ;
        RECT 314.400 294.600 315.450 295.950 ;
        RECT 320.400 295.050 321.450 332.400 ;
        RECT 328.950 328.950 331.050 333.000 ;
        RECT 335.400 331.050 336.450 361.950 ;
        RECT 347.400 343.200 348.450 403.950 ;
        RECT 350.400 397.050 351.450 416.100 ;
        RECT 356.400 415.350 357.600 416.100 ;
        RECT 362.400 415.350 363.600 417.600 ;
        RECT 367.950 415.950 370.050 418.050 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 358.950 412.950 361.050 415.050 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 352.950 409.950 355.050 412.050 ;
        RECT 359.400 410.400 360.600 412.650 ;
        RECT 349.950 394.950 352.050 397.050 ;
        RECT 353.400 391.050 354.450 409.950 ;
        RECT 359.400 406.050 360.450 410.400 ;
        RECT 367.950 409.950 370.050 412.050 ;
        RECT 358.950 403.950 361.050 406.050 ;
        RECT 358.950 394.950 361.050 397.050 ;
        RECT 352.950 388.950 355.050 391.050 ;
        RECT 359.400 388.050 360.450 394.950 ;
        RECT 358.950 385.950 361.050 388.050 ;
        RECT 364.950 379.950 367.050 382.050 ;
        RECT 365.400 373.200 366.450 379.950 ;
        RECT 356.400 372.450 357.600 372.600 ;
        RECT 353.400 371.400 357.600 372.450 ;
        RECT 353.400 352.050 354.450 371.400 ;
        RECT 356.400 370.350 357.600 371.400 ;
        RECT 364.950 371.100 367.050 373.200 ;
        RECT 365.400 370.350 366.600 371.100 ;
        RECT 356.100 367.950 358.200 370.050 ;
        RECT 359.400 367.950 361.500 370.050 ;
        RECT 364.800 367.950 366.900 370.050 ;
        RECT 359.400 365.400 360.600 367.650 ;
        RECT 355.950 361.950 358.050 364.050 ;
        RECT 352.950 349.950 355.050 352.050 ;
        RECT 352.950 343.950 355.050 346.050 ;
        RECT 337.950 340.950 340.050 343.050 ;
        RECT 346.950 341.100 349.050 343.200 ;
        RECT 338.400 333.900 339.450 340.950 ;
        RECT 346.950 337.950 349.050 340.050 ;
        RECT 353.400 339.600 354.450 343.950 ;
        RECT 356.400 340.050 357.450 361.950 ;
        RECT 347.400 337.350 348.600 337.950 ;
        RECT 353.400 337.350 354.600 339.600 ;
        RECT 355.950 337.950 358.050 340.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 344.400 333.900 345.600 334.650 ;
        RECT 337.950 331.800 340.050 333.900 ;
        RECT 343.950 331.800 346.050 333.900 ;
        RECT 350.400 332.400 351.600 334.650 ;
        RECT 334.950 328.950 337.050 331.050 ;
        RECT 340.950 328.950 343.050 331.050 ;
        RECT 325.950 313.950 328.050 316.050 ;
        RECT 322.950 295.950 325.050 298.050 ;
        RECT 308.400 292.350 309.600 293.100 ;
        RECT 314.400 292.350 315.600 294.600 ;
        RECT 319.950 292.950 322.050 295.050 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 311.400 288.900 312.600 289.650 ;
        RECT 301.950 286.800 304.050 288.900 ;
        RECT 310.950 286.800 313.050 288.900 ;
        RECT 317.400 288.000 318.600 289.650 ;
        RECT 298.950 268.950 301.050 271.050 ;
        RECT 283.950 265.950 286.050 268.050 ;
        RECT 295.950 265.950 298.050 268.050 ;
        RECT 286.950 260.100 289.050 262.200 ;
        RECT 287.400 259.350 288.600 260.100 ;
        RECT 284.100 256.950 286.200 259.050 ;
        RECT 287.400 256.950 289.500 259.050 ;
        RECT 292.800 256.950 294.900 259.050 ;
        RECT 284.400 254.400 285.600 256.650 ;
        RECT 293.400 254.400 294.600 256.650 ;
        RECT 296.400 256.050 297.450 265.950 ;
        RECT 280.950 247.950 283.050 250.050 ;
        RECT 284.400 247.050 285.450 254.400 ;
        RECT 286.950 250.950 289.050 253.050 ;
        RECT 283.950 244.950 286.050 247.050 ;
        RECT 277.950 241.950 280.050 244.050 ;
        RECT 287.400 243.450 288.450 250.950 ;
        RECT 284.400 242.400 288.450 243.450 ;
        RECT 274.950 217.950 277.050 220.050 ;
        RECT 272.400 214.350 273.600 216.600 ;
        RECT 277.950 216.000 280.050 220.050 ;
        RECT 278.400 214.350 279.600 216.000 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 275.400 210.900 276.600 211.650 ;
        RECT 274.950 208.800 277.050 210.900 ;
        RECT 265.950 202.950 268.050 205.050 ;
        RECT 274.950 202.950 277.050 205.050 ;
        RECT 268.950 193.950 271.050 196.050 ;
        RECT 259.950 184.950 262.050 187.050 ;
        RECT 269.400 184.200 270.450 193.950 ;
        RECT 256.950 181.950 259.050 184.050 ;
        RECT 262.950 182.100 265.050 184.200 ;
        RECT 268.950 182.100 271.050 184.200 ;
        RECT 263.400 181.350 264.600 182.100 ;
        RECT 269.400 181.350 270.600 182.100 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 256.800 175.950 258.900 178.050 ;
        RECT 260.400 177.900 261.600 178.650 ;
        RECT 253.950 160.950 256.050 163.050 ;
        RECT 253.950 154.950 256.050 157.050 ;
        RECT 244.950 143.400 249.450 144.450 ;
        RECT 244.950 142.950 247.050 143.400 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 238.950 137.100 241.050 139.200 ;
        RECT 245.400 138.600 246.450 142.950 ;
        RECT 239.400 136.350 240.600 137.100 ;
        RECT 245.400 136.350 246.600 138.600 ;
        RECT 247.950 136.950 250.050 141.900 ;
        RECT 250.950 139.950 253.050 142.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 236.400 131.400 237.600 133.650 ;
        RECT 242.400 132.900 243.600 133.650 ;
        RECT 251.400 132.900 252.450 139.950 ;
        RECT 254.400 138.450 255.450 154.950 ;
        RECT 257.400 142.050 258.450 175.950 ;
        RECT 259.950 175.800 262.050 177.900 ;
        RECT 266.400 177.000 267.600 178.650 ;
        RECT 260.400 160.050 261.450 175.800 ;
        RECT 265.950 172.950 268.050 177.000 ;
        RECT 271.950 175.950 274.050 178.050 ;
        RECT 259.950 157.950 262.050 160.050 ;
        RECT 268.950 148.950 271.050 151.050 ;
        RECT 256.950 139.950 259.050 142.050 ;
        RECT 257.400 138.450 258.600 138.600 ;
        RECT 254.400 137.400 258.600 138.450 ;
        RECT 262.950 138.000 265.050 142.050 ;
        RECT 269.400 138.450 270.450 148.950 ;
        RECT 272.400 142.050 273.450 175.950 ;
        RECT 275.400 175.050 276.450 202.950 ;
        RECT 284.400 202.050 285.450 242.400 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 283.950 199.950 286.050 202.050 ;
        RECT 287.400 190.050 288.450 235.950 ;
        RECT 293.400 235.050 294.450 254.400 ;
        RECT 295.950 253.950 298.050 256.050 ;
        RECT 299.400 244.050 300.450 268.950 ;
        RECT 302.400 253.050 303.450 286.800 ;
        RECT 316.950 283.950 319.050 288.000 ;
        RECT 319.950 286.950 322.050 289.050 ;
        RECT 307.950 274.950 310.050 277.050 ;
        RECT 308.400 261.600 309.450 274.950 ;
        RECT 308.400 259.350 309.600 261.600 ;
        RECT 320.400 261.450 321.450 286.950 ;
        RECT 317.400 260.400 321.450 261.450 ;
        RECT 323.400 261.600 324.450 295.950 ;
        RECT 326.400 286.050 327.450 313.950 ;
        RECT 328.950 301.950 331.050 304.050 ;
        RECT 329.400 295.050 330.450 301.950 ;
        RECT 328.950 292.950 331.050 295.050 ;
        RECT 334.950 294.000 337.050 298.050 ;
        RECT 341.400 295.200 342.450 328.950 ;
        RECT 350.400 310.050 351.450 332.400 ;
        RECT 359.400 319.050 360.450 365.400 ;
        RECT 368.400 358.050 369.450 409.950 ;
        RECT 374.400 403.050 375.450 463.950 ;
        RECT 377.400 433.050 378.450 484.650 ;
        RECT 379.950 457.950 382.050 460.050 ;
        RECT 380.400 451.050 381.450 457.950 ;
        RECT 383.400 457.050 384.450 505.950 ;
        RECT 386.400 505.050 387.450 511.950 ;
        RECT 392.400 508.050 393.450 523.950 ;
        RECT 400.950 520.800 403.050 522.900 ;
        RECT 401.400 511.050 402.450 520.800 ;
        RECT 404.400 517.050 405.450 547.950 ;
        RECT 409.950 541.950 415.050 544.050 ;
        RECT 409.950 535.950 412.050 538.050 ;
        RECT 406.950 529.950 409.050 532.050 ;
        RECT 403.950 514.950 406.050 517.050 ;
        RECT 400.950 508.950 403.050 511.050 ;
        RECT 391.950 505.950 394.050 508.050 ;
        RECT 385.950 502.950 388.050 505.050 ;
        RECT 403.950 502.950 406.050 505.050 ;
        RECT 385.950 493.950 388.050 496.050 ;
        RECT 394.950 494.100 397.050 496.200 ;
        RECT 386.400 489.900 387.450 493.950 ;
        RECT 395.400 493.350 396.600 494.100 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 385.950 487.800 388.050 489.900 ;
        RECT 392.400 489.000 393.600 490.650 ;
        RECT 398.400 489.900 399.600 490.650 ;
        RECT 391.950 484.950 394.050 489.000 ;
        RECT 397.950 487.800 400.050 489.900 ;
        RECT 398.400 487.050 399.450 487.800 ;
        RECT 394.950 485.400 399.450 487.050 ;
        RECT 394.950 484.950 399.000 485.400 ;
        RECT 392.400 481.050 393.450 484.950 ;
        RECT 391.950 478.950 394.050 481.050 ;
        RECT 385.950 460.950 388.050 463.050 ;
        RECT 386.400 457.050 387.450 460.950 ;
        RECT 382.800 454.950 384.900 457.050 ;
        RECT 385.950 454.950 388.050 457.050 ;
        RECT 379.950 448.950 382.050 451.050 ;
        RECT 386.400 450.600 387.450 454.950 ;
        RECT 404.400 451.200 405.450 502.950 ;
        RECT 407.400 484.050 408.450 529.950 ;
        RECT 410.400 529.050 411.450 535.950 ;
        RECT 412.950 530.100 415.050 535.050 ;
        RECT 416.400 532.050 417.450 553.950 ;
        RECT 418.950 541.950 421.050 544.050 ;
        RECT 419.400 532.050 420.450 541.950 ;
        RECT 425.400 541.050 426.450 556.950 ;
        RECT 431.400 556.050 432.450 565.950 ;
        RECT 430.950 553.950 433.050 556.050 ;
        RECT 437.400 553.050 438.450 566.400 ;
        RECT 436.950 550.950 439.050 553.050 ;
        RECT 443.400 550.050 444.450 566.400 ;
        RECT 449.400 556.050 450.450 610.950 ;
        RECT 455.400 610.050 456.450 619.950 ;
        RECT 454.950 607.950 457.050 610.050 ;
        RECT 452.100 604.950 454.200 607.050 ;
        RECT 452.400 603.900 453.600 604.650 ;
        RECT 451.950 601.800 454.050 603.900 ;
        RECT 454.950 598.950 457.050 601.050 ;
        RECT 455.400 592.050 456.450 598.950 ;
        RECT 454.950 589.950 457.050 592.050 ;
        RECT 458.400 589.050 459.450 634.950 ;
        RECT 473.400 622.050 474.450 658.950 ;
        RECT 479.400 655.050 480.450 706.950 ;
        RECT 485.400 702.450 486.450 718.950 ;
        RECT 488.400 706.050 489.450 721.800 ;
        RECT 506.400 720.450 507.450 721.800 ;
        RECT 503.400 719.400 507.450 720.450 ;
        RECT 496.800 709.950 498.900 712.050 ;
        RECT 487.950 703.950 490.050 706.050 ;
        RECT 485.400 701.400 489.450 702.450 ;
        RECT 484.800 682.950 486.900 685.050 ;
        RECT 485.400 680.400 486.600 682.650 ;
        RECT 485.400 676.050 486.450 680.400 ;
        RECT 484.950 673.950 487.050 676.050 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 478.950 652.950 481.050 655.050 ;
        RECT 481.950 650.100 484.050 652.200 ;
        RECT 482.400 649.350 483.600 650.100 ;
        RECT 476.100 646.950 478.200 649.050 ;
        RECT 481.500 646.950 483.600 649.050 ;
        RECT 476.400 645.900 477.600 646.650 ;
        RECT 485.400 646.050 486.450 667.950 ;
        RECT 475.950 643.800 478.050 645.900 ;
        RECT 484.950 643.950 487.050 646.050 ;
        RECT 488.400 643.050 489.450 701.400 ;
        RECT 493.800 682.950 495.900 685.050 ;
        RECT 494.400 681.450 495.600 682.650 ;
        RECT 497.400 681.450 498.450 709.950 ;
        RECT 499.950 682.950 502.050 685.050 ;
        RECT 494.400 680.400 498.450 681.450 ;
        RECT 500.400 661.050 501.450 682.950 ;
        RECT 503.400 670.050 504.450 719.400 ;
        RECT 509.400 679.050 510.450 722.400 ;
        RECT 514.950 721.800 517.050 723.900 ;
        RECT 520.950 721.800 523.050 723.900 ;
        RECT 526.950 721.800 529.050 723.900 ;
        RECT 529.950 712.950 532.050 715.050 ;
        RECT 530.400 703.050 531.450 712.950 ;
        RECT 536.400 712.050 537.450 727.800 ;
        RECT 539.400 723.900 540.450 739.950 ;
        RECT 542.400 730.050 543.450 784.800 ;
        RECT 548.400 784.050 549.450 793.950 ;
        RECT 547.950 781.950 550.050 784.050 ;
        RECT 545.700 774.300 547.800 776.400 ;
        RECT 546.300 769.500 547.800 774.300 ;
        RECT 545.700 767.400 547.800 769.500 ;
        RECT 546.300 749.700 547.800 767.400 ;
        RECT 545.700 747.600 547.800 749.700 ;
        RECT 548.700 771.300 550.800 776.400 ;
        RECT 551.700 774.300 553.800 776.400 ;
        RECT 570.600 774.300 572.700 776.400 ;
        RECT 573.600 774.300 576.600 776.400 ;
        RECT 548.700 749.700 549.900 771.300 ;
        RECT 551.700 769.500 553.200 774.300 ;
        RECT 554.100 771.300 556.200 773.400 ;
        RECT 551.100 767.400 553.200 769.500 ;
        RECT 551.700 749.700 553.200 767.400 ;
        RECT 554.700 764.100 555.900 771.300 ;
        RECT 559.500 769.800 561.600 771.900 ;
        RECT 568.200 771.300 570.300 773.400 ;
        RECT 554.100 762.000 556.200 764.100 ;
        RECT 560.700 763.200 561.600 769.800 ;
        RECT 554.700 749.700 555.900 762.000 ;
        RECT 559.500 761.100 561.600 763.200 ;
        RECT 556.800 754.500 558.900 756.600 ;
        RECT 560.700 750.600 561.600 761.100 ;
        RECT 562.950 758.100 565.050 760.200 ;
        RECT 563.400 757.350 564.600 758.100 ;
        RECT 563.100 754.950 565.200 757.050 ;
        RECT 548.700 747.600 550.800 749.700 ;
        RECT 551.700 747.600 553.800 749.700 ;
        RECT 554.700 747.600 556.800 749.700 ;
        RECT 560.100 748.500 562.200 750.600 ;
        RECT 569.100 749.700 570.300 771.300 ;
        RECT 571.500 768.300 572.700 774.300 ;
        RECT 571.500 766.200 573.600 768.300 ;
        RECT 571.500 749.700 572.700 766.200 ;
        RECT 575.100 755.400 576.600 774.300 ;
        RECT 574.500 753.300 576.600 755.400 ;
        RECT 574.500 749.700 575.700 753.300 ;
        RECT 568.200 747.600 570.300 749.700 ;
        RECT 571.200 747.600 573.300 749.700 ;
        RECT 574.200 747.600 576.300 749.700 ;
        RECT 578.400 748.050 579.450 796.800 ;
        RECT 581.400 793.050 582.450 833.400 ;
        RECT 586.950 829.950 589.050 834.000 ;
        RECT 604.950 829.950 607.050 834.000 ;
        RECT 611.400 826.050 612.450 838.950 ;
        RECT 620.400 838.350 621.600 839.100 ;
        RECT 628.800 838.950 630.900 841.050 ;
        RECT 634.800 838.950 636.900 841.050 ;
        RECT 637.950 838.950 640.050 841.050 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 617.400 835.050 618.600 835.650 ;
        RECT 613.950 833.400 618.600 835.050 ;
        RECT 623.400 834.000 624.600 835.650 ;
        RECT 613.950 832.950 618.000 833.400 ;
        RECT 622.950 829.950 625.050 834.000 ;
        RECT 610.950 823.950 613.050 826.050 ;
        RECT 628.950 820.950 631.050 823.050 ;
        RECT 613.950 811.950 616.050 814.050 ;
        RECT 583.950 806.100 586.050 811.050 ;
        RECT 614.400 808.200 615.450 811.950 ;
        RECT 584.400 805.350 585.600 806.100 ;
        RECT 592.950 805.950 595.050 808.050 ;
        RECT 607.950 806.100 610.050 808.200 ;
        RECT 613.950 806.100 616.050 808.200 ;
        RECT 629.400 807.600 630.450 820.950 ;
        RECT 623.400 807.450 624.600 807.600 ;
        RECT 617.400 806.400 624.600 807.450 ;
        RECT 584.400 802.950 586.500 805.050 ;
        RECT 589.800 802.950 591.900 805.050 ;
        RECT 590.400 801.900 591.600 802.650 ;
        RECT 589.950 799.800 592.050 801.900 ;
        RECT 580.950 790.950 583.050 793.050 ;
        RECT 580.950 784.950 583.050 787.050 ;
        RECT 581.400 778.050 582.450 784.950 ;
        RECT 583.950 778.950 586.050 781.050 ;
        RECT 580.950 775.950 583.050 778.050 ;
        RECT 584.400 775.050 585.450 778.950 ;
        RECT 583.950 772.950 586.050 775.050 ;
        RECT 587.400 765.450 588.600 765.600 ;
        RECT 590.400 765.450 591.450 799.800 ;
        RECT 587.400 764.400 591.450 765.450 ;
        RECT 587.400 763.350 588.600 764.400 ;
        RECT 581.100 760.950 583.200 763.050 ;
        RECT 587.100 760.950 589.200 763.050 ;
        RECT 577.950 745.950 580.050 748.050 ;
        RECT 574.950 742.950 577.050 745.050 ;
        RECT 556.950 741.450 559.050 742.050 ;
        RECT 551.400 740.400 559.050 741.450 ;
        RECT 551.400 736.050 552.450 740.400 ;
        RECT 556.950 739.950 559.050 740.400 ;
        RECT 553.950 736.950 556.050 739.050 ;
        RECT 550.950 733.950 553.050 736.050 ;
        RECT 554.400 733.050 555.450 736.950 ;
        RECT 553.950 730.950 556.050 733.050 ;
        RECT 541.950 727.950 544.050 730.050 ;
        RECT 547.950 728.100 550.050 730.200 ;
        RECT 554.400 729.600 555.450 730.950 ;
        RECT 548.400 727.350 549.600 728.100 ;
        RECT 554.400 727.350 555.600 729.600 ;
        RECT 559.950 727.950 562.050 730.050 ;
        RECT 565.950 728.100 568.050 730.200 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 538.950 721.800 541.050 723.900 ;
        RECT 541.950 721.950 544.050 724.050 ;
        RECT 545.400 723.900 546.600 724.650 ;
        RECT 551.400 723.900 552.600 724.650 ;
        RECT 542.400 715.050 543.450 721.950 ;
        RECT 544.950 721.800 547.050 723.900 ;
        RECT 550.950 721.800 553.050 723.900 ;
        RECT 560.400 715.050 561.450 727.950 ;
        RECT 566.400 727.350 567.600 728.100 ;
        RECT 566.400 724.950 568.500 727.050 ;
        RECT 571.800 724.950 573.900 727.050 ;
        RECT 575.400 726.450 576.450 742.950 ;
        RECT 578.400 730.200 579.450 745.950 ;
        RECT 593.400 738.450 594.450 805.950 ;
        RECT 608.400 805.350 609.600 806.100 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 602.100 802.950 604.200 805.050 ;
        RECT 607.500 802.950 609.600 805.050 ;
        RECT 596.400 790.050 597.450 802.950 ;
        RECT 602.400 800.400 603.600 802.650 ;
        RECT 595.950 787.950 598.050 790.050 ;
        RECT 602.400 778.050 603.450 800.400 ;
        RECT 610.950 793.950 613.050 796.050 ;
        RECT 601.950 775.950 604.050 778.050 ;
        RECT 595.950 766.950 598.050 769.050 ;
        RECT 604.950 766.950 607.050 769.050 ;
        RECT 596.400 748.050 597.450 766.950 ;
        RECT 605.400 762.600 606.450 766.950 ;
        RECT 607.950 763.950 610.050 769.050 ;
        RECT 605.400 760.350 606.600 762.600 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 602.400 756.450 603.600 757.650 ;
        RECT 599.400 755.400 603.600 756.450 ;
        RECT 595.950 745.950 598.050 748.050 ;
        RECT 599.400 745.050 600.450 755.400 ;
        RECT 601.950 751.950 604.050 754.050 ;
        RECT 607.950 753.450 610.050 757.050 ;
        RECT 605.400 753.000 610.050 753.450 ;
        RECT 605.400 752.400 609.450 753.000 ;
        RECT 598.950 742.950 601.050 745.050 ;
        RECT 593.400 737.400 597.450 738.450 ;
        RECT 577.950 728.100 580.050 730.200 ;
        RECT 592.950 729.000 595.050 733.050 ;
        RECT 596.400 730.200 597.450 737.400 ;
        RECT 593.400 727.350 594.600 729.000 ;
        RECT 595.950 728.100 598.050 730.200 ;
        RECT 575.400 725.400 579.450 726.450 ;
        RECT 562.950 721.950 565.050 724.050 ;
        RECT 572.400 723.900 573.600 724.650 ;
        RECT 541.950 712.950 544.050 715.050 ;
        RECT 559.950 712.950 562.050 715.050 ;
        RECT 535.950 709.950 538.050 712.050 ;
        RECT 523.950 700.950 526.050 703.050 ;
        RECT 529.950 700.950 532.050 703.050 ;
        RECT 514.950 683.100 517.050 685.200 ;
        RECT 515.400 682.350 516.600 683.100 ;
        RECT 515.100 679.950 517.200 682.050 ;
        RECT 508.950 676.950 511.050 679.050 ;
        RECT 509.400 673.050 510.450 676.950 ;
        RECT 511.950 673.950 514.050 676.050 ;
        RECT 508.950 670.950 511.050 673.050 ;
        RECT 502.950 667.950 505.050 670.050 ;
        RECT 508.950 661.950 511.050 664.050 ;
        RECT 499.950 658.950 502.050 661.050 ;
        RECT 505.950 655.950 508.050 658.050 ;
        RECT 490.950 652.950 493.050 655.050 ;
        RECT 478.950 640.950 481.050 643.050 ;
        RECT 487.950 640.950 490.050 643.050 ;
        RECT 461.700 618.300 463.800 620.400 ;
        RECT 462.300 613.500 463.800 618.300 ;
        RECT 461.700 611.400 463.800 613.500 ;
        RECT 462.300 593.700 463.800 611.400 ;
        RECT 461.700 591.600 463.800 593.700 ;
        RECT 464.700 615.300 466.800 620.400 ;
        RECT 467.700 618.300 469.800 620.400 ;
        RECT 472.950 619.950 475.050 622.050 ;
        RECT 464.700 593.700 465.900 615.300 ;
        RECT 467.700 613.500 469.200 618.300 ;
        RECT 470.100 615.300 472.200 617.400 ;
        RECT 467.100 611.400 469.200 613.500 ;
        RECT 467.700 593.700 469.200 611.400 ;
        RECT 470.700 608.100 471.900 615.300 ;
        RECT 475.500 613.800 477.600 615.900 ;
        RECT 470.100 606.000 472.200 608.100 ;
        RECT 476.700 607.200 477.600 613.800 ;
        RECT 479.400 612.450 480.450 640.950 ;
        RECT 491.400 640.050 492.450 652.950 ;
        RECT 499.950 651.000 502.050 655.050 ;
        RECT 506.400 652.050 507.450 655.950 ;
        RECT 500.400 649.350 501.600 651.000 ;
        RECT 505.950 649.950 508.050 652.050 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 493.950 643.950 496.050 646.050 ;
        RECT 497.400 645.900 498.600 646.650 ;
        RECT 490.950 637.950 493.050 640.050 ;
        RECT 494.400 634.050 495.450 643.950 ;
        RECT 496.950 643.800 499.050 645.900 ;
        RECT 503.400 644.400 504.600 646.650 ;
        RECT 493.950 631.950 496.050 634.050 ;
        RECT 503.400 625.050 504.450 644.400 ;
        RECT 502.950 622.950 505.050 625.050 ;
        RECT 486.600 618.300 488.700 620.400 ;
        RECT 489.600 618.300 492.600 620.400 ;
        RECT 484.200 615.300 486.300 617.400 ;
        RECT 479.400 611.400 483.450 612.450 ;
        RECT 470.700 593.700 471.900 606.000 ;
        RECT 475.500 605.100 477.600 607.200 ;
        RECT 472.800 598.500 474.900 600.600 ;
        RECT 476.700 594.600 477.600 605.100 ;
        RECT 478.800 602.100 480.900 604.200 ;
        RECT 482.400 604.050 483.450 611.400 ;
        RECT 479.400 601.350 480.600 602.100 ;
        RECT 481.950 601.950 484.050 604.050 ;
        RECT 479.100 598.950 481.200 601.050 ;
        RECT 464.700 591.600 466.800 593.700 ;
        RECT 467.700 591.600 469.800 593.700 ;
        RECT 470.700 591.600 472.800 593.700 ;
        RECT 476.100 592.500 478.200 594.600 ;
        RECT 485.100 593.700 486.300 615.300 ;
        RECT 487.500 612.300 488.700 618.300 ;
        RECT 487.500 610.200 489.600 612.300 ;
        RECT 487.500 593.700 488.700 610.200 ;
        RECT 491.100 599.400 492.600 618.300 ;
        RECT 509.400 610.200 510.450 661.950 ;
        RECT 512.400 652.050 513.450 673.950 ;
        RECT 517.950 658.950 520.050 661.050 ;
        RECT 511.950 649.950 514.050 652.050 ;
        RECT 518.400 651.600 519.450 658.950 ;
        RECT 524.400 652.200 525.450 700.950 ;
        RECT 538.950 682.950 541.050 685.050 ;
        RECT 553.950 683.100 556.050 685.200 ;
        RECT 533.100 679.950 535.200 682.050 ;
        RECT 539.400 676.050 540.450 682.950 ;
        RECT 554.400 682.350 555.600 683.100 ;
        RECT 554.100 679.950 556.200 682.050 ;
        RECT 538.950 673.950 541.050 676.050 ;
        RECT 535.950 658.950 538.050 661.050 ;
        RECT 529.950 655.950 532.050 658.050 ;
        RECT 518.400 649.350 519.600 651.600 ;
        RECT 523.950 650.100 526.050 652.200 ;
        RECT 524.400 649.350 525.600 650.100 ;
        RECT 530.400 649.200 531.450 655.950 ;
        RECT 514.950 646.950 517.050 649.050 ;
        RECT 517.950 646.950 520.050 649.050 ;
        RECT 520.950 646.950 523.050 649.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 529.950 647.100 532.050 649.200 ;
        RECT 511.950 643.950 514.050 646.050 ;
        RECT 515.400 644.400 516.600 646.650 ;
        RECT 521.400 644.400 522.600 646.650 ;
        RECT 530.400 646.350 531.600 647.100 ;
        RECT 512.400 613.050 513.450 643.950 ;
        RECT 515.400 640.050 516.450 644.400 ;
        RECT 517.950 640.950 520.050 643.050 ;
        RECT 514.950 637.950 517.050 640.050 ;
        RECT 511.950 610.950 514.050 613.050 ;
        RECT 502.950 608.100 505.050 610.200 ;
        RECT 508.950 608.100 511.050 610.200 ;
        RECT 503.400 607.350 504.600 608.100 ;
        RECT 497.100 604.950 499.200 607.050 ;
        RECT 503.100 604.950 505.200 607.050 ;
        RECT 512.100 604.950 514.200 607.050 ;
        RECT 490.500 597.300 492.600 599.400 ;
        RECT 512.400 602.400 513.600 604.650 ;
        RECT 490.500 593.700 491.700 597.300 ;
        RECT 484.200 591.600 486.300 593.700 ;
        RECT 487.200 591.600 489.300 593.700 ;
        RECT 490.200 591.600 492.300 593.700 ;
        RECT 457.950 586.950 460.050 589.050 ;
        RECT 466.950 586.950 469.050 589.050 ;
        RECT 454.950 580.950 457.050 583.050 ;
        RECT 463.950 580.950 466.050 583.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 452.400 559.050 453.450 568.950 ;
        RECT 451.950 556.950 454.050 559.050 ;
        RECT 448.950 553.950 451.050 556.050 ;
        RECT 442.950 547.950 445.050 550.050 ;
        RECT 430.950 544.950 433.050 547.050 ;
        RECT 424.950 538.950 427.050 541.050 ;
        RECT 415.800 529.950 417.900 532.050 ;
        RECT 409.950 526.950 412.050 529.050 ;
        RECT 412.950 526.950 415.050 529.050 ;
        RECT 418.950 528.000 421.050 532.050 ;
        RECT 425.400 531.600 426.450 538.950 ;
        RECT 431.400 535.050 432.450 544.950 ;
        RECT 433.950 541.950 436.050 544.050 ;
        RECT 430.950 532.950 433.050 535.050 ;
        RECT 425.400 529.350 426.600 531.600 ;
        RECT 434.400 529.050 435.450 541.950 ;
        RECT 437.400 540.300 440.400 542.400 ;
        RECT 441.300 540.300 443.400 542.400 ;
        RECT 452.400 541.050 453.450 556.950 ;
        RECT 455.400 544.050 456.450 580.950 ;
        RECT 464.400 573.600 465.450 580.950 ;
        RECT 464.400 571.350 465.600 573.600 ;
        RECT 467.400 571.050 468.450 586.950 ;
        RECT 512.400 586.050 513.450 602.400 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 511.950 583.950 514.050 586.050 ;
        RECT 482.700 579.300 484.800 581.400 ;
        RECT 485.700 579.300 487.800 581.400 ;
        RECT 488.700 579.300 490.800 581.400 ;
        RECT 472.950 574.950 475.050 577.050 ;
        RECT 483.300 575.700 484.500 579.300 ;
        RECT 458.100 568.950 460.200 571.050 ;
        RECT 463.500 568.950 465.600 571.050 ;
        RECT 466.950 568.950 469.050 571.050 ;
        RECT 473.400 570.900 474.450 574.950 ;
        RECT 478.950 571.950 481.050 574.050 ;
        RECT 482.400 573.600 484.500 575.700 ;
        RECT 472.950 568.800 475.050 570.900 ;
        RECT 458.400 567.900 459.600 568.650 ;
        RECT 457.950 565.800 460.050 567.900 ;
        RECT 469.800 565.950 471.900 568.050 ;
        RECT 475.800 565.950 477.900 568.050 ;
        RECT 470.400 564.450 471.600 565.650 ;
        RECT 467.400 563.400 471.600 564.450 ;
        RECT 467.400 559.050 468.450 563.400 ;
        RECT 469.950 559.950 472.050 562.050 ;
        RECT 475.950 559.950 478.050 562.050 ;
        RECT 466.950 556.950 469.050 559.050 ;
        RECT 467.400 553.050 468.450 556.950 ;
        RECT 466.950 550.950 469.050 553.050 ;
        RECT 454.950 541.950 457.050 544.050 ;
        RECT 413.400 526.350 414.600 526.950 ;
        RECT 419.400 526.350 420.600 528.000 ;
        RECT 424.800 526.950 426.900 529.050 ;
        RECT 430.800 526.950 432.900 529.050 ;
        RECT 433.950 526.950 436.050 529.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 427.950 523.950 430.050 526.050 ;
        RECT 409.950 520.950 412.050 523.050 ;
        RECT 416.400 521.400 417.600 523.650 ;
        RECT 410.400 505.050 411.450 520.950 ;
        RECT 416.400 517.050 417.450 521.400 ;
        RECT 421.950 520.950 424.050 523.050 ;
        RECT 415.950 514.950 418.050 517.050 ;
        RECT 412.950 511.950 415.050 514.050 ;
        RECT 409.950 502.950 412.050 505.050 ;
        RECT 413.400 495.600 414.450 511.950 ;
        RECT 413.400 495.450 414.600 495.600 ;
        RECT 410.400 494.400 414.600 495.450 ;
        RECT 406.950 481.950 409.050 484.050 ;
        RECT 410.400 466.050 411.450 494.400 ;
        RECT 413.400 493.350 414.600 494.400 ;
        RECT 413.400 490.950 415.500 493.050 ;
        RECT 418.800 490.950 420.900 493.050 ;
        RECT 419.400 489.000 420.600 490.650 ;
        RECT 422.400 489.900 423.450 520.950 ;
        RECT 428.400 496.200 429.450 523.950 ;
        RECT 433.950 520.950 436.050 523.050 ;
        RECT 437.400 521.400 438.900 540.300 ;
        RECT 441.300 534.300 442.500 540.300 ;
        RECT 440.400 532.200 442.500 534.300 ;
        RECT 434.400 508.050 435.450 520.950 ;
        RECT 437.400 519.300 439.500 521.400 ;
        RECT 438.300 515.700 439.500 519.300 ;
        RECT 441.300 515.700 442.500 532.200 ;
        RECT 443.700 537.300 445.800 539.400 ;
        RECT 451.950 538.950 454.050 541.050 ;
        RECT 460.200 540.300 462.300 542.400 ;
        RECT 443.700 515.700 444.900 537.300 ;
        RECT 448.950 535.950 451.050 538.050 ;
        RECT 449.400 525.600 450.450 535.950 ;
        RECT 452.400 535.800 454.500 537.900 ;
        RECT 457.800 537.300 459.900 539.400 ;
        RECT 452.400 529.200 453.300 535.800 ;
        RECT 458.100 530.100 459.300 537.300 ;
        RECT 460.800 535.500 462.300 540.300 ;
        RECT 463.200 537.300 465.300 542.400 ;
        RECT 460.800 533.400 462.900 535.500 ;
        RECT 452.400 527.100 454.500 529.200 ;
        RECT 457.800 528.000 459.900 530.100 ;
        RECT 449.400 523.350 450.600 525.600 ;
        RECT 448.800 520.950 450.900 523.050 ;
        RECT 452.400 516.600 453.300 527.100 ;
        RECT 455.100 520.500 457.200 522.600 ;
        RECT 437.700 513.600 439.800 515.700 ;
        RECT 440.700 513.600 442.800 515.700 ;
        RECT 443.700 513.600 445.800 515.700 ;
        RECT 451.800 514.500 453.900 516.600 ;
        RECT 458.100 515.700 459.300 528.000 ;
        RECT 460.800 515.700 462.300 533.400 ;
        RECT 464.100 515.700 465.300 537.300 ;
        RECT 457.200 513.600 459.300 515.700 ;
        RECT 460.200 513.600 462.300 515.700 ;
        RECT 463.200 513.600 465.300 515.700 ;
        RECT 466.200 540.300 468.300 542.400 ;
        RECT 470.400 541.050 471.450 559.950 ;
        RECT 472.950 556.950 475.050 559.050 ;
        RECT 473.400 547.050 474.450 556.950 ;
        RECT 472.950 544.950 475.050 547.050 ;
        RECT 466.200 535.500 467.700 540.300 ;
        RECT 469.950 538.950 472.050 541.050 ;
        RECT 466.200 533.400 468.300 535.500 ;
        RECT 476.400 535.050 477.450 559.950 ;
        RECT 466.200 515.700 467.700 533.400 ;
        RECT 475.950 532.950 478.050 535.050 ;
        RECT 475.800 526.950 477.900 529.050 ;
        RECT 476.400 525.900 477.600 526.650 ;
        RECT 475.950 523.800 478.050 525.900 ;
        RECT 466.200 513.600 468.300 515.700 ;
        RECT 479.400 514.050 480.450 571.950 ;
        RECT 482.400 554.700 483.900 573.600 ;
        RECT 486.300 562.800 487.500 579.300 ;
        RECT 485.400 560.700 487.500 562.800 ;
        RECT 486.300 554.700 487.500 560.700 ;
        RECT 488.700 557.700 489.900 579.300 ;
        RECT 496.800 578.400 498.900 580.500 ;
        RECT 502.200 579.300 504.300 581.400 ;
        RECT 505.200 579.300 507.300 581.400 ;
        RECT 508.200 579.300 510.300 581.400 ;
        RECT 493.800 571.950 495.900 574.050 ;
        RECT 494.400 570.900 495.600 571.650 ;
        RECT 493.950 568.800 496.050 570.900 ;
        RECT 497.400 567.900 498.300 578.400 ;
        RECT 500.100 572.400 502.200 574.500 ;
        RECT 497.400 565.800 499.500 567.900 ;
        RECT 503.100 567.000 504.300 579.300 ;
        RECT 497.400 559.200 498.300 565.800 ;
        RECT 502.800 564.900 504.900 567.000 ;
        RECT 488.700 555.600 490.800 557.700 ;
        RECT 497.400 557.100 499.500 559.200 ;
        RECT 503.100 557.700 504.300 564.900 ;
        RECT 505.800 561.600 507.300 579.300 ;
        RECT 505.800 559.500 507.900 561.600 ;
        RECT 502.800 555.600 504.900 557.700 ;
        RECT 505.800 554.700 507.300 559.500 ;
        RECT 509.100 557.700 510.300 579.300 ;
        RECT 482.400 552.600 485.400 554.700 ;
        RECT 486.300 552.600 488.400 554.700 ;
        RECT 493.950 550.950 496.050 553.050 ;
        RECT 505.200 552.600 507.300 554.700 ;
        RECT 508.200 552.600 510.300 557.700 ;
        RECT 511.200 579.300 513.300 581.400 ;
        RECT 511.200 561.600 512.700 579.300 ;
        RECT 511.200 559.500 513.300 561.600 ;
        RECT 511.200 554.700 512.700 559.500 ;
        RECT 511.200 552.600 513.300 554.700 ;
        RECT 487.950 547.950 490.050 550.050 ;
        RECT 484.800 526.950 486.900 529.050 ;
        RECT 485.400 525.000 486.600 526.650 ;
        RECT 484.950 520.950 487.050 525.000 ;
        RECT 481.950 514.950 484.050 517.050 ;
        RECT 478.950 511.950 481.050 514.050 ;
        RECT 482.400 508.050 483.450 514.950 ;
        RECT 433.950 505.950 436.050 508.050 ;
        RECT 442.950 505.950 445.050 508.050 ;
        RECT 448.950 505.950 451.050 508.050 ;
        RECT 481.950 505.950 484.050 508.050 ;
        RECT 427.950 494.100 430.050 496.200 ;
        RECT 439.950 494.100 442.050 496.200 ;
        RECT 440.400 493.350 441.600 494.100 ;
        RECT 434.100 490.950 436.200 493.050 ;
        RECT 439.500 490.950 441.600 493.050 ;
        RECT 418.950 484.950 421.050 489.000 ;
        RECT 421.950 487.800 424.050 489.900 ;
        RECT 434.400 488.400 435.600 490.650 ;
        RECT 409.950 463.950 412.050 466.050 ;
        RECT 415.950 463.950 418.050 466.050 ;
        RECT 412.950 454.950 415.050 457.050 ;
        RECT 409.950 451.950 412.050 454.050 ;
        RECT 386.400 448.350 387.600 450.600 ;
        RECT 391.950 449.100 394.050 451.200 ;
        RECT 397.950 449.100 400.050 451.200 ;
        RECT 403.950 449.100 406.050 451.200 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 383.400 444.900 384.600 445.650 ;
        RECT 382.950 442.800 385.050 444.900 ;
        RECT 379.950 439.950 382.050 442.050 ;
        RECT 376.950 430.950 379.050 433.050 ;
        RECT 376.950 424.950 379.050 427.050 ;
        RECT 373.950 400.950 376.050 403.050 ;
        RECT 370.950 388.950 373.050 391.050 ;
        RECT 367.950 355.950 370.050 358.050 ;
        RECT 364.950 352.950 367.050 355.050 ;
        RECT 365.400 349.050 366.450 352.950 ;
        RECT 364.950 346.950 367.050 349.050 ;
        RECT 361.950 343.950 364.050 346.050 ;
        RECT 362.400 340.200 363.450 343.950 ;
        RECT 371.400 343.050 372.450 388.950 ;
        RECT 373.950 382.950 376.050 385.050 ;
        RECT 361.950 338.100 364.050 340.200 ;
        RECT 364.950 339.000 367.050 343.050 ;
        RECT 370.950 340.950 373.050 343.050 ;
        RECT 365.400 337.350 366.600 339.000 ;
        RECT 365.400 334.950 367.500 337.050 ;
        RECT 370.800 334.950 372.900 337.050 ;
        RECT 371.400 332.400 372.600 334.650 ;
        RECT 358.950 316.950 361.050 319.050 ;
        RECT 361.950 313.950 364.050 316.050 ;
        RECT 349.950 307.950 352.050 310.050 ;
        RECT 362.400 304.050 363.450 313.950 ;
        RECT 371.400 307.050 372.450 332.400 ;
        RECT 370.950 304.950 373.050 307.050 ;
        RECT 361.950 301.950 364.050 304.050 ;
        RECT 374.400 303.450 375.450 382.950 ;
        RECT 371.400 302.400 375.450 303.450 ;
        RECT 349.950 295.950 352.050 298.050 ;
        RECT 335.400 292.350 336.600 294.000 ;
        RECT 340.950 293.100 343.050 295.200 ;
        RECT 346.950 293.100 349.050 295.200 ;
        RECT 341.400 292.350 342.600 293.100 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 332.400 287.400 333.600 289.650 ;
        RECT 338.400 288.900 339.600 289.650 ;
        RECT 325.950 283.950 328.050 286.050 ;
        RECT 332.400 274.050 333.450 287.400 ;
        RECT 337.950 286.800 340.050 288.900 ;
        RECT 331.950 271.950 334.050 274.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 311.400 255.000 312.600 256.650 ;
        RECT 301.950 250.950 304.050 253.050 ;
        RECT 310.950 250.950 313.050 255.000 ;
        RECT 298.950 241.950 301.050 244.050 ;
        RECT 310.950 241.950 313.050 244.050 ;
        RECT 295.950 240.900 300.000 241.050 ;
        RECT 295.950 238.950 301.050 240.900 ;
        RECT 301.950 238.950 304.050 241.050 ;
        RECT 304.950 238.950 307.050 241.050 ;
        RECT 298.950 238.800 301.050 238.950 ;
        RECT 292.950 232.950 295.050 235.050 ;
        RECT 298.950 232.950 301.050 235.050 ;
        RECT 293.400 226.050 294.450 232.950 ;
        RECT 292.950 223.950 295.050 226.050 ;
        RECT 292.950 215.100 295.050 220.050 ;
        RECT 299.400 216.600 300.450 232.950 ;
        RECT 302.400 222.450 303.450 238.950 ;
        RECT 305.400 232.050 306.450 238.950 ;
        RECT 304.950 229.950 307.050 232.050 ;
        RECT 307.950 229.950 310.050 232.050 ;
        RECT 304.950 222.450 307.050 223.050 ;
        RECT 302.400 221.400 307.050 222.450 ;
        RECT 304.950 220.950 307.050 221.400 ;
        RECT 305.400 217.050 306.450 220.950 ;
        RECT 293.400 214.350 294.600 215.100 ;
        RECT 299.400 214.350 300.600 216.600 ;
        RECT 304.950 214.950 307.050 217.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 289.950 208.950 292.050 211.050 ;
        RECT 296.400 209.400 297.600 211.650 ;
        RECT 302.400 210.900 303.600 211.650 ;
        RECT 290.400 196.050 291.450 208.950 ;
        RECT 292.950 205.950 295.050 208.050 ;
        RECT 289.950 193.950 292.050 196.050 ;
        RECT 277.950 187.950 280.050 190.050 ;
        RECT 286.950 187.950 289.050 190.050 ;
        RECT 274.950 172.950 277.050 175.050 ;
        RECT 274.950 169.800 277.050 171.900 ;
        RECT 275.400 166.050 276.450 169.800 ;
        RECT 274.950 163.950 277.050 166.050 ;
        RECT 275.400 154.050 276.450 163.950 ;
        RECT 278.400 160.050 279.450 187.950 ;
        RECT 286.950 182.100 289.050 184.200 ;
        RECT 293.400 184.050 294.450 205.950 ;
        RECT 296.400 205.050 297.450 209.400 ;
        RECT 301.950 208.800 304.050 210.900 ;
        RECT 304.950 208.950 307.050 211.050 ;
        RECT 296.400 203.400 301.050 205.050 ;
        RECT 297.000 202.950 301.050 203.400 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 301.950 199.950 304.050 202.050 ;
        RECT 287.400 181.350 288.600 182.100 ;
        RECT 292.950 181.950 295.050 184.050 ;
        RECT 283.950 178.950 286.050 181.050 ;
        RECT 286.950 178.950 289.050 181.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 284.400 176.400 285.600 178.650 ;
        RECT 290.400 177.900 291.600 178.650 ;
        RECT 280.950 172.950 283.050 175.050 ;
        RECT 281.400 168.450 282.450 172.950 ;
        RECT 284.400 172.050 285.450 176.400 ;
        RECT 289.950 175.800 292.050 177.900 ;
        RECT 283.950 169.950 286.050 172.050 ;
        RECT 289.950 169.950 292.050 174.750 ;
        RECT 296.400 172.050 297.450 199.950 ;
        RECT 298.950 196.950 301.050 199.050 ;
        RECT 299.400 184.050 300.450 196.950 ;
        RECT 302.400 187.050 303.450 199.950 ;
        RECT 305.400 190.050 306.450 208.950 ;
        RECT 308.400 205.050 309.450 229.950 ;
        RECT 311.400 210.450 312.450 241.950 ;
        RECT 317.400 232.050 318.450 260.400 ;
        RECT 323.400 259.350 324.600 261.600 ;
        RECT 328.950 260.100 331.050 262.200 ;
        RECT 337.800 260.100 339.900 262.200 ;
        RECT 340.950 260.100 343.050 262.200 ;
        RECT 347.400 261.600 348.450 293.100 ;
        RECT 350.400 289.050 351.450 295.950 ;
        RECT 355.950 294.000 358.050 298.050 ;
        RECT 356.400 292.350 357.600 294.000 ;
        RECT 361.950 293.100 364.050 295.200 ;
        RECT 362.400 292.350 363.600 293.100 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 349.950 286.950 352.050 289.050 ;
        RECT 359.400 287.400 360.600 289.650 ;
        RECT 365.400 288.900 366.600 289.650 ;
        RECT 371.400 289.050 372.450 302.400 ;
        RECT 377.400 300.450 378.450 424.950 ;
        RECT 380.400 418.200 381.450 439.950 ;
        RECT 383.400 427.050 384.450 442.800 ;
        RECT 382.950 424.950 385.050 427.050 ;
        RECT 379.950 416.100 382.050 418.200 ;
        RECT 380.400 415.350 381.600 416.100 ;
        RECT 380.400 412.950 382.500 415.050 ;
        RECT 385.800 412.950 387.900 415.050 ;
        RECT 386.400 410.400 387.600 412.650 ;
        RECT 379.950 397.950 382.050 400.050 ;
        RECT 380.400 391.050 381.450 397.950 ;
        RECT 379.950 388.950 382.050 391.050 ;
        RECT 380.400 372.600 381.450 388.950 ;
        RECT 386.400 388.050 387.450 410.400 ;
        RECT 392.400 409.050 393.450 449.100 ;
        RECT 398.400 448.350 399.600 449.100 ;
        RECT 404.400 448.350 405.600 449.100 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 400.950 445.950 403.050 448.050 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 401.400 443.400 402.600 445.650 ;
        RECT 394.950 439.950 397.050 442.050 ;
        RECT 391.950 406.950 394.050 409.050 ;
        RECT 385.950 385.950 388.050 388.050 ;
        RECT 380.400 370.350 381.600 372.600 ;
        RECT 388.950 372.000 391.050 376.050 ;
        RECT 389.400 370.350 390.600 372.000 ;
        RECT 380.100 367.950 382.200 370.050 ;
        RECT 385.500 367.950 387.600 370.050 ;
        RECT 388.800 367.950 390.900 370.050 ;
        RECT 386.400 366.000 387.600 367.650 ;
        RECT 385.950 361.950 388.050 366.000 ;
        RECT 392.400 360.450 393.450 406.950 ;
        RECT 395.400 366.900 396.450 439.950 ;
        RECT 401.400 439.050 402.450 443.400 ;
        RECT 406.950 442.950 409.050 445.050 ;
        RECT 400.950 436.950 403.050 439.050 ;
        RECT 401.400 417.600 402.450 436.950 ;
        RECT 407.400 421.050 408.450 442.950 ;
        RECT 406.950 418.950 409.050 421.050 ;
        RECT 401.400 415.350 402.600 417.600 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 404.400 411.900 405.600 412.650 ;
        RECT 403.950 409.800 406.050 411.900 ;
        RECT 410.400 406.050 411.450 451.950 ;
        RECT 413.400 451.050 414.450 454.950 ;
        RECT 416.400 454.050 417.450 463.950 ;
        RECT 412.950 448.950 415.050 451.050 ;
        RECT 415.950 450.000 418.050 454.050 ;
        RECT 421.950 450.000 424.050 454.050 ;
        RECT 434.400 451.200 435.450 488.400 ;
        RECT 443.400 481.050 444.450 505.950 ;
        RECT 442.950 478.950 445.050 481.050 ;
        RECT 449.400 466.050 450.450 505.950 ;
        RECT 484.950 502.950 487.050 505.050 ;
        RECT 451.950 499.950 454.050 502.050 ;
        RECT 448.950 463.950 451.050 466.050 ;
        RECT 436.950 451.950 439.050 454.050 ;
        RECT 416.400 448.350 417.600 450.000 ;
        RECT 422.400 448.350 423.600 450.000 ;
        RECT 427.950 449.100 430.050 451.200 ;
        RECT 433.950 449.100 436.050 451.200 ;
        RECT 428.400 448.350 429.600 449.100 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 424.950 445.950 427.050 448.050 ;
        RECT 427.950 445.950 430.050 448.050 ;
        RECT 419.400 444.900 420.600 445.650 ;
        RECT 418.950 439.950 421.050 444.900 ;
        RECT 425.400 443.400 426.600 445.650 ;
        RECT 412.950 433.950 415.050 436.050 ;
        RECT 400.950 403.950 403.050 406.050 ;
        RECT 409.950 403.950 412.050 406.050 ;
        RECT 401.400 372.600 402.450 403.950 ;
        RECT 401.400 372.450 402.600 372.600 ;
        RECT 398.400 371.400 402.600 372.450 ;
        RECT 394.950 364.800 397.050 366.900 ;
        RECT 392.400 359.400 396.450 360.450 ;
        RECT 391.950 355.950 394.050 358.050 ;
        RECT 382.950 346.950 385.050 349.050 ;
        RECT 379.950 340.950 382.050 343.050 ;
        RECT 374.400 299.400 378.450 300.450 ;
        RECT 359.400 268.050 360.450 287.400 ;
        RECT 364.950 286.800 367.050 288.900 ;
        RECT 370.950 286.950 373.050 289.050 ;
        RECT 361.950 283.950 364.050 286.050 ;
        RECT 358.950 265.950 361.050 268.050 ;
        RECT 329.400 259.350 330.600 260.100 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 319.950 253.950 322.050 256.050 ;
        RECT 326.400 255.000 327.600 256.650 ;
        RECT 313.950 230.400 318.450 232.050 ;
        RECT 313.950 229.950 318.000 230.400 ;
        RECT 316.950 223.950 319.050 226.050 ;
        RECT 313.950 217.950 316.050 220.050 ;
        RECT 314.400 214.050 315.450 217.950 ;
        RECT 317.400 216.600 318.450 223.950 ;
        RECT 320.400 219.450 321.450 253.950 ;
        RECT 325.950 250.950 328.050 255.000 ;
        RECT 332.400 254.400 333.600 256.650 ;
        RECT 332.400 253.050 333.450 254.400 ;
        RECT 334.950 253.950 337.050 256.050 ;
        RECT 331.950 250.950 334.050 253.050 ;
        RECT 332.400 243.450 333.450 250.950 ;
        RECT 329.400 242.400 333.450 243.450 ;
        RECT 322.950 232.950 325.050 235.050 ;
        RECT 323.400 226.050 324.450 232.950 ;
        RECT 322.950 223.950 325.050 226.050 ;
        RECT 324.000 222.450 328.050 223.050 ;
        RECT 323.400 222.000 328.050 222.450 ;
        RECT 322.950 220.950 328.050 222.000 ;
        RECT 322.950 219.450 325.050 220.950 ;
        RECT 320.400 218.400 325.050 219.450 ;
        RECT 322.950 217.950 325.050 218.400 ;
        RECT 317.400 214.350 318.600 216.600 ;
        RECT 325.950 215.100 328.050 217.200 ;
        RECT 326.400 214.350 327.600 215.100 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 317.100 211.950 319.200 214.050 ;
        RECT 322.500 211.950 324.600 214.050 ;
        RECT 325.800 211.950 327.900 214.050 ;
        RECT 323.400 210.900 324.600 211.650 ;
        RECT 311.400 209.400 315.450 210.450 ;
        RECT 310.950 205.950 313.050 208.050 ;
        RECT 307.950 202.950 310.050 205.050 ;
        RECT 304.950 187.950 307.050 190.050 ;
        RECT 301.950 184.950 304.050 187.050 ;
        RECT 298.950 181.950 301.050 184.050 ;
        RECT 304.950 182.100 307.050 184.200 ;
        RECT 311.400 184.050 312.450 205.950 ;
        RECT 305.400 181.350 306.600 182.100 ;
        RECT 310.950 181.950 313.050 184.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 302.400 177.900 303.600 178.650 ;
        RECT 308.400 177.900 309.600 178.650 ;
        RECT 301.950 175.800 304.050 177.900 ;
        RECT 307.950 175.800 310.050 177.900 ;
        RECT 295.950 169.950 298.050 172.050 ;
        RECT 302.400 169.050 303.450 175.800 ;
        RECT 304.950 172.950 307.050 175.050 ;
        RECT 281.400 167.400 285.450 168.450 ;
        RECT 284.400 163.050 285.450 167.400 ;
        RECT 301.950 166.950 304.050 169.050 ;
        RECT 305.400 163.050 306.450 172.950 ;
        RECT 283.950 160.950 286.050 163.050 ;
        RECT 304.950 160.950 307.050 163.050 ;
        RECT 277.950 157.950 280.050 160.050 ;
        RECT 274.950 151.950 277.050 154.050 ;
        RECT 271.950 139.950 274.050 142.050 ;
        RECT 274.950 139.950 277.050 142.050 ;
        RECT 257.400 136.350 258.600 137.400 ;
        RECT 263.400 136.350 264.600 138.000 ;
        RECT 269.400 137.400 273.450 138.450 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 260.400 132.900 261.600 133.650 ;
        RECT 266.400 132.900 267.600 133.650 ;
        RECT 229.950 121.950 232.050 124.050 ;
        RECT 236.400 121.050 237.450 131.400 ;
        RECT 241.950 130.800 244.050 132.900 ;
        RECT 250.950 130.800 253.050 132.900 ;
        RECT 259.950 130.800 262.050 132.900 ;
        RECT 265.950 130.800 268.050 132.900 ;
        RECT 272.400 132.450 273.450 137.400 ;
        RECT 269.400 131.400 273.450 132.450 ;
        RECT 238.950 127.950 241.050 130.050 ;
        RECT 235.950 120.450 238.050 121.050 ;
        RECT 233.400 119.400 238.050 120.450 ;
        RECT 226.950 112.950 229.050 115.050 ;
        RECT 233.400 111.450 234.450 119.400 ;
        RECT 235.950 118.950 238.050 119.400 ;
        RECT 239.400 118.050 240.450 127.950 ;
        RECT 265.950 121.950 268.050 124.050 ;
        RECT 244.950 118.950 247.050 121.050 ;
        RECT 259.950 118.950 262.050 121.050 ;
        RECT 238.950 115.950 241.050 118.050 ;
        RECT 235.950 114.450 238.050 115.050 ;
        RECT 241.950 114.450 244.050 115.050 ;
        RECT 235.950 113.400 244.050 114.450 ;
        RECT 235.950 112.950 238.050 113.400 ;
        RECT 241.950 112.950 244.050 113.400 ;
        RECT 245.400 111.450 246.450 118.950 ;
        RECT 253.950 112.950 256.050 115.050 ;
        RECT 233.400 110.400 246.450 111.450 ;
        RECT 229.950 106.950 232.050 109.050 ;
        RECT 218.400 103.350 219.600 105.000 ;
        RECT 224.400 103.350 225.600 105.600 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 220.950 100.950 223.050 103.050 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 211.950 97.950 214.050 100.050 ;
        RECT 221.400 98.400 222.600 100.650 ;
        RECT 221.400 91.050 222.450 98.400 ;
        RECT 220.950 88.950 223.050 91.050 ;
        RECT 230.400 85.050 231.450 106.950 ;
        RECT 238.950 104.100 241.050 106.200 ;
        RECT 244.950 104.100 247.050 106.200 ;
        RECT 239.400 103.350 240.600 104.100 ;
        RECT 245.400 103.350 246.600 104.100 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 242.400 98.400 243.600 100.650 ;
        RECT 248.400 99.900 249.600 100.650 ;
        RECT 229.950 82.950 232.050 85.050 ;
        RECT 211.950 73.950 214.050 76.050 ;
        RECT 206.400 68.400 210.450 69.450 ;
        RECT 191.400 58.350 192.600 59.100 ;
        RECT 197.400 58.350 198.600 59.100 ;
        RECT 202.950 58.950 205.050 61.050 ;
        RECT 181.950 57.000 186.450 57.450 ;
        RECT 182.400 56.400 186.450 57.000 ;
        RECT 143.400 49.050 144.450 53.400 ;
        RECT 148.950 52.800 151.050 54.900 ;
        RECT 160.950 52.800 163.050 54.900 ;
        RECT 167.400 53.400 168.600 55.650 ;
        RECT 173.400 54.900 174.600 55.650 ;
        RECT 142.950 46.950 145.050 49.050 ;
        RECT 167.400 46.050 168.450 53.400 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 178.950 52.950 184.050 55.050 ;
        RECT 185.400 52.050 186.450 56.400 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 187.950 52.950 190.050 55.050 ;
        RECT 194.400 54.000 195.600 55.650 ;
        RECT 200.400 54.900 201.600 55.650 ;
        RECT 206.400 54.900 207.450 68.400 ;
        RECT 208.950 64.950 211.050 67.050 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 178.950 46.950 181.050 49.050 ;
        RECT 166.950 43.950 169.050 46.050 ;
        RECT 127.950 37.950 130.050 40.050 ;
        RECT 136.950 37.950 139.050 40.050 ;
        RECT 121.950 34.950 124.050 37.050 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 97.950 22.950 100.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 118.950 22.950 121.050 25.050 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 83.400 21.900 84.600 22.650 ;
        RECT 89.400 21.900 90.600 22.650 ;
        RECT 82.950 19.800 85.050 21.900 ;
        RECT 88.950 19.800 91.050 21.900 ;
        RECT 100.950 19.950 103.050 22.050 ;
        RECT 104.400 20.400 105.600 22.650 ;
        RECT 110.400 21.900 111.600 22.650 ;
        RECT 73.950 16.950 76.050 19.050 ;
        RECT 101.400 16.050 102.450 19.950 ;
        RECT 100.950 13.950 103.050 16.050 ;
        RECT 52.950 10.950 55.050 13.050 ;
        RECT 104.400 10.050 105.450 20.400 ;
        RECT 109.950 19.800 112.050 21.900 ;
        RECT 122.400 16.050 123.450 34.950 ;
        RECT 128.400 28.200 129.450 37.950 ;
        RECT 169.950 34.950 172.050 37.050 ;
        RECT 166.950 31.950 169.050 34.050 ;
        RECT 157.950 28.950 160.050 31.050 ;
        RECT 127.950 26.100 130.050 28.200 ;
        RECT 143.400 27.450 144.600 27.600 ;
        RECT 137.400 26.400 144.600 27.450 ;
        RECT 128.400 25.350 129.600 26.100 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 131.400 21.900 132.600 22.650 ;
        RECT 121.950 13.950 124.050 16.050 ;
        RECT 125.400 10.050 126.450 19.950 ;
        RECT 130.950 19.800 133.050 21.900 ;
        RECT 137.400 13.050 138.450 26.400 ;
        RECT 143.400 25.350 144.600 26.400 ;
        RECT 148.950 26.100 151.050 28.200 ;
        RECT 149.400 25.350 150.600 26.100 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 146.400 21.000 147.600 22.650 ;
        RECT 152.400 21.900 153.600 22.650 ;
        RECT 145.950 16.950 148.050 21.000 ;
        RECT 151.950 19.800 154.050 21.900 ;
        RECT 158.400 19.050 159.450 28.950 ;
        RECT 167.400 28.200 168.450 31.950 ;
        RECT 170.400 31.050 171.450 34.950 ;
        RECT 169.950 28.950 172.050 31.050 ;
        RECT 166.950 26.100 169.050 28.200 ;
        RECT 174.000 27.600 178.050 28.050 ;
        RECT 167.400 25.350 168.600 26.100 ;
        RECT 173.400 25.950 178.050 27.600 ;
        RECT 173.400 25.350 174.600 25.950 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 164.400 21.900 165.600 22.650 ;
        RECT 170.400 21.900 171.600 22.650 ;
        RECT 179.400 22.050 180.450 46.950 ;
        RECT 188.400 34.050 189.450 52.950 ;
        RECT 193.950 49.950 196.050 54.000 ;
        RECT 199.950 52.800 202.050 54.900 ;
        RECT 205.950 52.800 208.050 54.900 ;
        RECT 196.950 40.950 199.050 43.050 ;
        RECT 187.950 31.950 190.050 34.050 ;
        RECT 181.950 26.100 184.050 28.200 ;
        RECT 190.950 26.100 193.050 28.200 ;
        RECT 197.400 27.600 198.450 40.950 ;
        RECT 200.400 31.050 201.450 52.800 ;
        RECT 209.400 37.050 210.450 64.950 ;
        RECT 212.400 61.050 213.450 73.950 ;
        RECT 217.950 64.950 220.050 67.050 ;
        RECT 211.950 58.950 214.050 61.050 ;
        RECT 218.400 60.600 219.450 64.950 ;
        RECT 218.400 58.350 219.600 60.600 ;
        RECT 223.950 59.100 226.050 61.200 ;
        RECT 229.950 59.100 232.050 61.200 ;
        RECT 235.950 59.100 238.050 61.200 ;
        RECT 242.400 61.050 243.450 98.400 ;
        RECT 247.950 97.800 250.050 99.900 ;
        RECT 244.950 88.950 247.050 91.050 ;
        RECT 224.400 58.350 225.600 59.100 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 220.950 55.950 223.050 58.050 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 215.400 54.900 216.600 55.650 ;
        RECT 214.950 52.800 217.050 54.900 ;
        RECT 221.400 53.400 222.600 55.650 ;
        RECT 221.400 49.050 222.450 53.400 ;
        RECT 220.950 46.950 223.050 49.050 ;
        RECT 217.950 40.950 220.050 43.050 ;
        RECT 218.400 37.050 219.450 40.950 ;
        RECT 221.400 40.050 222.450 46.950 ;
        RECT 220.950 37.950 223.050 40.050 ;
        RECT 208.950 34.950 211.050 37.050 ;
        RECT 217.950 34.950 220.050 37.050 ;
        RECT 199.950 28.950 202.050 31.050 ;
        RECT 163.950 19.800 166.050 21.900 ;
        RECT 169.950 19.800 172.050 21.900 ;
        RECT 178.950 19.950 181.050 22.050 ;
        RECT 157.950 16.950 160.050 19.050 ;
        RECT 136.950 10.950 139.050 13.050 ;
        RECT 103.950 7.950 106.050 10.050 ;
        RECT 124.950 7.950 127.050 10.050 ;
        RECT 164.400 7.050 165.450 19.800 ;
        RECT 182.400 16.050 183.450 26.100 ;
        RECT 191.400 25.350 192.600 26.100 ;
        RECT 197.400 25.350 198.600 27.600 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 202.950 22.950 205.050 28.200 ;
        RECT 211.950 26.100 214.050 28.200 ;
        RECT 217.950 26.100 220.050 28.200 ;
        RECT 230.400 28.050 231.450 59.100 ;
        RECT 236.400 58.350 237.600 59.100 ;
        RECT 241.950 58.950 244.050 61.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 239.400 54.000 240.600 55.650 ;
        RECT 245.400 55.050 246.450 88.950 ;
        RECT 248.400 67.050 249.450 97.800 ;
        RECT 254.400 97.050 255.450 112.950 ;
        RECT 256.950 103.950 259.050 106.050 ;
        RECT 260.400 105.450 261.450 118.950 ;
        RECT 262.950 115.950 265.050 118.050 ;
        RECT 263.400 109.050 264.450 115.950 ;
        RECT 266.400 115.050 267.450 121.950 ;
        RECT 265.950 112.950 268.050 115.050 ;
        RECT 262.950 106.950 265.050 109.050 ;
        RECT 269.400 105.600 270.450 131.400 ;
        RECT 271.950 124.950 274.050 127.050 ;
        RECT 272.400 109.050 273.450 124.950 ;
        RECT 271.950 106.950 274.050 109.050 ;
        RECT 275.400 106.050 276.450 139.950 ;
        RECT 277.950 138.450 280.050 145.050 ;
        RECT 283.800 142.200 285.900 144.300 ;
        RECT 292.800 142.500 294.900 144.600 ;
        RECT 307.950 142.950 310.050 145.050 ;
        RECT 281.400 138.450 282.600 138.600 ;
        RECT 277.950 138.000 282.600 138.450 ;
        RECT 278.400 137.400 282.600 138.000 ;
        RECT 281.400 136.350 282.600 137.400 ;
        RECT 281.100 133.950 283.200 136.050 ;
        RECT 284.100 129.600 285.000 142.200 ;
        RECT 290.400 139.350 291.600 141.600 ;
        RECT 290.100 136.950 292.200 139.050 ;
        RECT 285.900 135.900 288.000 136.200 ;
        RECT 294.000 135.900 294.900 142.500 ;
        RECT 298.950 136.950 301.050 139.050 ;
        RECT 308.400 138.600 309.450 142.950 ;
        RECT 314.400 142.200 315.450 209.400 ;
        RECT 322.950 208.800 325.050 210.900 ;
        RECT 329.400 208.050 330.450 242.400 ;
        RECT 335.400 241.050 336.450 253.950 ;
        RECT 334.950 238.950 337.050 241.050 ;
        RECT 338.400 235.050 339.450 260.100 ;
        RECT 341.400 253.050 342.450 260.100 ;
        RECT 347.400 259.350 348.600 261.600 ;
        RECT 352.950 260.100 355.050 262.200 ;
        RECT 353.400 259.350 354.600 260.100 ;
        RECT 362.400 259.050 363.450 283.950 ;
        RECT 370.950 283.800 373.050 285.900 ;
        RECT 367.950 280.950 370.050 283.050 ;
        RECT 364.950 277.950 367.050 280.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 350.400 255.000 351.600 256.650 ;
        RECT 356.400 255.450 357.600 256.650 ;
        RECT 365.400 256.050 366.450 277.950 ;
        RECT 368.400 262.050 369.450 280.950 ;
        RECT 367.950 259.950 370.050 262.050 ;
        RECT 371.400 261.600 372.450 283.800 ;
        RECT 374.400 280.050 375.450 299.400 ;
        RECT 380.400 298.050 381.450 340.950 ;
        RECT 383.400 339.600 384.450 346.950 ;
        RECT 383.400 337.350 384.600 339.600 ;
        RECT 383.400 334.950 385.500 337.050 ;
        RECT 388.800 334.950 390.900 337.050 ;
        RECT 389.400 332.400 390.600 334.650 ;
        RECT 389.400 310.050 390.450 332.400 ;
        RECT 388.950 307.950 391.050 310.050 ;
        RECT 382.950 298.950 385.050 301.050 ;
        RECT 379.950 295.950 382.050 298.050 ;
        RECT 383.400 294.600 384.450 298.950 ;
        RECT 383.400 292.350 384.600 294.600 ;
        RECT 388.950 293.100 391.050 295.200 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 380.400 288.900 381.600 289.650 ;
        RECT 379.950 286.800 382.050 288.900 ;
        RECT 376.950 280.950 379.050 283.050 ;
        RECT 373.950 277.950 376.050 280.050 ;
        RECT 377.400 271.050 378.450 280.950 ;
        RECT 376.950 268.950 379.050 271.050 ;
        RECT 371.400 259.350 372.600 261.600 ;
        RECT 371.400 256.950 373.500 259.050 ;
        RECT 376.800 256.950 378.900 259.050 ;
        RECT 340.950 250.950 343.050 253.050 ;
        RECT 349.950 250.950 352.050 255.000 ;
        RECT 356.400 254.400 360.450 255.450 ;
        RECT 349.950 244.950 352.050 247.050 ;
        RECT 343.950 238.950 346.050 241.050 ;
        RECT 337.950 232.950 340.050 235.050 ;
        RECT 331.950 226.950 334.050 229.050 ;
        RECT 337.950 226.950 340.050 229.050 ;
        RECT 328.950 205.950 331.050 208.050 ;
        RECT 332.400 199.050 333.450 226.950 ;
        RECT 338.400 217.200 339.450 226.950 ;
        RECT 337.950 215.100 340.050 217.200 ;
        RECT 344.400 216.600 345.450 238.950 ;
        RECT 338.400 214.350 339.600 215.100 ;
        RECT 344.400 214.350 345.600 216.600 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 341.400 210.900 342.600 211.650 ;
        RECT 340.950 208.800 343.050 210.900 ;
        RECT 346.950 208.950 349.050 211.050 ;
        RECT 337.950 205.950 340.050 208.050 ;
        RECT 331.950 196.950 334.050 199.050 ;
        RECT 334.950 193.950 337.050 196.050 ;
        RECT 331.950 187.950 334.050 190.050 ;
        RECT 316.950 181.950 319.050 184.050 ;
        RECT 325.950 182.100 328.050 184.200 ;
        RECT 332.400 184.050 333.450 187.950 ;
        RECT 335.400 187.050 336.450 193.950 ;
        RECT 334.950 184.950 337.050 187.050 ;
        RECT 332.400 183.900 336.000 184.050 ;
        RECT 317.400 169.050 318.450 181.950 ;
        RECT 326.400 181.350 327.600 182.100 ;
        RECT 332.400 181.950 337.050 183.900 ;
        RECT 332.400 181.350 333.600 181.950 ;
        RECT 334.950 181.800 337.050 181.950 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 319.950 175.800 322.050 177.900 ;
        RECT 323.400 176.400 324.600 178.650 ;
        RECT 329.400 176.400 330.600 178.650 ;
        RECT 338.400 178.050 339.450 205.950 ;
        RECT 340.950 202.950 343.050 205.050 ;
        RECT 316.950 166.950 319.050 169.050 ;
        RECT 320.400 166.050 321.450 175.800 ;
        RECT 319.950 163.950 322.050 166.050 ;
        RECT 323.400 163.050 324.450 176.400 ;
        RECT 322.950 160.950 325.050 163.050 ;
        RECT 329.400 160.050 330.450 176.400 ;
        RECT 337.950 175.950 340.050 178.050 ;
        RECT 337.950 160.950 340.050 163.050 ;
        RECT 328.950 157.950 331.050 160.050 ;
        RECT 322.950 154.950 325.050 157.050 ;
        RECT 334.950 154.950 337.050 157.050 ;
        RECT 319.950 142.950 322.050 145.050 ;
        RECT 313.950 140.100 316.050 142.200 ;
        RECT 285.900 135.000 294.900 135.900 ;
        RECT 285.900 134.100 288.000 135.000 ;
        RECT 291.000 133.200 293.100 134.100 ;
        RECT 285.900 132.000 293.100 133.200 ;
        RECT 285.900 131.100 288.000 132.000 ;
        RECT 283.500 127.500 285.600 129.600 ;
        RECT 290.100 128.100 292.200 130.200 ;
        RECT 294.000 129.900 294.900 135.000 ;
        RECT 295.800 133.950 297.900 136.050 ;
        RECT 296.400 132.450 297.600 133.650 ;
        RECT 299.400 132.450 300.450 136.950 ;
        RECT 308.400 136.350 309.600 138.600 ;
        RECT 313.950 136.950 316.050 139.050 ;
        RECT 314.400 136.350 315.600 136.950 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 296.400 131.400 300.450 132.450 ;
        RECT 304.950 130.950 307.050 133.050 ;
        RECT 311.400 131.400 312.600 133.650 ;
        RECT 320.400 133.050 321.450 142.950 ;
        RECT 323.400 133.050 324.450 154.950 ;
        RECT 335.400 142.050 336.450 154.950 ;
        RECT 334.950 139.950 337.050 142.050 ;
        RECT 331.950 137.100 334.050 139.200 ;
        RECT 338.400 139.050 339.450 160.950 ;
        RECT 341.400 157.050 342.450 202.950 ;
        RECT 343.950 196.950 346.050 199.050 ;
        RECT 344.400 190.050 345.450 196.950 ;
        RECT 343.950 187.950 346.050 190.050 ;
        RECT 347.400 186.450 348.450 208.950 ;
        RECT 350.400 205.050 351.450 244.950 ;
        RECT 355.950 235.950 358.050 238.050 ;
        RECT 352.950 220.950 355.050 223.050 ;
        RECT 353.400 217.050 354.450 220.950 ;
        RECT 356.400 219.450 357.450 235.950 ;
        RECT 359.400 235.050 360.450 254.400 ;
        RECT 364.950 253.950 367.050 256.050 ;
        RECT 377.400 255.000 378.600 256.650 ;
        RECT 370.950 250.950 373.050 253.050 ;
        RECT 376.950 250.950 379.050 255.000 ;
        RECT 358.800 232.950 360.900 235.050 ;
        RECT 361.950 232.950 364.050 235.050 ;
        RECT 359.400 223.050 360.450 232.950 ;
        RECT 362.400 226.050 363.450 232.950 ;
        RECT 364.950 226.950 367.050 229.050 ;
        RECT 361.950 223.950 364.050 226.050 ;
        RECT 358.950 220.950 361.050 223.050 ;
        RECT 356.400 218.400 360.450 219.450 ;
        RECT 352.950 214.950 355.050 217.050 ;
        RECT 359.400 216.600 360.450 218.400 ;
        RECT 365.400 216.600 366.450 226.950 ;
        RECT 359.400 214.350 360.600 216.600 ;
        RECT 365.400 214.350 366.600 216.600 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 352.950 208.950 355.050 211.050 ;
        RECT 356.400 209.400 357.600 211.650 ;
        RECT 362.400 209.400 363.600 211.650 ;
        RECT 371.400 211.050 372.450 250.950 ;
        RECT 380.400 250.050 381.450 286.800 ;
        RECT 382.950 283.950 385.050 286.050 ;
        RECT 379.950 247.950 382.050 250.050 ;
        RECT 373.950 244.950 376.050 247.050 ;
        RECT 349.950 202.950 352.050 205.050 ;
        RECT 353.400 202.050 354.450 208.950 ;
        RECT 352.950 199.950 355.050 202.050 ;
        RECT 356.400 199.050 357.450 209.400 ;
        RECT 362.400 199.050 363.450 209.400 ;
        RECT 370.950 208.950 373.050 211.050 ;
        RECT 374.400 208.050 375.450 244.950 ;
        RECT 379.950 238.950 382.050 241.050 ;
        RECT 380.400 232.050 381.450 238.950 ;
        RECT 379.950 229.950 382.050 232.050 ;
        RECT 380.400 216.600 381.450 229.950 ;
        RECT 383.400 220.050 384.450 283.950 ;
        RECT 389.400 268.050 390.450 293.100 ;
        RECT 392.400 286.050 393.450 355.950 ;
        RECT 395.400 316.050 396.450 359.400 ;
        RECT 398.400 349.050 399.450 371.400 ;
        RECT 401.400 370.350 402.600 371.400 ;
        RECT 409.950 371.100 412.050 373.200 ;
        RECT 410.400 370.350 411.600 371.100 ;
        RECT 401.100 367.950 403.200 370.050 ;
        RECT 406.500 367.950 408.600 370.050 ;
        RECT 409.800 367.950 411.900 370.050 ;
        RECT 407.400 366.900 408.600 367.650 ;
        RECT 406.950 364.800 409.050 366.900 ;
        RECT 397.950 346.950 400.050 349.050 ;
        RECT 413.400 345.450 414.450 433.950 ;
        RECT 418.950 424.950 421.050 427.050 ;
        RECT 419.400 417.600 420.450 424.950 ;
        RECT 425.400 424.050 426.450 443.400 ;
        RECT 424.950 421.950 427.050 424.050 ;
        RECT 419.400 415.350 420.600 417.600 ;
        RECT 424.950 416.100 427.050 418.200 ;
        RECT 425.400 415.350 426.600 416.100 ;
        RECT 418.950 412.950 421.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 422.400 411.900 423.600 412.650 ;
        RECT 421.950 406.950 424.050 411.900 ;
        RECT 428.400 410.400 429.600 412.650 ;
        RECT 434.400 411.450 435.450 449.100 ;
        RECT 437.400 444.900 438.450 451.950 ;
        RECT 439.950 448.950 442.050 454.050 ;
        RECT 445.950 449.100 448.050 451.200 ;
        RECT 446.400 448.350 447.600 449.100 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 436.950 442.800 439.050 444.900 ;
        RECT 439.950 442.950 442.050 445.050 ;
        RECT 443.400 444.900 444.600 445.650 ;
        RECT 436.950 427.950 439.050 430.050 ;
        RECT 431.400 410.400 435.450 411.450 ;
        RECT 428.400 406.050 429.450 410.400 ;
        RECT 427.950 403.950 430.050 406.050 ;
        RECT 431.400 391.050 432.450 410.400 ;
        RECT 433.950 403.950 436.050 406.050 ;
        RECT 430.950 388.950 433.050 391.050 ;
        RECT 418.950 379.950 421.050 382.050 ;
        RECT 430.950 381.600 433.050 382.050 ;
        RECT 425.400 380.550 433.050 381.600 ;
        RECT 419.400 358.050 420.450 379.950 ;
        RECT 425.400 373.200 426.450 380.550 ;
        RECT 430.950 379.950 433.050 380.550 ;
        RECT 430.950 376.800 433.050 378.900 ;
        RECT 424.950 371.100 427.050 373.200 ;
        RECT 431.400 372.600 432.450 376.800 ;
        RECT 434.400 373.050 435.450 403.950 ;
        RECT 437.400 379.050 438.450 427.950 ;
        RECT 440.400 418.200 441.450 442.950 ;
        RECT 442.950 442.800 445.050 444.900 ;
        RECT 443.400 433.050 444.450 442.800 ;
        RECT 452.400 436.050 453.450 499.950 ;
        RECT 485.400 499.050 486.450 502.950 ;
        RECT 488.400 502.050 489.450 547.950 ;
        RECT 490.950 538.950 493.050 541.050 ;
        RECT 491.400 532.050 492.450 538.950 ;
        RECT 490.950 529.950 493.050 532.050 ;
        RECT 494.400 531.600 495.450 550.950 ;
        RECT 515.400 550.050 516.450 601.950 ;
        RECT 518.400 574.050 519.450 640.950 ;
        RECT 521.400 625.050 522.450 644.400 ;
        RECT 526.950 642.450 529.050 646.050 ;
        RECT 530.100 643.950 532.200 646.050 ;
        RECT 524.400 642.000 529.050 642.450 ;
        RECT 524.400 641.400 528.450 642.000 ;
        RECT 520.950 622.950 523.050 625.050 ;
        RECT 524.400 610.050 525.450 641.400 ;
        RECT 536.400 637.050 537.450 658.950 ;
        RECT 539.400 648.600 540.450 673.950 ;
        RECT 563.400 664.050 564.450 721.950 ;
        RECT 571.950 721.800 574.050 723.900 ;
        RECT 568.950 709.950 571.050 712.050 ;
        RECT 565.950 676.950 568.050 679.050 ;
        RECT 566.400 667.050 567.450 676.950 ;
        RECT 569.400 676.050 570.450 709.950 ;
        RECT 572.100 679.950 574.200 682.050 ;
        RECT 568.950 673.950 571.050 676.050 ;
        RECT 578.400 673.050 579.450 725.400 ;
        RECT 587.400 724.950 589.500 727.050 ;
        RECT 592.500 724.950 594.600 727.050 ;
        RECT 596.400 709.050 597.450 728.100 ;
        RECT 595.950 706.950 598.050 709.050 ;
        RECT 580.950 700.800 583.050 702.900 ;
        RECT 581.400 678.900 582.450 700.800 ;
        RECT 602.400 700.050 603.450 751.950 ;
        RECT 598.950 697.950 603.450 700.050 ;
        RECT 589.950 683.100 592.050 685.200 ;
        RECT 595.800 683.100 597.900 685.200 ;
        RECT 602.400 685.050 603.450 697.950 ;
        RECT 605.400 688.050 606.450 752.400 ;
        RECT 611.400 745.050 612.450 793.950 ;
        RECT 614.400 763.050 615.450 806.100 ;
        RECT 617.400 769.050 618.450 806.400 ;
        RECT 623.400 805.350 624.600 806.400 ;
        RECT 629.400 805.350 630.600 807.600 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 626.400 801.000 627.600 802.650 ;
        RECT 625.950 796.950 628.050 801.000 ;
        RECT 632.400 800.400 633.600 802.650 ;
        RECT 616.950 766.950 619.050 769.050 ;
        RECT 613.950 760.950 616.050 763.050 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 622.950 762.000 625.050 766.050 ;
        RECT 617.400 760.350 618.600 761.100 ;
        RECT 623.400 760.350 624.600 762.000 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 625.950 757.950 628.050 760.050 ;
        RECT 613.950 751.950 616.050 757.050 ;
        RECT 620.400 756.900 621.600 757.650 ;
        RECT 619.950 754.800 622.050 756.900 ;
        RECT 626.400 755.400 627.600 757.650 ;
        RECT 619.950 748.950 622.050 751.050 ;
        RECT 610.950 742.950 613.050 745.050 ;
        RECT 616.950 739.950 619.050 742.050 ;
        RECT 617.400 733.050 618.450 739.950 ;
        RECT 616.950 730.950 619.050 733.050 ;
        RECT 607.950 728.100 610.050 730.200 ;
        RECT 608.400 727.350 609.600 728.100 ;
        RECT 620.400 727.200 621.450 748.950 ;
        RECT 626.400 747.450 627.450 755.400 ;
        RECT 628.950 754.950 631.050 757.050 ;
        RECT 623.400 747.000 627.450 747.450 ;
        RECT 622.950 746.400 627.450 747.000 ;
        RECT 622.950 742.950 625.050 746.400 ;
        RECT 629.400 744.450 630.450 754.950 ;
        RECT 626.400 743.400 630.450 744.450 ;
        RECT 608.400 724.950 610.500 727.050 ;
        RECT 613.800 724.950 615.900 727.050 ;
        RECT 619.950 725.100 622.050 727.200 ;
        RECT 614.400 722.400 615.600 724.650 ;
        RECT 620.400 724.350 621.600 725.100 ;
        RECT 614.400 706.050 615.450 722.400 ;
        RECT 620.100 721.950 622.200 724.050 ;
        RECT 613.950 703.950 616.050 706.050 ;
        RECT 626.400 697.050 627.450 743.400 ;
        RECT 628.950 739.950 631.050 742.050 ;
        RECT 629.400 726.600 630.450 739.950 ;
        RECT 632.400 736.050 633.450 800.400 ;
        RECT 638.400 796.050 639.450 838.950 ;
        RECT 641.400 833.400 642.900 852.300 ;
        RECT 645.300 846.300 646.500 852.300 ;
        RECT 644.400 844.200 646.500 846.300 ;
        RECT 641.400 831.300 643.500 833.400 ;
        RECT 642.300 827.700 643.500 831.300 ;
        RECT 645.300 827.700 646.500 844.200 ;
        RECT 647.700 849.300 649.800 851.400 ;
        RECT 647.700 827.700 648.900 849.300 ;
        RECT 656.400 847.800 658.500 849.900 ;
        RECT 661.800 849.300 663.900 851.400 ;
        RECT 656.400 841.200 657.300 847.800 ;
        RECT 662.100 842.100 663.300 849.300 ;
        RECT 664.800 847.500 666.300 852.300 ;
        RECT 667.200 849.300 669.300 854.400 ;
        RECT 664.800 845.400 666.900 847.500 ;
        RECT 652.950 837.000 655.050 841.050 ;
        RECT 656.400 839.100 658.500 841.200 ;
        RECT 661.800 840.000 663.900 842.100 ;
        RECT 653.400 835.350 654.600 837.000 ;
        RECT 652.800 832.950 654.900 835.050 ;
        RECT 656.400 828.600 657.300 839.100 ;
        RECT 659.100 832.500 661.200 834.600 ;
        RECT 641.700 825.600 643.800 827.700 ;
        RECT 644.700 825.600 646.800 827.700 ;
        RECT 647.700 825.600 649.800 827.700 ;
        RECT 655.800 826.500 657.900 828.600 ;
        RECT 662.100 827.700 663.300 840.000 ;
        RECT 664.800 827.700 666.300 845.400 ;
        RECT 668.100 827.700 669.300 849.300 ;
        RECT 661.200 825.600 663.300 827.700 ;
        RECT 664.200 825.600 666.300 827.700 ;
        RECT 667.200 825.600 669.300 827.700 ;
        RECT 670.200 852.300 672.300 854.400 ;
        RECT 670.200 847.500 671.700 852.300 ;
        RECT 670.200 845.400 672.300 847.500 ;
        RECT 670.200 827.700 671.700 845.400 ;
        RECT 670.200 825.600 672.300 827.700 ;
        RECT 674.400 823.050 675.450 859.950 ;
        RECT 679.800 838.950 681.900 841.050 ;
        RECT 680.400 836.400 681.600 838.650 ;
        RECT 680.400 823.050 681.450 836.400 ;
        RECT 658.950 820.950 661.050 823.050 ;
        RECT 673.950 820.950 676.050 823.050 ;
        RECT 679.950 820.950 682.050 823.050 ;
        RECT 659.400 817.050 660.450 820.950 ;
        RECT 658.950 814.950 661.050 817.050 ;
        RECT 649.950 811.950 652.050 814.050 ;
        RECT 642.000 807.450 646.050 808.050 ;
        RECT 641.400 805.950 646.050 807.450 ;
        RECT 650.400 807.600 651.450 811.950 ;
        RECT 637.950 793.950 640.050 796.050 ;
        RECT 641.400 766.050 642.450 805.950 ;
        RECT 650.400 805.350 651.600 807.600 ;
        RECT 655.950 805.950 658.050 811.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 652.950 802.950 655.050 805.050 ;
        RECT 647.400 801.000 648.600 802.650 ;
        RECT 653.400 801.900 654.600 802.650 ;
        RECT 659.400 801.900 660.450 814.950 ;
        RECT 661.950 811.950 664.050 814.050 ;
        RECT 673.950 811.950 676.050 814.050 ;
        RECT 662.400 808.050 663.450 811.950 ;
        RECT 661.950 805.950 664.050 808.050 ;
        RECT 667.950 806.100 670.050 808.200 ;
        RECT 674.400 807.600 675.450 811.950 ;
        RECT 668.400 805.350 669.600 806.100 ;
        RECT 674.400 805.350 675.600 807.600 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 646.950 796.950 649.050 801.000 ;
        RECT 652.950 799.800 655.050 801.900 ;
        RECT 658.800 799.800 660.900 801.900 ;
        RECT 661.950 799.950 664.050 802.050 ;
        RECT 665.400 800.400 666.600 802.650 ;
        RECT 671.400 800.400 672.600 802.650 ;
        RECT 677.400 801.900 678.600 802.650 ;
        RECT 662.400 790.050 663.450 799.950 ;
        RECT 665.400 790.050 666.450 800.400 ;
        RECT 671.400 796.050 672.450 800.400 ;
        RECT 676.950 799.800 679.050 801.900 ;
        RECT 679.950 796.950 682.050 799.050 ;
        RECT 670.950 793.950 673.050 796.050 ;
        RECT 661.800 787.950 663.900 790.050 ;
        RECT 664.950 787.950 667.050 790.050 ;
        RECT 643.950 775.950 646.050 778.050 ;
        RECT 661.950 775.950 664.050 778.050 ;
        RECT 640.950 763.950 643.050 766.050 ;
        RECT 644.400 763.200 645.450 775.950 ;
        RECT 649.950 769.950 652.050 772.050 ;
        RECT 634.950 762.600 639.000 763.050 ;
        RECT 634.950 760.950 639.600 762.600 ;
        RECT 643.950 761.100 646.050 763.200 ;
        RECT 638.400 760.350 639.600 760.950 ;
        RECT 644.400 760.350 645.600 761.100 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 634.950 754.950 637.050 757.050 ;
        RECT 641.400 756.900 642.600 757.650 ;
        RECT 635.400 751.050 636.450 754.950 ;
        RECT 640.950 754.800 643.050 756.900 ;
        RECT 634.950 748.950 637.050 751.050 ;
        RECT 650.400 742.050 651.450 769.950 ;
        RECT 652.950 763.950 655.050 766.050 ;
        RECT 653.400 757.050 654.450 763.950 ;
        RECT 662.400 762.600 663.450 775.950 ;
        RECT 662.400 760.350 663.600 762.600 ;
        RECT 667.950 762.000 670.050 766.050 ;
        RECT 680.400 763.050 681.450 796.950 ;
        RECT 683.400 766.050 684.450 868.950 ;
        RECT 686.400 844.050 687.450 874.950 ;
        RECT 695.400 871.050 696.450 916.950 ;
        RECT 697.950 913.800 700.050 915.900 ;
        RECT 707.400 913.950 709.500 916.050 ;
        RECT 712.800 913.950 714.900 916.050 ;
        RECT 719.400 915.900 720.600 916.650 ;
        RECT 718.950 913.800 721.050 915.900 ;
        RECT 728.400 914.400 729.600 916.650 ;
        RECT 698.400 886.200 699.450 913.800 ;
        RECT 707.400 912.000 708.600 913.650 ;
        RECT 706.950 907.950 709.050 912.000 ;
        RECT 718.950 901.950 721.050 904.050 ;
        RECT 700.950 898.950 703.050 901.050 ;
        RECT 697.950 884.100 700.050 886.200 ;
        RECT 694.950 868.950 697.050 871.050 ;
        RECT 694.950 862.950 697.050 865.050 ;
        RECT 695.400 853.050 696.450 862.950 ;
        RECT 694.950 850.950 697.050 853.050 ;
        RECT 685.950 841.950 688.050 844.050 ;
        RECT 694.950 841.950 697.050 847.050 ;
        RECT 698.400 841.200 699.450 884.100 ;
        RECT 701.400 850.050 702.450 898.950 ;
        RECT 709.950 889.950 712.050 892.050 ;
        RECT 710.400 885.600 711.450 889.950 ;
        RECT 710.400 883.350 711.600 885.600 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 712.950 880.950 715.050 883.050 ;
        RECT 707.400 878.400 708.600 880.650 ;
        RECT 713.400 879.900 714.600 880.650 ;
        RECT 719.400 879.900 720.450 901.950 ;
        RECT 728.400 901.050 729.450 914.400 ;
        RECT 738.300 905.700 739.800 923.400 ;
        RECT 737.700 903.600 739.800 905.700 ;
        RECT 740.700 927.300 742.800 932.400 ;
        RECT 743.700 930.300 745.800 932.400 ;
        RECT 762.600 930.300 764.700 932.400 ;
        RECT 765.600 930.300 768.600 932.400 ;
        RECT 740.700 905.700 741.900 927.300 ;
        RECT 743.700 925.500 745.200 930.300 ;
        RECT 746.100 927.300 748.200 929.400 ;
        RECT 743.100 923.400 745.200 925.500 ;
        RECT 743.700 905.700 745.200 923.400 ;
        RECT 746.700 920.100 747.900 927.300 ;
        RECT 751.500 925.800 753.600 927.900 ;
        RECT 760.200 927.300 762.300 929.400 ;
        RECT 746.100 918.000 748.200 920.100 ;
        RECT 752.700 919.200 753.600 925.800 ;
        RECT 754.950 922.800 757.050 924.900 ;
        RECT 746.700 905.700 747.900 918.000 ;
        RECT 751.500 917.100 753.600 919.200 ;
        RECT 748.800 910.500 750.900 912.600 ;
        RECT 752.700 906.600 753.600 917.100 ;
        RECT 755.400 915.600 756.450 922.800 ;
        RECT 755.400 913.350 756.600 915.600 ;
        RECT 755.100 910.950 757.200 913.050 ;
        RECT 740.700 903.600 742.800 905.700 ;
        RECT 743.700 903.600 745.800 905.700 ;
        RECT 746.700 903.600 748.800 905.700 ;
        RECT 752.100 904.500 754.200 906.600 ;
        RECT 761.100 905.700 762.300 927.300 ;
        RECT 763.500 924.300 764.700 930.300 ;
        RECT 763.500 922.200 765.600 924.300 ;
        RECT 763.500 905.700 764.700 922.200 ;
        RECT 767.100 911.400 768.600 930.300 ;
        RECT 793.950 922.950 796.050 925.050 ;
        RECT 898.950 922.950 901.050 925.050 ;
        RECT 922.950 922.950 925.050 925.050 ;
        RECT 779.400 921.450 780.600 921.600 ;
        RECT 779.400 920.400 786.450 921.450 ;
        RECT 779.400 919.350 780.600 920.400 ;
        RECT 773.100 916.950 775.200 919.050 ;
        RECT 779.100 916.950 781.200 919.050 ;
        RECT 766.500 909.300 768.600 911.400 ;
        RECT 766.500 905.700 767.700 909.300 ;
        RECT 760.200 903.600 762.300 905.700 ;
        RECT 763.200 903.600 765.300 905.700 ;
        RECT 766.200 903.600 768.300 905.700 ;
        RECT 724.950 899.400 729.450 901.050 ;
        RECT 724.950 898.950 729.000 899.400 ;
        RECT 727.950 895.950 730.050 898.050 ;
        RECT 728.400 885.600 729.450 895.950 ;
        RECT 733.950 892.950 736.050 895.050 ;
        RECT 745.950 892.950 748.050 895.050 ;
        RECT 734.400 885.600 735.450 892.950 ;
        RECT 728.400 883.350 729.600 885.600 ;
        RECT 734.400 883.350 735.600 885.600 ;
        RECT 742.950 883.950 745.050 886.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 733.950 880.950 736.050 883.050 ;
        RECT 736.950 880.950 739.050 883.050 ;
        RECT 707.400 871.050 708.450 878.400 ;
        RECT 712.950 877.800 715.050 879.900 ;
        RECT 718.950 877.800 721.050 879.900 ;
        RECT 725.400 879.450 726.600 880.650 ;
        RECT 722.400 878.400 726.600 879.450 ;
        RECT 731.400 878.400 732.600 880.650 ;
        RECT 737.400 879.450 738.600 880.650 ;
        RECT 743.400 879.450 744.450 883.950 ;
        RECT 746.400 879.900 747.450 892.950 ;
        RECT 760.950 889.950 763.050 892.050 ;
        RECT 775.950 889.950 778.050 892.050 ;
        RECT 754.950 884.100 757.050 886.200 ;
        RECT 761.400 885.600 762.450 889.950 ;
        RECT 776.400 885.600 777.450 889.950 ;
        RECT 755.400 883.350 756.600 884.100 ;
        RECT 761.400 883.350 762.600 885.600 ;
        RECT 776.400 883.350 777.600 885.600 ;
        RECT 781.950 884.100 784.050 886.200 ;
        RECT 785.400 886.050 786.450 920.400 ;
        RECT 794.400 918.600 795.450 922.950 ;
        RECT 794.400 916.350 795.600 918.600 ;
        RECT 802.950 917.100 805.050 919.200 ;
        RECT 803.400 916.350 804.600 917.100 ;
        RECT 805.950 916.950 808.050 919.050 ;
        RECT 808.950 917.100 811.050 919.200 ;
        RECT 811.950 918.600 816.000 919.050 ;
        RECT 794.100 913.950 796.200 916.050 ;
        RECT 799.500 913.950 801.600 916.050 ;
        RECT 802.800 913.950 804.900 916.050 ;
        RECT 800.400 911.400 801.600 913.650 ;
        RECT 800.400 909.450 801.450 911.400 ;
        RECT 800.400 908.400 804.450 909.450 ;
        RECT 803.400 901.050 804.450 908.400 ;
        RECT 806.400 906.450 807.450 916.950 ;
        RECT 809.400 913.050 810.450 917.100 ;
        RECT 811.950 916.950 816.600 918.600 ;
        RECT 820.950 917.100 823.050 919.200 ;
        RECT 832.950 917.100 835.050 919.200 ;
        RECT 838.950 917.100 841.050 919.200 ;
        RECT 865.950 918.000 868.050 922.050 ;
        RECT 871.950 919.950 874.050 922.050 ;
        RECT 877.950 921.450 882.000 922.050 ;
        RECT 877.950 919.950 882.450 921.450 ;
        RECT 889.950 919.950 892.050 922.050 ;
        RECT 815.400 916.350 816.600 916.950 ;
        RECT 821.400 916.350 822.600 917.100 ;
        RECT 814.950 913.950 817.050 916.050 ;
        RECT 817.950 913.950 820.050 916.050 ;
        RECT 820.950 913.950 823.050 916.050 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 808.950 910.950 811.050 913.050 ;
        RECT 818.400 912.900 819.600 913.650 ;
        RECT 817.950 910.800 820.050 912.900 ;
        RECT 824.400 911.400 825.600 913.650 ;
        RECT 806.400 905.400 810.450 906.450 ;
        RECT 802.950 898.950 805.050 901.050 ;
        RECT 787.950 889.950 790.050 892.050 ;
        RECT 782.400 883.350 783.600 884.100 ;
        RECT 784.950 883.950 787.050 886.050 ;
        RECT 751.950 880.950 754.050 883.050 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 757.950 880.950 760.050 883.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 778.950 880.950 781.050 883.050 ;
        RECT 781.950 880.950 784.050 883.050 ;
        RECT 737.400 878.400 744.450 879.450 ;
        RECT 706.950 868.950 709.050 871.050 ;
        RECT 718.950 853.950 721.050 856.050 ;
        RECT 700.950 847.950 703.050 850.050 ;
        RECT 719.400 844.050 720.450 853.950 ;
        RECT 700.950 841.950 703.050 844.050 ;
        RECT 688.800 838.950 690.900 841.050 ;
        RECT 697.950 839.100 700.050 841.200 ;
        RECT 689.400 838.050 690.600 838.650 ;
        RECT 685.950 836.400 690.600 838.050 ;
        RECT 685.950 835.950 690.450 836.400 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 689.400 828.450 690.450 835.950 ;
        RECT 692.400 832.050 693.450 835.950 ;
        RECT 691.950 829.950 694.050 832.050 ;
        RECT 689.400 827.400 693.450 828.450 ;
        RECT 692.400 807.600 693.450 827.400 ;
        RECT 692.400 805.350 693.600 807.600 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 689.400 801.900 690.600 802.650 ;
        RECT 688.950 799.800 691.050 801.900 ;
        RECT 698.400 799.050 699.450 839.100 ;
        RECT 701.400 801.450 702.450 841.950 ;
        RECT 706.950 840.000 709.050 844.050 ;
        RECT 718.950 841.950 721.050 844.050 ;
        RECT 707.400 838.350 708.600 840.000 ;
        RECT 712.950 839.100 715.050 841.200 ;
        RECT 713.400 838.350 714.600 839.100 ;
        RECT 706.950 835.950 709.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 710.400 834.900 711.600 835.650 ;
        RECT 709.950 832.800 712.050 834.900 ;
        RECT 712.950 820.950 715.050 823.050 ;
        RECT 709.950 811.950 712.050 814.050 ;
        RECT 710.400 808.200 711.450 811.950 ;
        RECT 709.950 806.100 712.050 808.200 ;
        RECT 710.400 805.350 711.600 806.100 ;
        RECT 704.400 802.950 706.500 805.050 ;
        RECT 709.500 802.950 711.600 805.050 ;
        RECT 704.400 801.450 705.600 802.650 ;
        RECT 701.400 800.400 705.600 801.450 ;
        RECT 713.400 799.050 714.450 820.950 ;
        RECT 697.950 796.950 700.050 799.050 ;
        RECT 703.950 796.950 706.050 799.050 ;
        RECT 712.950 796.950 715.050 799.050 ;
        RECT 697.950 790.950 700.050 793.050 ;
        RECT 691.950 781.950 694.050 784.050 ;
        RECT 682.950 763.950 685.050 766.050 ;
        RECT 688.950 763.950 691.050 766.050 ;
        RECT 668.400 760.350 669.600 762.000 ;
        RECT 679.950 760.950 682.050 763.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 685.800 757.950 687.900 760.050 ;
        RECT 652.950 754.950 655.050 757.050 ;
        RECT 659.400 755.400 660.600 757.650 ;
        RECT 665.400 755.400 666.600 757.650 ;
        RECT 659.400 742.050 660.450 755.400 ;
        RECT 661.950 751.950 664.050 754.050 ;
        RECT 662.400 745.050 663.450 751.950 ;
        RECT 665.400 751.050 666.450 755.400 ;
        RECT 664.950 748.950 667.050 751.050 ;
        RECT 670.950 748.950 673.050 751.050 ;
        RECT 661.950 742.950 664.050 745.050 ;
        RECT 634.950 739.950 637.050 742.050 ;
        RECT 649.950 739.950 652.050 742.050 ;
        RECT 658.950 739.950 661.050 742.050 ;
        RECT 631.950 733.950 634.050 736.050 ;
        RECT 629.400 724.350 630.600 726.600 ;
        RECT 629.100 721.950 631.200 724.050 ;
        RECT 635.400 712.050 636.450 739.950 ;
        RECT 638.700 735.300 640.800 737.400 ;
        RECT 639.300 717.600 640.800 735.300 ;
        RECT 638.700 715.500 640.800 717.600 ;
        RECT 634.950 709.950 637.050 712.050 ;
        RECT 639.300 710.700 640.800 715.500 ;
        RECT 638.700 708.600 640.800 710.700 ;
        RECT 641.700 735.300 643.800 737.400 ;
        RECT 644.700 735.300 646.800 737.400 ;
        RECT 647.700 735.300 649.800 737.400 ;
        RECT 641.700 713.700 642.900 735.300 ;
        RECT 644.700 717.600 646.200 735.300 ;
        RECT 647.700 723.000 648.900 735.300 ;
        RECT 653.100 734.400 655.200 736.500 ;
        RECT 661.200 735.300 663.300 737.400 ;
        RECT 664.200 735.300 666.300 737.400 ;
        RECT 667.200 735.300 669.300 737.400 ;
        RECT 649.800 728.400 651.900 730.500 ;
        RECT 653.700 723.900 654.600 734.400 ;
        RECT 656.100 727.950 658.200 730.050 ;
        RECT 656.400 727.050 657.600 727.650 ;
        RECT 656.400 725.400 661.050 727.050 ;
        RECT 657.000 724.950 661.050 725.400 ;
        RECT 647.100 720.900 649.200 723.000 ;
        RECT 652.500 721.800 654.600 723.900 ;
        RECT 655.950 721.950 658.050 724.050 ;
        RECT 644.100 715.500 646.200 717.600 ;
        RECT 641.700 708.600 643.800 713.700 ;
        RECT 644.700 710.700 646.200 715.500 ;
        RECT 647.700 713.700 648.900 720.900 ;
        RECT 653.700 715.200 654.600 721.800 ;
        RECT 647.100 711.600 649.200 713.700 ;
        RECT 652.500 713.100 654.600 715.200 ;
        RECT 644.700 708.600 646.800 710.700 ;
        RECT 634.950 703.950 637.050 706.050 ;
        RECT 607.950 694.950 610.050 697.050 ;
        RECT 625.950 694.950 628.050 697.050 ;
        RECT 604.950 685.950 607.050 688.050 ;
        RECT 590.400 682.350 591.600 683.100 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 587.400 678.900 588.600 679.650 ;
        RECT 596.400 679.050 597.450 683.100 ;
        RECT 598.950 682.950 601.050 685.050 ;
        RECT 601.950 682.950 604.050 685.050 ;
        RECT 608.400 684.600 609.450 694.950 ;
        RECT 580.950 676.800 583.050 678.900 ;
        RECT 586.950 676.800 589.050 678.900 ;
        RECT 595.950 676.950 598.050 679.050 ;
        RECT 595.950 673.800 598.050 675.900 ;
        RECT 577.950 670.950 580.050 673.050 ;
        RECT 586.950 670.950 589.050 673.050 ;
        RECT 565.950 664.950 568.050 667.050 ;
        RECT 544.950 661.950 547.050 664.050 ;
        RECT 562.950 661.950 565.050 664.050 ;
        RECT 541.950 652.950 544.050 655.050 ;
        RECT 542.400 649.050 543.450 652.950 ;
        RECT 539.400 646.350 540.600 648.600 ;
        RECT 541.800 646.950 543.900 649.050 ;
        RECT 539.100 643.950 541.200 646.050 ;
        RECT 545.400 643.050 546.450 661.950 ;
        RECT 548.700 657.300 550.800 659.400 ;
        RECT 541.800 640.950 543.900 643.050 ;
        RECT 544.950 640.950 547.050 643.050 ;
        RECT 535.950 634.950 538.050 637.050 ;
        RECT 542.400 622.050 543.450 640.950 ;
        RECT 549.300 639.600 550.800 657.300 ;
        RECT 548.700 637.500 550.800 639.600 ;
        RECT 549.300 632.700 550.800 637.500 ;
        RECT 548.700 630.600 550.800 632.700 ;
        RECT 551.700 657.300 553.800 659.400 ;
        RECT 554.700 657.300 556.800 659.400 ;
        RECT 557.700 657.300 559.800 659.400 ;
        RECT 551.700 635.700 552.900 657.300 ;
        RECT 554.700 639.600 556.200 657.300 ;
        RECT 557.700 645.000 558.900 657.300 ;
        RECT 563.100 656.400 565.200 658.500 ;
        RECT 571.200 657.300 573.300 659.400 ;
        RECT 574.200 657.300 576.300 659.400 ;
        RECT 577.200 657.300 579.300 659.400 ;
        RECT 559.800 650.400 561.900 652.500 ;
        RECT 563.700 645.900 564.600 656.400 ;
        RECT 566.100 649.950 568.200 652.050 ;
        RECT 557.100 642.900 559.200 645.000 ;
        RECT 562.500 643.800 564.600 645.900 ;
        RECT 554.100 637.500 556.200 639.600 ;
        RECT 551.700 630.600 553.800 635.700 ;
        RECT 554.700 632.700 556.200 637.500 ;
        RECT 557.700 635.700 558.900 642.900 ;
        RECT 563.700 637.200 564.600 643.800 ;
        RECT 557.100 633.600 559.200 635.700 ;
        RECT 562.500 635.100 564.600 637.200 ;
        RECT 566.400 647.400 567.600 649.650 ;
        RECT 566.400 637.050 567.450 647.400 ;
        RECT 568.950 646.950 571.050 649.050 ;
        RECT 569.400 640.050 570.450 646.950 ;
        RECT 568.950 637.950 571.050 640.050 ;
        RECT 565.950 634.950 568.050 637.050 ;
        RECT 572.100 635.700 573.300 657.300 ;
        RECT 571.200 633.600 573.300 635.700 ;
        RECT 574.500 640.800 575.700 657.300 ;
        RECT 577.500 653.700 578.700 657.300 ;
        RECT 577.500 651.600 579.600 653.700 ;
        RECT 574.500 638.700 576.600 640.800 ;
        RECT 574.500 632.700 575.700 638.700 ;
        RECT 578.100 632.700 579.600 651.600 ;
        RECT 587.400 649.050 588.450 670.950 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 584.100 643.950 586.200 646.050 ;
        RECT 590.100 643.950 592.200 646.050 ;
        RECT 590.400 642.900 591.600 643.650 ;
        RECT 596.400 643.050 597.450 673.800 ;
        RECT 599.400 673.050 600.450 682.950 ;
        RECT 608.400 682.350 609.600 684.600 ;
        RECT 613.950 684.000 616.050 688.050 ;
        RECT 625.950 685.950 628.050 688.050 ;
        RECT 614.400 682.350 615.600 684.000 ;
        RECT 620.100 682.950 622.200 685.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 607.950 679.950 610.050 682.050 ;
        RECT 610.950 679.950 613.050 682.050 ;
        RECT 613.950 679.950 616.050 682.050 ;
        RECT 620.400 680.400 621.600 682.650 ;
        RECT 601.950 676.950 604.050 679.050 ;
        RECT 605.400 678.900 606.600 679.650 ;
        RECT 598.950 670.950 601.050 673.050 ;
        RECT 602.400 669.450 603.450 676.950 ;
        RECT 604.950 676.800 607.050 678.900 ;
        RECT 611.400 677.400 612.600 679.650 ;
        RECT 605.400 675.450 606.450 676.800 ;
        RECT 605.400 674.400 609.450 675.450 ;
        RECT 599.400 668.400 603.450 669.450 ;
        RECT 599.400 649.050 600.450 668.400 ;
        RECT 601.950 661.950 604.050 664.050 ;
        RECT 598.950 646.950 601.050 649.050 ;
        RECT 602.400 646.050 603.450 661.950 ;
        RECT 608.400 651.600 609.450 674.400 ;
        RECT 611.400 673.050 612.450 677.400 ;
        RECT 610.800 670.950 612.900 673.050 ;
        RECT 613.950 670.950 616.050 673.050 ;
        RECT 614.400 667.050 615.450 670.950 ;
        RECT 620.400 667.050 621.450 680.400 ;
        RECT 613.950 664.950 616.050 667.050 ;
        RECT 619.950 664.950 622.050 667.050 ;
        RECT 626.400 664.050 627.450 685.950 ;
        RECT 629.100 682.950 631.200 685.050 ;
        RECT 629.400 680.400 630.600 682.650 ;
        RECT 629.400 676.050 630.450 680.400 ;
        RECT 628.950 673.950 631.050 676.050 ;
        RECT 625.950 661.950 628.050 664.050 ;
        RECT 635.400 658.050 636.450 703.950 ;
        RECT 638.700 696.300 640.800 698.400 ;
        RECT 639.300 691.500 640.800 696.300 ;
        RECT 638.700 689.400 640.800 691.500 ;
        RECT 639.300 671.700 640.800 689.400 ;
        RECT 638.700 669.600 640.800 671.700 ;
        RECT 641.700 693.300 643.800 698.400 ;
        RECT 644.700 696.300 646.800 698.400 ;
        RECT 656.400 697.050 657.450 721.950 ;
        RECT 662.100 713.700 663.300 735.300 ;
        RECT 661.200 711.600 663.300 713.700 ;
        RECT 664.500 718.800 665.700 735.300 ;
        RECT 667.500 731.700 668.700 735.300 ;
        RECT 667.500 729.600 669.600 731.700 ;
        RECT 664.500 716.700 666.600 718.800 ;
        RECT 664.500 710.700 665.700 716.700 ;
        RECT 668.100 710.700 669.600 729.600 ;
        RECT 671.400 727.050 672.450 748.950 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 674.100 721.950 676.200 724.050 ;
        RECT 680.100 721.950 682.200 724.050 ;
        RECT 680.400 719.400 681.600 721.650 ;
        RECT 663.600 708.600 665.700 710.700 ;
        RECT 666.600 708.600 669.600 710.700 ;
        RECT 670.950 709.950 673.050 712.050 ;
        RECT 641.700 671.700 642.900 693.300 ;
        RECT 644.700 691.500 646.200 696.300 ;
        RECT 647.100 693.300 649.200 695.400 ;
        RECT 655.950 694.950 658.050 697.050 ;
        RECT 663.600 696.300 665.700 698.400 ;
        RECT 666.600 696.300 669.600 698.400 ;
        RECT 644.100 689.400 646.200 691.500 ;
        RECT 644.700 671.700 646.200 689.400 ;
        RECT 647.700 686.100 648.900 693.300 ;
        RECT 652.500 691.800 654.600 693.900 ;
        RECT 661.200 693.300 663.300 695.400 ;
        RECT 647.100 684.000 649.200 686.100 ;
        RECT 653.700 685.200 654.600 691.800 ;
        RECT 647.700 671.700 648.900 684.000 ;
        RECT 652.500 683.100 654.600 685.200 ;
        RECT 649.800 676.500 651.900 678.600 ;
        RECT 653.700 672.600 654.600 683.100 ;
        RECT 655.950 681.000 658.050 685.050 ;
        RECT 656.400 679.350 657.600 681.000 ;
        RECT 656.100 676.950 658.200 679.050 ;
        RECT 641.700 669.600 643.800 671.700 ;
        RECT 644.700 669.600 646.800 671.700 ;
        RECT 647.700 669.600 649.800 671.700 ;
        RECT 653.100 670.500 655.200 672.600 ;
        RECT 662.100 671.700 663.300 693.300 ;
        RECT 664.500 690.300 665.700 696.300 ;
        RECT 664.500 688.200 666.600 690.300 ;
        RECT 664.500 671.700 665.700 688.200 ;
        RECT 668.100 677.400 669.600 696.300 ;
        RECT 667.500 675.300 669.600 677.400 ;
        RECT 671.400 676.050 672.450 709.950 ;
        RECT 680.400 706.050 681.450 719.400 ;
        RECT 689.400 712.050 690.450 763.950 ;
        RECT 692.400 745.050 693.450 781.950 ;
        RECT 698.400 751.050 699.450 790.950 ;
        RECT 704.400 772.050 705.450 796.950 ;
        RECT 719.400 781.050 720.450 841.950 ;
        RECT 722.400 808.050 723.450 878.400 ;
        RECT 731.400 871.050 732.450 878.400 ;
        RECT 745.950 877.800 748.050 879.900 ;
        RECT 752.400 878.400 753.600 880.650 ;
        RECT 758.400 878.400 759.600 880.650 ;
        RECT 773.400 879.900 774.600 880.650 ;
        RECT 752.400 871.050 753.450 878.400 ;
        RECT 730.950 868.950 733.050 871.050 ;
        RECT 751.950 868.950 754.050 871.050 ;
        RECT 758.400 868.050 759.450 878.400 ;
        RECT 772.950 877.800 775.050 879.900 ;
        RECT 779.400 878.400 780.600 880.650 ;
        RECT 788.400 880.050 789.450 889.950 ;
        RECT 805.950 884.100 808.050 886.200 ;
        RECT 796.950 880.950 799.050 883.050 ;
        RECT 799.950 880.950 802.050 883.050 ;
        RECT 757.950 865.950 760.050 868.050 ;
        RECT 751.950 853.950 754.050 856.050 ;
        RECT 772.950 853.950 775.050 856.050 ;
        RECT 724.950 847.950 727.050 850.050 ;
        RECT 725.400 820.050 726.450 847.950 ;
        RECT 739.950 839.100 742.050 841.200 ;
        RECT 752.400 840.600 753.450 853.950 ;
        RECT 760.950 850.950 763.050 853.050 ;
        RECT 728.100 835.950 730.200 838.050 ;
        RECT 733.500 835.950 735.600 838.050 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 734.400 833.400 735.600 835.650 ;
        RECT 727.950 826.950 730.050 829.050 ;
        RECT 724.950 817.950 727.050 820.050 ;
        RECT 721.950 805.950 724.050 808.050 ;
        RECT 724.800 802.950 726.900 805.050 ;
        RECT 718.950 778.950 721.050 781.050 ;
        RECT 728.400 778.050 729.450 826.950 ;
        RECT 734.400 811.050 735.450 833.400 ;
        RECT 737.400 826.050 738.450 835.950 ;
        RECT 736.950 823.950 739.050 826.050 ;
        RECT 740.400 822.450 741.450 839.100 ;
        RECT 752.400 838.350 753.600 840.600 ;
        RECT 748.950 835.950 751.050 838.050 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 749.400 834.900 750.600 835.650 ;
        RECT 748.950 832.800 751.050 834.900 ;
        RECT 761.400 829.050 762.450 850.950 ;
        RECT 766.950 839.100 769.050 841.200 ;
        RECT 773.400 840.600 774.450 853.950 ;
        RECT 779.400 847.050 780.450 878.400 ;
        RECT 784.950 877.950 787.050 880.050 ;
        RECT 787.950 877.950 790.050 880.050 ;
        RECT 797.400 879.900 798.600 880.650 ;
        RECT 785.400 874.050 786.450 877.950 ;
        RECT 796.950 877.800 799.050 879.900 ;
        RECT 784.950 871.950 787.050 874.050 ;
        RECT 796.950 868.950 799.050 871.050 ;
        RECT 784.950 856.950 787.050 859.050 ;
        RECT 785.400 853.050 786.450 856.950 ;
        RECT 784.950 850.950 787.050 853.050 ;
        RECT 787.950 847.950 790.050 850.050 ;
        RECT 778.950 844.950 781.050 847.050 ;
        RECT 767.400 838.350 768.600 839.100 ;
        RECT 773.400 838.350 774.600 840.600 ;
        RECT 782.100 838.950 784.200 841.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 772.950 835.950 775.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 782.400 836.400 783.600 838.650 ;
        RECT 770.400 833.400 771.600 835.650 ;
        RECT 776.400 834.900 777.600 835.650 ;
        RECT 770.400 829.050 771.450 833.400 ;
        RECT 775.950 832.800 778.050 834.900 ;
        RECT 760.950 826.950 763.050 829.050 ;
        RECT 769.950 826.950 772.050 829.050 ;
        RECT 737.400 821.400 741.450 822.450 ;
        RECT 733.950 808.950 736.050 811.050 ;
        RECT 730.950 806.100 733.050 808.200 ;
        RECT 727.950 775.950 730.050 778.050 ;
        RECT 703.950 769.950 706.050 772.050 ;
        RECT 704.400 762.600 705.450 769.950 ;
        RECT 715.950 766.950 718.050 769.050 ;
        RECT 704.400 760.350 705.600 762.600 ;
        RECT 703.800 757.950 705.900 760.050 ;
        RECT 716.400 754.050 717.450 766.950 ;
        RECT 724.950 761.100 727.050 763.200 ;
        RECT 731.400 763.050 732.450 806.100 ;
        RECT 737.400 793.050 738.450 821.400 ;
        RECT 745.950 817.950 748.050 820.050 ;
        RECT 742.800 802.950 744.900 805.050 ;
        RECT 743.400 801.450 744.600 802.650 ;
        RECT 746.400 801.450 747.450 817.950 ;
        RECT 770.400 817.050 771.450 826.950 ;
        RECT 782.400 826.050 783.450 836.400 ;
        RECT 788.400 835.050 789.450 847.950 ;
        RECT 791.100 838.950 793.200 841.050 ;
        RECT 791.400 836.400 792.600 838.650 ;
        RECT 787.950 832.950 790.050 835.050 ;
        RECT 781.950 823.950 784.050 826.050 ;
        RECT 791.400 820.050 792.450 836.400 ;
        RECT 797.400 823.050 798.450 868.950 ;
        RECT 806.400 865.050 807.450 884.100 ;
        RECT 809.400 868.050 810.450 905.400 ;
        RECT 824.400 901.050 825.450 911.400 ;
        RECT 820.800 898.950 822.900 901.050 ;
        RECT 823.950 898.950 826.050 901.050 ;
        RECT 814.950 884.100 817.050 886.200 ;
        RECT 821.400 885.600 822.450 898.950 ;
        RECT 826.950 889.950 829.050 892.050 ;
        RECT 827.400 885.600 828.450 889.950 ;
        RECT 815.400 883.350 816.600 884.100 ;
        RECT 821.400 883.350 822.600 885.600 ;
        RECT 827.400 883.350 828.600 885.600 ;
        RECT 829.950 883.950 832.050 889.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 817.950 880.950 820.050 883.050 ;
        RECT 820.950 880.950 823.050 883.050 ;
        RECT 823.950 880.950 826.050 883.050 ;
        RECT 826.950 880.950 829.050 883.050 ;
        RECT 811.950 877.950 814.050 880.050 ;
        RECT 818.400 879.900 819.600 880.650 ;
        RECT 812.400 871.050 813.450 877.950 ;
        RECT 817.950 877.800 820.050 879.900 ;
        RECT 824.400 878.400 825.600 880.650 ;
        RECT 811.950 868.950 814.050 871.050 ;
        RECT 808.950 865.950 811.050 868.050 ;
        RECT 805.950 862.950 808.050 865.050 ;
        RECT 824.400 859.050 825.450 878.400 ;
        RECT 823.950 856.950 826.050 859.050 ;
        RECT 800.700 852.300 802.800 854.400 ;
        RECT 801.300 847.500 802.800 852.300 ;
        RECT 800.700 845.400 802.800 847.500 ;
        RECT 801.300 827.700 802.800 845.400 ;
        RECT 800.700 825.600 802.800 827.700 ;
        RECT 803.700 849.300 805.800 854.400 ;
        RECT 806.700 852.300 808.800 854.400 ;
        RECT 803.700 827.700 804.900 849.300 ;
        RECT 806.700 847.500 808.200 852.300 ;
        RECT 809.100 849.300 811.200 851.400 ;
        RECT 817.950 850.950 820.050 853.050 ;
        RECT 825.600 852.300 827.700 854.400 ;
        RECT 828.600 852.300 831.600 854.400 ;
        RECT 806.100 845.400 808.200 847.500 ;
        RECT 806.700 827.700 808.200 845.400 ;
        RECT 809.700 842.100 810.900 849.300 ;
        RECT 814.500 847.800 816.600 849.900 ;
        RECT 809.100 840.000 811.200 842.100 ;
        RECT 815.700 841.200 816.600 847.800 ;
        RECT 809.700 827.700 810.900 840.000 ;
        RECT 814.500 839.100 816.600 841.200 ;
        RECT 811.800 832.500 813.900 834.600 ;
        RECT 815.700 828.600 816.600 839.100 ;
        RECT 818.400 837.600 819.450 850.950 ;
        RECT 823.200 849.300 825.300 851.400 ;
        RECT 818.400 835.350 819.600 837.600 ;
        RECT 818.100 832.950 820.200 835.050 ;
        RECT 803.700 825.600 805.800 827.700 ;
        RECT 806.700 825.600 808.800 827.700 ;
        RECT 809.700 825.600 811.800 827.700 ;
        RECT 815.100 826.500 817.200 828.600 ;
        RECT 824.100 827.700 825.300 849.300 ;
        RECT 826.500 846.300 827.700 852.300 ;
        RECT 826.500 844.200 828.600 846.300 ;
        RECT 826.500 827.700 827.700 844.200 ;
        RECT 830.100 833.400 831.600 852.300 ;
        RECT 833.400 850.050 834.450 917.100 ;
        RECT 839.400 916.350 840.600 917.100 ;
        RECT 866.400 916.350 867.600 918.000 ;
        RECT 838.950 913.950 841.050 916.050 ;
        RECT 841.950 913.950 844.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 859.950 913.950 862.050 916.050 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 865.950 913.950 868.050 916.050 ;
        RECT 835.950 910.950 838.050 913.050 ;
        RECT 863.400 911.400 864.600 913.650 ;
        RECT 836.400 895.050 837.450 910.950 ;
        RECT 863.400 901.050 864.450 911.400 ;
        RECT 838.950 900.450 841.050 901.050 ;
        RECT 844.950 900.450 847.050 901.050 ;
        RECT 838.950 899.400 847.050 900.450 ;
        RECT 838.950 898.950 841.050 899.400 ;
        RECT 844.950 898.950 847.050 899.400 ;
        RECT 862.950 898.950 865.050 901.050 ;
        RECT 835.950 892.950 838.050 895.050 ;
        RECT 872.400 892.050 873.450 919.950 ;
        RECT 881.400 918.600 882.450 919.950 ;
        RECT 881.400 916.350 882.600 918.600 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 880.950 913.950 883.050 916.050 ;
        RECT 883.950 913.950 886.050 916.050 ;
        RECT 884.400 912.900 885.600 913.650 ;
        RECT 890.400 912.900 891.450 919.950 ;
        RECT 899.400 918.600 900.450 922.950 ;
        RECT 913.950 919.950 916.050 922.050 ;
        RECT 899.400 916.350 900.600 918.600 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 901.950 913.950 904.050 916.050 ;
        RECT 904.950 913.950 907.050 916.050 ;
        RECT 883.950 910.800 886.050 912.900 ;
        RECT 889.950 910.800 892.050 912.900 ;
        RECT 896.400 911.400 897.600 913.650 ;
        RECT 902.400 911.400 903.600 913.650 ;
        RECT 896.400 904.050 897.450 911.400 ;
        RECT 902.400 907.050 903.450 911.400 ;
        RECT 901.800 904.950 903.900 907.050 ;
        RECT 904.950 904.950 907.050 907.050 ;
        RECT 877.950 901.950 880.050 904.050 ;
        RECT 895.950 901.950 898.050 904.050 ;
        RECT 871.950 889.950 874.050 892.050 ;
        RECT 841.950 889.050 844.050 889.200 ;
        RECT 844.950 889.050 847.050 889.200 ;
        RECT 841.950 887.100 847.050 889.050 ;
        RECT 843.000 886.950 846.000 887.100 ;
        RECT 835.950 883.950 838.050 886.050 ;
        RECT 841.950 883.950 844.050 886.050 ;
        RECT 853.950 884.100 856.050 886.200 ;
        RECT 862.950 884.100 865.050 886.200 ;
        RECT 836.400 865.050 837.450 883.950 ;
        RECT 842.400 883.350 843.600 883.950 ;
        RECT 841.950 880.950 844.050 883.050 ;
        RECT 844.950 880.950 847.050 883.050 ;
        RECT 845.400 879.900 846.600 880.650 ;
        RECT 844.950 877.800 847.050 879.900 ;
        RECT 841.950 871.950 844.050 874.050 ;
        RECT 835.950 862.950 838.050 865.050 ;
        RECT 832.950 847.950 835.050 850.050 ;
        RECT 842.400 844.200 843.450 871.950 ;
        RECT 854.400 871.050 855.450 884.100 ;
        RECT 863.400 883.350 864.600 884.100 ;
        RECT 860.100 880.950 862.200 883.050 ;
        RECT 863.400 880.950 865.500 883.050 ;
        RECT 868.800 880.950 870.900 883.050 ;
        RECT 860.400 878.400 861.600 880.650 ;
        RECT 869.400 878.400 870.600 880.650 ;
        RECT 878.400 880.050 879.450 901.950 ;
        RECT 892.950 889.950 895.050 892.050 ;
        RECT 886.950 884.100 889.050 889.050 ;
        RECT 893.400 885.600 894.450 889.950 ;
        RECT 901.950 886.950 904.050 889.050 ;
        RECT 887.400 883.350 888.600 884.100 ;
        RECT 893.400 883.350 894.600 885.600 ;
        RECT 883.950 880.950 886.050 883.050 ;
        RECT 886.950 880.950 889.050 883.050 ;
        RECT 889.950 880.950 892.050 883.050 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 853.950 868.950 856.050 871.050 ;
        RECT 850.950 850.950 853.050 853.050 ;
        RECT 832.950 841.950 835.050 844.050 ;
        RECT 841.950 842.100 844.050 844.200 ;
        RECT 829.500 831.300 831.600 833.400 ;
        RECT 829.500 827.700 830.700 831.300 ;
        RECT 823.200 825.600 825.300 827.700 ;
        RECT 826.200 825.600 828.300 827.700 ;
        RECT 829.200 825.600 831.300 827.700 ;
        RECT 796.950 820.950 799.050 823.050 ;
        RECT 775.950 817.950 778.050 820.050 ;
        RECT 790.950 817.950 793.050 820.050 ;
        RECT 769.950 814.950 772.050 817.050 ;
        RECT 757.950 807.000 760.050 811.050 ;
        RECT 766.950 808.950 769.050 811.050 ;
        RECT 758.400 805.350 759.600 807.000 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 767.400 804.600 768.450 808.950 ;
        RECT 776.400 804.600 777.450 817.950 ;
        RECT 785.700 813.300 787.800 815.400 ;
        RECT 743.400 800.400 747.450 801.450 ;
        RECT 761.400 800.400 762.600 802.650 ;
        RECT 767.400 802.350 768.600 804.600 ;
        RECT 776.400 802.350 777.600 804.600 ;
        RECT 736.950 790.950 739.050 793.050 ;
        RECT 742.950 781.950 745.050 784.050 ;
        RECT 739.950 778.950 742.050 781.050 ;
        RECT 725.400 760.350 726.600 761.100 ;
        RECT 730.950 760.950 733.050 763.050 ;
        RECT 740.400 762.600 741.450 778.950 ;
        RECT 743.400 778.050 744.450 781.950 ;
        RECT 742.950 775.950 745.050 778.050 ;
        RECT 761.400 775.050 762.450 800.400 ;
        RECT 767.100 799.950 769.200 802.050 ;
        RECT 776.100 799.950 778.200 802.050 ;
        RECT 786.300 795.600 787.800 813.300 ;
        RECT 785.700 793.500 787.800 795.600 ;
        RECT 766.950 787.950 769.050 790.050 ;
        RECT 786.300 788.700 787.800 793.500 ;
        RECT 760.950 772.950 763.050 775.050 ;
        RECT 740.400 760.350 741.600 762.600 ;
        RECT 748.950 760.950 751.050 763.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 736.950 757.950 739.050 760.050 ;
        RECT 739.950 757.950 742.050 760.050 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 722.400 755.400 723.600 757.650 ;
        RECT 737.400 756.900 738.600 757.650 ;
        RECT 743.400 756.900 744.600 757.650 ;
        RECT 749.400 756.900 750.450 760.950 ;
        RECT 758.100 757.950 760.200 760.050 ;
        RECT 763.500 757.950 765.600 760.050 ;
        RECT 764.400 756.900 765.600 757.650 ;
        RECT 767.400 757.050 768.450 787.950 ;
        RECT 785.700 786.600 787.800 788.700 ;
        RECT 788.700 813.300 790.800 815.400 ;
        RECT 791.700 813.300 793.800 815.400 ;
        RECT 794.700 813.300 796.800 815.400 ;
        RECT 788.700 791.700 789.900 813.300 ;
        RECT 791.700 795.600 793.200 813.300 ;
        RECT 794.700 801.000 795.900 813.300 ;
        RECT 800.100 812.400 802.200 814.500 ;
        RECT 808.200 813.300 810.300 815.400 ;
        RECT 811.200 813.300 813.300 815.400 ;
        RECT 814.200 813.300 816.300 815.400 ;
        RECT 796.800 806.400 798.900 808.500 ;
        RECT 800.700 801.900 801.600 812.400 ;
        RECT 803.100 805.950 805.200 808.050 ;
        RECT 794.100 798.900 796.200 801.000 ;
        RECT 799.500 799.800 801.600 801.900 ;
        RECT 791.100 793.500 793.200 795.600 ;
        RECT 788.700 786.600 790.800 791.700 ;
        RECT 791.700 788.700 793.200 793.500 ;
        RECT 794.700 791.700 795.900 798.900 ;
        RECT 800.700 793.200 801.600 799.800 ;
        RECT 794.100 789.600 796.200 791.700 ;
        RECT 799.500 791.100 801.600 793.200 ;
        RECT 803.400 803.400 804.600 805.650 ;
        RECT 791.700 786.600 793.800 788.700 ;
        RECT 803.400 784.050 804.450 803.400 ;
        RECT 809.100 791.700 810.300 813.300 ;
        RECT 808.200 789.600 810.300 791.700 ;
        RECT 811.500 796.800 812.700 813.300 ;
        RECT 814.500 809.700 815.700 813.300 ;
        RECT 814.500 807.600 816.600 809.700 ;
        RECT 811.500 794.700 813.600 796.800 ;
        RECT 811.500 788.700 812.700 794.700 ;
        RECT 815.100 788.700 816.600 807.600 ;
        RECT 833.400 805.050 834.450 841.950 ;
        RECT 842.400 841.350 843.600 842.100 ;
        RECT 836.100 838.950 838.200 841.050 ;
        RECT 842.100 838.950 844.200 841.050 ;
        RECT 851.400 834.900 852.450 850.950 ;
        RECT 860.400 843.450 861.450 878.400 ;
        RECT 869.400 874.050 870.450 878.400 ;
        RECT 877.950 877.950 880.050 880.050 ;
        RECT 884.400 879.900 885.600 880.650 ;
        RECT 883.950 877.800 886.050 879.900 ;
        RECT 890.400 878.400 891.600 880.650 ;
        RECT 896.400 878.400 897.600 880.650 ;
        RECT 890.400 874.050 891.450 878.400 ;
        RECT 868.950 871.950 871.050 874.050 ;
        RECT 889.950 871.950 892.050 874.050 ;
        RECT 874.950 856.950 877.050 859.050 ;
        RECT 862.950 847.950 865.050 850.050 ;
        RECT 857.400 842.400 861.450 843.450 ;
        RECT 857.400 840.600 858.450 842.400 ;
        RECT 863.400 840.600 864.450 847.950 ;
        RECT 857.400 838.350 858.600 840.600 ;
        RECT 863.400 838.350 864.600 840.600 ;
        RECT 871.950 838.950 874.050 841.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 860.400 834.900 861.600 835.650 ;
        RECT 866.400 834.900 867.600 835.650 ;
        RECT 872.400 834.900 873.450 838.950 ;
        RECT 875.400 834.900 876.450 856.950 ;
        RECT 883.950 850.950 886.050 853.050 ;
        RECT 884.400 840.600 885.450 850.950 ;
        RECT 896.400 844.050 897.450 878.400 ;
        RECT 895.950 841.950 898.050 844.050 ;
        RECT 902.400 841.200 903.450 886.950 ;
        RECT 905.400 850.050 906.450 904.950 ;
        RECT 914.400 889.050 915.450 919.950 ;
        RECT 923.400 918.600 924.450 922.950 ;
        RECT 923.400 916.350 924.600 918.600 ;
        RECT 937.950 918.000 940.050 922.050 ;
        RECT 938.400 916.350 939.600 918.000 ;
        RECT 919.950 913.950 922.050 916.050 ;
        RECT 922.950 913.950 925.050 916.050 ;
        RECT 925.950 913.950 928.050 916.050 ;
        RECT 937.950 913.950 940.050 916.050 ;
        RECT 940.950 913.950 943.050 916.050 ;
        RECT 920.400 911.400 921.600 913.650 ;
        RECT 920.400 907.050 921.450 911.400 ;
        RECT 919.950 904.950 922.050 907.050 ;
        RECT 913.950 888.450 916.050 889.050 ;
        RECT 913.950 887.400 918.450 888.450 ;
        RECT 913.950 886.950 916.050 887.400 ;
        RECT 917.400 885.600 918.450 887.400 ;
        RECT 917.400 883.350 918.600 885.600 ;
        RECT 922.950 883.950 925.050 886.050 ;
        RECT 928.950 884.100 931.050 886.200 ;
        RECT 910.950 880.950 913.050 883.050 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 914.400 879.900 915.600 880.650 ;
        RECT 913.950 877.800 916.050 879.900 ;
        RECT 923.400 853.050 924.450 883.950 ;
        RECT 929.400 883.350 930.600 884.100 ;
        RECT 929.400 880.950 931.500 883.050 ;
        RECT 934.800 880.950 936.900 883.050 ;
        RECT 922.950 850.950 925.050 853.050 ;
        RECT 904.950 847.950 907.050 850.050 ;
        RECT 884.400 838.350 885.600 840.600 ;
        RECT 889.950 839.100 892.050 841.200 ;
        RECT 901.950 839.100 904.050 841.200 ;
        RECT 904.950 840.000 907.050 844.050 ;
        RECT 923.400 843.450 924.450 850.950 ;
        RECT 920.400 842.400 924.450 843.450 ;
        RECT 890.400 838.350 891.600 839.100 ;
        RECT 905.400 838.350 906.600 840.000 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 907.950 835.950 910.050 838.050 ;
        RECT 850.950 832.800 853.050 834.900 ;
        RECT 859.950 832.800 862.050 834.900 ;
        RECT 865.950 832.800 868.050 834.900 ;
        RECT 871.800 832.800 873.900 834.900 ;
        RECT 874.950 832.800 877.050 834.900 ;
        RECT 881.400 833.400 882.600 835.650 ;
        RECT 887.400 833.400 888.600 835.650 ;
        RECT 908.400 834.900 909.600 835.650 ;
        RECT 881.400 829.050 882.450 833.400 ;
        RECT 880.950 826.950 883.050 829.050 ;
        RECT 887.400 823.050 888.450 833.400 ;
        RECT 907.950 832.800 910.050 834.900 ;
        RECT 920.400 834.450 921.450 842.400 ;
        RECT 923.400 835.950 925.500 838.050 ;
        RECT 928.800 835.950 930.900 838.050 ;
        RECT 923.400 834.450 924.600 835.650 ;
        RECT 920.400 833.400 924.600 834.450 ;
        RECT 886.950 820.950 889.050 823.050 ;
        RECT 848.700 813.300 850.800 815.400 ;
        RECT 851.700 813.300 853.800 815.400 ;
        RECT 854.700 813.300 856.800 815.400 ;
        RECT 849.300 809.700 850.500 813.300 ;
        RECT 848.400 807.600 850.500 809.700 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 821.100 799.950 823.200 802.050 ;
        RECT 827.100 799.950 829.200 802.050 ;
        RECT 835.800 799.950 837.900 802.050 ;
        RECT 841.800 799.950 843.900 802.050 ;
        RECT 827.400 798.900 828.600 799.650 ;
        RECT 836.400 798.900 837.600 799.650 ;
        RECT 826.950 796.800 829.050 798.900 ;
        RECT 835.950 796.800 838.050 798.900 ;
        RECT 810.600 786.600 812.700 788.700 ;
        RECT 813.600 786.600 816.600 788.700 ;
        RECT 848.400 788.700 849.900 807.600 ;
        RECT 852.300 796.800 853.500 813.300 ;
        RECT 851.400 794.700 853.500 796.800 ;
        RECT 852.300 788.700 853.500 794.700 ;
        RECT 854.700 791.700 855.900 813.300 ;
        RECT 862.800 812.400 864.900 814.500 ;
        RECT 868.200 813.300 870.300 815.400 ;
        RECT 871.200 813.300 873.300 815.400 ;
        RECT 874.200 813.300 876.300 815.400 ;
        RECT 859.800 805.950 861.900 808.050 ;
        RECT 860.400 804.900 861.600 805.650 ;
        RECT 859.950 802.800 862.050 804.900 ;
        RECT 863.400 801.900 864.300 812.400 ;
        RECT 866.100 806.400 868.200 808.500 ;
        RECT 863.400 799.800 865.500 801.900 ;
        RECT 869.100 801.000 870.300 813.300 ;
        RECT 863.400 793.200 864.300 799.800 ;
        RECT 868.800 798.900 870.900 801.000 ;
        RECT 854.700 789.600 856.800 791.700 ;
        RECT 863.400 791.100 865.500 793.200 ;
        RECT 869.100 791.700 870.300 798.900 ;
        RECT 871.800 795.600 873.300 813.300 ;
        RECT 871.800 793.500 873.900 795.600 ;
        RECT 868.800 789.600 870.900 791.700 ;
        RECT 871.800 788.700 873.300 793.500 ;
        RECT 875.100 791.700 876.300 813.300 ;
        RECT 848.400 786.600 851.400 788.700 ;
        RECT 852.300 786.600 854.400 788.700 ;
        RECT 871.200 786.600 873.300 788.700 ;
        RECT 874.200 786.600 876.300 791.700 ;
        RECT 877.200 813.300 879.300 815.400 ;
        RECT 886.950 814.950 889.050 817.050 ;
        RECT 877.200 795.600 878.700 813.300 ;
        RECT 880.950 802.800 883.050 804.900 ;
        RECT 887.400 804.600 888.450 814.950 ;
        RECT 895.950 811.950 898.050 814.050 ;
        RECT 925.950 811.950 928.050 814.050 ;
        RECT 896.400 804.600 897.450 811.950 ;
        RECT 898.950 806.100 901.050 808.200 ;
        RECT 913.950 806.100 916.050 808.200 ;
        RECT 926.400 807.450 927.450 811.950 ;
        RECT 929.400 807.450 930.600 807.600 ;
        RECT 926.400 806.400 930.600 807.450 ;
        RECT 877.200 793.500 879.300 795.600 ;
        RECT 877.200 788.700 878.700 793.500 ;
        RECT 877.200 786.600 879.300 788.700 ;
        RECT 802.950 781.950 805.050 784.050 ;
        RECT 808.950 781.950 811.050 784.050 ;
        RECT 799.950 772.950 802.050 775.050 ;
        RECT 796.950 769.950 799.050 772.050 ;
        RECT 783.000 768.450 787.050 769.050 ;
        RECT 782.400 768.000 787.050 768.450 ;
        RECT 781.950 766.950 787.050 768.000 ;
        RECT 772.950 763.950 775.050 766.050 ;
        RECT 781.950 764.100 784.050 766.950 ;
        RECT 793.950 763.950 796.050 769.050 ;
        RECT 715.950 751.950 718.050 754.050 ;
        RECT 722.400 751.050 723.450 755.400 ;
        RECT 736.950 754.800 739.050 756.900 ;
        RECT 742.950 754.800 745.050 756.900 ;
        RECT 748.950 754.800 751.050 756.900 ;
        RECT 754.950 754.800 757.050 756.900 ;
        RECT 763.950 754.800 766.050 756.900 ;
        RECT 766.950 754.950 769.050 757.050 ;
        RECT 697.950 748.950 700.050 751.050 ;
        RECT 721.950 748.950 724.050 751.050 ;
        RECT 691.950 742.950 694.050 745.050 ;
        RECT 698.400 732.450 699.450 748.950 ;
        RECT 706.950 739.950 709.050 742.050 ;
        RECT 698.400 731.400 702.450 732.450 ;
        RECT 701.400 729.600 702.450 731.400 ;
        RECT 707.400 729.600 708.450 739.950 ;
        RECT 712.950 733.950 715.050 736.050 ;
        RECT 733.950 733.950 736.050 739.050 ;
        RECT 736.950 736.950 739.050 739.050 ;
        RECT 701.400 727.350 702.600 729.600 ;
        RECT 707.400 727.350 708.600 729.600 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 698.400 723.000 699.600 724.650 ;
        RECT 704.400 723.900 705.600 724.650 ;
        RECT 713.400 723.900 714.450 733.950 ;
        RECT 721.950 728.100 724.050 730.200 ;
        RECT 727.950 728.100 730.050 733.050 ;
        RECT 722.400 727.350 723.600 728.100 ;
        RECT 728.400 727.350 729.600 728.100 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 724.950 724.950 727.050 727.050 ;
        RECT 727.950 724.950 730.050 727.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 719.400 723.900 720.600 724.650 ;
        RECT 697.950 718.950 700.050 723.000 ;
        RECT 703.950 721.800 706.050 723.900 ;
        RECT 712.950 721.800 715.050 723.900 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 725.400 722.400 726.600 724.650 ;
        RECT 731.400 723.900 732.600 724.650 ;
        RECT 688.950 709.950 691.050 712.050 ;
        RECT 679.950 703.950 682.050 706.050 ;
        RECT 680.400 688.200 681.450 703.950 ;
        RECT 725.400 703.050 726.450 722.400 ;
        RECT 730.950 721.800 733.050 723.900 ;
        RECT 737.400 723.450 738.450 736.950 ;
        RECT 743.400 733.050 744.450 754.800 ;
        RECT 745.950 735.600 748.050 736.050 ;
        RECT 751.950 735.600 754.050 736.050 ;
        RECT 745.950 734.550 754.050 735.600 ;
        RECT 745.950 733.950 748.050 734.550 ;
        RECT 751.950 733.950 754.050 734.550 ;
        RECT 755.400 733.050 756.450 754.800 ;
        RECT 773.400 742.050 774.450 763.950 ;
        RECT 781.950 760.950 784.050 763.050 ;
        RECT 782.400 760.350 783.600 760.950 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 775.950 754.950 778.050 757.050 ;
        RECT 779.400 756.900 780.600 757.650 ;
        RECT 776.400 750.450 777.450 754.950 ;
        RECT 778.950 754.800 781.050 756.900 ;
        RECT 785.400 755.400 786.600 757.650 ;
        RECT 797.400 756.900 798.450 769.950 ;
        RECT 800.400 762.450 801.450 772.950 ;
        RECT 805.950 763.950 808.050 769.050 ;
        RECT 809.400 762.600 810.450 781.950 ;
        RECT 814.950 778.950 817.050 781.050 ;
        RECT 815.400 775.050 816.450 778.950 ;
        RECT 826.950 775.950 829.050 778.050 ;
        RECT 847.950 775.950 850.050 778.050 ;
        RECT 814.950 772.950 817.050 775.050 ;
        RECT 823.950 772.950 826.050 775.050 ;
        RECT 803.400 762.450 804.600 762.600 ;
        RECT 800.400 761.400 804.600 762.450 ;
        RECT 803.400 760.350 804.600 761.400 ;
        RECT 809.400 760.350 810.600 762.600 ;
        RECT 814.950 761.100 817.050 763.200 ;
        RECT 820.950 761.100 823.050 763.200 ;
        RECT 815.400 760.350 816.600 761.100 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 776.400 749.400 783.450 750.450 ;
        RECT 772.950 739.950 775.050 742.050 ;
        RECT 760.950 736.950 763.050 739.050 ;
        RECT 757.950 733.950 760.050 736.050 ;
        RECT 742.950 730.950 745.050 733.050 ;
        RECT 745.950 729.000 748.050 732.900 ;
        RECT 754.950 730.950 757.050 733.050 ;
        RECT 746.400 727.350 747.600 729.000 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 749.400 723.900 750.600 724.650 ;
        RECT 734.400 722.400 738.450 723.450 ;
        RECT 712.950 700.950 715.050 703.050 ;
        RECT 724.950 700.950 727.050 703.050 ;
        RECT 697.950 694.950 700.050 697.050 ;
        RECT 701.400 696.300 704.400 698.400 ;
        RECT 705.300 696.300 707.400 698.400 ;
        RECT 679.950 686.100 682.050 688.200 ;
        RECT 688.950 686.100 691.050 688.200 ;
        RECT 680.400 685.350 681.600 686.100 ;
        RECT 689.400 685.350 690.600 686.100 ;
        RECT 674.100 682.950 676.200 685.050 ;
        RECT 680.100 682.950 682.200 685.050 ;
        RECT 688.800 682.950 690.900 685.050 ;
        RECT 694.800 682.950 696.900 685.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 667.500 671.700 668.700 675.300 ;
        RECT 670.950 673.950 673.050 676.050 ;
        RECT 661.200 669.600 663.300 671.700 ;
        RECT 664.200 669.600 666.300 671.700 ;
        RECT 667.200 669.600 669.300 671.700 ;
        RECT 670.950 670.800 673.050 672.900 ;
        RECT 640.950 664.950 643.050 667.050 ;
        RECT 622.950 655.950 625.050 658.050 ;
        RECT 634.950 655.950 637.050 658.050 ;
        RECT 608.400 649.350 609.600 651.600 ;
        RECT 613.950 651.000 616.050 655.050 ;
        RECT 614.400 649.350 615.600 651.000 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 601.950 645.450 604.050 646.050 ;
        RECT 599.400 644.400 604.050 645.450 ;
        RECT 589.950 640.800 592.050 642.900 ;
        RECT 595.950 640.950 598.050 643.050 ;
        RECT 554.700 630.600 556.800 632.700 ;
        RECT 573.600 630.600 575.700 632.700 ;
        RECT 576.600 630.600 579.600 632.700 ;
        RECT 586.950 631.950 589.050 634.050 ;
        RECT 587.400 622.050 588.450 631.950 ;
        RECT 530.700 618.300 532.800 620.400 ;
        RECT 531.300 613.500 532.800 618.300 ;
        RECT 526.950 610.950 529.050 613.050 ;
        RECT 530.700 611.400 532.800 613.500 ;
        RECT 523.950 607.950 526.050 610.050 ;
        RECT 521.100 604.950 523.200 607.050 ;
        RECT 521.400 603.000 522.600 604.650 ;
        RECT 520.950 598.950 523.050 603.000 ;
        RECT 523.950 601.950 526.050 604.050 ;
        RECT 517.950 571.950 520.050 574.050 ;
        RECT 521.400 570.600 522.450 598.950 ;
        RECT 524.400 589.050 525.450 601.950 ;
        RECT 527.400 601.050 528.450 610.950 ;
        RECT 526.950 598.950 529.050 601.050 ;
        RECT 531.300 593.700 532.800 611.400 ;
        RECT 530.700 591.600 532.800 593.700 ;
        RECT 533.700 615.300 535.800 620.400 ;
        RECT 536.700 618.300 538.800 620.400 ;
        RECT 541.950 619.950 544.050 622.050 ;
        RECT 547.950 619.950 550.050 622.050 ;
        RECT 533.700 593.700 534.900 615.300 ;
        RECT 536.700 613.500 538.200 618.300 ;
        RECT 539.100 615.300 541.200 617.400 ;
        RECT 536.100 611.400 538.200 613.500 ;
        RECT 536.700 593.700 538.200 611.400 ;
        RECT 539.700 608.100 540.900 615.300 ;
        RECT 544.500 613.800 546.600 615.900 ;
        RECT 539.100 606.000 541.200 608.100 ;
        RECT 545.700 607.200 546.600 613.800 ;
        RECT 539.700 593.700 540.900 606.000 ;
        RECT 544.500 605.100 546.600 607.200 ;
        RECT 541.800 598.500 543.900 600.600 ;
        RECT 545.700 594.600 546.600 605.100 ;
        RECT 548.400 603.600 549.450 619.950 ;
        RECT 555.600 618.300 557.700 620.400 ;
        RECT 558.600 618.300 561.600 620.400 ;
        RECT 577.950 619.950 580.050 622.050 ;
        RECT 586.950 619.950 589.050 622.050 ;
        RECT 553.200 615.300 555.300 617.400 ;
        RECT 548.400 601.350 549.600 603.600 ;
        RECT 548.100 598.950 550.200 601.050 ;
        RECT 533.700 591.600 535.800 593.700 ;
        RECT 536.700 591.600 538.800 593.700 ;
        RECT 539.700 591.600 541.800 593.700 ;
        RECT 545.100 592.500 547.200 594.600 ;
        RECT 554.100 593.700 555.300 615.300 ;
        RECT 556.500 612.300 557.700 618.300 ;
        RECT 556.500 610.200 558.600 612.300 ;
        RECT 556.500 593.700 557.700 610.200 ;
        RECT 560.100 599.400 561.600 618.300 ;
        RECT 562.950 616.950 565.050 619.050 ;
        RECT 559.500 597.300 561.600 599.400 ;
        RECT 559.500 593.700 560.700 597.300 ;
        RECT 553.200 591.600 555.300 593.700 ;
        RECT 556.200 591.600 558.300 593.700 ;
        RECT 559.200 591.600 561.300 593.700 ;
        RECT 523.950 586.950 526.050 589.050 ;
        RECT 544.950 586.950 547.050 589.050 ;
        RECT 559.950 586.950 562.050 589.050 ;
        RECT 538.950 577.950 541.050 580.050 ;
        RECT 535.950 571.950 538.050 574.050 ;
        RECT 521.400 570.450 522.600 570.600 ;
        RECT 530.400 570.450 531.600 570.600 ;
        RECT 521.400 569.400 525.450 570.450 ;
        RECT 521.400 568.350 522.600 569.400 ;
        RECT 520.800 565.950 522.900 568.050 ;
        RECT 517.950 562.950 520.050 565.050 ;
        RECT 514.950 547.950 517.050 550.050 ;
        RECT 502.950 541.950 505.050 544.050 ;
        RECT 494.400 529.350 495.600 531.600 ;
        RECT 493.800 526.950 495.900 529.050 ;
        RECT 499.800 526.950 501.900 529.050 ;
        RECT 503.400 525.900 504.450 541.950 ;
        RECT 506.400 540.300 509.400 542.400 ;
        RECT 510.300 540.300 512.400 542.400 ;
        RECT 502.950 523.800 505.050 525.900 ;
        RECT 506.400 521.400 507.900 540.300 ;
        RECT 510.300 534.300 511.500 540.300 ;
        RECT 509.400 532.200 511.500 534.300 ;
        RECT 493.950 517.950 496.050 520.050 ;
        RECT 506.400 519.300 508.500 521.400 ;
        RECT 487.950 499.950 490.050 502.050 ;
        RECT 494.400 499.050 495.450 517.950 ;
        RECT 507.300 515.700 508.500 519.300 ;
        RECT 510.300 515.700 511.500 532.200 ;
        RECT 512.700 537.300 514.800 539.400 ;
        RECT 512.700 515.700 513.900 537.300 ;
        RECT 518.400 525.600 519.450 562.950 ;
        RECT 524.400 553.050 525.450 569.400 ;
        RECT 530.400 569.400 534.450 570.450 ;
        RECT 530.400 568.350 531.600 569.400 ;
        RECT 529.800 565.950 531.900 568.050 ;
        RECT 533.400 562.050 534.450 569.400 ;
        RECT 536.400 568.050 537.450 571.950 ;
        RECT 535.950 565.950 538.050 568.050 ;
        RECT 532.950 559.950 535.050 562.050 ;
        RECT 539.400 559.050 540.450 577.950 ;
        RECT 545.400 573.600 546.450 586.950 ;
        RECT 560.400 580.050 561.450 586.950 ;
        RECT 559.950 577.950 562.050 580.050 ;
        RECT 559.950 574.800 562.050 576.900 ;
        RECT 545.400 571.350 546.600 573.600 ;
        RECT 550.950 572.100 553.050 574.200 ;
        RECT 551.400 571.350 552.600 572.100 ;
        RECT 544.950 568.950 547.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 548.400 567.000 549.600 568.650 ;
        RECT 554.400 567.900 555.600 568.650 ;
        RECT 547.950 562.950 550.050 567.000 ;
        RECT 553.950 565.800 556.050 567.900 ;
        RECT 538.950 556.950 541.050 559.050 ;
        RECT 523.950 550.950 526.050 553.050 ;
        RECT 547.950 550.950 550.050 553.050 ;
        RECT 524.400 544.050 525.450 550.950 ;
        RECT 523.950 541.950 526.050 544.050 ;
        RECT 529.200 540.300 531.300 542.400 ;
        RECT 521.400 535.800 523.500 537.900 ;
        RECT 526.800 537.300 528.900 539.400 ;
        RECT 521.400 529.200 522.300 535.800 ;
        RECT 527.100 530.100 528.300 537.300 ;
        RECT 529.800 535.500 531.300 540.300 ;
        RECT 532.200 537.300 534.300 542.400 ;
        RECT 529.800 533.400 531.900 535.500 ;
        RECT 521.400 527.100 523.500 529.200 ;
        RECT 526.800 528.000 528.900 530.100 ;
        RECT 518.400 523.350 519.600 525.600 ;
        RECT 517.800 520.950 519.900 523.050 ;
        RECT 521.400 516.600 522.300 527.100 ;
        RECT 524.100 520.500 526.200 522.600 ;
        RECT 502.950 511.950 505.050 514.050 ;
        RECT 506.700 513.600 508.800 515.700 ;
        RECT 509.700 513.600 511.800 515.700 ;
        RECT 512.700 513.600 514.800 515.700 ;
        RECT 520.800 514.500 522.900 516.600 ;
        RECT 527.100 515.700 528.300 528.000 ;
        RECT 529.800 515.700 531.300 533.400 ;
        RECT 533.100 515.700 534.300 537.300 ;
        RECT 526.200 513.600 528.300 515.700 ;
        RECT 529.200 513.600 531.300 515.700 ;
        RECT 532.200 513.600 534.300 515.700 ;
        RECT 535.200 540.300 537.300 542.400 ;
        RECT 535.200 535.500 536.700 540.300 ;
        RECT 535.200 533.400 537.300 535.500 ;
        RECT 535.200 515.700 536.700 533.400 ;
        RECT 538.950 532.800 541.050 534.900 ;
        RECT 535.200 513.600 537.300 515.700 ;
        RECT 496.950 508.950 499.050 511.050 ;
        RECT 481.950 496.950 484.050 499.050 ;
        RECT 484.950 496.950 487.050 499.050 ;
        RECT 493.950 496.950 496.050 499.050 ;
        RECT 454.950 494.100 457.050 496.200 ;
        RECT 472.950 494.100 475.050 496.200 ;
        RECT 455.400 493.350 456.600 494.100 ;
        RECT 473.400 493.350 474.600 494.100 ;
        RECT 455.400 490.950 457.500 493.050 ;
        RECT 460.800 490.950 462.900 493.050 ;
        RECT 473.400 490.950 475.500 493.050 ;
        RECT 478.800 490.950 480.900 493.050 ;
        RECT 461.400 488.400 462.600 490.650 ;
        RECT 479.400 488.400 480.600 490.650 ;
        RECT 461.400 484.050 462.450 488.400 ;
        RECT 472.950 484.950 475.050 487.050 ;
        RECT 460.950 481.950 463.050 484.050 ;
        RECT 466.950 481.950 469.050 484.050 ;
        RECT 460.950 475.950 463.050 478.050 ;
        RECT 461.400 450.600 462.450 475.950 ;
        RECT 463.950 472.950 466.050 475.050 ;
        RECT 464.400 460.050 465.450 472.950 ;
        RECT 463.950 457.950 466.050 460.050 ;
        RECT 467.400 453.450 468.450 481.950 ;
        RECT 469.950 469.950 472.050 472.050 ;
        RECT 470.400 460.050 471.450 469.950 ;
        RECT 469.950 457.950 472.050 460.050 ;
        RECT 467.400 452.400 471.450 453.450 ;
        RECT 470.400 450.600 471.450 452.400 ;
        RECT 461.400 450.450 462.600 450.600 ;
        RECT 458.400 449.400 462.600 450.450 ;
        RECT 458.400 438.450 459.450 449.400 ;
        RECT 461.400 448.350 462.600 449.400 ;
        RECT 470.400 448.350 471.600 450.600 ;
        RECT 473.400 448.050 474.450 484.950 ;
        RECT 475.950 463.950 478.050 466.050 ;
        RECT 461.100 445.950 463.200 448.050 ;
        RECT 464.400 445.950 466.500 448.050 ;
        RECT 469.800 445.950 471.900 448.050 ;
        RECT 472.950 445.950 475.050 448.050 ;
        RECT 464.400 444.900 465.600 445.650 ;
        RECT 463.950 442.800 466.050 444.900 ;
        RECT 472.950 442.800 475.050 444.900 ;
        RECT 458.400 437.400 462.450 438.450 ;
        RECT 451.950 433.950 454.050 436.050 ;
        RECT 457.950 433.950 460.050 436.050 ;
        RECT 442.950 430.950 445.050 433.050 ;
        RECT 439.950 416.100 442.050 418.200 ;
        RECT 445.950 416.100 448.050 418.200 ;
        RECT 451.950 416.100 454.050 418.200 ;
        RECT 446.400 415.350 447.600 416.100 ;
        RECT 452.400 415.350 453.600 416.100 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 439.950 409.950 442.050 412.050 ;
        RECT 443.400 411.000 444.600 412.650 ;
        RECT 436.950 376.950 439.050 379.050 ;
        RECT 436.950 373.800 439.050 375.900 ;
        RECT 425.400 370.350 426.600 371.100 ;
        RECT 431.400 370.350 432.600 372.600 ;
        RECT 433.950 370.950 436.050 373.050 ;
        RECT 424.950 367.950 427.050 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 428.400 366.900 429.600 367.650 ;
        RECT 427.950 364.800 430.050 366.900 ;
        RECT 433.950 364.950 436.050 367.050 ;
        RECT 418.950 355.950 421.050 358.050 ;
        RECT 424.950 355.950 427.050 358.050 ;
        RECT 406.500 341.400 408.600 343.500 ;
        RECT 413.400 343.200 414.600 345.450 ;
        RECT 404.100 334.950 406.200 337.050 ;
        RECT 404.400 333.450 405.600 334.650 ;
        RECT 401.400 332.400 405.600 333.450 ;
        RECT 394.950 313.950 397.050 316.050 ;
        RECT 401.400 298.050 402.450 332.400 ;
        RECT 407.100 328.800 408.000 341.400 ;
        RECT 413.100 340.800 415.200 342.900 ;
        RECT 416.400 341.100 418.500 343.200 ;
        RECT 408.900 339.000 411.000 339.900 ;
        RECT 408.900 337.800 416.100 339.000 ;
        RECT 414.000 336.900 416.100 337.800 ;
        RECT 408.900 336.000 411.000 336.900 ;
        RECT 417.000 336.000 417.900 341.100 ;
        RECT 418.950 339.450 421.050 340.200 ;
        RECT 418.950 338.400 423.450 339.450 ;
        RECT 418.950 338.100 421.050 338.400 ;
        RECT 419.400 337.350 420.600 338.100 ;
        RECT 408.900 335.100 417.900 336.000 ;
        RECT 408.900 334.800 411.000 335.100 ;
        RECT 413.100 331.950 415.200 334.050 ;
        RECT 413.400 329.400 414.600 331.650 ;
        RECT 406.800 326.700 408.900 328.800 ;
        RECT 417.000 328.500 417.900 335.100 ;
        RECT 418.800 334.950 420.900 337.050 ;
        RECT 422.400 333.900 423.450 338.400 ;
        RECT 421.950 331.800 424.050 333.900 ;
        RECT 409.950 325.950 412.050 328.050 ;
        RECT 415.800 326.400 417.900 328.500 ;
        RECT 403.950 322.950 406.050 325.050 ;
        RECT 404.400 301.050 405.450 322.950 ;
        RECT 403.950 298.950 406.050 301.050 ;
        RECT 400.950 295.950 403.050 298.050 ;
        RECT 397.950 293.100 400.050 295.200 ;
        RECT 404.400 294.600 405.450 298.950 ;
        RECT 398.400 292.350 399.600 293.100 ;
        RECT 404.400 292.350 405.600 294.600 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 401.400 288.900 402.600 289.650 ;
        RECT 400.950 286.800 403.050 288.900 ;
        RECT 391.950 283.950 394.050 286.050 ;
        RECT 394.950 274.950 397.050 277.050 ;
        RECT 395.400 268.050 396.450 274.950 ;
        RECT 388.950 265.950 391.050 268.050 ;
        RECT 394.950 265.950 397.050 268.050 ;
        RECT 389.400 247.050 390.450 265.950 ;
        RECT 395.400 261.600 396.450 265.950 ;
        RECT 395.400 259.350 396.600 261.600 ;
        RECT 406.950 259.950 409.050 262.050 ;
        RECT 392.100 256.950 394.200 259.050 ;
        RECT 395.400 256.950 397.500 259.050 ;
        RECT 400.800 256.950 402.900 259.050 ;
        RECT 392.400 254.400 393.600 256.650 ;
        RECT 401.400 255.000 402.600 256.650 ;
        RECT 388.950 244.950 391.050 247.050 ;
        RECT 392.400 232.050 393.450 254.400 ;
        RECT 400.950 252.450 403.050 255.000 ;
        RECT 400.950 251.400 405.450 252.450 ;
        RECT 400.950 250.950 403.050 251.400 ;
        RECT 397.950 247.950 400.050 250.050 ;
        RECT 391.950 229.950 394.050 232.050 ;
        RECT 391.950 226.800 394.050 228.900 ;
        RECT 382.950 217.950 385.050 220.050 ;
        RECT 380.400 214.350 381.600 216.600 ;
        RECT 385.950 216.000 388.050 220.050 ;
        RECT 392.400 217.050 393.450 226.800 ;
        RECT 394.950 217.950 397.050 220.050 ;
        RECT 386.400 214.350 387.600 216.000 ;
        RECT 391.950 214.950 394.050 217.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 383.400 209.400 384.600 211.650 ;
        RECT 389.400 210.900 390.600 211.650 ;
        RECT 373.950 205.950 376.050 208.050 ;
        RECT 355.950 196.950 358.050 199.050 ;
        RECT 361.950 196.950 364.050 199.050 ;
        RECT 373.950 196.950 376.050 199.050 ;
        RECT 361.950 193.800 364.050 195.900 ;
        RECT 349.950 187.950 352.050 190.050 ;
        RECT 344.400 186.000 348.450 186.450 ;
        RECT 343.950 185.400 348.450 186.000 ;
        RECT 343.950 181.950 346.050 185.400 ;
        RECT 350.400 183.600 351.450 187.950 ;
        RECT 358.950 184.950 361.050 190.050 ;
        RECT 350.400 181.350 351.600 183.600 ;
        RECT 355.950 182.100 358.050 184.200 ;
        RECT 356.400 181.350 357.600 182.100 ;
        RECT 362.400 181.050 363.450 193.800 ;
        RECT 364.950 187.950 367.050 190.050 ;
        RECT 367.950 187.950 370.050 190.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 343.950 175.950 346.050 178.050 ;
        RECT 347.400 176.400 348.600 178.650 ;
        RECT 353.400 177.900 354.600 178.650 ;
        RECT 340.950 154.950 343.050 157.050 ;
        RECT 340.950 148.950 343.050 151.050 ;
        RECT 332.400 136.350 333.600 137.100 ;
        RECT 337.950 136.950 340.050 139.050 ;
        RECT 328.950 133.950 331.050 136.050 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 329.400 133.050 330.600 133.650 ;
        RECT 293.400 127.800 295.500 129.900 ;
        RECT 290.400 125.550 291.600 127.800 ;
        RECT 283.950 121.950 286.050 124.050 ;
        RECT 284.400 118.050 285.450 121.950 ;
        RECT 290.400 118.050 291.450 125.550 ;
        RECT 283.950 115.950 286.050 118.050 ;
        RECT 289.950 115.950 292.050 118.050 ;
        RECT 301.950 115.950 304.050 118.050 ;
        RECT 286.950 114.450 289.050 115.050 ;
        RECT 286.950 114.000 294.450 114.450 ;
        RECT 286.950 113.400 295.050 114.000 ;
        RECT 286.950 112.950 289.050 113.400 ;
        RECT 289.800 109.950 291.900 112.050 ;
        RECT 292.950 109.950 295.050 113.400 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 290.400 106.200 291.450 109.950 ;
        RECT 263.400 105.450 264.600 105.600 ;
        RECT 260.400 104.400 264.600 105.450 ;
        RECT 253.950 94.950 256.050 97.050 ;
        RECT 257.400 94.050 258.450 103.950 ;
        RECT 263.400 103.350 264.600 104.400 ;
        RECT 269.400 103.350 270.600 105.600 ;
        RECT 274.950 103.950 277.050 106.050 ;
        RECT 280.950 103.950 283.050 106.050 ;
        RECT 289.950 104.100 292.050 106.200 ;
        RECT 296.400 105.600 297.450 112.950 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 277.950 100.950 280.050 103.050 ;
        RECT 266.400 99.900 267.600 100.650 ;
        RECT 272.400 99.900 273.600 100.650 ;
        RECT 265.950 97.800 268.050 99.900 ;
        RECT 271.950 97.800 274.050 99.900 ;
        RECT 265.950 96.300 268.050 96.750 ;
        RECT 271.950 96.300 274.050 96.750 ;
        RECT 265.950 95.250 274.050 96.300 ;
        RECT 265.950 94.650 268.050 95.250 ;
        RECT 271.950 94.650 274.050 95.250 ;
        RECT 256.950 91.950 259.050 94.050 ;
        RECT 278.400 91.050 279.450 100.950 ;
        RECT 277.950 88.950 280.050 91.050 ;
        RECT 281.400 85.050 282.450 103.950 ;
        RECT 290.400 103.350 291.600 104.100 ;
        RECT 296.400 103.350 297.600 105.600 ;
        RECT 298.950 103.950 301.050 109.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 287.400 99.900 288.600 100.650 ;
        RECT 286.950 97.800 289.050 99.900 ;
        RECT 293.400 99.000 294.600 100.650 ;
        RECT 292.950 94.950 295.050 99.000 ;
        RECT 298.950 94.950 301.050 99.900 ;
        RECT 280.950 82.950 283.050 85.050 ;
        RECT 268.950 70.950 271.050 73.050 ;
        RECT 247.950 64.950 250.050 67.050 ;
        RECT 247.950 58.950 250.050 61.050 ;
        RECT 253.950 60.000 256.050 64.050 ;
        RECT 238.950 49.950 241.050 54.000 ;
        RECT 244.950 52.950 247.050 55.050 ;
        RECT 248.400 49.050 249.450 58.950 ;
        RECT 254.400 58.350 255.600 60.000 ;
        RECT 259.950 59.100 262.050 61.200 ;
        RECT 260.400 58.350 261.600 59.100 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 257.400 53.400 258.600 55.650 ;
        RECT 263.400 54.900 264.600 55.650 ;
        RECT 247.950 46.950 250.050 49.050 ;
        RECT 257.400 40.050 258.450 53.400 ;
        RECT 262.950 52.800 265.050 54.900 ;
        RECT 265.950 52.950 268.050 55.050 ;
        RECT 256.950 37.950 259.050 40.050 ;
        RECT 232.950 34.950 235.050 37.050 ;
        RECT 233.400 31.050 234.450 34.950 ;
        RECT 235.950 31.950 238.050 34.050 ;
        RECT 247.950 31.950 250.050 34.050 ;
        RECT 262.950 31.950 265.050 34.050 ;
        RECT 232.950 28.950 235.050 31.050 ;
        RECT 212.400 25.350 213.600 26.100 ;
        RECT 218.400 25.350 219.600 26.100 ;
        RECT 223.950 25.950 226.050 28.050 ;
        RECT 226.950 25.950 229.050 28.050 ;
        RECT 229.950 25.950 232.050 28.050 ;
        RECT 236.400 27.600 237.450 31.950 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 184.950 16.950 187.050 22.050 ;
        RECT 188.400 20.400 189.600 22.650 ;
        RECT 194.400 21.900 195.600 22.650 ;
        RECT 181.950 13.950 184.050 16.050 ;
        RECT 188.400 10.050 189.450 20.400 ;
        RECT 193.950 19.800 196.050 21.900 ;
        RECT 205.950 19.950 208.050 22.050 ;
        RECT 209.400 21.900 210.600 22.650 ;
        RECT 202.950 16.950 205.050 19.050 ;
        RECT 187.950 7.950 190.050 10.050 ;
        RECT 203.400 7.050 204.450 16.950 ;
        RECT 206.400 10.050 207.450 19.950 ;
        RECT 208.950 19.800 211.050 21.900 ;
        RECT 215.400 20.400 216.600 22.650 ;
        RECT 205.950 7.950 208.050 10.050 ;
        RECT 209.400 7.050 210.450 19.800 ;
        RECT 211.950 16.950 214.050 19.050 ;
        RECT 163.950 4.950 166.050 7.050 ;
        RECT 202.950 4.950 205.050 7.050 ;
        RECT 208.950 4.950 211.050 7.050 ;
        RECT 212.400 6.450 213.450 16.950 ;
        RECT 215.400 16.050 216.450 20.400 ;
        RECT 220.950 16.950 223.050 19.050 ;
        RECT 214.950 13.950 217.050 16.050 ;
        RECT 221.400 13.050 222.450 16.950 ;
        RECT 220.950 10.950 223.050 13.050 ;
        RECT 224.400 12.450 225.450 25.950 ;
        RECT 227.400 19.050 228.450 25.950 ;
        RECT 236.400 25.350 237.600 27.600 ;
        RECT 241.950 26.100 244.050 28.200 ;
        RECT 242.400 25.350 243.600 26.100 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 233.400 21.900 234.600 22.650 ;
        RECT 232.950 19.800 235.050 21.900 ;
        RECT 239.400 21.000 240.600 22.650 ;
        RECT 248.400 22.050 249.450 31.950 ;
        RECT 256.950 27.000 259.050 31.050 ;
        RECT 257.400 25.350 258.600 27.000 ;
        RECT 259.950 25.950 262.050 31.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 226.950 16.950 229.050 19.050 ;
        RECT 238.950 13.950 241.050 21.000 ;
        RECT 247.950 19.950 250.050 22.050 ;
        RECT 254.400 21.900 255.600 22.650 ;
        RECT 253.950 19.800 256.050 21.900 ;
        RECT 235.950 12.450 238.050 13.050 ;
        RECT 241.950 12.450 244.050 13.050 ;
        RECT 224.400 11.400 228.450 12.450 ;
        RECT 217.950 9.450 220.050 10.050 ;
        RECT 223.950 9.450 226.050 10.050 ;
        RECT 217.950 8.400 226.050 9.450 ;
        RECT 217.950 7.950 220.050 8.400 ;
        RECT 223.950 7.950 226.050 8.400 ;
        RECT 227.400 7.050 228.450 11.400 ;
        RECT 235.950 11.400 244.050 12.450 ;
        RECT 235.950 10.950 238.050 11.400 ;
        RECT 241.950 10.950 244.050 11.400 ;
        RECT 232.950 9.450 235.050 10.050 ;
        RECT 244.950 9.450 247.050 10.050 ;
        RECT 232.950 8.400 247.050 9.450 ;
        RECT 232.950 7.950 235.050 8.400 ;
        RECT 244.950 7.950 247.050 8.400 ;
        RECT 263.400 7.050 264.450 31.950 ;
        RECT 266.400 22.050 267.450 52.950 ;
        RECT 269.400 28.050 270.450 70.950 ;
        RECT 302.400 64.050 303.450 115.950 ;
        RECT 305.400 94.050 306.450 130.950 ;
        RECT 311.400 118.050 312.450 131.400 ;
        RECT 319.950 130.950 322.050 133.050 ;
        RECT 322.950 130.950 325.050 133.050 ;
        RECT 325.950 131.400 330.600 133.050 ;
        RECT 335.400 132.000 336.600 133.650 ;
        RECT 325.950 130.950 330.000 131.400 ;
        RECT 319.950 127.800 322.050 129.900 ;
        RECT 334.950 127.950 337.050 132.000 ;
        RECT 310.950 115.950 313.050 118.050 ;
        RECT 316.950 115.950 319.050 118.050 ;
        RECT 317.400 109.050 318.450 115.950 ;
        RECT 320.400 115.050 321.450 127.800 ;
        RECT 325.950 124.950 328.050 127.050 ;
        RECT 319.950 112.950 322.050 115.050 ;
        RECT 316.950 106.950 319.050 109.050 ;
        RECT 313.950 104.100 316.050 106.200 ;
        RECT 320.400 105.600 321.450 112.950 ;
        RECT 326.400 106.050 327.450 124.950 ;
        RECT 334.950 124.800 337.050 126.900 ;
        RECT 328.950 118.950 331.050 121.050 ;
        RECT 314.400 103.350 315.600 104.100 ;
        RECT 320.400 103.350 321.600 105.600 ;
        RECT 325.950 103.950 328.050 106.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 313.950 100.950 316.050 103.050 ;
        RECT 316.950 100.950 319.050 103.050 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 311.400 98.400 312.600 100.650 ;
        RECT 317.400 98.400 318.600 100.650 ;
        RECT 323.400 99.900 324.600 100.650 ;
        RECT 304.950 91.950 307.050 94.050 ;
        RECT 271.950 59.100 274.050 61.200 ;
        RECT 277.950 59.100 280.050 61.200 ;
        RECT 283.950 59.100 286.050 64.050 ;
        RECT 272.400 49.050 273.450 59.100 ;
        RECT 278.400 58.350 279.600 59.100 ;
        RECT 284.400 58.350 285.600 59.100 ;
        RECT 289.950 58.950 292.050 64.050 ;
        RECT 292.950 61.950 295.050 64.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 274.950 52.950 277.050 55.050 ;
        RECT 281.400 53.400 282.600 55.650 ;
        RECT 287.400 53.400 288.600 55.650 ;
        RECT 271.950 46.950 274.050 49.050 ;
        RECT 275.400 40.050 276.450 52.950 ;
        RECT 281.400 51.450 282.450 53.400 ;
        RECT 281.400 51.000 285.450 51.450 ;
        RECT 280.950 50.400 285.450 51.000 ;
        RECT 280.950 46.950 283.050 50.400 ;
        RECT 284.400 46.050 285.450 50.400 ;
        RECT 287.400 49.050 288.450 53.400 ;
        RECT 286.950 46.950 289.050 49.050 ;
        RECT 283.950 43.950 286.050 46.050 ;
        RECT 280.950 40.950 283.050 43.050 ;
        RECT 274.950 37.950 277.050 40.050 ;
        RECT 274.950 31.950 277.050 34.050 ;
        RECT 268.950 25.950 271.050 28.050 ;
        RECT 275.400 27.600 276.450 31.950 ;
        RECT 281.400 27.600 282.450 40.950 ;
        RECT 286.950 31.950 289.050 34.050 ;
        RECT 275.400 25.350 276.600 27.600 ;
        RECT 281.400 25.350 282.600 27.600 ;
        RECT 287.400 25.050 288.450 31.950 ;
        RECT 293.400 31.050 294.450 61.950 ;
        RECT 298.950 60.000 301.050 64.050 ;
        RECT 301.950 61.950 304.050 64.050 ;
        RECT 304.950 60.000 307.050 64.050 ;
        RECT 311.400 61.050 312.450 98.400 ;
        RECT 313.950 88.950 316.050 91.050 ;
        RECT 299.400 58.350 300.600 60.000 ;
        RECT 305.400 58.350 306.600 60.000 ;
        RECT 310.950 58.950 313.050 61.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 302.400 54.900 303.600 55.650 ;
        RECT 301.950 52.800 304.050 54.900 ;
        RECT 308.400 54.450 309.600 55.650 ;
        RECT 308.400 53.400 312.450 54.450 ;
        RECT 301.950 37.950 304.050 40.050 ;
        RECT 295.950 31.950 298.050 34.050 ;
        RECT 292.950 28.950 295.050 31.050 ;
        RECT 289.950 25.950 292.050 28.050 ;
        RECT 296.400 27.600 297.450 31.950 ;
        RECT 302.400 27.600 303.450 37.950 ;
        RECT 311.400 34.050 312.450 53.400 ;
        RECT 314.400 49.050 315.450 88.950 ;
        RECT 317.400 85.050 318.450 98.400 ;
        RECT 322.950 97.800 325.050 99.900 ;
        RECT 323.400 94.050 324.450 97.800 ;
        RECT 329.400 94.050 330.450 118.950 ;
        RECT 335.400 115.050 336.450 124.800 ;
        RECT 341.400 121.050 342.450 148.950 ;
        RECT 344.400 130.050 345.450 175.950 ;
        RECT 347.400 169.050 348.450 176.400 ;
        RECT 352.950 175.800 355.050 177.900 ;
        RECT 358.950 172.950 361.050 178.050 ;
        RECT 365.400 177.900 366.450 187.950 ;
        RECT 368.400 184.050 369.450 187.950 ;
        RECT 367.950 181.950 370.050 184.050 ;
        RECT 374.400 183.600 375.450 196.950 ;
        RECT 383.400 196.050 384.450 209.400 ;
        RECT 388.950 208.800 391.050 210.900 ;
        RECT 385.950 202.950 388.050 205.050 ;
        RECT 382.950 193.950 385.050 196.050 ;
        RECT 381.000 183.600 385.050 184.050 ;
        RECT 374.400 181.350 375.600 183.600 ;
        RECT 380.400 181.950 385.050 183.600 ;
        RECT 380.400 181.350 381.600 181.950 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 371.400 177.900 372.600 178.650 ;
        RECT 377.400 177.900 378.600 178.650 ;
        RECT 364.950 175.800 367.050 177.900 ;
        RECT 370.950 175.800 373.050 177.900 ;
        RECT 376.950 175.800 379.050 177.900 ;
        RECT 382.950 175.950 385.050 178.050 ;
        RECT 373.950 172.950 376.050 175.050 ;
        RECT 370.950 169.950 373.050 172.050 ;
        RECT 346.950 166.950 349.050 169.050 ;
        RECT 347.400 157.050 348.450 166.950 ;
        RECT 361.950 160.950 364.050 163.050 ;
        RECT 346.950 154.950 349.050 157.050 ;
        RECT 362.400 151.050 363.450 160.950 ;
        RECT 358.800 148.950 360.900 151.050 ;
        RECT 361.950 148.950 364.050 151.050 ;
        RECT 352.950 137.100 355.050 139.200 ;
        RECT 359.400 138.600 360.450 148.950 ;
        RECT 367.950 142.950 370.050 145.050 ;
        RECT 353.400 136.350 354.600 137.100 ;
        RECT 359.400 136.350 360.600 138.600 ;
        RECT 364.950 137.100 367.050 139.200 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 352.950 133.950 355.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 350.400 132.000 351.600 133.650 ;
        RECT 343.950 127.950 346.050 130.050 ;
        RECT 349.950 127.950 352.050 132.000 ;
        RECT 356.400 131.400 357.600 133.650 ;
        RECT 346.950 124.950 349.050 127.050 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 340.950 118.950 343.050 121.050 ;
        RECT 334.950 112.950 337.050 115.050 ;
        RECT 337.950 109.950 340.050 112.050 ;
        RECT 338.400 106.200 339.450 109.950 ;
        RECT 337.950 104.100 340.050 106.200 ;
        RECT 338.400 103.350 339.600 104.100 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 335.400 100.050 336.600 100.650 ;
        RECT 331.950 98.400 336.600 100.050 ;
        RECT 344.400 99.900 345.450 121.950 ;
        RECT 347.400 121.050 348.450 124.950 ;
        RECT 356.400 121.050 357.450 131.400 ;
        RECT 365.400 130.050 366.450 137.100 ;
        RECT 364.950 127.950 367.050 130.050 ;
        RECT 368.400 127.050 369.450 142.950 ;
        RECT 371.400 139.050 372.450 169.950 ;
        RECT 374.400 139.200 375.450 172.950 ;
        RECT 383.400 139.200 384.450 175.950 ;
        RECT 370.950 136.950 373.050 139.050 ;
        RECT 373.950 137.100 376.050 139.200 ;
        RECT 380.400 138.450 381.600 138.600 ;
        RECT 382.950 138.450 385.050 139.200 ;
        RECT 380.400 137.400 385.050 138.450 ;
        RECT 374.400 136.350 375.600 137.100 ;
        RECT 380.400 136.350 381.600 137.400 ;
        RECT 382.950 137.100 385.050 137.400 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 370.950 127.950 373.050 133.050 ;
        RECT 377.400 131.400 378.600 133.650 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 367.950 124.950 370.050 127.050 ;
        RECT 346.950 118.950 349.050 121.050 ;
        RECT 355.950 118.950 358.050 121.050 ;
        RECT 364.950 118.950 367.050 121.050 ;
        RECT 361.950 115.950 364.050 118.050 ;
        RECT 355.950 112.950 358.050 115.050 ;
        RECT 349.950 104.100 352.050 106.200 ;
        RECT 356.400 105.600 357.450 112.950 ;
        RECT 362.400 109.050 363.450 115.950 ;
        RECT 361.950 106.950 364.050 109.050 ;
        RECT 350.400 103.350 351.600 104.100 ;
        RECT 356.400 103.350 357.600 105.600 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 352.950 100.950 355.050 103.050 ;
        RECT 355.950 100.950 358.050 103.050 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 353.400 99.900 354.600 100.650 ;
        RECT 331.950 97.950 336.000 98.400 ;
        RECT 343.950 97.800 346.050 99.900 ;
        RECT 352.950 97.800 355.050 99.900 ;
        RECT 359.400 98.400 360.600 100.650 ;
        RECT 322.950 91.950 325.050 94.050 ;
        RECT 328.950 91.950 331.050 94.050 ;
        RECT 334.800 91.950 336.900 94.050 ;
        RECT 337.950 91.950 340.050 94.050 ;
        RECT 335.400 88.050 336.450 91.950 ;
        RECT 334.950 85.950 337.050 88.050 ;
        RECT 316.950 82.950 319.050 85.050 ;
        RECT 319.950 76.950 322.050 79.050 ;
        RECT 316.950 61.950 319.050 64.050 ;
        RECT 317.400 52.050 318.450 61.950 ;
        RECT 320.400 61.050 321.450 76.950 ;
        RECT 331.950 67.050 334.050 70.050 ;
        RECT 331.950 66.000 337.050 67.050 ;
        RECT 332.400 65.400 337.050 66.000 ;
        RECT 333.000 64.950 337.050 65.400 ;
        RECT 319.950 58.950 322.050 61.050 ;
        RECT 325.950 59.100 328.050 64.050 ;
        RECT 331.950 60.000 334.050 64.050 ;
        RECT 326.400 58.350 327.600 59.100 ;
        RECT 332.400 58.350 333.600 60.000 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 323.400 53.400 324.600 55.650 ;
        RECT 329.400 54.900 330.600 55.650 ;
        RECT 338.400 55.050 339.450 91.950 ;
        RECT 359.400 88.050 360.450 98.400 ;
        RECT 358.950 85.950 361.050 88.050 ;
        RECT 340.950 67.950 343.050 70.050 ;
        RECT 346.950 67.950 349.050 70.050 ;
        RECT 355.950 67.950 358.050 70.050 ;
        RECT 341.400 61.200 342.450 67.950 ;
        RECT 340.950 59.100 343.050 61.200 ;
        RECT 347.400 60.600 348.450 67.950 ;
        RECT 356.400 63.450 357.450 67.950 ;
        RECT 365.400 63.450 366.450 118.950 ;
        RECT 374.400 105.600 375.450 127.950 ;
        RECT 377.400 108.450 378.450 131.400 ;
        RECT 386.400 124.050 387.450 202.950 ;
        RECT 395.400 193.050 396.450 217.950 ;
        RECT 398.400 205.050 399.450 247.950 ;
        RECT 404.400 232.050 405.450 251.400 ;
        RECT 407.400 250.050 408.450 259.950 ;
        RECT 410.400 253.050 411.450 325.950 ;
        RECT 418.950 310.950 421.050 313.050 ;
        RECT 412.950 307.950 415.050 310.050 ;
        RECT 413.400 277.050 414.450 307.950 ;
        RECT 419.400 294.600 420.450 310.950 ;
        RECT 425.400 304.050 426.450 355.950 ;
        RECT 434.400 339.600 435.450 364.950 ;
        RECT 437.400 343.050 438.450 373.800 ;
        RECT 440.400 367.050 441.450 409.950 ;
        RECT 442.950 406.950 445.050 411.000 ;
        RECT 449.400 410.400 450.600 412.650 ;
        RECT 458.400 412.050 459.450 433.950 ;
        RECT 461.400 430.050 462.450 437.400 ;
        RECT 460.950 427.950 463.050 430.050 ;
        RECT 464.400 424.050 465.450 442.800 ;
        RECT 469.950 439.950 472.050 442.050 ;
        RECT 470.400 436.050 471.450 439.950 ;
        RECT 469.950 433.950 472.050 436.050 ;
        RECT 463.950 421.950 466.050 424.050 ;
        RECT 469.950 421.950 472.050 424.050 ;
        RECT 460.950 415.950 463.050 418.050 ;
        RECT 470.400 417.600 471.450 421.950 ;
        RECT 473.400 421.050 474.450 442.800 ;
        RECT 476.400 442.050 477.450 463.950 ;
        RECT 479.400 448.050 480.450 488.400 ;
        RECT 482.400 451.050 483.450 496.950 ;
        RECT 485.400 469.050 486.450 496.950 ;
        RECT 497.400 495.600 498.450 508.950 ;
        RECT 503.400 499.050 504.450 511.950 ;
        RECT 514.950 505.950 517.050 508.050 ;
        RECT 502.950 496.950 505.050 499.050 ;
        RECT 497.400 493.350 498.600 495.600 ;
        RECT 505.950 493.950 508.050 496.050 ;
        RECT 515.400 495.600 516.450 505.950 ;
        RECT 539.400 505.050 540.450 532.800 ;
        RECT 544.800 526.950 546.900 529.050 ;
        RECT 541.950 523.800 544.050 525.900 ;
        RECT 545.400 525.450 546.600 526.650 ;
        RECT 548.400 525.450 549.450 550.950 ;
        RECT 556.950 547.950 559.050 550.050 ;
        RECT 550.950 535.950 553.050 538.050 ;
        RECT 551.400 532.050 552.450 535.950 ;
        RECT 550.950 529.950 553.050 532.050 ;
        RECT 553.800 526.950 555.900 529.050 ;
        RECT 554.400 525.900 555.600 526.650 ;
        RECT 545.400 524.400 549.450 525.450 ;
        RECT 553.950 523.800 556.050 525.900 ;
        RECT 542.400 520.050 543.450 523.800 ;
        RECT 541.950 517.950 544.050 520.050 ;
        RECT 544.950 514.950 547.050 517.050 ;
        RECT 526.950 502.950 529.050 505.050 ;
        RECT 538.950 502.950 541.050 505.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 487.950 487.950 490.050 490.050 ;
        RECT 494.400 488.400 495.600 490.650 ;
        RECT 484.950 466.950 487.050 469.050 ;
        RECT 488.400 460.050 489.450 487.950 ;
        RECT 494.400 484.050 495.450 488.400 ;
        RECT 506.400 484.050 507.450 493.950 ;
        RECT 515.400 493.350 516.600 495.600 ;
        RECT 523.950 493.950 526.050 496.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 512.400 489.000 513.600 490.650 ;
        RECT 518.400 489.900 519.600 490.650 ;
        RECT 511.950 484.950 514.050 489.000 ;
        RECT 517.950 487.800 520.050 489.900 ;
        RECT 493.950 481.950 496.050 484.050 ;
        RECT 505.950 481.950 508.050 484.050 ;
        RECT 490.950 466.950 493.050 469.050 ;
        RECT 487.950 457.950 490.050 460.050 ;
        RECT 488.400 453.450 489.450 457.950 ;
        RECT 485.400 452.400 489.450 453.450 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 485.400 450.600 486.450 452.400 ;
        RECT 491.400 450.600 492.450 466.950 ;
        RECT 508.950 463.950 511.050 466.050 ;
        RECT 509.400 457.050 510.450 463.950 ;
        RECT 512.400 463.050 513.450 484.950 ;
        RECT 514.950 475.950 517.050 478.050 ;
        RECT 515.400 466.050 516.450 475.950 ;
        RECT 518.400 475.050 519.450 487.800 ;
        RECT 520.950 484.950 523.050 487.050 ;
        RECT 517.950 472.950 520.050 475.050 ;
        RECT 521.400 471.450 522.450 484.950 ;
        RECT 524.400 481.050 525.450 493.950 ;
        RECT 527.400 487.050 528.450 502.950 ;
        RECT 535.950 495.000 538.050 499.050 ;
        RECT 536.400 493.350 537.600 495.000 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 533.400 489.000 534.600 490.650 ;
        RECT 526.950 484.950 529.050 487.050 ;
        RECT 532.950 484.950 535.050 489.000 ;
        RECT 539.400 488.400 540.600 490.650 ;
        RECT 539.400 481.050 540.450 488.400 ;
        RECT 545.400 484.050 546.450 514.950 ;
        RECT 557.400 514.050 558.450 547.950 ;
        RECT 560.400 526.050 561.450 574.800 ;
        RECT 563.400 567.900 564.450 616.950 ;
        RECT 571.950 608.100 574.050 610.200 ;
        RECT 572.400 607.350 573.600 608.100 ;
        RECT 566.100 604.950 568.200 607.050 ;
        RECT 572.100 604.950 574.200 607.050 ;
        RECT 568.950 598.950 571.050 601.050 ;
        RECT 565.950 580.950 568.050 583.050 ;
        RECT 566.400 577.050 567.450 580.950 ;
        RECT 569.400 577.050 570.450 598.950 ;
        RECT 578.400 580.050 579.450 619.950 ;
        RECT 580.950 610.950 583.050 613.050 ;
        RECT 581.400 601.050 582.450 610.950 ;
        RECT 590.400 610.200 591.450 640.800 ;
        RECT 595.950 634.950 598.050 637.050 ;
        RECT 592.950 628.950 595.050 631.050 ;
        RECT 589.950 608.100 592.050 610.200 ;
        RECT 593.400 606.600 594.450 628.950 ;
        RECT 596.400 613.050 597.450 634.950 ;
        RECT 599.400 619.050 600.450 644.400 ;
        RECT 601.950 643.950 604.050 644.400 ;
        RECT 604.950 643.950 607.050 646.050 ;
        RECT 611.400 645.900 612.600 646.650 ;
        RECT 617.400 645.900 618.600 646.650 ;
        RECT 601.950 640.800 604.050 642.900 ;
        RECT 598.950 616.950 601.050 619.050 ;
        RECT 595.950 610.950 598.050 613.050 ;
        RECT 593.400 604.350 594.600 606.600 ;
        RECT 598.950 606.000 601.050 610.050 ;
        RECT 602.400 607.050 603.450 640.800 ;
        RECT 605.400 634.050 606.450 643.950 ;
        RECT 610.950 643.800 613.050 645.900 ;
        RECT 616.950 643.800 619.050 645.900 ;
        RECT 611.400 640.050 612.450 643.800 ;
        RECT 623.400 642.900 624.450 655.950 ;
        RECT 631.950 650.100 634.050 652.200 ;
        RECT 632.400 649.350 633.600 650.100 ;
        RECT 628.950 646.950 631.050 649.050 ;
        RECT 631.950 646.950 634.050 649.050 ;
        RECT 634.950 646.950 637.050 649.050 ;
        RECT 629.400 644.400 630.600 646.650 ;
        RECT 635.400 644.400 636.600 646.650 ;
        RECT 622.950 640.800 625.050 642.900 ;
        RECT 629.400 640.050 630.450 644.400 ;
        RECT 631.950 640.950 634.050 643.050 ;
        RECT 610.950 637.950 613.050 640.050 ;
        RECT 628.950 637.950 631.050 640.050 ;
        RECT 607.950 634.950 610.050 637.050 ;
        RECT 604.950 631.950 607.050 634.050 ;
        RECT 604.950 613.950 607.050 616.050 ;
        RECT 599.400 604.350 600.600 606.000 ;
        RECT 601.950 604.950 604.050 607.050 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 580.950 598.950 583.050 601.050 ;
        RECT 586.950 598.950 589.050 601.050 ;
        RECT 590.400 599.400 591.600 601.650 ;
        RECT 596.400 600.900 597.600 601.650 ;
        RECT 587.400 592.050 588.450 598.950 ;
        RECT 590.400 595.050 591.450 599.400 ;
        RECT 595.950 598.800 598.050 600.900 ;
        RECT 589.950 592.950 592.050 595.050 ;
        RECT 601.950 592.950 604.050 595.050 ;
        RECT 586.950 589.950 589.050 592.050 ;
        RECT 598.950 586.950 601.050 589.050 ;
        RECT 577.950 577.950 580.050 580.050 ;
        RECT 589.950 577.950 592.050 580.050 ;
        RECT 565.950 574.950 568.050 577.050 ;
        RECT 568.950 574.950 571.050 577.050 ;
        RECT 590.400 574.200 591.450 577.950 ;
        RECT 571.950 572.100 574.050 574.200 ;
        RECT 589.950 572.100 592.050 574.200 ;
        RECT 572.400 571.350 573.600 572.100 ;
        RECT 590.400 571.350 591.600 572.100 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 580.950 568.950 583.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 562.950 565.800 565.050 567.900 ;
        RECT 569.400 566.400 570.600 568.650 ;
        RECT 575.400 567.900 576.600 568.650 ;
        RECT 562.950 550.950 565.050 553.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 560.400 517.050 561.450 523.950 ;
        RECT 559.950 514.950 562.050 517.050 ;
        RECT 556.950 511.950 559.050 514.050 ;
        RECT 563.400 513.450 564.450 550.950 ;
        RECT 569.400 538.050 570.450 566.400 ;
        RECT 574.950 565.800 577.050 567.900 ;
        RECT 581.400 565.050 582.450 568.950 ;
        RECT 593.400 566.400 594.600 568.650 ;
        RECT 580.950 562.950 583.050 565.050 ;
        RECT 589.950 562.950 592.050 565.050 ;
        RECT 583.950 556.950 586.050 559.050 ;
        RECT 568.950 535.950 571.050 538.050 ;
        RECT 569.400 528.600 570.450 535.950 ;
        RECT 574.950 532.950 577.050 535.050 ;
        RECT 575.400 528.600 576.450 532.950 ;
        RECT 569.400 526.350 570.600 528.600 ;
        RECT 575.400 526.350 576.600 528.600 ;
        RECT 580.950 527.100 583.050 529.200 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 572.400 522.900 573.600 523.650 ;
        RECT 571.950 520.800 574.050 522.900 ;
        RECT 581.400 520.050 582.450 527.100 ;
        RECT 580.950 517.950 583.050 520.050 ;
        RECT 574.950 514.950 577.050 517.050 ;
        RECT 560.400 512.400 564.450 513.450 ;
        RECT 553.950 499.950 556.050 502.050 ;
        RECT 554.400 495.600 555.450 499.950 ;
        RECT 560.400 496.050 561.450 512.400 ;
        RECT 562.950 508.950 565.050 511.050 ;
        RECT 554.400 493.350 555.600 495.600 ;
        RECT 559.950 493.950 562.050 496.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 551.400 488.400 552.600 490.650 ;
        RECT 557.400 488.400 558.600 490.650 ;
        RECT 544.950 481.950 547.050 484.050 ;
        RECT 523.950 478.950 526.050 481.050 ;
        RECT 538.950 480.450 541.050 481.050 ;
        RECT 538.950 479.400 543.450 480.450 ;
        RECT 538.950 478.950 541.050 479.400 ;
        RECT 518.400 470.400 522.450 471.450 ;
        RECT 514.950 463.950 517.050 466.050 ;
        RECT 511.950 460.950 514.050 463.050 ;
        RECT 514.950 457.950 517.050 460.050 ;
        RECT 508.950 454.950 511.050 457.050 ;
        RECT 485.400 448.350 486.600 450.600 ;
        RECT 491.400 448.350 492.600 450.600 ;
        RECT 505.950 449.100 508.050 451.200 ;
        RECT 512.400 450.450 513.600 450.600 ;
        RECT 515.400 450.450 516.450 457.950 ;
        RECT 512.400 449.400 516.450 450.450 ;
        RECT 506.400 448.350 507.600 449.100 ;
        RECT 512.400 448.350 513.600 449.400 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 490.950 445.950 493.050 448.050 ;
        RECT 496.950 445.950 499.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 488.400 443.400 489.600 445.650 ;
        RECT 475.950 439.950 478.050 442.050 ;
        RECT 475.950 436.800 478.050 438.900 ;
        RECT 472.950 418.950 475.050 421.050 ;
        RECT 476.400 417.600 477.450 436.800 ;
        RECT 488.400 436.050 489.450 443.400 ;
        RECT 487.950 435.450 490.050 436.050 ;
        RECT 485.400 434.400 490.050 435.450 ;
        RECT 478.950 430.950 481.050 433.050 ;
        RECT 479.400 418.050 480.450 430.950 ;
        RECT 481.950 421.950 484.050 424.050 ;
        RECT 449.400 406.050 450.450 410.400 ;
        RECT 457.950 409.950 460.050 412.050 ;
        RECT 457.950 406.800 460.050 408.900 ;
        RECT 448.950 403.950 451.050 406.050 ;
        RECT 442.950 379.950 445.050 382.050 ;
        RECT 443.400 372.450 444.450 379.950 ;
        RECT 446.400 372.450 447.600 372.600 ;
        RECT 443.400 371.400 447.600 372.450 ;
        RECT 446.400 370.350 447.600 371.400 ;
        RECT 451.950 371.100 454.050 373.200 ;
        RECT 458.400 373.050 459.450 406.800 ;
        RECT 461.400 400.050 462.450 415.950 ;
        RECT 470.400 415.350 471.600 417.600 ;
        RECT 476.400 415.350 477.600 417.600 ;
        RECT 478.950 415.950 481.050 418.050 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 472.950 412.950 475.050 415.050 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 467.400 410.400 468.600 412.650 ;
        RECT 473.400 411.000 474.600 412.650 ;
        RECT 467.400 406.050 468.450 410.400 ;
        RECT 472.950 406.950 475.050 411.000 ;
        RECT 478.950 409.950 481.050 412.050 ;
        RECT 479.400 406.050 480.450 409.950 ;
        RECT 466.950 403.950 469.050 406.050 ;
        RECT 478.950 403.950 481.050 406.050 ;
        RECT 471.000 402.450 475.050 403.050 ;
        RECT 470.400 402.000 475.050 402.450 ;
        RECT 469.950 400.950 475.050 402.000 ;
        RECT 460.950 397.950 463.050 400.050 ;
        RECT 469.950 397.950 472.050 400.950 ;
        RECT 469.950 388.950 472.050 391.050 ;
        RECT 460.950 385.950 463.050 388.050 ;
        RECT 452.400 370.350 453.600 371.100 ;
        RECT 457.950 370.950 460.050 373.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 439.950 364.950 442.050 367.050 ;
        RECT 449.400 366.000 450.600 367.650 ;
        RECT 448.950 361.950 451.050 366.000 ;
        RECT 455.400 365.400 456.600 367.650 ;
        RECT 442.950 349.950 445.050 352.050 ;
        RECT 436.950 340.950 439.050 343.050 ;
        RECT 434.400 337.350 435.600 339.600 ;
        RECT 439.950 338.100 442.050 340.200 ;
        RECT 443.400 340.050 444.450 349.950 ;
        RECT 445.950 346.950 448.050 349.050 ;
        RECT 451.950 346.950 454.050 349.050 ;
        RECT 440.400 337.350 441.600 338.100 ;
        RECT 442.950 337.950 445.050 340.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 431.400 332.400 432.600 334.650 ;
        RECT 437.400 333.900 438.600 334.650 ;
        RECT 431.400 325.050 432.450 332.400 ;
        RECT 436.950 331.800 439.050 333.900 ;
        RECT 442.950 331.950 445.050 334.050 ;
        RECT 443.400 328.050 444.450 331.950 ;
        RECT 442.950 325.950 445.050 328.050 ;
        RECT 446.400 325.050 447.450 346.950 ;
        RECT 448.950 340.950 451.050 343.050 ;
        RECT 452.400 342.450 453.450 346.950 ;
        RECT 455.400 346.050 456.450 365.400 ;
        RECT 461.400 352.050 462.450 385.950 ;
        RECT 470.400 384.450 471.450 388.950 ;
        RECT 482.400 388.050 483.450 421.950 ;
        RECT 485.400 418.050 486.450 434.400 ;
        RECT 487.950 433.950 490.050 434.400 ;
        RECT 490.950 429.450 493.050 433.050 ;
        RECT 488.400 429.000 493.050 429.450 ;
        RECT 488.400 428.400 492.450 429.000 ;
        RECT 488.400 418.050 489.450 428.400 ;
        RECT 497.400 427.050 498.450 445.950 ;
        RECT 503.400 443.400 504.600 445.650 ;
        RECT 509.400 443.400 510.600 445.650 ;
        RECT 518.400 444.450 519.450 470.400 ;
        RECT 526.800 463.950 528.900 466.050 ;
        RECT 529.950 463.950 532.050 466.050 ;
        RECT 538.950 463.950 541.050 466.050 ;
        RECT 527.400 454.050 528.450 463.950 ;
        RECT 526.950 451.950 529.050 454.050 ;
        RECT 523.950 449.100 526.050 451.200 ;
        RECT 530.400 450.600 531.450 463.950 ;
        RECT 535.950 457.950 538.050 460.050 ;
        RECT 536.400 451.050 537.450 457.950 ;
        RECT 524.400 448.350 525.600 449.100 ;
        RECT 530.400 448.350 531.600 450.600 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 515.400 443.400 519.450 444.450 ;
        RECT 503.400 433.050 504.450 443.400 ;
        RECT 509.400 433.050 510.450 443.400 ;
        RECT 502.950 430.950 505.050 433.050 ;
        RECT 508.950 430.950 511.050 433.050 ;
        RECT 490.950 424.950 493.050 427.050 ;
        RECT 496.950 424.950 499.050 427.050 ;
        RECT 505.950 424.950 508.050 427.050 ;
        RECT 484.950 415.950 487.050 418.050 ;
        RECT 487.950 415.950 490.050 418.050 ;
        RECT 491.400 417.600 492.450 424.950 ;
        RECT 496.950 421.800 499.050 423.900 ;
        RECT 497.400 417.600 498.450 421.800 ;
        RECT 491.400 415.350 492.600 417.600 ;
        RECT 497.400 415.350 498.600 417.600 ;
        RECT 502.950 416.100 505.050 418.200 ;
        RECT 506.400 418.050 507.450 424.950 ;
        RECT 503.400 415.350 504.600 416.100 ;
        RECT 505.950 415.950 508.050 418.050 ;
        RECT 484.950 409.800 487.050 414.900 ;
        RECT 490.950 412.950 493.050 415.050 ;
        RECT 493.950 412.950 496.050 415.050 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 494.400 411.900 495.600 412.650 ;
        RECT 500.400 411.900 501.600 412.650 ;
        RECT 493.950 409.800 496.050 411.900 ;
        RECT 499.950 409.800 502.050 411.900 ;
        RECT 505.950 409.950 508.050 412.050 ;
        RECT 487.950 403.950 490.050 406.050 ;
        RECT 481.950 385.950 484.050 388.050 ;
        RECT 478.950 384.450 481.050 385.050 ;
        RECT 470.400 383.400 481.050 384.450 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 469.950 379.950 472.050 382.050 ;
        RECT 475.950 379.950 478.050 382.050 ;
        RECT 463.950 373.950 466.050 376.050 ;
        RECT 464.400 364.050 465.450 373.950 ;
        RECT 470.400 373.200 471.450 379.950 ;
        RECT 469.950 371.100 472.050 373.200 ;
        RECT 476.400 372.600 477.450 379.950 ;
        RECT 481.950 376.950 484.050 379.050 ;
        RECT 482.400 372.600 483.450 376.950 ;
        RECT 470.400 370.350 471.600 371.100 ;
        RECT 476.400 370.350 477.600 372.600 ;
        RECT 482.400 370.350 483.600 372.600 ;
        RECT 469.950 367.950 472.050 370.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 466.950 364.950 469.050 367.050 ;
        RECT 473.400 365.400 474.600 367.650 ;
        RECT 479.400 365.400 480.600 367.650 ;
        RECT 488.400 367.050 489.450 403.950 ;
        RECT 490.950 391.950 493.050 394.050 ;
        RECT 491.400 367.050 492.450 391.950 ;
        RECT 502.950 382.950 505.050 385.050 ;
        RECT 503.400 376.050 504.450 382.950 ;
        RECT 506.400 379.050 507.450 409.950 ;
        RECT 505.950 376.950 508.050 379.050 ;
        RECT 502.950 373.950 505.050 376.050 ;
        RECT 496.950 371.100 499.050 373.200 ;
        RECT 506.400 373.050 507.450 376.950 ;
        RECT 509.400 376.050 510.450 430.950 ;
        RECT 511.950 421.950 514.050 424.050 ;
        RECT 508.950 373.950 511.050 376.050 ;
        RECT 503.400 372.450 504.600 372.600 ;
        RECT 505.950 372.450 508.050 373.050 ;
        RECT 512.400 372.450 513.450 421.950 ;
        RECT 515.400 418.050 516.450 443.400 ;
        RECT 520.950 442.950 523.050 445.050 ;
        RECT 527.400 444.900 528.600 445.650 ;
        RECT 521.400 439.050 522.450 442.950 ;
        RECT 526.950 442.800 529.050 444.900 ;
        RECT 533.400 443.400 534.600 445.650 ;
        RECT 520.950 436.950 523.050 439.050 ;
        RECT 517.950 433.950 520.050 436.050 ;
        RECT 514.950 415.950 517.050 418.050 ;
        RECT 518.400 417.600 519.450 433.950 ;
        RECT 533.400 427.050 534.450 443.400 ;
        RECT 539.400 433.050 540.450 463.950 ;
        RECT 542.400 439.050 543.450 479.400 ;
        RECT 551.400 463.050 552.450 488.400 ;
        RECT 557.400 484.050 558.450 488.400 ;
        RECT 559.950 487.950 562.050 490.050 ;
        RECT 556.950 481.950 559.050 484.050 ;
        RECT 560.400 475.050 561.450 487.950 ;
        RECT 559.950 472.950 562.050 475.050 ;
        RECT 553.950 466.950 556.050 469.050 ;
        RECT 550.950 460.950 553.050 463.050 ;
        RECT 547.950 450.000 550.050 454.050 ;
        RECT 554.400 450.600 555.450 466.950 ;
        RECT 548.400 448.350 549.600 450.000 ;
        RECT 554.400 448.350 555.600 450.600 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 556.950 445.950 559.050 448.050 ;
        RECT 551.400 444.900 552.600 445.650 ;
        RECT 550.950 442.800 553.050 444.900 ;
        RECT 557.400 443.400 558.600 445.650 ;
        RECT 541.950 436.950 544.050 439.050 ;
        RECT 547.950 436.950 550.050 439.050 ;
        RECT 538.950 430.950 541.050 433.050 ;
        RECT 532.950 424.950 535.050 427.050 ;
        RECT 523.950 421.950 526.050 424.050 ;
        RECT 524.400 418.200 525.450 421.950 ;
        RECT 518.400 415.350 519.600 417.600 ;
        RECT 523.950 416.100 526.050 418.200 ;
        RECT 529.950 416.100 532.050 418.200 ;
        RECT 524.400 415.350 525.600 416.100 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 514.950 409.950 517.050 412.050 ;
        RECT 521.400 410.400 522.600 412.650 ;
        RECT 515.400 400.050 516.450 409.950 ;
        RECT 521.400 409.050 522.450 410.400 ;
        RECT 521.400 407.400 526.050 409.050 ;
        RECT 522.000 406.950 526.050 407.400 ;
        RECT 517.950 403.950 520.050 406.050 ;
        RECT 526.950 403.950 529.050 406.050 ;
        RECT 514.950 397.950 517.050 400.050 ;
        RECT 503.400 371.400 508.050 372.450 ;
        RECT 497.400 370.350 498.600 371.100 ;
        RECT 503.400 370.350 504.600 371.400 ;
        RECT 505.950 370.950 508.050 371.400 ;
        RECT 509.400 371.400 513.450 372.450 ;
        RECT 514.950 372.000 517.050 376.050 ;
        RECT 518.400 375.450 519.450 403.950 ;
        RECT 518.400 374.400 522.450 375.450 ;
        RECT 521.400 372.600 522.450 374.400 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 463.950 361.950 466.050 364.050 ;
        RECT 461.400 350.400 466.050 352.050 ;
        RECT 462.000 349.950 466.050 350.400 ;
        RECT 454.950 343.950 457.050 346.050 ;
        RECT 463.950 343.950 466.050 346.050 ;
        RECT 452.400 341.400 456.450 342.450 ;
        RECT 449.400 337.050 450.450 340.950 ;
        RECT 455.400 339.600 456.450 341.400 ;
        RECT 464.400 340.050 465.450 343.950 ;
        RECT 467.400 342.450 468.450 364.950 ;
        RECT 473.400 361.050 474.450 365.400 ;
        RECT 472.950 358.950 475.050 361.050 ;
        RECT 469.950 342.450 472.050 343.050 ;
        RECT 467.400 341.400 472.050 342.450 ;
        RECT 469.950 340.950 472.050 341.400 ;
        RECT 455.400 337.350 456.600 339.600 ;
        RECT 463.950 337.950 466.050 340.050 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 452.100 334.950 454.200 337.050 ;
        RECT 455.400 334.950 457.500 337.050 ;
        RECT 460.800 334.950 462.900 337.050 ;
        RECT 448.950 328.950 451.050 333.900 ;
        RECT 452.400 332.400 453.600 334.650 ;
        RECT 461.400 332.400 462.600 334.650 ;
        RECT 430.950 322.950 433.050 325.050 ;
        RECT 439.950 322.950 442.050 325.050 ;
        RECT 430.950 316.950 433.050 319.050 ;
        RECT 431.400 310.050 432.450 316.950 ;
        RECT 430.950 307.950 433.050 310.050 ;
        RECT 424.950 301.950 427.050 304.050 ;
        RECT 424.950 298.800 427.050 300.900 ;
        RECT 425.400 294.600 426.450 298.800 ;
        RECT 419.400 292.350 420.600 294.600 ;
        RECT 425.400 292.350 426.600 294.600 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 422.400 287.400 423.600 289.650 ;
        RECT 415.950 280.950 418.050 283.050 ;
        RECT 412.950 274.950 415.050 277.050 ;
        RECT 416.400 274.050 417.450 280.950 ;
        RECT 415.950 271.950 418.050 274.050 ;
        RECT 418.950 260.100 421.050 262.200 ;
        RECT 422.400 261.450 423.450 287.400 ;
        RECT 431.400 271.050 432.450 307.950 ;
        RECT 433.950 301.950 436.050 304.050 ;
        RECT 434.400 280.050 435.450 301.950 ;
        RECT 440.400 294.600 441.450 322.950 ;
        RECT 442.950 322.800 445.050 324.900 ;
        RECT 445.950 322.950 448.050 325.050 ;
        RECT 448.950 322.950 451.050 327.900 ;
        RECT 443.400 310.050 444.450 322.800 ;
        RECT 452.400 316.050 453.450 332.400 ;
        RECT 461.400 322.050 462.450 332.400 ;
        RECT 460.950 319.950 463.050 322.050 ;
        RECT 451.950 313.950 454.050 316.050 ;
        RECT 445.950 310.950 448.050 313.050 ;
        RECT 442.950 307.950 445.050 310.050 ;
        RECT 446.400 307.050 447.450 310.950 ;
        RECT 452.400 309.450 453.450 313.950 ;
        RECT 449.400 308.400 453.450 309.450 ;
        RECT 445.950 304.950 448.050 307.050 ;
        RECT 446.400 294.600 447.450 304.950 ;
        RECT 449.400 301.050 450.450 308.400 ;
        RECT 451.950 304.950 454.050 307.050 ;
        RECT 448.950 298.950 451.050 301.050 ;
        RECT 440.400 292.350 441.600 294.600 ;
        RECT 446.400 292.350 447.600 294.600 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 443.400 288.900 444.600 289.650 ;
        RECT 442.950 286.800 445.050 288.900 ;
        RECT 448.950 286.950 451.050 289.050 ;
        RECT 433.950 277.950 436.050 280.050 ;
        RECT 430.950 268.950 433.050 271.050 ;
        RECT 431.400 262.200 432.450 268.950 ;
        RECT 443.400 268.050 444.450 286.800 ;
        RECT 445.950 277.950 448.050 280.050 ;
        RECT 436.950 265.950 439.050 268.050 ;
        RECT 442.950 265.950 445.050 268.050 ;
        RECT 437.400 262.200 438.450 265.950 ;
        RECT 422.400 260.400 426.450 261.450 ;
        RECT 419.400 259.350 420.600 260.100 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 416.400 254.400 417.600 256.650 ;
        RECT 409.950 250.950 412.050 253.050 ;
        RECT 416.400 250.050 417.450 254.400 ;
        RECT 421.950 253.950 424.050 256.050 ;
        RECT 418.950 250.950 421.050 253.050 ;
        RECT 406.950 247.950 409.050 250.050 ;
        RECT 415.950 247.950 418.050 250.050 ;
        RECT 403.950 229.950 406.050 232.050 ;
        RECT 400.950 220.950 403.050 223.050 ;
        RECT 397.950 202.950 400.050 205.050 ;
        RECT 394.950 190.950 397.050 193.050 ;
        RECT 391.950 187.950 394.050 190.050 ;
        RECT 392.400 184.200 393.450 187.950 ;
        RECT 391.950 182.100 394.050 184.200 ;
        RECT 392.400 181.350 393.600 182.100 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 394.950 178.950 397.050 181.050 ;
        RECT 395.400 178.050 396.600 178.650 ;
        RECT 395.400 177.900 400.050 178.050 ;
        RECT 394.950 175.950 400.050 177.900 ;
        RECT 394.950 175.800 397.050 175.950 ;
        RECT 401.400 175.050 402.450 220.950 ;
        RECT 404.400 216.600 405.450 229.950 ;
        RECT 404.400 214.350 405.600 216.600 ;
        RECT 413.400 216.450 414.600 216.600 ;
        RECT 413.400 215.400 417.450 216.450 ;
        RECT 413.400 214.350 414.600 215.400 ;
        RECT 404.100 211.950 406.200 214.050 ;
        RECT 409.500 211.950 411.600 214.050 ;
        RECT 412.800 211.950 414.900 214.050 ;
        RECT 410.400 210.900 411.600 211.650 ;
        RECT 409.950 208.800 412.050 210.900 ;
        RECT 403.950 205.950 406.050 208.050 ;
        RECT 404.400 178.050 405.450 205.950 ;
        RECT 410.400 205.050 411.450 208.800 ;
        RECT 409.950 202.950 412.050 205.050 ;
        RECT 406.950 193.950 409.050 196.050 ;
        RECT 407.400 184.050 408.450 193.950 ;
        RECT 416.400 187.050 417.450 215.400 ;
        RECT 419.400 211.050 420.450 250.950 ;
        RECT 422.400 244.050 423.450 253.950 ;
        RECT 421.950 241.950 424.050 244.050 ;
        RECT 425.400 216.450 426.450 260.400 ;
        RECT 430.950 260.100 433.050 262.200 ;
        RECT 436.950 260.100 439.050 262.200 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 428.400 253.050 429.450 256.950 ;
        RECT 427.950 250.950 430.050 253.050 ;
        RECT 427.950 226.950 430.050 229.050 ;
        RECT 431.400 228.450 432.450 260.100 ;
        RECT 437.400 259.350 438.600 260.100 ;
        RECT 434.100 256.950 436.200 259.050 ;
        RECT 437.400 256.950 439.500 259.050 ;
        RECT 442.800 256.950 444.900 259.050 ;
        RECT 434.400 254.400 435.600 256.650 ;
        RECT 443.400 255.450 444.600 256.650 ;
        RECT 446.400 255.900 447.450 277.950 ;
        RECT 445.950 255.450 448.050 255.900 ;
        RECT 443.400 254.400 448.050 255.450 ;
        RECT 434.400 232.050 435.450 254.400 ;
        RECT 445.950 253.800 448.050 254.400 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 433.950 229.950 436.050 232.050 ;
        RECT 442.950 229.950 445.050 232.050 ;
        RECT 431.400 227.400 435.450 228.450 ;
        RECT 428.400 223.050 429.450 226.950 ;
        RECT 427.950 220.950 430.050 223.050 ;
        RECT 422.400 215.400 426.450 216.450 ;
        RECT 427.950 216.000 430.050 219.900 ;
        RECT 434.400 217.200 435.450 227.400 ;
        RECT 439.950 220.950 442.050 223.050 ;
        RECT 418.950 208.950 421.050 211.050 ;
        RECT 418.950 202.950 421.050 205.050 ;
        RECT 415.950 184.950 418.050 187.050 ;
        RECT 406.950 181.950 409.050 184.050 ;
        RECT 412.950 182.100 415.050 184.200 ;
        RECT 419.400 184.050 420.450 202.950 ;
        RECT 413.400 181.350 414.600 182.100 ;
        RECT 418.950 181.950 421.050 184.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 415.950 178.950 418.050 181.050 ;
        RECT 403.950 175.950 406.050 178.050 ;
        RECT 410.400 176.400 411.600 178.650 ;
        RECT 416.400 176.400 417.600 178.650 ;
        RECT 400.950 172.950 403.050 175.050 ;
        RECT 406.950 172.950 409.050 175.050 ;
        RECT 388.950 169.950 391.050 172.050 ;
        RECT 385.950 121.950 388.050 124.050 ;
        RECT 389.400 112.050 390.450 169.950 ;
        RECT 391.950 137.100 394.050 139.200 ;
        RECT 401.400 138.450 402.600 138.600 ;
        RECT 401.400 137.400 405.450 138.450 ;
        RECT 392.400 136.350 393.600 137.100 ;
        RECT 401.400 136.350 402.600 137.400 ;
        RECT 392.100 133.950 394.200 136.050 ;
        RECT 397.500 133.950 399.600 136.050 ;
        RECT 400.800 133.950 402.900 136.050 ;
        RECT 398.400 132.900 399.600 133.650 ;
        RECT 397.950 130.800 400.050 132.900 ;
        RECT 391.950 127.950 394.050 130.050 ;
        RECT 388.950 109.950 391.050 112.050 ;
        RECT 377.400 107.400 381.450 108.450 ;
        RECT 374.400 103.350 375.600 105.600 ;
        RECT 380.400 105.450 381.450 107.400 ;
        RECT 380.400 104.400 384.450 105.450 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 373.950 100.950 376.050 103.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 371.400 99.900 372.600 100.650 ;
        RECT 370.950 97.800 373.050 99.900 ;
        RECT 377.400 98.400 378.600 100.650 ;
        RECT 371.400 94.050 372.450 97.800 ;
        RECT 370.950 91.950 373.050 94.050 ;
        RECT 377.400 91.050 378.450 98.400 ;
        RECT 376.950 88.950 379.050 91.050 ;
        RECT 383.400 76.050 384.450 104.400 ;
        RECT 385.950 104.100 388.050 106.200 ;
        RECT 392.400 105.600 393.450 127.950 ;
        RECT 386.400 91.050 387.450 104.100 ;
        RECT 392.400 103.350 393.600 105.600 ;
        RECT 397.950 104.100 400.050 106.200 ;
        RECT 404.400 106.050 405.450 137.400 ;
        RECT 398.400 103.350 399.600 104.100 ;
        RECT 403.950 103.950 406.050 106.050 ;
        RECT 407.400 103.050 408.450 172.950 ;
        RECT 410.400 154.050 411.450 176.400 ;
        RECT 416.400 172.050 417.450 176.400 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 415.950 169.950 418.050 172.050 ;
        RECT 419.400 166.050 420.450 175.950 ;
        RECT 418.950 163.950 421.050 166.050 ;
        RECT 422.400 163.050 423.450 215.400 ;
        RECT 428.400 214.350 429.600 216.000 ;
        RECT 433.950 215.100 436.050 217.200 ;
        RECT 434.400 214.350 435.600 215.100 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 430.950 211.950 433.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 424.950 208.950 427.050 211.050 ;
        RECT 431.400 210.000 432.600 211.650 ;
        RECT 425.400 169.050 426.450 208.950 ;
        RECT 430.950 205.950 433.050 210.000 ;
        RECT 433.950 193.950 436.050 196.050 ;
        RECT 427.950 181.950 430.050 187.050 ;
        RECT 434.400 183.600 435.450 193.950 ;
        RECT 440.400 190.050 441.450 220.950 ;
        RECT 439.950 187.950 442.050 190.050 ;
        RECT 443.400 186.450 444.450 229.950 ;
        RECT 446.400 229.050 447.450 235.950 ;
        RECT 445.950 226.950 448.050 229.050 ;
        RECT 446.400 216.600 447.450 226.950 ;
        RECT 449.400 223.050 450.450 286.950 ;
        RECT 452.400 250.050 453.450 304.950 ;
        RECT 457.950 293.100 460.050 295.200 ;
        RECT 464.400 294.600 465.450 337.950 ;
        RECT 466.950 337.800 469.050 339.900 ;
        RECT 467.400 328.050 468.450 337.800 ;
        RECT 466.950 325.950 469.050 328.050 ;
        RECT 470.400 295.050 471.450 340.950 ;
        RECT 473.400 340.050 474.450 358.950 ;
        RECT 479.400 352.050 480.450 365.400 ;
        RECT 487.950 364.950 490.050 367.050 ;
        RECT 490.950 364.950 493.050 367.050 ;
        RECT 500.400 366.900 501.600 367.650 ;
        RECT 499.950 364.800 502.050 366.900 ;
        RECT 481.950 358.950 484.050 364.050 ;
        RECT 493.950 358.950 496.050 361.050 ;
        RECT 478.950 349.950 481.050 352.050 ;
        RECT 481.950 343.950 484.050 346.050 ;
        RECT 490.950 343.950 493.050 346.050 ;
        RECT 472.950 337.950 475.050 340.050 ;
        RECT 475.950 339.000 478.050 343.050 ;
        RECT 482.400 339.600 483.450 343.950 ;
        RECT 476.400 337.350 477.600 339.000 ;
        RECT 482.400 337.350 483.600 339.600 ;
        RECT 487.950 337.950 490.050 343.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 479.400 332.400 480.600 334.650 ;
        RECT 485.400 333.900 486.600 334.650 ;
        RECT 479.400 307.050 480.450 332.400 ;
        RECT 484.950 331.800 487.050 333.900 ;
        RECT 491.400 328.050 492.450 343.950 ;
        RECT 494.400 340.050 495.450 358.950 ;
        RECT 499.950 349.950 502.050 352.050 ;
        RECT 493.950 337.950 496.050 340.050 ;
        RECT 500.400 339.600 501.450 349.950 ;
        RECT 500.400 337.350 501.600 339.600 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 497.400 333.900 498.600 334.650 ;
        RECT 496.950 331.800 499.050 333.900 ;
        RECT 503.400 333.000 504.600 334.650 ;
        RECT 502.950 328.950 505.050 333.000 ;
        RECT 490.950 325.950 493.050 328.050 ;
        RECT 496.950 322.950 499.050 325.050 ;
        RECT 493.950 319.950 496.050 322.050 ;
        RECT 494.400 310.050 495.450 319.950 ;
        RECT 493.950 307.950 496.050 310.050 ;
        RECT 478.950 304.950 481.050 307.050 ;
        RECT 487.950 298.950 490.050 301.050 ;
        RECT 458.400 292.350 459.600 293.100 ;
        RECT 464.400 292.350 465.600 294.600 ;
        RECT 469.800 292.950 471.900 295.050 ;
        RECT 472.950 292.950 475.050 295.050 ;
        RECT 478.950 293.100 481.050 295.200 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 461.400 287.400 462.600 289.650 ;
        RECT 467.400 288.900 468.600 289.650 ;
        RECT 473.400 288.900 474.450 292.950 ;
        RECT 479.400 292.350 480.600 293.100 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 482.400 288.900 483.600 289.650 ;
        RECT 461.400 280.050 462.450 287.400 ;
        RECT 466.950 286.800 469.050 288.900 ;
        RECT 472.950 286.800 475.050 288.900 ;
        RECT 481.950 286.800 484.050 288.900 ;
        RECT 460.950 277.950 463.050 280.050 ;
        RECT 469.950 277.950 472.050 280.050 ;
        RECT 457.950 271.950 460.050 274.050 ;
        RECT 454.950 268.950 457.050 271.050 ;
        RECT 455.400 265.050 456.450 268.950 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 458.400 261.600 459.450 271.950 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 464.400 261.600 465.450 265.950 ;
        RECT 458.400 259.350 459.600 261.600 ;
        RECT 464.400 259.350 465.600 261.600 ;
        RECT 457.950 256.950 460.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 461.400 254.400 462.600 256.650 ;
        RECT 457.950 250.950 460.050 253.050 ;
        RECT 451.950 247.950 454.050 250.050 ;
        RECT 448.950 220.950 451.050 223.050 ;
        RECT 446.400 214.350 447.600 216.600 ;
        RECT 454.950 215.100 457.050 217.200 ;
        RECT 455.400 214.350 456.600 215.100 ;
        RECT 446.100 211.950 448.200 214.050 ;
        RECT 451.500 211.950 453.600 214.050 ;
        RECT 454.800 211.950 456.900 214.050 ;
        RECT 452.400 210.900 453.600 211.650 ;
        RECT 451.950 208.800 454.050 210.900 ;
        RECT 448.950 205.950 451.050 208.050 ;
        RECT 458.400 207.450 459.450 250.950 ;
        RECT 455.400 206.400 459.450 207.450 ;
        RECT 440.400 185.400 444.450 186.450 ;
        RECT 440.400 183.600 441.450 185.400 ;
        RECT 434.400 181.350 435.600 183.600 ;
        RECT 440.400 181.350 441.600 183.600 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 431.400 176.400 432.600 178.650 ;
        RECT 437.400 176.400 438.600 178.650 ;
        RECT 443.400 177.900 444.600 178.650 ;
        RECT 431.400 174.450 432.450 176.400 ;
        RECT 431.400 173.400 435.450 174.450 ;
        RECT 424.950 166.950 427.050 169.050 ;
        RECT 430.950 166.950 433.050 169.050 ;
        RECT 427.950 163.950 430.050 166.050 ;
        RECT 421.950 160.950 424.050 163.050 ;
        RECT 409.950 151.950 412.050 154.050 ;
        RECT 422.400 145.050 423.450 160.950 ;
        RECT 415.950 142.950 418.050 145.050 ;
        RECT 421.950 142.950 424.050 145.050 ;
        RECT 416.400 138.600 417.450 142.950 ;
        RECT 428.400 142.050 429.450 163.950 ;
        RECT 416.400 136.350 417.600 138.600 ;
        RECT 421.950 138.000 424.050 141.900 ;
        RECT 427.950 139.950 430.050 142.050 ;
        RECT 422.400 136.350 423.600 138.000 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 413.400 131.400 414.600 133.650 ;
        RECT 419.400 132.900 420.600 133.650 ;
        RECT 428.400 133.050 429.450 139.950 ;
        RECT 413.400 121.050 414.450 131.400 ;
        RECT 418.950 130.800 421.050 132.900 ;
        RECT 427.950 130.800 430.050 133.050 ;
        RECT 431.400 130.050 432.450 166.950 ;
        RECT 434.400 157.050 435.450 173.400 ;
        RECT 433.950 154.950 436.050 157.050 ;
        RECT 437.400 148.050 438.450 176.400 ;
        RECT 442.950 175.800 445.050 177.900 ;
        RECT 445.950 169.950 448.050 172.050 ;
        RECT 446.400 157.050 447.450 169.950 ;
        RECT 449.400 166.050 450.450 205.950 ;
        RECT 455.400 184.050 456.450 206.400 ;
        RECT 461.400 196.050 462.450 254.400 ;
        RECT 470.400 220.050 471.450 277.950 ;
        RECT 482.400 277.050 483.450 286.800 ;
        RECT 488.400 286.050 489.450 298.950 ;
        RECT 494.400 295.200 495.450 307.950 ;
        RECT 497.400 304.050 498.450 322.950 ;
        RECT 505.950 310.950 508.050 313.050 ;
        RECT 496.950 301.950 499.050 304.050 ;
        RECT 497.400 298.050 498.450 301.950 ;
        RECT 496.950 295.950 499.050 298.050 ;
        RECT 493.950 293.100 496.050 295.200 ;
        RECT 499.950 293.100 502.050 295.200 ;
        RECT 506.400 294.600 507.450 310.950 ;
        RECT 494.400 292.350 495.600 293.100 ;
        RECT 500.400 292.350 501.600 293.100 ;
        RECT 506.400 292.350 507.600 294.600 ;
        RECT 509.400 294.450 510.450 371.400 ;
        RECT 515.400 370.350 516.600 372.000 ;
        RECT 521.400 370.350 522.600 372.600 ;
        RECT 514.950 367.950 517.050 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 511.950 364.950 514.050 367.050 ;
        RECT 518.400 366.900 519.600 367.650 ;
        RECT 512.400 340.050 513.450 364.950 ;
        RECT 517.950 364.800 520.050 366.900 ;
        RECT 523.950 358.950 526.050 361.050 ;
        RECT 511.950 337.950 514.050 340.050 ;
        RECT 517.950 338.100 520.050 340.200 ;
        RECT 524.400 339.600 525.450 358.950 ;
        RECT 518.400 337.350 519.600 338.100 ;
        RECT 524.400 337.350 525.600 339.600 ;
        RECT 527.400 339.450 528.450 403.950 ;
        RECT 530.400 403.050 531.450 416.100 ;
        RECT 532.950 415.950 535.050 421.050 ;
        RECT 538.950 416.100 541.050 418.200 ;
        RECT 544.950 417.000 547.050 421.050 ;
        RECT 548.400 418.050 549.450 436.950 ;
        RECT 557.400 430.050 558.450 443.400 ;
        RECT 563.400 436.050 564.450 508.950 ;
        RECT 568.950 499.950 571.050 502.050 ;
        RECT 565.950 496.950 568.050 499.050 ;
        RECT 566.400 481.050 567.450 496.950 ;
        RECT 569.400 489.450 570.450 499.950 ;
        RECT 575.400 495.600 576.450 514.950 ;
        RECT 575.400 493.350 576.600 495.600 ;
        RECT 572.100 490.950 574.200 493.050 ;
        RECT 575.400 490.950 577.500 493.050 ;
        RECT 580.800 490.950 582.900 493.050 ;
        RECT 572.400 489.450 573.600 490.650 ;
        RECT 569.400 488.400 573.600 489.450 ;
        RECT 581.400 488.400 582.600 490.650 ;
        RECT 584.400 490.050 585.450 556.950 ;
        RECT 590.400 553.050 591.450 562.950 ;
        RECT 593.400 562.050 594.450 566.400 ;
        RECT 595.950 565.950 598.050 568.050 ;
        RECT 592.950 559.950 595.050 562.050 ;
        RECT 589.950 550.950 592.050 553.050 ;
        RECT 590.400 528.600 591.450 550.950 ;
        RECT 596.400 535.050 597.450 565.950 ;
        RECT 599.400 562.050 600.450 586.950 ;
        RECT 598.950 559.950 601.050 562.050 ;
        RECT 598.950 550.950 601.050 553.050 ;
        RECT 595.950 532.950 598.050 535.050 ;
        RECT 590.400 526.350 591.600 528.600 ;
        RECT 595.950 528.450 598.050 529.200 ;
        RECT 599.400 528.450 600.450 550.950 ;
        RECT 602.400 544.050 603.450 592.950 ;
        RECT 605.400 556.050 606.450 613.950 ;
        RECT 608.400 598.050 609.450 634.950 ;
        RECT 610.950 631.950 613.050 634.050 ;
        RECT 622.950 631.950 625.050 634.050 ;
        RECT 611.400 607.050 612.450 631.950 ;
        RECT 610.950 604.950 613.050 607.050 ;
        RECT 616.950 606.000 619.050 610.050 ;
        RECT 623.400 607.050 624.450 631.950 ;
        RECT 632.400 613.050 633.450 640.950 ;
        RECT 635.400 628.050 636.450 644.400 ;
        RECT 641.400 637.050 642.450 664.950 ;
        RECT 652.950 661.950 655.050 664.050 ;
        RECT 643.950 652.950 646.050 655.050 ;
        RECT 640.950 634.950 643.050 637.050 ;
        RECT 644.400 634.050 645.450 652.950 ;
        RECT 653.400 651.600 654.450 661.950 ;
        RECT 671.400 654.450 672.450 670.800 ;
        RECT 683.400 667.050 684.450 679.950 ;
        RECT 698.400 673.050 699.450 694.950 ;
        RECT 701.400 677.400 702.900 696.300 ;
        RECT 705.300 690.300 706.500 696.300 ;
        RECT 704.400 688.200 706.500 690.300 ;
        RECT 701.400 675.300 703.500 677.400 ;
        RECT 688.950 670.950 691.050 673.050 ;
        RECT 697.950 670.950 700.050 673.050 ;
        RECT 702.300 671.700 703.500 675.300 ;
        RECT 705.300 671.700 706.500 688.200 ;
        RECT 707.700 693.300 709.800 695.400 ;
        RECT 707.700 671.700 708.900 693.300 ;
        RECT 713.400 681.600 714.450 700.950 ;
        RECT 724.200 696.300 726.300 698.400 ;
        RECT 716.400 691.800 718.500 693.900 ;
        RECT 721.800 693.300 723.900 695.400 ;
        RECT 716.400 685.200 717.300 691.800 ;
        RECT 722.100 686.100 723.300 693.300 ;
        RECT 724.800 691.500 726.300 696.300 ;
        RECT 727.200 693.300 729.300 698.400 ;
        RECT 724.800 689.400 726.900 691.500 ;
        RECT 716.400 683.100 718.500 685.200 ;
        RECT 721.800 684.000 723.900 686.100 ;
        RECT 713.400 679.350 714.600 681.600 ;
        RECT 712.800 676.950 714.900 679.050 ;
        RECT 716.400 672.600 717.300 683.100 ;
        RECT 719.100 676.500 721.200 678.600 ;
        RECT 682.950 664.950 685.050 667.050 ;
        RECT 676.950 661.950 679.050 664.050 ;
        RECT 677.400 655.050 678.450 661.950 ;
        RECT 671.400 653.400 675.450 654.450 ;
        RECT 674.400 651.600 675.450 653.400 ;
        RECT 676.950 652.950 679.050 655.050 ;
        RECT 653.400 649.350 654.600 651.600 ;
        RECT 674.400 649.350 675.600 651.600 ;
        RECT 679.950 650.100 682.050 652.200 ;
        RECT 689.400 652.050 690.450 670.950 ;
        RECT 701.700 669.600 703.800 671.700 ;
        RECT 704.700 669.600 706.800 671.700 ;
        RECT 707.700 669.600 709.800 671.700 ;
        RECT 715.800 670.500 717.900 672.600 ;
        RECT 722.100 671.700 723.300 684.000 ;
        RECT 724.800 671.700 726.300 689.400 ;
        RECT 728.100 671.700 729.300 693.300 ;
        RECT 721.200 669.600 723.300 671.700 ;
        RECT 724.200 669.600 726.300 671.700 ;
        RECT 727.200 669.600 729.300 671.700 ;
        RECT 730.200 696.300 732.300 698.400 ;
        RECT 730.200 691.500 731.700 696.300 ;
        RECT 730.200 689.400 732.300 691.500 ;
        RECT 730.200 671.700 731.700 689.400 ;
        RECT 730.200 669.600 732.300 671.700 ;
        RECT 734.400 667.050 735.450 722.400 ;
        RECT 748.950 721.800 751.050 723.900 ;
        RECT 742.950 688.950 745.050 691.050 ;
        RECT 739.800 682.950 741.900 685.050 ;
        RECT 740.400 680.400 741.600 682.650 ;
        RECT 740.400 676.050 741.450 680.400 ;
        RECT 739.950 673.950 742.050 676.050 ;
        RECT 706.950 664.950 709.050 667.050 ;
        RECT 718.950 664.950 721.050 667.050 ;
        RECT 733.950 664.950 736.050 667.050 ;
        RECT 680.400 649.350 681.600 650.100 ;
        RECT 685.950 649.950 688.050 652.050 ;
        RECT 688.950 649.950 691.050 652.050 ;
        RECT 694.950 650.100 697.050 652.200 ;
        RECT 700.950 650.100 703.050 652.200 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 650.400 644.400 651.600 646.650 ;
        RECT 656.400 644.400 657.600 646.650 ;
        RECT 671.400 645.000 672.600 646.650 ;
        RECT 677.400 645.900 678.600 646.650 ;
        RECT 650.400 637.050 651.450 644.400 ;
        RECT 649.950 634.950 652.050 637.050 ;
        RECT 643.950 631.950 646.050 634.050 ;
        RECT 640.950 628.950 643.050 631.050 ;
        RECT 634.950 625.950 637.050 628.050 ;
        RECT 631.950 610.950 634.050 613.050 ;
        RECT 625.950 607.950 628.050 610.050 ;
        RECT 617.400 604.350 618.600 606.000 ;
        RECT 622.950 604.950 625.050 607.050 ;
        RECT 613.950 601.950 616.050 604.050 ;
        RECT 616.950 601.950 619.050 604.050 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 610.950 598.950 613.050 601.050 ;
        RECT 614.400 599.400 615.600 601.650 ;
        RECT 620.400 599.400 621.600 601.650 ;
        RECT 626.400 600.450 627.450 607.950 ;
        RECT 634.950 606.000 637.050 610.050 ;
        RECT 641.400 607.200 642.450 628.950 ;
        RECT 652.950 625.950 655.050 628.050 ;
        RECT 635.400 604.350 636.600 606.000 ;
        RECT 640.950 605.100 643.050 607.200 ;
        RECT 649.950 605.100 652.050 607.200 ;
        RECT 641.400 604.350 642.600 605.100 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 623.400 599.400 627.450 600.450 ;
        RECT 607.950 595.950 610.050 598.050 ;
        RECT 611.400 594.450 612.450 598.950 ;
        RECT 608.400 593.400 612.450 594.450 ;
        RECT 608.400 573.600 609.450 593.400 ;
        RECT 614.400 589.050 615.450 599.400 ;
        RECT 616.950 595.950 619.050 598.050 ;
        RECT 620.400 597.450 621.450 599.400 ;
        RECT 623.400 597.450 624.450 599.400 ;
        RECT 628.950 598.950 631.050 601.050 ;
        RECT 632.400 599.400 633.600 601.650 ;
        RECT 638.400 600.900 639.600 601.650 ;
        RECT 620.400 596.400 624.450 597.450 ;
        RECT 613.950 586.950 616.050 589.050 ;
        RECT 608.400 571.350 609.600 573.600 ;
        RECT 608.400 568.950 610.500 571.050 ;
        RECT 613.800 568.950 615.900 571.050 ;
        RECT 614.400 566.400 615.600 568.650 ;
        RECT 614.400 562.050 615.450 566.400 ;
        RECT 613.950 559.950 616.050 562.050 ;
        RECT 604.950 553.950 607.050 556.050 ;
        RECT 617.400 550.050 618.450 595.950 ;
        RECT 619.950 580.950 622.050 583.050 ;
        RECT 616.950 547.950 619.050 550.050 ;
        RECT 601.950 541.950 604.050 544.050 ;
        RECT 595.950 527.400 600.450 528.450 ;
        RECT 595.950 527.100 598.050 527.400 ;
        RECT 596.400 526.350 597.600 527.100 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 593.400 521.400 594.600 523.650 ;
        RECT 589.950 517.950 592.050 520.050 ;
        RECT 590.400 511.050 591.450 517.950 ;
        RECT 593.400 517.050 594.450 521.400 ;
        RECT 592.950 514.950 595.050 517.050 ;
        RECT 589.950 508.950 592.050 511.050 ;
        RECT 586.950 505.950 589.050 508.050 ;
        RECT 581.400 484.050 582.450 488.400 ;
        RECT 583.950 487.950 586.050 490.050 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 580.950 481.950 583.050 484.050 ;
        RECT 565.950 478.950 568.050 481.050 ;
        RECT 568.950 469.950 571.050 472.050 ;
        RECT 565.950 460.950 568.050 463.050 ;
        RECT 566.400 444.900 567.450 460.950 ;
        RECT 569.400 457.050 570.450 469.950 ;
        RECT 568.950 454.950 571.050 457.050 ;
        RECT 572.400 451.200 573.450 481.950 ;
        RECT 583.950 472.950 586.050 475.050 ;
        RECT 577.950 454.950 580.050 457.050 ;
        RECT 571.950 449.100 574.050 451.200 ;
        RECT 578.400 450.600 579.450 454.950 ;
        RECT 584.400 451.050 585.450 472.950 ;
        RECT 587.400 460.050 588.450 505.950 ;
        RECT 602.400 505.050 603.450 541.950 ;
        RECT 607.950 527.100 610.050 529.200 ;
        RECT 608.400 526.350 609.600 527.100 ;
        RECT 607.950 523.950 610.050 526.050 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 611.400 521.400 612.600 523.650 ;
        RECT 607.950 508.950 610.050 511.050 ;
        RECT 592.950 502.950 595.050 505.050 ;
        RECT 601.950 502.950 604.050 505.050 ;
        RECT 593.400 495.600 594.450 502.950 ;
        RECT 593.400 493.350 594.600 495.600 ;
        RECT 598.950 494.100 601.050 496.200 ;
        RECT 599.400 493.350 600.600 494.100 ;
        RECT 604.950 493.950 607.050 499.050 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 589.950 487.950 592.050 490.050 ;
        RECT 596.400 489.900 597.600 490.650 ;
        RECT 586.950 457.950 589.050 460.050 ;
        RECT 572.400 448.350 573.600 449.100 ;
        RECT 578.400 448.350 579.600 450.600 ;
        RECT 584.400 448.950 589.050 451.050 ;
        RECT 584.400 448.350 585.600 448.950 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 577.950 445.950 580.050 448.050 ;
        RECT 580.950 445.950 583.050 448.050 ;
        RECT 583.950 445.950 586.050 448.050 ;
        RECT 575.400 444.900 576.600 445.650 ;
        RECT 581.400 444.900 582.600 445.650 ;
        RECT 565.950 442.800 568.050 444.900 ;
        RECT 574.950 442.800 577.050 444.900 ;
        RECT 580.950 442.800 583.050 444.900 ;
        RECT 586.950 442.950 589.050 445.050 ;
        RECT 581.400 439.050 582.450 442.800 ;
        RECT 574.950 436.950 577.050 439.050 ;
        RECT 580.950 436.950 583.050 439.050 ;
        RECT 562.950 433.950 565.050 436.050 ;
        RECT 571.950 433.950 574.050 436.050 ;
        RECT 562.950 430.800 565.050 432.900 ;
        RECT 556.950 427.950 559.050 430.050 ;
        RECT 550.950 424.950 553.050 427.050 ;
        RECT 539.400 415.350 540.600 416.100 ;
        RECT 545.400 415.350 546.600 417.000 ;
        RECT 547.950 415.950 550.050 418.050 ;
        RECT 535.950 412.950 538.050 415.050 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 532.950 409.950 535.050 412.050 ;
        RECT 536.400 411.000 537.600 412.650 ;
        RECT 542.400 411.900 543.600 412.650 ;
        RECT 551.400 412.050 552.450 424.950 ;
        RECT 553.950 421.950 556.050 424.050 ;
        RECT 529.950 400.950 532.050 403.050 ;
        RECT 533.400 372.450 534.450 409.950 ;
        RECT 535.950 406.950 538.050 411.000 ;
        RECT 541.950 409.800 544.050 411.900 ;
        RECT 550.950 409.950 553.050 412.050 ;
        RECT 550.950 406.800 553.050 408.900 ;
        RECT 554.400 408.450 555.450 421.950 ;
        RECT 563.400 417.600 564.450 430.800 ;
        RECT 563.400 415.350 564.600 417.600 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 560.400 412.050 561.600 412.650 ;
        RECT 556.950 410.400 561.600 412.050 ;
        RECT 566.400 411.000 567.600 412.650 ;
        RECT 556.950 409.950 561.000 410.400 ;
        RECT 554.400 407.400 558.450 408.450 ;
        RECT 538.950 391.950 541.050 394.050 ;
        RECT 547.950 391.950 550.050 394.050 ;
        RECT 530.400 371.400 534.450 372.450 ;
        RECT 539.400 372.600 540.450 391.950 ;
        RECT 548.400 388.050 549.450 391.950 ;
        RECT 547.950 385.950 550.050 388.050 ;
        RECT 551.400 385.050 552.450 406.800 ;
        RECT 550.950 382.950 553.050 385.050 ;
        RECT 544.950 379.950 547.050 382.050 ;
        RECT 553.950 379.950 556.050 382.050 ;
        RECT 545.400 372.600 546.450 379.950 ;
        RECT 530.400 343.050 531.450 371.400 ;
        RECT 539.400 370.350 540.600 372.600 ;
        RECT 545.400 370.350 546.600 372.600 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 536.400 366.900 537.600 367.650 ;
        RECT 535.950 364.800 538.050 366.900 ;
        RECT 542.400 365.400 543.600 367.650 ;
        RECT 548.400 365.400 549.600 367.650 ;
        RECT 554.400 366.900 555.450 379.950 ;
        RECT 542.400 355.050 543.450 365.400 ;
        RECT 544.950 355.950 547.050 358.050 ;
        RECT 541.950 352.950 544.050 355.050 ;
        RECT 538.950 351.450 541.050 352.050 ;
        RECT 545.400 351.450 546.450 355.950 ;
        RECT 538.950 350.400 546.450 351.450 ;
        RECT 538.950 349.950 541.050 350.400 ;
        RECT 544.950 346.950 547.050 349.050 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 527.400 338.400 531.450 339.450 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 511.950 331.950 514.050 334.050 ;
        RECT 515.400 333.000 516.600 334.650 ;
        RECT 521.400 333.000 522.600 334.650 ;
        RECT 512.400 301.050 513.450 331.950 ;
        RECT 514.950 328.950 517.050 333.000 ;
        RECT 520.950 328.950 523.050 333.000 ;
        RECT 520.950 322.950 523.050 325.050 ;
        RECT 521.400 316.050 522.450 322.950 ;
        RECT 520.950 313.950 523.050 316.050 ;
        RECT 511.950 298.950 514.050 301.050 ;
        RECT 521.400 294.600 522.450 313.950 ;
        RECT 526.950 310.950 529.050 313.050 ;
        RECT 527.400 294.600 528.450 310.950 ;
        RECT 530.400 301.050 531.450 338.400 ;
        RECT 538.950 338.100 541.050 340.200 ;
        RECT 545.400 339.600 546.450 346.950 ;
        RECT 548.400 346.050 549.450 365.400 ;
        RECT 553.950 364.800 556.050 366.900 ;
        RECT 557.400 352.050 558.450 407.400 ;
        RECT 565.950 406.950 568.050 411.000 ;
        RECT 559.950 397.950 562.050 400.050 ;
        RECT 572.400 399.450 573.450 433.950 ;
        RECT 575.400 418.050 576.450 436.950 ;
        RECT 580.950 424.950 583.050 427.050 ;
        RECT 574.950 415.950 577.050 418.050 ;
        RECT 581.400 417.600 582.450 424.950 ;
        RECT 587.400 421.050 588.450 442.950 ;
        RECT 586.950 418.950 589.050 421.050 ;
        RECT 581.400 415.350 582.600 417.600 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 580.950 412.950 583.050 415.050 ;
        RECT 583.950 412.950 586.050 415.050 ;
        RECT 578.400 410.400 579.600 412.650 ;
        RECT 584.400 411.900 585.600 412.650 ;
        RECT 578.400 406.050 579.450 410.400 ;
        RECT 583.950 409.800 586.050 411.900 ;
        RECT 580.950 408.750 585.000 409.050 ;
        RECT 580.950 406.950 586.050 408.750 ;
        RECT 583.950 406.650 586.050 406.950 ;
        RECT 577.950 403.950 580.050 406.050 ;
        RECT 582.000 402.450 586.050 403.050 ;
        RECT 581.400 400.950 586.050 402.450 ;
        RECT 586.950 400.950 589.050 403.050 ;
        RECT 572.400 398.400 576.450 399.450 ;
        RECT 560.400 388.050 561.450 397.950 ;
        RECT 571.950 394.950 574.050 397.050 ;
        RECT 559.950 385.950 562.050 388.050 ;
        RECT 568.950 385.950 571.050 388.050 ;
        RECT 565.950 371.100 568.050 373.200 ;
        RECT 569.400 373.050 570.450 385.950 ;
        RECT 566.400 370.350 567.600 371.100 ;
        RECT 568.950 370.950 571.050 373.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 563.400 366.900 564.600 367.650 ;
        RECT 562.950 364.800 565.050 366.900 ;
        RECT 572.400 366.450 573.450 394.950 ;
        RECT 569.400 365.400 573.450 366.450 ;
        RECT 550.950 349.950 553.050 352.050 ;
        RECT 556.950 349.950 559.050 352.050 ;
        RECT 547.950 343.950 550.050 346.050 ;
        RECT 548.400 340.050 549.450 343.950 ;
        RECT 539.400 337.350 540.600 338.100 ;
        RECT 545.400 337.350 546.600 339.600 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 535.950 334.950 538.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 536.400 333.900 537.600 334.650 ;
        RECT 535.950 331.800 538.050 333.900 ;
        RECT 542.400 332.400 543.600 334.650 ;
        RECT 532.950 328.950 535.050 331.050 ;
        RECT 538.950 328.950 541.050 331.050 ;
        RECT 529.950 298.950 532.050 301.050 ;
        RECT 509.400 293.400 513.450 294.450 ;
        RECT 493.950 289.950 496.050 292.050 ;
        RECT 496.950 289.950 499.050 292.050 ;
        RECT 499.950 289.950 502.050 292.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 497.400 288.000 498.600 289.650 ;
        RECT 503.400 288.900 504.600 289.650 ;
        RECT 487.950 283.950 490.050 286.050 ;
        RECT 496.950 283.950 499.050 288.000 ;
        RECT 502.950 286.800 505.050 288.900 ;
        RECT 508.950 286.950 511.050 289.050 ;
        RECT 481.950 274.950 484.050 277.050 ;
        RECT 509.400 274.050 510.450 286.950 ;
        RECT 493.950 271.950 496.050 274.050 ;
        RECT 508.950 271.950 511.050 274.050 ;
        RECT 484.950 265.950 487.050 268.050 ;
        RECT 478.950 261.000 481.050 265.050 ;
        RECT 485.400 262.200 486.450 265.950 ;
        RECT 479.400 259.350 480.600 261.000 ;
        RECT 484.950 260.100 487.050 262.200 ;
        RECT 485.400 259.350 486.600 260.100 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 476.400 254.400 477.600 256.650 ;
        RECT 482.400 254.400 483.600 256.650 ;
        RECT 488.400 255.900 489.600 256.650 ;
        RECT 476.400 238.050 477.450 254.400 ;
        RECT 478.950 241.950 481.050 244.050 ;
        RECT 475.950 235.950 478.050 238.050 ;
        RECT 472.950 232.950 475.050 235.050 ;
        RECT 473.400 220.050 474.450 232.950 ;
        RECT 475.950 229.950 478.050 232.050 ;
        RECT 463.950 217.950 466.050 220.050 ;
        RECT 469.800 217.950 471.900 220.050 ;
        RECT 472.950 217.950 475.050 220.050 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 464.400 190.050 465.450 217.950 ;
        RECT 476.400 217.200 477.450 229.950 ;
        RECT 466.950 216.600 471.000 217.050 ;
        RECT 466.950 214.950 471.600 216.600 ;
        RECT 475.950 215.100 478.050 217.200 ;
        RECT 479.400 216.450 480.450 241.950 ;
        RECT 482.400 229.050 483.450 254.400 ;
        RECT 487.950 253.800 490.050 255.900 ;
        RECT 494.400 253.050 495.450 271.950 ;
        RECT 502.950 260.100 505.050 262.200 ;
        RECT 503.400 259.350 504.600 260.100 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 496.950 253.950 499.050 256.050 ;
        RECT 500.400 254.400 501.600 256.650 ;
        RECT 506.400 256.050 507.600 256.650 ;
        RECT 506.400 254.400 511.050 256.050 ;
        RECT 493.950 250.950 496.050 253.050 ;
        RECT 493.950 247.800 496.050 249.900 ;
        RECT 481.950 226.950 484.050 229.050 ;
        RECT 479.400 215.400 483.450 216.450 ;
        RECT 470.400 214.350 471.600 214.950 ;
        RECT 476.400 214.350 477.600 215.100 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 472.950 211.950 475.050 214.050 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 466.950 208.950 469.050 211.050 ;
        RECT 473.400 209.400 474.600 211.650 ;
        RECT 482.400 210.900 483.450 215.400 ;
        RECT 487.950 215.100 490.050 217.200 ;
        RECT 494.400 216.600 495.450 247.800 ;
        RECT 497.400 244.050 498.450 253.950 ;
        RECT 496.950 241.950 499.050 244.050 ;
        RECT 500.400 232.050 501.450 254.400 ;
        RECT 507.000 253.950 511.050 254.400 ;
        RECT 502.800 250.950 504.900 253.050 ;
        RECT 505.950 250.950 508.050 253.050 ;
        RECT 499.950 229.950 502.050 232.050 ;
        RECT 500.400 223.050 501.450 229.950 ;
        RECT 499.950 220.950 502.050 223.050 ;
        RECT 488.400 214.350 489.600 215.100 ;
        RECT 494.400 214.350 495.600 216.600 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 467.400 199.050 468.450 208.950 ;
        RECT 473.400 205.050 474.450 209.400 ;
        RECT 481.950 208.800 484.050 210.900 ;
        RECT 491.400 209.400 492.600 211.650 ;
        RECT 497.400 210.900 498.600 211.650 ;
        RECT 472.950 202.950 475.050 205.050 ;
        RECT 466.950 196.950 469.050 199.050 ;
        RECT 472.950 196.950 475.050 199.050 ;
        RECT 457.950 187.950 460.050 190.050 ;
        RECT 463.950 187.950 466.050 190.050 ;
        RECT 469.950 187.950 472.050 190.050 ;
        RECT 451.950 181.950 454.050 184.050 ;
        RECT 454.950 181.950 457.050 184.050 ;
        RECT 458.400 183.600 459.450 187.950 ;
        RECT 452.400 172.050 453.450 181.950 ;
        RECT 458.400 181.350 459.600 183.600 ;
        RECT 463.950 182.100 466.050 184.200 ;
        RECT 470.400 184.050 471.450 187.950 ;
        RECT 464.400 181.350 465.600 182.100 ;
        RECT 469.950 181.950 472.050 184.050 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 463.950 178.950 466.050 181.050 ;
        RECT 466.950 178.950 469.050 181.050 ;
        RECT 454.950 175.950 457.050 178.050 ;
        RECT 461.400 176.400 462.600 178.650 ;
        RECT 467.400 177.000 468.600 178.650 ;
        RECT 451.950 169.950 454.050 172.050 ;
        RECT 455.400 169.050 456.450 175.950 ;
        RECT 454.950 166.950 457.050 169.050 ;
        RECT 448.950 163.950 451.050 166.050 ;
        RECT 461.400 160.050 462.450 176.400 ;
        RECT 466.950 172.950 469.050 177.000 ;
        RECT 469.950 175.950 472.050 178.050 ;
        RECT 466.950 166.950 469.050 169.050 ;
        RECT 460.800 157.950 462.900 160.050 ;
        RECT 463.950 157.950 466.050 160.050 ;
        RECT 445.950 154.950 448.050 157.050 ;
        RECT 464.400 151.050 465.450 157.950 ;
        RECT 463.950 148.950 466.050 151.050 ;
        RECT 436.950 145.950 439.050 148.050 ;
        RECT 433.950 136.950 436.050 142.050 ;
        RECT 441.000 138.600 445.050 139.050 ;
        RECT 440.400 136.950 445.050 138.600 ;
        RECT 451.950 138.600 456.000 139.050 ;
        RECT 451.950 138.450 456.600 138.600 ;
        RECT 449.400 137.400 456.600 138.450 ;
        RECT 460.950 138.000 463.050 142.050 ;
        RECT 467.400 139.050 468.450 166.950 ;
        RECT 470.400 139.050 471.450 175.950 ;
        RECT 473.400 175.050 474.450 196.950 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 472.950 172.950 475.050 175.050 ;
        RECT 476.400 145.050 477.450 193.950 ;
        RECT 491.400 186.450 492.450 209.400 ;
        RECT 496.950 208.800 499.050 210.900 ;
        RECT 493.950 196.950 496.050 199.050 ;
        RECT 488.400 185.400 492.450 186.450 ;
        RECT 481.950 182.100 484.050 184.200 ;
        RECT 488.400 183.600 489.450 185.400 ;
        RECT 494.400 184.050 495.450 196.950 ;
        RECT 499.950 193.950 502.050 196.050 ;
        RECT 496.950 187.950 499.050 190.050 ;
        RECT 482.400 181.350 483.600 182.100 ;
        RECT 488.400 181.350 489.600 183.600 ;
        RECT 493.950 181.950 496.050 184.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 484.950 178.950 487.050 181.050 ;
        RECT 487.950 178.950 490.050 181.050 ;
        RECT 490.950 178.950 493.050 181.050 ;
        RECT 478.950 175.950 481.050 178.050 ;
        RECT 485.400 176.400 486.600 178.650 ;
        RECT 491.400 177.900 492.600 178.650 ;
        RECT 479.400 151.050 480.450 175.950 ;
        RECT 485.400 172.050 486.450 176.400 ;
        RECT 490.950 175.800 493.050 177.900 ;
        RECT 493.950 175.950 496.050 178.050 ;
        RECT 497.400 177.900 498.450 187.950 ;
        RECT 500.400 184.050 501.450 193.950 ;
        RECT 503.400 187.050 504.450 250.950 ;
        RECT 506.400 226.050 507.450 250.950 ;
        RECT 512.400 238.050 513.450 293.400 ;
        RECT 521.400 292.350 522.600 294.600 ;
        RECT 527.400 292.350 528.600 294.600 ;
        RECT 517.950 289.950 520.050 292.050 ;
        RECT 520.950 289.950 523.050 292.050 ;
        RECT 523.950 289.950 526.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 518.400 287.400 519.600 289.650 ;
        RECT 524.400 288.900 525.600 289.650 ;
        RECT 514.950 283.950 517.050 286.050 ;
        RECT 515.400 256.050 516.450 283.950 ;
        RECT 518.400 280.050 519.450 287.400 ;
        RECT 523.950 286.800 526.050 288.900 ;
        RECT 533.400 288.450 534.450 328.950 ;
        RECT 539.400 319.050 540.450 328.950 ;
        RECT 542.400 328.050 543.450 332.400 ;
        RECT 541.950 325.950 544.050 328.050 ;
        RECT 551.400 325.050 552.450 349.950 ;
        RECT 565.950 346.950 568.050 349.050 ;
        RECT 559.950 343.950 562.050 346.050 ;
        RECT 560.400 339.600 561.450 343.950 ;
        RECT 566.400 340.050 567.450 346.950 ;
        RECT 560.400 337.350 561.600 339.600 ;
        RECT 565.950 337.950 568.050 340.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 557.400 332.400 558.600 334.650 ;
        RECT 563.400 332.400 564.600 334.650 ;
        RECT 569.400 333.450 570.450 365.400 ;
        RECT 575.400 364.050 576.450 398.400 ;
        RECT 581.400 388.050 582.450 400.950 ;
        RECT 583.950 391.950 586.050 394.050 ;
        RECT 580.950 385.950 583.050 388.050 ;
        RECT 584.400 382.050 585.450 391.950 ;
        RECT 587.400 391.050 588.450 400.950 ;
        RECT 590.400 397.050 591.450 487.950 ;
        RECT 595.950 487.800 598.050 489.900 ;
        RECT 602.400 488.400 603.600 490.650 ;
        RECT 602.400 484.050 603.450 488.400 ;
        RECT 601.950 481.950 604.050 484.050 ;
        RECT 608.400 474.450 609.450 508.950 ;
        RECT 611.400 505.050 612.450 521.400 ;
        RECT 610.950 502.950 613.050 505.050 ;
        RECT 617.400 499.050 618.450 547.950 ;
        RECT 620.400 538.050 621.450 580.950 ;
        RECT 623.400 568.050 624.450 596.400 ;
        RECT 625.950 592.950 628.050 595.050 ;
        RECT 626.400 577.050 627.450 592.950 ;
        RECT 629.400 583.050 630.450 598.950 ;
        RECT 632.400 592.050 633.450 599.400 ;
        RECT 637.950 598.800 640.050 600.900 ;
        RECT 644.400 599.400 645.600 601.650 ;
        RECT 650.400 601.050 651.450 605.100 ;
        RECT 634.950 595.950 637.050 598.050 ;
        RECT 631.950 589.950 634.050 592.050 ;
        RECT 635.400 588.450 636.450 595.950 ;
        RECT 632.400 587.400 636.450 588.450 ;
        RECT 628.950 580.950 631.050 583.050 ;
        RECT 625.950 574.950 628.050 577.050 ;
        RECT 632.400 574.200 633.450 587.400 ;
        RECT 644.400 586.050 645.450 599.400 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 653.400 595.050 654.450 625.950 ;
        RECT 656.400 625.050 657.450 644.400 ;
        RECT 658.950 640.950 664.050 643.050 ;
        RECT 670.950 640.950 673.050 645.000 ;
        RECT 676.950 643.800 679.050 645.900 ;
        RECT 682.950 643.950 685.050 646.050 ;
        RECT 667.950 637.950 670.050 640.050 ;
        RECT 655.950 622.950 658.050 625.050 ;
        RECT 656.400 607.050 657.450 622.950 ;
        RECT 668.400 621.450 669.450 637.950 ;
        RECT 665.400 620.400 669.450 621.450 ;
        RECT 655.950 604.950 658.050 607.050 ;
        RECT 658.950 605.100 661.050 607.200 ;
        RECT 665.400 606.600 666.450 620.400 ;
        RECT 677.400 613.050 678.450 643.800 ;
        RECT 676.950 610.950 679.050 613.050 ;
        RECT 683.400 610.200 684.450 643.950 ;
        RECT 686.400 640.050 687.450 649.950 ;
        RECT 695.400 649.350 696.600 650.100 ;
        RECT 701.400 649.350 702.600 650.100 ;
        RECT 691.950 646.950 694.050 649.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 692.400 645.900 693.600 646.650 ;
        RECT 691.950 643.800 694.050 645.900 ;
        RECT 698.400 644.400 699.600 646.650 ;
        RECT 698.400 642.450 699.450 644.400 ;
        RECT 695.400 641.400 699.450 642.450 ;
        RECT 685.950 637.950 688.050 640.050 ;
        RECT 695.400 631.050 696.450 641.400 ;
        RECT 694.950 628.950 697.050 631.050 ;
        RECT 670.950 607.950 673.050 610.050 ;
        RECT 682.950 608.100 685.050 610.200 ;
        RECT 659.400 604.350 660.600 605.100 ;
        RECT 665.400 604.350 666.600 606.600 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 655.950 598.950 658.050 601.050 ;
        RECT 662.400 599.400 663.600 601.650 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 643.950 583.950 646.050 586.050 ;
        RECT 631.950 572.100 634.050 574.200 ;
        RECT 637.950 572.100 640.050 574.200 ;
        RECT 643.950 572.100 646.050 574.200 ;
        RECT 632.400 571.350 633.600 572.100 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 622.950 565.950 625.050 568.050 ;
        RECT 629.400 567.900 630.600 568.650 ;
        RECT 628.950 565.800 631.050 567.900 ;
        RECT 619.950 535.950 622.050 538.050 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 629.400 528.600 630.450 565.800 ;
        RECT 638.400 553.050 639.450 572.100 ;
        RECT 644.400 571.350 645.600 572.100 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 647.400 567.900 648.600 568.650 ;
        RECT 646.950 565.800 649.050 567.900 ;
        RECT 637.800 550.950 639.900 553.050 ;
        RECT 640.950 550.950 643.050 553.050 ;
        RECT 610.950 496.950 613.050 499.050 ;
        RECT 616.950 496.950 619.050 499.050 ;
        RECT 620.400 498.450 621.450 527.100 ;
        RECT 629.400 526.350 630.600 528.600 ;
        RECT 634.950 527.100 637.050 529.200 ;
        RECT 635.400 526.350 636.600 527.100 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 631.950 523.950 634.050 526.050 ;
        RECT 634.950 523.950 637.050 526.050 ;
        RECT 626.400 521.400 627.600 523.650 ;
        RECT 632.400 522.900 633.600 523.650 ;
        RECT 641.400 523.050 642.450 550.950 ;
        RECT 643.950 541.950 646.050 544.050 ;
        RECT 622.950 514.950 625.050 517.050 ;
        RECT 623.400 501.450 624.450 514.950 ;
        RECT 626.400 514.050 627.450 521.400 ;
        RECT 631.950 520.800 634.050 522.900 ;
        RECT 640.950 520.950 643.050 523.050 ;
        RECT 644.400 522.450 645.450 541.950 ;
        RECT 647.400 529.200 648.450 565.800 ;
        RECT 653.400 565.050 654.450 592.950 ;
        RECT 652.950 562.950 655.050 565.050 ;
        RECT 656.400 562.050 657.450 598.950 ;
        RECT 662.400 595.050 663.450 599.400 ;
        RECT 671.400 598.050 672.450 607.950 ;
        RECT 673.950 604.950 676.050 607.050 ;
        RECT 682.950 604.950 685.050 607.050 ;
        RECT 688.950 605.100 691.050 607.200 ;
        RECT 670.950 595.950 673.050 598.050 ;
        RECT 674.400 595.050 675.450 604.950 ;
        RECT 683.400 604.350 684.600 604.950 ;
        RECT 689.400 604.350 690.600 605.100 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 680.400 599.400 681.600 601.650 ;
        RECT 686.400 600.900 687.600 601.650 ;
        RECT 695.400 601.050 696.450 628.950 ;
        RECT 707.400 625.050 708.450 664.950 ;
        RECT 719.400 651.600 720.450 664.950 ;
        RECT 743.400 657.450 744.450 688.950 ;
        RECT 748.800 682.950 750.900 685.050 ;
        RECT 749.400 681.900 750.600 682.650 ;
        RECT 755.400 681.900 756.450 730.950 ;
        RECT 758.400 730.050 759.450 733.950 ;
        RECT 757.950 727.950 760.050 730.050 ;
        RECT 761.400 729.600 762.450 736.950 ;
        RECT 761.400 727.350 762.600 729.600 ;
        RECT 766.950 728.100 769.050 730.200 ;
        RECT 775.950 728.100 778.050 730.200 ;
        RECT 782.400 729.600 783.450 749.400 ;
        RECT 785.400 739.050 786.450 755.400 ;
        RECT 796.950 754.800 799.050 756.900 ;
        RECT 806.400 756.000 807.600 757.650 ;
        RECT 812.400 756.900 813.600 757.650 ;
        RECT 787.950 751.950 793.050 754.050 ;
        RECT 805.950 748.950 808.050 756.000 ;
        RECT 811.950 754.800 814.050 756.900 ;
        RECT 821.400 754.050 822.450 761.100 ;
        RECT 814.950 751.950 817.050 754.050 ;
        RECT 820.950 751.950 823.050 754.050 ;
        RECT 784.950 736.950 787.050 739.050 ;
        RECT 805.950 736.950 808.050 739.050 ;
        RECT 767.400 727.350 768.600 728.100 ;
        RECT 760.950 724.950 763.050 727.050 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 764.400 722.400 765.600 724.650 ;
        RECT 770.400 723.000 771.600 724.650 ;
        RECT 760.950 685.950 763.050 688.050 ;
        RECT 748.950 679.800 751.050 681.900 ;
        RECT 754.950 679.800 757.050 681.900 ;
        RECT 761.400 664.050 762.450 685.950 ;
        RECT 764.400 685.050 765.450 722.400 ;
        RECT 769.950 718.950 772.050 723.000 ;
        RECT 776.400 709.050 777.450 728.100 ;
        RECT 782.400 727.350 783.600 729.600 ;
        RECT 787.950 728.100 790.050 730.200 ;
        RECT 788.400 727.350 789.600 728.100 ;
        RECT 799.950 727.950 802.050 730.050 ;
        RECT 806.400 729.600 807.450 736.950 ;
        RECT 811.950 733.950 814.050 736.050 ;
        RECT 812.400 730.050 813.450 733.950 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 787.950 724.950 790.050 727.050 ;
        RECT 790.950 724.950 793.050 727.050 ;
        RECT 785.400 723.900 786.600 724.650 ;
        RECT 784.950 721.800 787.050 723.900 ;
        RECT 791.400 723.000 792.600 724.650 ;
        RECT 781.950 720.750 786.000 721.050 ;
        RECT 781.950 718.950 787.050 720.750 ;
        RECT 790.950 718.950 793.050 723.000 ;
        RECT 784.950 718.650 787.050 718.950 ;
        RECT 775.950 706.950 778.050 709.050 ;
        RECT 784.950 706.950 787.050 709.050 ;
        RECT 769.950 697.950 772.050 700.050 ;
        RECT 781.950 697.950 784.050 700.050 ;
        RECT 770.400 691.050 771.450 697.950 ;
        RECT 775.950 691.950 778.050 694.050 ;
        RECT 769.950 688.950 772.050 691.050 ;
        RECT 763.950 682.950 766.050 685.050 ;
        RECT 770.400 684.600 771.450 688.950 ;
        RECT 776.400 688.050 777.450 691.950 ;
        RECT 770.400 682.350 771.600 684.600 ;
        RECT 775.950 684.000 778.050 688.050 ;
        RECT 776.400 682.350 777.600 684.000 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 767.400 678.900 768.600 679.650 ;
        RECT 773.400 678.900 774.600 679.650 ;
        RECT 766.950 676.800 769.050 678.900 ;
        RECT 772.950 676.800 775.050 678.900 ;
        RECT 778.950 676.800 781.050 678.900 ;
        RECT 779.400 667.050 780.450 676.800 ;
        RECT 778.950 664.950 781.050 667.050 ;
        RECT 751.950 661.950 754.050 664.050 ;
        RECT 760.950 661.950 763.050 664.050 ;
        RECT 743.400 655.200 744.600 657.450 ;
        RECT 738.900 651.900 741.000 653.700 ;
        RECT 742.800 652.800 744.900 654.900 ;
        RECT 746.100 654.300 748.200 656.400 ;
        RECT 719.400 649.350 720.600 651.600 ;
        RECT 737.400 650.700 746.100 651.900 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 734.100 646.950 736.200 649.050 ;
        RECT 716.400 645.900 717.600 646.650 ;
        RECT 715.950 643.800 718.050 645.900 ;
        RECT 722.400 644.400 723.600 646.650 ;
        RECT 734.400 645.450 735.600 646.650 ;
        RECT 731.400 644.400 735.600 645.450 ;
        RECT 722.400 640.050 723.450 644.400 ;
        RECT 721.950 637.950 724.050 640.050 ;
        RECT 731.400 631.050 732.450 644.400 ;
        RECT 737.400 641.700 738.300 650.700 ;
        RECT 744.000 649.800 746.100 650.700 ;
        RECT 747.000 648.900 747.900 654.300 ;
        RECT 749.400 651.450 750.600 651.600 ;
        RECT 752.400 651.450 753.450 661.950 ;
        RECT 772.950 655.950 775.050 658.050 ;
        RECT 773.400 655.200 774.600 655.950 ;
        RECT 768.900 651.900 771.000 653.700 ;
        RECT 772.800 652.800 774.900 654.900 ;
        RECT 776.100 654.300 778.200 656.400 ;
        RECT 782.400 655.050 783.450 697.950 ;
        RECT 785.400 676.050 786.450 706.950 ;
        RECT 800.400 706.050 801.450 727.950 ;
        RECT 806.400 727.350 807.600 729.600 ;
        RECT 811.950 727.950 814.050 730.050 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 809.400 722.400 810.600 724.650 ;
        RECT 802.950 718.950 805.050 721.050 ;
        RECT 803.400 714.450 804.450 718.950 ;
        RECT 805.950 717.450 808.050 721.050 ;
        RECT 809.400 718.050 810.450 722.400 ;
        RECT 815.400 721.050 816.450 751.950 ;
        RECT 820.950 739.950 823.050 742.050 ;
        RECT 821.400 733.050 822.450 739.950 ;
        RECT 824.400 733.050 825.450 772.950 ;
        RECT 827.400 763.050 828.450 775.950 ;
        RECT 826.950 760.950 829.050 763.050 ;
        RECT 832.950 761.100 835.050 763.200 ;
        RECT 838.950 761.100 841.050 763.200 ;
        RECT 844.950 761.100 847.050 763.200 ;
        RECT 833.400 760.350 834.600 761.100 ;
        RECT 839.400 760.350 840.600 761.100 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 838.950 757.950 841.050 760.050 ;
        RECT 826.950 754.950 829.050 757.050 ;
        RECT 830.400 755.400 831.600 757.650 ;
        RECT 836.400 755.400 837.600 757.650 ;
        RECT 827.400 751.050 828.450 754.950 ;
        RECT 826.950 748.950 829.050 751.050 ;
        RECT 830.400 747.450 831.450 755.400 ;
        RECT 827.400 746.400 831.450 747.450 ;
        RECT 827.400 736.050 828.450 746.400 ;
        RECT 836.400 745.050 837.450 755.400 ;
        RECT 838.950 751.950 841.050 754.050 ;
        RECT 835.950 742.950 838.050 745.050 ;
        RECT 829.950 739.950 832.050 742.050 ;
        RECT 826.950 733.950 829.050 736.050 ;
        RECT 820.800 730.950 822.900 733.050 ;
        RECT 823.950 730.950 826.050 733.050 ;
        RECT 830.400 729.600 831.450 739.950 ;
        RECT 835.950 736.950 838.050 739.050 ;
        RECT 836.400 730.050 837.450 736.950 ;
        RECT 824.400 729.450 825.600 729.600 ;
        RECT 818.400 728.400 825.600 729.450 ;
        RECT 814.950 718.950 817.050 721.050 ;
        RECT 808.950 717.450 811.050 718.050 ;
        RECT 805.950 717.000 811.050 717.450 ;
        RECT 806.400 716.400 811.050 717.000 ;
        RECT 808.950 715.950 811.050 716.400 ;
        RECT 803.400 713.400 807.450 714.450 ;
        RECT 799.950 703.950 802.050 706.050 ;
        RECT 799.950 697.950 802.050 700.050 ;
        RECT 793.950 691.950 796.050 694.050 ;
        RECT 794.400 684.600 795.450 691.950 ;
        RECT 800.400 684.600 801.450 697.950 ;
        RECT 794.400 682.350 795.600 684.600 ;
        RECT 800.400 682.350 801.600 684.600 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 791.400 678.000 792.600 679.650 ;
        RECT 797.400 678.900 798.600 679.650 ;
        RECT 784.950 673.950 787.050 676.050 ;
        RECT 790.950 673.950 793.050 678.000 ;
        RECT 796.950 676.800 799.050 678.900 ;
        RECT 797.400 667.050 798.450 676.800 ;
        RECT 806.400 673.050 807.450 713.400 ;
        RECT 818.400 712.050 819.450 728.400 ;
        RECT 824.400 727.350 825.600 728.400 ;
        RECT 830.400 727.350 831.600 729.600 ;
        RECT 835.950 727.950 838.050 730.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 832.950 724.950 835.050 727.050 ;
        RECT 820.950 721.950 823.050 724.050 ;
        RECT 827.400 723.900 828.600 724.650 ;
        RECT 833.400 723.900 834.600 724.650 ;
        RECT 821.400 715.050 822.450 721.950 ;
        RECT 826.950 721.800 829.050 723.900 ;
        RECT 832.950 721.800 835.050 723.900 ;
        RECT 828.000 720.750 831.000 721.050 ;
        RECT 826.950 720.300 831.000 720.750 ;
        RECT 826.950 718.950 831.450 720.300 ;
        RECT 826.950 718.650 829.050 718.950 ;
        RECT 830.400 718.050 831.450 718.950 ;
        RECT 830.400 716.400 835.050 718.050 ;
        RECT 831.000 715.950 835.050 716.400 ;
        RECT 820.950 712.950 823.050 715.050 ;
        RECT 839.400 712.050 840.450 751.950 ;
        RECT 845.400 751.050 846.450 761.100 ;
        RECT 844.950 748.950 847.050 751.050 ;
        RECT 848.400 745.050 849.450 775.950 ;
        RECT 859.950 772.950 862.050 775.050 ;
        RECT 853.950 761.100 856.050 763.200 ;
        RECT 860.400 762.600 861.450 772.950 ;
        RECT 868.950 766.950 871.050 769.050 ;
        RECT 854.400 760.350 855.600 761.100 ;
        RECT 860.400 760.350 861.600 762.600 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 856.950 757.950 859.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 862.950 757.950 865.050 760.050 ;
        RECT 850.950 754.950 853.050 757.050 ;
        RECT 857.400 755.400 858.600 757.650 ;
        RECT 863.400 755.400 864.600 757.650 ;
        RECT 847.950 742.950 850.050 745.050 ;
        RECT 851.400 739.050 852.450 754.950 ;
        RECT 857.400 751.050 858.450 755.400 ;
        RECT 859.950 751.950 862.050 754.050 ;
        RECT 856.950 748.950 859.050 751.050 ;
        RECT 860.400 745.050 861.450 751.950 ;
        RECT 863.400 748.050 864.450 755.400 ;
        RECT 869.400 754.050 870.450 766.950 ;
        RECT 874.950 761.100 877.050 763.200 ;
        RECT 881.400 762.600 882.450 802.800 ;
        RECT 887.400 802.350 888.600 804.600 ;
        RECT 896.400 802.350 897.600 804.600 ;
        RECT 886.800 799.950 888.900 802.050 ;
        RECT 895.800 799.950 897.900 802.050 ;
        RECT 899.400 795.450 900.450 806.100 ;
        RECT 914.400 805.350 915.600 806.100 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 896.400 794.400 900.450 795.450 ;
        RECT 917.400 800.400 918.600 802.650 ;
        RECT 892.950 790.950 895.050 793.050 ;
        RECT 889.950 766.950 892.050 769.050 ;
        RECT 875.400 760.350 876.600 761.100 ;
        RECT 881.400 760.350 882.600 762.600 ;
        RECT 887.400 762.450 888.600 762.600 ;
        RECT 890.400 762.450 891.450 766.950 ;
        RECT 887.400 761.400 891.450 762.450 ;
        RECT 887.400 760.350 888.600 761.400 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 880.950 757.950 883.050 760.050 ;
        RECT 883.950 757.950 886.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 878.400 756.000 879.600 757.650 ;
        RECT 868.950 751.950 871.050 754.050 ;
        RECT 874.950 751.950 877.050 754.050 ;
        RECT 877.950 751.950 880.050 756.000 ;
        RECT 884.400 755.400 885.600 757.650 ;
        RECT 862.950 745.950 865.050 748.050 ;
        RECT 859.950 742.950 862.050 745.050 ;
        RECT 865.950 742.950 868.050 745.050 ;
        RECT 850.950 736.950 853.050 739.050 ;
        RECT 862.950 733.950 865.050 736.050 ;
        RECT 841.950 727.950 844.050 730.050 ;
        RECT 850.950 729.000 853.050 733.050 ;
        RECT 842.400 718.050 843.450 727.950 ;
        RECT 851.400 727.350 852.600 729.000 ;
        RECT 856.950 728.100 859.050 730.200 ;
        RECT 857.400 727.350 858.600 728.100 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 856.950 724.950 859.050 727.050 ;
        RECT 848.400 722.400 849.600 724.650 ;
        RECT 854.400 723.000 855.600 724.650 ;
        RECT 848.400 718.050 849.450 722.400 ;
        RECT 853.950 718.950 856.050 723.000 ;
        RECT 859.950 721.950 862.050 724.050 ;
        RECT 841.950 715.950 844.050 718.050 ;
        RECT 847.950 715.950 850.050 718.050 ;
        RECT 817.950 709.950 820.050 712.050 ;
        RECT 823.950 709.950 826.050 712.050 ;
        RECT 838.950 709.950 841.050 712.050 ;
        RECT 820.950 703.950 823.050 706.050 ;
        RECT 811.950 683.100 814.050 685.200 ;
        RECT 812.400 682.350 813.600 683.100 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 815.400 678.900 816.600 679.650 ;
        RECT 814.950 676.800 817.050 678.900 ;
        RECT 817.950 676.950 820.050 679.050 ;
        RECT 805.950 670.950 808.050 673.050 ;
        RECT 811.950 670.950 814.050 673.050 ;
        RECT 796.950 664.950 799.050 667.050 ;
        RECT 802.950 664.950 805.050 667.050 ;
        RECT 749.400 650.400 753.450 651.450 ;
        RECT 767.400 650.700 776.100 651.900 ;
        RECT 749.400 649.350 750.600 650.400 ;
        RECT 741.000 647.700 747.900 648.900 ;
        RECT 741.000 645.300 741.900 647.700 ;
        RECT 739.800 643.200 741.900 645.300 ;
        RECT 742.800 643.950 744.900 646.050 ;
        RECT 736.500 639.600 738.600 641.700 ;
        RECT 743.400 641.400 744.600 643.650 ;
        RECT 746.700 640.500 747.900 647.700 ;
        RECT 748.800 646.950 750.900 649.050 ;
        RECT 764.100 646.950 766.200 649.050 ;
        RECT 764.400 645.450 765.600 646.650 ;
        RECT 761.400 644.400 765.600 645.450 ;
        RECT 746.100 638.400 748.200 640.500 ;
        RECT 761.400 637.050 762.450 644.400 ;
        RECT 767.400 641.700 768.300 650.700 ;
        RECT 774.000 649.800 776.100 650.700 ;
        RECT 777.000 648.900 777.900 654.300 ;
        RECT 781.950 652.950 784.050 655.050 ;
        RECT 779.400 651.450 780.600 651.600 ;
        RECT 779.400 650.400 783.450 651.450 ;
        RECT 790.950 651.000 793.050 655.050 ;
        RECT 779.400 649.350 780.600 650.400 ;
        RECT 771.000 647.700 777.900 648.900 ;
        RECT 771.000 645.300 771.900 647.700 ;
        RECT 769.800 643.200 771.900 645.300 ;
        RECT 772.800 643.950 774.900 646.050 ;
        RECT 766.500 639.600 768.600 641.700 ;
        RECT 773.400 641.400 774.600 643.650 ;
        RECT 776.700 640.500 777.900 647.700 ;
        RECT 778.800 646.950 780.900 649.050 ;
        RECT 776.100 638.400 778.200 640.500 ;
        RECT 748.950 634.950 751.050 637.050 ;
        RECT 760.950 634.950 763.050 637.050 ;
        RECT 730.950 628.950 733.050 631.050 ;
        RECT 715.950 625.950 718.050 628.050 ;
        RECT 706.950 622.950 709.050 625.050 ;
        RECT 716.400 610.050 717.450 625.950 ;
        RECT 730.950 622.950 733.050 625.050 ;
        RECT 700.950 606.000 703.050 610.050 ;
        RECT 715.950 607.950 718.050 610.050 ;
        RECT 701.400 604.350 702.600 606.000 ;
        RECT 706.950 605.100 709.050 607.200 ;
        RECT 707.400 604.350 708.600 605.100 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 661.950 592.950 664.050 595.050 ;
        RECT 673.950 592.950 676.050 595.050 ;
        RECT 661.950 583.950 664.050 586.050 ;
        RECT 662.400 573.600 663.450 583.950 ;
        RECT 667.950 580.950 670.050 583.050 ;
        RECT 668.400 573.600 669.450 580.950 ;
        RECT 676.950 574.950 679.050 577.050 ;
        RECT 662.400 571.350 663.600 573.600 ;
        RECT 668.400 571.350 669.600 573.600 ;
        RECT 661.950 568.950 664.050 571.050 ;
        RECT 664.950 568.950 667.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 665.400 567.900 666.600 568.650 ;
        RECT 671.400 567.900 672.600 568.650 ;
        RECT 677.400 567.900 678.450 574.950 ;
        RECT 680.400 574.050 681.450 599.400 ;
        RECT 685.950 598.800 688.050 600.900 ;
        RECT 694.950 598.950 697.050 601.050 ;
        RECT 704.400 600.900 705.600 601.650 ;
        RECT 703.950 598.800 706.050 600.900 ;
        RECT 716.400 600.450 717.450 607.950 ;
        RECT 724.950 605.100 727.050 607.200 ;
        RECT 725.400 604.350 726.600 605.100 ;
        RECT 721.950 601.950 724.050 604.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 722.400 600.900 723.600 601.650 ;
        RECT 716.400 599.400 720.450 600.450 ;
        RECT 697.950 592.950 700.050 595.050 ;
        RECT 694.950 580.950 697.050 583.050 ;
        RECT 679.950 571.950 682.050 574.050 ;
        RECT 685.950 573.000 688.050 577.050 ;
        RECT 686.400 571.350 687.600 573.000 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 685.950 568.950 688.050 571.050 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 664.950 565.800 667.050 567.900 ;
        RECT 670.950 565.800 673.050 567.900 ;
        RECT 676.950 565.800 679.050 567.900 ;
        RECT 683.400 566.400 684.600 568.650 ;
        RECT 689.400 566.400 690.600 568.650 ;
        RECT 661.950 562.950 664.050 565.050 ;
        RECT 655.950 559.950 658.050 562.050 ;
        RECT 646.950 527.100 649.050 529.200 ;
        RECT 652.950 527.100 655.050 529.200 ;
        RECT 658.950 527.100 661.050 529.200 ;
        RECT 662.400 529.050 663.450 562.950 ;
        RECT 683.400 553.050 684.450 566.400 ;
        RECT 682.950 550.950 685.050 553.050 ;
        RECT 664.950 535.950 667.050 538.050 ;
        RECT 653.400 526.350 654.600 527.100 ;
        RECT 659.400 526.350 660.600 527.100 ;
        RECT 661.950 526.950 664.050 529.050 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 650.400 522.450 651.600 523.650 ;
        RECT 644.400 521.400 651.600 522.450 ;
        RECT 656.400 521.400 657.600 523.650 ;
        RECT 628.950 517.950 631.050 520.050 ;
        RECT 625.950 511.950 628.050 514.050 ;
        RECT 629.400 508.050 630.450 517.950 ;
        RECT 634.950 511.950 637.050 514.050 ;
        RECT 628.950 505.950 631.050 508.050 ;
        RECT 628.950 501.450 631.050 502.050 ;
        RECT 623.400 500.400 631.050 501.450 ;
        RECT 628.950 499.950 631.050 500.400 ;
        RECT 620.400 497.400 630.450 498.450 ;
        RECT 611.400 478.050 612.450 496.950 ;
        RECT 620.400 495.600 621.450 497.400 ;
        RECT 620.400 493.350 621.600 495.600 ;
        RECT 625.950 494.100 628.050 496.200 ;
        RECT 629.400 495.450 630.450 497.400 ;
        RECT 629.400 494.400 633.450 495.450 ;
        RECT 626.400 493.350 627.600 494.100 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 625.950 490.950 628.050 493.050 ;
        RECT 617.400 490.050 618.600 490.650 ;
        RECT 613.950 488.400 618.600 490.050 ;
        RECT 623.400 489.900 624.600 490.650 ;
        RECT 613.950 487.950 618.000 488.400 ;
        RECT 622.950 487.800 625.050 489.900 ;
        RECT 628.950 487.950 631.050 490.050 ;
        RECT 623.400 484.050 624.450 487.800 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 629.400 481.050 630.450 487.950 ;
        RECT 632.400 484.050 633.450 494.400 ;
        RECT 631.950 481.950 634.050 484.050 ;
        RECT 628.950 478.950 631.050 481.050 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 608.400 473.400 612.450 474.450 ;
        RECT 607.950 463.950 610.050 466.050 ;
        RECT 592.950 456.450 595.050 457.050 ;
        RECT 598.950 456.450 601.050 457.050 ;
        RECT 592.950 455.400 601.050 456.450 ;
        RECT 592.950 454.950 595.050 455.400 ;
        RECT 598.950 454.950 601.050 455.400 ;
        RECT 595.950 449.100 598.050 451.200 ;
        RECT 601.950 449.100 604.050 451.200 ;
        RECT 596.400 448.350 597.600 449.100 ;
        RECT 602.400 448.350 603.600 449.100 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 598.950 445.950 601.050 448.050 ;
        RECT 601.950 445.950 604.050 448.050 ;
        RECT 599.400 444.000 600.600 445.650 ;
        RECT 598.950 439.950 601.050 444.000 ;
        RECT 592.950 436.950 595.050 439.050 ;
        RECT 593.400 409.050 594.450 436.950 ;
        RECT 604.950 430.950 607.050 433.050 ;
        RECT 605.400 424.050 606.450 430.950 ;
        RECT 608.400 430.050 609.450 463.950 ;
        RECT 611.400 439.050 612.450 473.400 ;
        RECT 619.950 457.950 622.050 460.050 ;
        RECT 628.950 459.450 631.050 460.050 ;
        RECT 623.400 458.400 631.050 459.450 ;
        RECT 620.400 450.600 621.450 457.950 ;
        RECT 623.400 454.050 624.450 458.400 ;
        RECT 628.950 457.950 631.050 458.400 ;
        RECT 625.950 454.950 628.050 457.050 ;
        RECT 622.950 451.950 625.050 454.050 ;
        RECT 626.400 451.200 627.450 454.950 ;
        RECT 620.400 448.350 621.600 450.600 ;
        RECT 625.950 449.100 628.050 451.200 ;
        RECT 626.400 448.350 627.600 449.100 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 617.400 444.900 618.600 445.650 ;
        RECT 623.400 444.900 624.600 445.650 ;
        RECT 629.400 444.900 630.600 445.650 ;
        RECT 616.950 439.950 619.050 444.900 ;
        RECT 622.950 442.800 625.050 444.900 ;
        RECT 628.950 442.800 631.050 444.900 ;
        RECT 628.950 439.650 631.050 441.750 ;
        RECT 610.950 436.950 613.050 439.050 ;
        RECT 607.950 427.950 610.050 430.050 ;
        RECT 604.950 421.950 607.050 424.050 ;
        RECT 610.950 418.950 613.050 421.050 ;
        RECT 601.950 416.100 604.050 418.200 ;
        RECT 602.400 415.350 603.600 416.100 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 595.950 409.800 598.050 411.900 ;
        RECT 599.400 410.400 600.600 412.650 ;
        RECT 605.400 411.900 606.600 412.650 ;
        RECT 592.950 406.950 595.050 409.050 ;
        RECT 589.950 394.950 592.050 397.050 ;
        RECT 586.950 388.950 589.050 391.050 ;
        RECT 583.950 379.950 586.050 382.050 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 580.950 376.950 583.050 379.050 ;
        RECT 577.950 370.950 580.050 373.050 ;
        RECT 581.400 372.600 582.450 376.950 ;
        RECT 590.400 373.200 591.450 379.950 ;
        RECT 574.950 361.950 577.050 364.050 ;
        RECT 574.950 358.800 577.050 360.900 ;
        RECT 571.950 352.950 574.050 355.050 ;
        RECT 572.400 343.050 573.450 352.950 ;
        RECT 575.400 343.200 576.450 358.800 ;
        RECT 578.400 349.050 579.450 370.950 ;
        RECT 581.400 370.350 582.600 372.600 ;
        RECT 589.950 371.100 592.050 373.200 ;
        RECT 590.400 370.350 591.600 371.100 ;
        RECT 593.400 370.050 594.450 406.950 ;
        RECT 596.400 403.050 597.450 409.800 ;
        RECT 599.400 409.050 600.450 410.400 ;
        RECT 604.950 409.800 607.050 411.900 ;
        RECT 598.950 406.950 601.050 409.050 ;
        RECT 595.950 400.950 598.050 403.050 ;
        RECT 595.950 391.950 598.050 394.050 ;
        RECT 581.100 367.950 583.200 370.050 ;
        RECT 584.400 367.950 586.500 370.050 ;
        RECT 589.800 367.950 591.900 370.050 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 584.400 365.400 585.600 367.650 ;
        RECT 584.400 364.050 585.450 365.400 ;
        RECT 583.950 361.950 586.050 364.050 ;
        RECT 580.950 352.950 583.050 355.050 ;
        RECT 577.950 346.950 580.050 349.050 ;
        RECT 581.400 346.050 582.450 352.950 ;
        RECT 580.950 343.950 583.050 346.050 ;
        RECT 571.950 340.950 574.050 343.050 ;
        RECT 574.950 341.100 577.050 343.200 ;
        RECT 574.950 337.950 577.050 340.050 ;
        RECT 580.800 338.100 582.900 340.200 ;
        RECT 584.400 340.050 585.450 361.950 ;
        RECT 586.950 355.950 589.050 358.050 ;
        RECT 593.400 357.450 594.450 367.950 ;
        RECT 596.400 361.050 597.450 391.950 ;
        RECT 599.400 382.050 600.450 406.950 ;
        RECT 605.400 406.050 606.450 409.800 ;
        RECT 604.950 403.950 607.050 406.050 ;
        RECT 611.400 400.050 612.450 418.950 ;
        RECT 613.950 415.950 616.050 418.050 ;
        RECT 619.950 416.100 622.050 418.200 ;
        RECT 610.950 397.950 613.050 400.050 ;
        RECT 614.400 388.050 615.450 415.950 ;
        RECT 620.400 415.350 621.600 416.100 ;
        RECT 617.100 412.950 619.200 415.050 ;
        RECT 620.400 412.950 622.500 415.050 ;
        RECT 625.800 412.950 627.900 415.050 ;
        RECT 617.400 411.000 618.600 412.650 ;
        RECT 616.950 406.950 619.050 411.000 ;
        RECT 626.400 410.400 627.600 412.650 ;
        RECT 626.400 406.050 627.450 410.400 ;
        RECT 616.950 403.800 619.050 405.900 ;
        RECT 625.950 403.950 628.050 406.050 ;
        RECT 613.950 385.950 616.050 388.050 ;
        RECT 598.950 379.950 601.050 382.050 ;
        RECT 604.950 372.000 607.050 376.050 ;
        RECT 610.950 373.950 613.050 379.050 ;
        RECT 613.950 373.950 616.050 376.050 ;
        RECT 605.400 370.350 606.600 372.000 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 602.400 367.050 603.600 367.650 ;
        RECT 598.950 365.400 603.600 367.050 ;
        RECT 608.400 366.000 609.600 367.650 ;
        RECT 598.950 364.950 603.000 365.400 ;
        RECT 607.950 361.950 610.050 366.000 ;
        RECT 614.400 361.050 615.450 373.950 ;
        RECT 617.400 364.050 618.450 403.800 ;
        RECT 622.950 397.950 625.050 400.050 ;
        RECT 623.400 376.050 624.450 397.950 ;
        RECT 629.400 394.050 630.450 439.650 ;
        RECT 635.400 436.050 636.450 511.950 ;
        RECT 637.950 498.450 642.000 499.050 ;
        RECT 637.950 496.950 642.450 498.450 ;
        RECT 641.400 495.600 642.450 496.950 ;
        RECT 641.400 493.350 642.600 495.600 ;
        RECT 638.100 490.950 640.200 493.050 ;
        RECT 641.400 490.950 643.500 493.050 ;
        RECT 646.800 490.950 648.900 493.050 ;
        RECT 638.400 488.400 639.600 490.650 ;
        RECT 647.400 488.400 648.600 490.650 ;
        RECT 638.400 484.050 639.450 488.400 ;
        RECT 637.950 481.950 640.050 484.050 ;
        RECT 647.400 478.050 648.450 488.400 ;
        RECT 637.950 475.950 640.050 478.050 ;
        RECT 646.950 475.950 649.050 478.050 ;
        RECT 638.400 442.050 639.450 475.950 ;
        RECT 650.400 466.050 651.450 521.400 ;
        RECT 652.950 517.950 655.050 520.050 ;
        RECT 649.950 463.950 652.050 466.050 ;
        RECT 653.400 463.050 654.450 517.950 ;
        RECT 656.400 516.450 657.450 521.400 ;
        RECT 656.400 515.400 660.450 516.450 ;
        RECT 655.950 511.950 658.050 514.050 ;
        RECT 656.400 478.050 657.450 511.950 ;
        RECT 659.400 499.050 660.450 515.400 ;
        RECT 665.400 511.050 666.450 535.950 ;
        RECT 675.000 531.450 679.050 532.050 ;
        RECT 674.400 529.950 679.050 531.450 ;
        RECT 674.400 528.600 675.450 529.950 ;
        RECT 674.400 526.350 675.600 528.600 ;
        RECT 679.950 527.100 682.050 529.200 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 667.950 520.950 670.050 523.050 ;
        RECT 671.400 521.400 672.600 523.650 ;
        RECT 664.950 508.950 667.050 511.050 ;
        RECT 658.950 496.950 661.050 499.050 ;
        RECT 664.950 495.000 667.050 499.050 ;
        RECT 668.400 498.450 669.450 520.950 ;
        RECT 671.400 502.050 672.450 521.400 ;
        RECT 680.400 514.050 681.450 527.100 ;
        RECT 683.400 522.900 684.450 550.950 ;
        RECT 689.400 550.050 690.450 566.400 ;
        RECT 695.400 553.050 696.450 580.950 ;
        RECT 698.400 573.450 699.450 592.950 ;
        RECT 706.950 589.950 709.050 592.050 ;
        RECT 707.400 579.450 708.450 589.950 ;
        RECT 707.400 577.200 708.600 579.450 ;
        RECT 703.500 575.100 705.600 577.200 ;
        RECT 701.400 573.450 702.600 573.600 ;
        RECT 698.400 572.400 702.600 573.450 ;
        RECT 701.400 571.350 702.600 572.400 ;
        RECT 701.100 568.950 703.200 571.050 ;
        RECT 704.100 570.000 705.000 575.100 ;
        RECT 706.800 574.800 708.900 576.900 ;
        RECT 713.400 575.400 715.500 577.500 ;
        RECT 711.000 573.000 713.100 573.900 ;
        RECT 705.900 571.800 713.100 573.000 ;
        RECT 705.900 570.900 708.000 571.800 ;
        RECT 711.000 570.000 713.100 570.900 ;
        RECT 704.100 569.100 713.100 570.000 ;
        RECT 704.100 562.500 705.000 569.100 ;
        RECT 711.000 568.800 713.100 569.100 ;
        RECT 706.800 565.950 708.900 568.050 ;
        RECT 707.400 563.400 708.600 565.650 ;
        RECT 714.000 562.800 714.900 575.400 ;
        RECT 715.800 568.950 717.900 571.050 ;
        RECT 716.400 567.900 717.600 568.650 ;
        RECT 715.950 565.800 718.050 567.900 ;
        RECT 704.100 560.400 706.200 562.500 ;
        RECT 713.100 560.700 715.200 562.800 ;
        RECT 719.400 559.050 720.450 599.400 ;
        RECT 721.950 598.800 724.050 600.900 ;
        RECT 722.400 592.050 723.450 598.800 ;
        RECT 724.950 592.950 727.050 595.050 ;
        RECT 721.950 589.950 724.050 592.050 ;
        RECT 706.950 556.950 709.050 559.050 ;
        RECT 718.950 556.950 721.050 559.050 ;
        RECT 694.950 550.950 697.050 553.050 ;
        RECT 688.950 547.950 691.050 550.050 ;
        RECT 694.950 547.800 697.050 549.900 ;
        RECT 703.950 547.950 706.050 550.050 ;
        RECT 688.950 528.000 691.050 532.050 ;
        RECT 695.400 529.200 696.450 547.800 ;
        RECT 689.400 526.350 690.600 528.000 ;
        RECT 694.950 527.100 697.050 529.200 ;
        RECT 695.400 526.350 696.600 527.100 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 694.950 523.950 697.050 526.050 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 692.400 522.900 693.600 523.650 ;
        RECT 682.950 520.800 685.050 522.900 ;
        RECT 691.950 520.800 694.050 522.900 ;
        RECT 698.400 522.450 699.600 523.650 ;
        RECT 704.400 522.450 705.450 547.950 ;
        RECT 698.400 521.400 705.450 522.450 ;
        RECT 703.950 517.950 706.050 520.050 ;
        RECT 679.950 511.950 682.050 514.050 ;
        RECT 685.950 511.950 688.050 514.050 ;
        RECT 676.950 508.950 679.050 511.050 ;
        RECT 670.950 499.950 673.050 502.050 ;
        RECT 668.400 497.400 672.450 498.450 ;
        RECT 665.400 493.350 666.600 495.000 ;
        RECT 659.100 490.950 661.200 493.050 ;
        RECT 664.500 490.950 666.600 493.050 ;
        RECT 667.800 490.950 669.900 493.050 ;
        RECT 659.400 489.900 660.600 490.650 ;
        RECT 658.950 487.800 661.050 489.900 ;
        RECT 668.400 488.400 669.600 490.650 ;
        RECT 668.400 484.050 669.450 488.400 ;
        RECT 667.950 481.950 670.050 484.050 ;
        RECT 671.400 481.050 672.450 497.400 ;
        RECT 673.950 493.950 676.050 496.050 ;
        RECT 677.400 495.450 678.450 508.950 ;
        RECT 686.400 495.600 687.450 511.950 ;
        RECT 704.400 508.050 705.450 517.950 ;
        RECT 707.400 514.050 708.450 556.950 ;
        RECT 725.400 544.050 726.450 592.950 ;
        RECT 731.400 589.050 732.450 622.950 ;
        RECT 739.950 605.100 742.050 607.200 ;
        RECT 740.400 604.350 741.600 605.100 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 737.400 599.400 738.600 601.650 ;
        RECT 749.400 601.050 750.450 634.950 ;
        RECT 782.400 628.050 783.450 650.400 ;
        RECT 791.400 649.350 792.600 651.000 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 794.400 646.050 795.600 646.650 ;
        RECT 803.400 646.050 804.450 664.950 ;
        RECT 812.400 651.600 813.450 670.950 ;
        RECT 818.400 651.600 819.450 676.950 ;
        RECT 821.400 667.050 822.450 703.950 ;
        RECT 820.950 664.950 823.050 667.050 ;
        RECT 812.400 649.350 813.600 651.600 ;
        RECT 818.400 649.350 819.600 651.600 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 809.400 646.050 810.600 646.650 ;
        RECT 787.950 643.950 790.050 646.050 ;
        RECT 794.400 644.400 799.050 646.050 ;
        RECT 795.000 643.950 799.050 644.400 ;
        RECT 802.950 643.950 805.050 646.050 ;
        RECT 805.950 644.400 810.600 646.050 ;
        RECT 815.400 645.900 816.600 646.650 ;
        RECT 805.950 643.950 810.000 644.400 ;
        RECT 781.950 625.950 784.050 628.050 ;
        RECT 763.950 613.950 766.050 616.050 ;
        RECT 757.950 610.950 760.050 613.050 ;
        RECT 758.400 606.600 759.450 610.950 ;
        RECT 758.400 604.350 759.600 606.600 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 737.400 595.050 738.450 599.400 ;
        RECT 748.950 598.950 751.050 601.050 ;
        RECT 755.400 599.400 756.600 601.650 ;
        RECT 764.400 601.050 765.450 613.950 ;
        RECT 775.950 610.950 778.050 613.050 ;
        RECT 769.950 605.100 772.050 607.200 ;
        RECT 776.400 606.600 777.450 610.950 ;
        RECT 784.950 607.950 787.050 610.050 ;
        RECT 770.400 604.350 771.600 605.100 ;
        RECT 776.400 604.350 777.600 606.600 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 755.400 595.050 756.450 599.400 ;
        RECT 763.950 598.950 766.050 601.050 ;
        RECT 773.400 600.900 774.600 601.650 ;
        RECT 772.950 598.800 775.050 600.900 ;
        RECT 779.400 600.450 780.600 601.650 ;
        RECT 785.400 600.450 786.450 607.950 ;
        RECT 779.400 599.400 786.450 600.450 ;
        RECT 736.950 592.950 739.050 595.050 ;
        RECT 754.950 592.950 757.050 595.050 ;
        RECT 730.950 586.950 733.050 589.050 ;
        RECT 733.950 572.100 736.050 574.200 ;
        RECT 734.400 571.350 735.600 572.100 ;
        RECT 745.950 571.950 748.050 574.050 ;
        RECT 755.400 573.600 756.450 592.950 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 733.950 568.950 736.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 731.400 567.900 732.600 568.650 ;
        RECT 730.950 565.800 733.050 567.900 ;
        RECT 737.400 566.400 738.600 568.650 ;
        RECT 746.400 567.900 747.450 571.950 ;
        RECT 755.400 571.350 756.600 573.600 ;
        RECT 760.950 571.950 763.050 577.050 ;
        RECT 769.950 573.000 772.050 577.050 ;
        RECT 770.400 571.350 771.600 573.000 ;
        RECT 775.950 572.100 778.050 574.200 ;
        RECT 776.400 571.350 777.600 572.100 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 752.400 567.900 753.600 568.650 ;
        RECT 731.400 550.050 732.450 565.800 ;
        RECT 737.400 553.050 738.450 566.400 ;
        RECT 745.950 565.800 748.050 567.900 ;
        RECT 751.950 565.800 754.050 567.900 ;
        RECT 758.400 567.000 759.600 568.650 ;
        RECT 752.400 559.050 753.450 565.800 ;
        RECT 757.950 562.950 760.050 567.000 ;
        RECT 764.400 565.050 765.450 568.950 ;
        RECT 773.400 567.900 774.600 568.650 ;
        RECT 782.400 568.050 783.450 599.400 ;
        RECT 784.950 595.950 787.050 598.050 ;
        RECT 772.950 565.800 775.050 567.900 ;
        RECT 781.950 565.950 784.050 568.050 ;
        RECT 763.950 562.950 766.050 565.050 ;
        RECT 769.950 562.950 772.050 565.050 ;
        RECT 751.950 556.950 754.050 559.050 ;
        RECT 748.950 553.950 751.050 556.050 ;
        RECT 736.950 550.950 739.050 553.050 ;
        RECT 730.950 547.950 733.050 550.050 ;
        RECT 724.950 541.950 727.050 544.050 ;
        RECT 715.950 528.000 718.050 532.050 ;
        RECT 716.400 526.350 717.600 528.000 ;
        RECT 721.950 527.100 724.050 529.200 ;
        RECT 725.400 529.050 726.450 541.950 ;
        RECT 727.950 529.950 730.050 532.050 ;
        RECT 722.400 526.350 723.600 527.100 ;
        RECT 724.950 526.950 727.050 529.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 718.950 523.950 721.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 713.400 522.000 714.600 523.650 ;
        RECT 719.400 522.900 720.600 523.650 ;
        RECT 712.950 517.950 715.050 522.000 ;
        RECT 718.950 520.800 721.050 522.900 ;
        RECT 724.950 517.950 727.050 523.050 ;
        RECT 706.950 511.950 709.050 514.050 ;
        RECT 728.400 511.050 729.450 529.950 ;
        RECT 730.950 527.100 733.050 529.200 ;
        RECT 736.950 527.100 739.050 529.200 ;
        RECT 742.950 528.000 745.050 532.050 ;
        RECT 749.400 529.050 750.450 553.950 ;
        RECT 766.950 547.950 769.050 550.050 ;
        RECT 731.400 520.050 732.450 527.100 ;
        RECT 737.400 526.350 738.600 527.100 ;
        RECT 743.400 526.350 744.600 528.000 ;
        RECT 748.950 526.950 751.050 529.050 ;
        RECT 757.950 528.000 760.050 532.050 ;
        RECT 767.400 529.200 768.450 547.950 ;
        RECT 758.400 526.350 759.600 528.000 ;
        RECT 766.950 527.100 769.050 529.200 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 751.950 523.950 754.050 526.050 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 733.950 520.950 736.050 523.050 ;
        RECT 740.400 521.400 741.600 523.650 ;
        RECT 746.400 521.400 747.600 523.650 ;
        RECT 730.800 517.950 732.900 520.050 ;
        RECT 712.950 508.950 715.050 511.050 ;
        RECT 727.950 508.950 730.050 511.050 ;
        RECT 703.950 505.950 706.050 508.050 ;
        RECT 704.400 495.600 705.450 505.950 ;
        RECT 680.400 495.450 681.600 495.600 ;
        RECT 677.400 494.400 681.600 495.450 ;
        RECT 670.950 478.950 673.050 481.050 ;
        RECT 655.950 475.950 658.050 478.050 ;
        RECT 646.950 460.950 649.050 463.050 ;
        RECT 652.950 460.950 655.050 463.050 ;
        RECT 674.400 462.450 675.450 493.950 ;
        RECT 680.400 493.350 681.600 494.400 ;
        RECT 686.400 493.350 687.600 495.600 ;
        RECT 704.400 493.350 705.600 495.600 ;
        RECT 679.950 490.950 682.050 493.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 683.400 489.900 684.600 490.650 ;
        RECT 682.950 487.800 685.050 489.900 ;
        RECT 689.400 488.400 690.600 490.650 ;
        RECT 707.400 488.400 708.600 490.650 ;
        RECT 689.400 478.050 690.450 488.400 ;
        RECT 691.950 478.950 694.050 481.050 ;
        RECT 688.950 475.950 691.050 478.050 ;
        RECT 674.400 461.400 678.450 462.450 ;
        RECT 647.400 450.600 648.450 460.950 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 673.950 457.950 676.050 460.050 ;
        RECT 647.400 448.350 648.600 450.600 ;
        RECT 652.950 449.100 655.050 451.200 ;
        RECT 653.400 448.350 654.600 449.100 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 644.400 444.900 645.600 445.650 ;
        RECT 643.950 442.800 646.050 444.900 ;
        RECT 650.400 443.400 651.600 445.650 ;
        RECT 637.950 439.950 640.050 442.050 ;
        RECT 646.950 439.950 649.050 442.050 ;
        RECT 634.950 433.950 637.050 436.050 ;
        RECT 631.950 424.950 634.050 427.050 ;
        RECT 632.400 415.050 633.450 424.950 ;
        RECT 634.950 421.950 637.050 424.050 ;
        RECT 643.950 421.950 646.050 424.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 628.950 391.950 631.050 394.050 ;
        RECT 622.950 373.950 625.050 376.050 ;
        RECT 625.950 372.000 628.050 376.050 ;
        RECT 632.400 372.600 633.450 412.950 ;
        RECT 635.400 400.050 636.450 421.950 ;
        RECT 644.400 421.200 645.600 421.950 ;
        RECT 640.500 419.100 642.600 421.200 ;
        RECT 647.400 421.050 648.450 439.950 ;
        RECT 650.400 427.050 651.450 443.400 ;
        RECT 659.400 442.050 660.450 457.950 ;
        RECT 667.950 449.100 670.050 451.200 ;
        RECT 668.400 448.350 669.600 449.100 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 665.400 444.900 666.600 445.650 ;
        RECT 664.950 442.800 667.050 444.900 ;
        RECT 674.400 444.450 675.450 457.950 ;
        RECT 677.400 451.050 678.450 461.400 ;
        RECT 676.950 448.950 679.050 451.050 ;
        RECT 682.950 449.100 685.050 451.200 ;
        RECT 683.400 448.350 684.600 449.100 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 671.400 443.400 675.450 444.450 ;
        RECT 680.400 443.400 681.600 445.650 ;
        RECT 686.400 444.900 687.600 445.650 ;
        RECT 658.950 439.950 661.050 442.050 ;
        RECT 649.950 424.950 652.050 427.050 ;
        RECT 655.950 424.950 658.050 427.050 ;
        RECT 637.950 416.100 640.050 418.200 ;
        RECT 638.400 415.350 639.600 416.100 ;
        RECT 638.100 412.950 640.200 415.050 ;
        RECT 641.100 414.000 642.000 419.100 ;
        RECT 643.800 418.800 645.900 420.900 ;
        RECT 646.950 418.950 649.050 421.050 ;
        RECT 650.400 419.400 652.500 421.500 ;
        RECT 648.000 417.000 650.100 417.900 ;
        RECT 642.900 415.800 650.100 417.000 ;
        RECT 642.900 414.900 645.000 415.800 ;
        RECT 648.000 414.000 650.100 414.900 ;
        RECT 641.100 413.100 650.100 414.000 ;
        RECT 641.100 406.500 642.000 413.100 ;
        RECT 648.000 412.800 650.100 413.100 ;
        RECT 643.800 409.950 645.900 412.050 ;
        RECT 644.400 407.400 645.600 409.650 ;
        RECT 651.000 406.800 651.900 419.400 ;
        RECT 652.800 412.950 654.900 415.050 ;
        RECT 653.400 411.450 654.600 412.650 ;
        RECT 656.400 411.450 657.450 424.950 ;
        RECT 664.950 416.100 667.050 418.200 ;
        RECT 671.400 417.600 672.450 443.400 ;
        RECT 680.400 436.050 681.450 443.400 ;
        RECT 685.950 442.800 688.050 444.900 ;
        RECT 679.950 433.950 682.050 436.050 ;
        RECT 679.950 427.950 682.050 430.050 ;
        RECT 665.400 415.350 666.600 416.100 ;
        RECT 671.400 415.350 672.600 417.600 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 653.400 410.400 657.450 411.450 ;
        RECT 668.400 410.400 669.600 412.650 ;
        RECT 674.400 411.900 675.600 412.650 ;
        RECT 641.100 404.400 643.200 406.500 ;
        RECT 650.100 404.700 652.200 406.800 ;
        RECT 634.950 397.950 637.050 400.050 ;
        RECT 637.950 397.950 640.050 400.050 ;
        RECT 646.950 397.950 649.050 400.050 ;
        RECT 634.950 388.950 637.050 391.050 ;
        RECT 635.400 373.050 636.450 388.950 ;
        RECT 626.400 370.350 627.600 372.000 ;
        RECT 632.400 370.350 633.600 372.600 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 623.400 365.400 624.600 367.650 ;
        RECT 629.400 366.900 630.600 367.650 ;
        RECT 638.400 366.900 639.450 397.950 ;
        RECT 640.950 391.950 643.050 394.050 ;
        RECT 616.950 361.950 619.050 364.050 ;
        RECT 623.400 361.050 624.450 365.400 ;
        RECT 628.950 364.800 631.050 366.900 ;
        RECT 637.950 364.800 640.050 366.900 ;
        RECT 625.950 361.950 628.050 364.050 ;
        RECT 595.950 358.950 598.050 361.050 ;
        RECT 604.950 358.950 607.050 361.050 ;
        RECT 613.950 358.950 616.050 361.050 ;
        RECT 622.950 358.950 625.050 361.050 ;
        RECT 593.400 356.400 597.450 357.450 ;
        RECT 575.400 337.350 576.600 337.950 ;
        RECT 581.400 337.350 582.600 338.100 ;
        RECT 583.950 337.950 586.050 340.050 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 566.400 333.000 570.450 333.450 ;
        RECT 565.950 332.400 570.450 333.000 ;
        RECT 557.400 325.050 558.450 332.400 ;
        RECT 559.950 328.950 562.050 331.050 ;
        RECT 550.950 322.950 553.050 325.050 ;
        RECT 556.950 322.950 559.050 325.050 ;
        RECT 538.950 316.950 541.050 319.050 ;
        RECT 556.950 313.950 559.050 316.050 ;
        RECT 541.800 310.950 543.900 313.050 ;
        RECT 544.950 310.950 547.050 313.050 ;
        RECT 535.950 298.950 538.050 301.050 ;
        RECT 530.400 287.400 534.450 288.450 ;
        RECT 517.950 277.950 520.050 280.050 ;
        RECT 530.400 265.050 531.450 287.400 ;
        RECT 532.950 274.950 535.050 277.050 ;
        RECT 529.950 262.950 532.050 265.050 ;
        RECT 523.950 260.100 526.050 262.200 ;
        RECT 524.400 259.350 525.600 260.100 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 514.950 253.950 517.050 256.050 ;
        RECT 521.400 255.450 522.600 256.650 ;
        RECT 518.400 254.400 522.600 255.450 ;
        RECT 527.400 256.050 528.600 256.650 ;
        RECT 527.400 254.400 532.050 256.050 ;
        RECT 518.400 249.450 519.450 254.400 ;
        RECT 528.000 253.950 532.050 254.400 ;
        RECT 533.400 253.050 534.450 274.950 ;
        RECT 536.400 268.050 537.450 298.950 ;
        RECT 542.400 294.600 543.450 310.950 ;
        RECT 545.400 298.050 546.450 310.950 ;
        RECT 553.950 307.950 556.050 310.050 ;
        RECT 544.800 295.950 546.900 298.050 ;
        RECT 542.400 292.350 543.600 294.600 ;
        RECT 547.950 294.000 550.050 298.050 ;
        RECT 554.400 295.200 555.450 307.950 ;
        RECT 557.400 301.050 558.450 313.950 ;
        RECT 556.950 298.950 559.050 301.050 ;
        RECT 548.400 292.350 549.600 294.000 ;
        RECT 553.950 293.100 556.050 295.200 ;
        RECT 554.400 292.350 555.600 293.100 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 545.400 288.900 546.600 289.650 ;
        RECT 544.950 286.800 547.050 288.900 ;
        RECT 551.400 288.000 552.600 289.650 ;
        RECT 550.950 283.950 553.050 288.000 ;
        RECT 556.950 286.950 559.050 289.050 ;
        RECT 557.400 277.050 558.450 286.950 ;
        RECT 556.950 274.950 559.050 277.050 ;
        RECT 560.400 274.050 561.450 328.950 ;
        RECT 563.400 316.050 564.450 332.400 ;
        RECT 565.950 331.050 568.050 332.400 ;
        RECT 571.950 331.950 574.050 334.050 ;
        RECT 578.400 333.900 579.600 334.650 ;
        RECT 565.800 330.000 568.050 331.050 ;
        RECT 565.800 328.950 567.900 330.000 ;
        RECT 568.950 328.950 571.050 331.050 ;
        RECT 565.950 322.950 568.050 325.050 ;
        RECT 562.950 313.950 565.050 316.050 ;
        RECT 562.950 301.950 565.050 304.050 ;
        RECT 563.400 286.050 564.450 301.950 ;
        RECT 566.400 295.050 567.450 322.950 ;
        RECT 569.400 310.050 570.450 328.950 ;
        RECT 572.400 319.050 573.450 331.950 ;
        RECT 577.950 331.800 580.050 333.900 ;
        RECT 574.950 328.950 577.050 331.050 ;
        RECT 583.950 328.950 586.050 331.050 ;
        RECT 571.950 316.950 574.050 319.050 ;
        RECT 575.400 315.450 576.450 328.950 ;
        RECT 584.400 325.050 585.450 328.950 ;
        RECT 587.400 325.050 588.450 355.950 ;
        RECT 589.950 352.950 592.050 355.050 ;
        RECT 590.400 343.050 591.450 352.950 ;
        RECT 592.950 343.950 595.050 346.050 ;
        RECT 589.950 340.950 592.050 343.050 ;
        RECT 589.950 337.800 592.050 339.900 ;
        RECT 593.400 339.450 594.450 343.950 ;
        RECT 596.400 343.050 597.450 356.400 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 596.400 339.450 597.600 339.600 ;
        RECT 593.400 338.400 597.600 339.450 ;
        RECT 590.400 334.050 591.450 337.800 ;
        RECT 596.400 337.350 597.600 338.400 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 589.950 331.950 592.050 334.050 ;
        RECT 599.400 333.900 600.600 334.650 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 601.950 325.950 604.050 328.050 ;
        RECT 583.800 322.950 585.900 325.050 ;
        RECT 586.950 322.950 589.050 325.050 ;
        RECT 595.950 319.950 598.050 322.050 ;
        RECT 580.950 316.950 583.050 319.050 ;
        RECT 572.400 314.400 576.450 315.450 ;
        RECT 568.950 307.950 571.050 310.050 ;
        RECT 572.400 307.050 573.450 314.400 ;
        RECT 574.950 310.950 577.050 313.050 ;
        RECT 571.950 304.950 574.050 307.050 ;
        RECT 565.950 292.950 568.050 295.050 ;
        RECT 568.950 293.100 571.050 295.200 ;
        RECT 575.400 294.600 576.450 310.950 ;
        RECT 569.400 292.350 570.600 293.100 ;
        RECT 575.400 292.350 576.600 294.600 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 572.400 288.900 573.600 289.650 ;
        RECT 571.950 286.800 574.050 288.900 ;
        RECT 581.400 288.450 582.450 316.950 ;
        RECT 596.400 316.050 597.450 319.950 ;
        RECT 595.800 313.950 597.900 316.050 ;
        RECT 598.950 313.950 601.050 316.050 ;
        RECT 583.950 301.950 586.050 304.050 ;
        RECT 584.400 294.450 585.450 301.950 ;
        RECT 599.400 295.200 600.450 313.950 ;
        RECT 602.400 313.050 603.450 325.950 ;
        RECT 605.400 316.050 606.450 358.950 ;
        RECT 616.950 352.950 619.050 355.050 ;
        RECT 613.950 346.950 616.050 349.050 ;
        RECT 614.400 339.600 615.450 346.950 ;
        RECT 617.400 343.050 618.450 352.950 ;
        RECT 616.950 340.950 619.050 343.050 ;
        RECT 614.400 337.350 615.600 339.600 ;
        RECT 619.950 338.100 622.050 340.200 ;
        RECT 620.400 337.350 621.600 338.100 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 611.400 333.900 612.600 334.650 ;
        RECT 610.950 331.800 613.050 333.900 ;
        RECT 617.400 332.400 618.600 334.650 ;
        RECT 617.400 325.050 618.450 332.400 ;
        RECT 622.950 331.950 625.050 334.050 ;
        RECT 616.950 322.950 619.050 325.050 ;
        RECT 604.950 313.950 607.050 316.050 ;
        RECT 601.950 310.950 604.050 313.050 ;
        RECT 604.950 298.950 607.050 301.050 ;
        RECT 601.950 295.950 604.050 298.050 ;
        RECT 587.400 294.450 588.600 294.600 ;
        RECT 584.400 293.400 588.600 294.450 ;
        RECT 587.400 292.350 588.600 293.400 ;
        RECT 592.950 293.100 595.050 295.200 ;
        RECT 598.950 293.100 601.050 295.200 ;
        RECT 593.400 292.350 594.600 293.100 ;
        RECT 586.950 289.950 589.050 292.050 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 578.400 287.400 582.450 288.450 ;
        RECT 590.400 287.400 591.600 289.650 ;
        RECT 562.950 283.950 565.050 286.050 ;
        RECT 550.950 271.950 553.050 274.050 ;
        RECT 559.950 271.950 562.050 274.050 ;
        RECT 535.950 265.950 538.050 268.050 ;
        RECT 535.950 260.100 538.050 262.200 ;
        RECT 541.950 260.100 544.050 262.200 ;
        RECT 520.800 250.950 522.900 253.050 ;
        RECT 523.950 250.950 526.050 253.050 ;
        RECT 532.950 250.950 535.050 253.050 ;
        RECT 515.400 248.400 519.450 249.450 ;
        RECT 511.950 235.950 514.050 238.050 ;
        RECT 505.950 223.950 508.050 226.050 ;
        RECT 505.950 220.800 508.050 222.900 ;
        RECT 511.950 220.950 514.050 223.050 ;
        RECT 506.400 217.050 507.450 220.800 ;
        RECT 505.950 214.950 508.050 217.050 ;
        RECT 512.400 216.600 513.450 220.950 ;
        RECT 515.400 217.050 516.450 248.400 ;
        RECT 517.950 238.950 520.050 241.050 ;
        RECT 518.400 232.050 519.450 238.950 ;
        RECT 517.950 229.950 520.050 232.050 ;
        RECT 512.400 214.350 513.600 216.600 ;
        RECT 514.800 214.950 516.900 217.050 ;
        RECT 517.950 215.100 520.050 217.200 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 509.400 210.900 510.600 211.650 ;
        RECT 508.950 208.800 511.050 210.900 ;
        RECT 509.400 196.050 510.450 208.800 ;
        RECT 514.950 207.450 517.050 211.050 ;
        RECT 512.400 207.000 517.050 207.450 ;
        RECT 512.400 206.400 516.450 207.000 ;
        RECT 508.950 193.950 511.050 196.050 ;
        RECT 505.950 187.950 508.050 190.050 ;
        RECT 502.950 184.950 505.050 187.050 ;
        RECT 499.950 181.950 502.050 184.050 ;
        RECT 506.400 183.600 507.450 187.950 ;
        RECT 512.400 184.050 513.450 206.400 ;
        RECT 518.400 205.050 519.450 215.100 ;
        RECT 517.950 202.950 520.050 205.050 ;
        RECT 514.950 184.950 517.050 187.050 ;
        RECT 506.400 181.350 507.600 183.600 ;
        RECT 511.950 181.950 514.050 184.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 505.950 178.950 508.050 181.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 503.400 177.900 504.600 178.650 ;
        RECT 509.400 177.900 510.600 178.650 ;
        RECT 484.950 169.950 487.050 172.050 ;
        RECT 481.950 160.950 484.050 163.050 ;
        RECT 478.950 148.950 481.050 151.050 ;
        RECT 475.950 140.100 478.050 145.050 ;
        RECT 440.400 136.350 441.600 136.950 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 437.400 133.050 438.600 133.650 ;
        RECT 433.950 131.400 438.600 133.050 ;
        RECT 449.400 132.900 450.450 137.400 ;
        RECT 451.950 136.950 456.600 137.400 ;
        RECT 455.400 136.350 456.600 136.950 ;
        RECT 461.400 136.350 462.600 138.000 ;
        RECT 466.950 136.950 469.050 139.050 ;
        RECT 469.950 136.950 472.050 139.050 ;
        RECT 475.950 136.950 478.050 139.050 ;
        RECT 482.400 138.600 483.450 160.950 ;
        RECT 494.400 154.050 495.450 175.950 ;
        RECT 496.950 175.800 499.050 177.900 ;
        RECT 502.950 175.800 505.050 177.900 ;
        RECT 508.950 175.800 511.050 177.900 ;
        RECT 509.400 157.050 510.450 175.800 ;
        RECT 508.950 154.950 511.050 157.050 ;
        RECT 493.950 151.950 496.050 154.050 ;
        RECT 502.950 142.950 505.050 145.050 ;
        RECT 503.400 139.200 504.450 142.950 ;
        RECT 476.400 136.350 477.600 136.950 ;
        RECT 482.400 136.350 483.600 138.600 ;
        RECT 496.950 137.100 499.050 139.200 ;
        RECT 502.950 137.100 505.050 139.200 ;
        RECT 497.400 136.350 498.600 137.100 ;
        RECT 503.400 136.350 504.600 137.100 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 457.950 133.950 460.050 136.050 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 469.950 133.800 472.050 135.900 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 478.950 133.950 481.050 136.050 ;
        RECT 481.950 133.950 484.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 499.950 133.950 502.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 433.950 130.950 438.000 131.400 ;
        RECT 448.950 130.800 451.050 132.900 ;
        RECT 458.400 131.400 459.600 133.650 ;
        RECT 464.400 131.400 465.600 133.650 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 436.950 127.950 439.050 130.050 ;
        RECT 412.950 118.950 415.050 121.050 ;
        RECT 437.400 115.050 438.450 127.950 ;
        RECT 430.950 112.950 433.050 115.050 ;
        RECT 436.950 112.950 439.050 115.050 ;
        RECT 409.950 104.100 412.050 106.200 ;
        RECT 418.950 104.100 421.050 106.200 ;
        RECT 424.950 104.100 427.050 106.200 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 394.950 100.950 397.050 103.050 ;
        RECT 397.950 100.950 400.050 103.050 ;
        RECT 400.950 100.950 403.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 395.400 99.000 396.600 100.650 ;
        RECT 401.400 99.900 402.600 100.650 ;
        RECT 410.400 100.050 411.450 104.100 ;
        RECT 419.400 103.350 420.600 104.100 ;
        RECT 425.400 103.350 426.600 104.100 ;
        RECT 415.950 100.950 418.050 103.050 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 394.950 94.950 397.050 99.000 ;
        RECT 400.950 97.800 403.050 99.900 ;
        RECT 406.950 97.800 409.050 99.900 ;
        RECT 409.800 97.950 411.900 100.050 ;
        RECT 385.950 88.950 388.050 91.050 ;
        RECT 382.950 75.450 385.050 76.050 ;
        RECT 380.400 74.400 385.050 75.450 ;
        RECT 367.950 64.950 370.050 67.050 ;
        RECT 356.400 62.400 360.450 63.450 ;
        RECT 362.400 63.000 366.450 63.450 ;
        RECT 347.400 58.350 348.600 60.600 ;
        RECT 352.950 59.100 355.050 61.200 ;
        RECT 353.400 58.350 354.600 59.100 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 346.950 55.950 349.050 58.050 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 316.950 49.950 319.050 52.050 ;
        RECT 313.950 46.950 316.050 49.050 ;
        RECT 310.950 31.950 313.050 34.050 ;
        RECT 271.950 22.950 274.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 265.950 19.950 268.050 22.050 ;
        RECT 268.950 18.300 271.050 22.050 ;
        RECT 272.400 21.900 273.600 22.650 ;
        RECT 278.400 21.900 279.600 22.650 ;
        RECT 271.950 19.800 274.050 21.900 ;
        RECT 277.950 19.800 280.050 21.900 ;
        RECT 290.400 19.050 291.450 25.950 ;
        RECT 296.400 25.350 297.600 27.600 ;
        RECT 302.400 25.350 303.600 27.600 ;
        RECT 307.950 25.950 310.050 31.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 299.400 20.400 300.600 22.650 ;
        RECT 305.400 21.900 306.600 22.650 ;
        RECT 299.400 19.050 300.450 20.400 ;
        RECT 304.950 19.800 307.050 21.900 ;
        RECT 277.950 18.300 280.050 18.750 ;
        RECT 268.950 18.000 280.050 18.300 ;
        RECT 269.400 17.250 280.050 18.000 ;
        RECT 277.950 16.650 280.050 17.250 ;
        RECT 289.950 16.950 292.050 19.050 ;
        RECT 298.950 16.950 301.050 19.050 ;
        RECT 299.400 13.050 300.450 16.950 ;
        RECT 311.400 16.050 312.450 31.950 ;
        RECT 320.400 28.200 321.450 52.950 ;
        RECT 323.400 34.050 324.450 53.400 ;
        RECT 328.950 52.800 331.050 54.900 ;
        RECT 337.800 52.950 339.900 55.050 ;
        RECT 340.950 52.950 343.050 55.050 ;
        RECT 344.400 54.000 345.600 55.650 ;
        RECT 331.950 37.950 334.050 40.050 ;
        RECT 322.950 31.950 325.050 34.050 ;
        RECT 319.950 26.100 322.050 28.200 ;
        RECT 325.950 26.100 328.050 28.200 ;
        RECT 320.400 25.350 321.600 26.100 ;
        RECT 326.400 25.350 327.600 26.100 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 313.950 19.950 316.050 22.050 ;
        RECT 317.400 21.900 318.600 22.650 ;
        RECT 314.400 16.050 315.450 19.950 ;
        RECT 316.950 19.800 319.050 21.900 ;
        RECT 323.400 21.000 324.600 22.650 ;
        RECT 322.950 16.950 325.050 21.000 ;
        RECT 328.950 19.950 331.050 22.050 ;
        RECT 332.400 21.900 333.450 37.950 ;
        RECT 341.400 30.450 342.450 52.950 ;
        RECT 343.950 49.950 346.050 54.000 ;
        RECT 350.400 53.400 351.600 55.650 ;
        RECT 341.400 29.400 345.450 30.450 ;
        RECT 334.950 27.600 339.000 28.050 ;
        RECT 344.400 27.600 345.450 29.400 ;
        RECT 334.950 25.950 339.600 27.600 ;
        RECT 338.400 25.350 339.600 25.950 ;
        RECT 344.400 25.350 345.600 27.600 ;
        RECT 350.400 27.450 351.450 53.400 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 356.400 40.050 357.450 52.950 ;
        RECT 359.400 49.050 360.450 62.400 ;
        RECT 361.950 62.400 366.450 63.000 ;
        RECT 361.950 58.950 364.050 62.400 ;
        RECT 368.400 60.600 369.450 64.950 ;
        RECT 368.400 58.350 369.600 60.600 ;
        RECT 373.950 59.100 376.050 61.200 ;
        RECT 374.400 58.350 375.600 59.100 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 365.400 54.900 366.600 55.650 ;
        RECT 364.950 52.800 367.050 54.900 ;
        RECT 371.400 53.400 372.600 55.650 ;
        RECT 358.950 46.950 361.050 49.050 ;
        RECT 365.400 46.050 366.450 52.800 ;
        RECT 364.950 43.950 367.050 46.050 ;
        RECT 358.950 40.950 361.050 43.050 ;
        RECT 355.950 37.950 358.050 40.050 ;
        RECT 355.950 31.950 358.050 34.050 ;
        RECT 350.400 26.400 354.450 27.450 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 341.400 21.900 342.600 22.650 ;
        RECT 310.950 13.950 313.050 16.050 ;
        RECT 314.400 14.400 319.050 16.050 ;
        RECT 315.000 13.950 319.050 14.400 ;
        RECT 298.950 10.950 301.050 13.050 ;
        RECT 329.400 10.050 330.450 19.950 ;
        RECT 331.950 19.800 334.050 21.900 ;
        RECT 340.950 19.800 343.050 21.900 ;
        RECT 347.400 21.000 348.600 22.650 ;
        RECT 341.400 16.050 342.450 19.800 ;
        RECT 346.950 16.950 349.050 21.000 ;
        RECT 334.950 13.950 337.050 16.050 ;
        RECT 340.950 13.950 343.050 16.050 ;
        RECT 335.400 10.050 336.450 13.950 ;
        RECT 353.400 13.050 354.450 26.400 ;
        RECT 356.400 19.050 357.450 31.950 ;
        RECT 359.400 28.050 360.450 40.950 ;
        RECT 371.400 40.050 372.450 53.400 ;
        RECT 376.950 52.950 379.050 55.050 ;
        RECT 373.950 45.450 376.050 46.050 ;
        RECT 377.400 45.450 378.450 52.950 ;
        RECT 373.950 44.400 378.450 45.450 ;
        RECT 373.950 43.950 376.050 44.400 ;
        RECT 370.950 37.950 373.050 40.050 ;
        RECT 361.950 31.950 364.050 34.050 ;
        RECT 367.950 31.950 370.050 34.050 ;
        RECT 358.950 25.950 361.050 28.050 ;
        RECT 362.400 27.600 363.450 31.950 ;
        RECT 368.400 27.600 369.450 31.950 ;
        RECT 374.400 28.050 375.450 43.950 ;
        RECT 376.950 31.950 379.050 34.050 ;
        RECT 362.400 25.350 363.600 27.600 ;
        RECT 368.400 25.350 369.600 27.600 ;
        RECT 373.950 25.950 376.050 28.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 370.950 22.950 373.050 25.050 ;
        RECT 365.400 21.900 366.600 22.650 ;
        RECT 371.400 21.900 372.600 22.650 ;
        RECT 364.950 19.800 367.050 21.900 ;
        RECT 370.950 19.800 373.050 21.900 ;
        RECT 377.400 19.050 378.450 31.950 ;
        RECT 355.950 16.950 358.050 19.050 ;
        RECT 366.000 18.750 369.000 19.050 ;
        RECT 364.950 18.300 369.000 18.750 ;
        RECT 364.950 16.950 369.450 18.300 ;
        RECT 376.950 16.950 379.050 19.050 ;
        RECT 364.950 16.650 367.050 16.950 ;
        RECT 368.400 16.050 369.450 16.950 ;
        RECT 380.400 16.050 381.450 74.400 ;
        RECT 382.950 73.950 385.050 74.400 ;
        RECT 407.400 70.050 408.450 97.800 ;
        RECT 412.950 94.950 415.050 100.050 ;
        RECT 416.400 98.400 417.600 100.650 ;
        RECT 422.400 99.900 423.600 100.650 ;
        RECT 431.400 99.900 432.450 112.950 ;
        RECT 436.950 109.800 439.050 111.900 ;
        RECT 437.400 105.600 438.450 109.800 ;
        RECT 437.400 103.350 438.600 105.600 ;
        RECT 442.950 105.000 445.050 109.050 ;
        RECT 443.400 103.350 444.600 105.000 ;
        RECT 451.950 103.950 454.050 106.050 ;
        RECT 458.400 105.450 459.450 131.400 ;
        RECT 464.400 124.050 465.450 131.400 ;
        RECT 470.400 127.050 471.450 133.800 ;
        RECT 479.400 132.900 480.600 133.650 ;
        RECT 478.950 130.800 481.050 132.900 ;
        RECT 485.400 131.400 486.600 133.650 ;
        RECT 500.400 132.900 501.600 133.650 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 460.800 121.950 462.900 124.050 ;
        RECT 463.950 121.950 466.050 124.050 ;
        RECT 455.400 104.400 459.450 105.450 ;
        RECT 461.400 105.600 462.450 121.950 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 416.400 91.050 417.450 98.400 ;
        RECT 421.950 97.800 424.050 99.900 ;
        RECT 430.950 97.800 433.050 99.900 ;
        RECT 440.400 98.400 441.600 100.650 ;
        RECT 446.400 99.900 447.600 100.650 ;
        RECT 452.400 99.900 453.450 103.950 ;
        RECT 415.950 88.950 418.050 91.050 ;
        RECT 421.950 88.950 424.050 91.050 ;
        RECT 422.400 85.050 423.450 88.950 ;
        RECT 440.400 85.050 441.450 98.400 ;
        RECT 445.950 97.800 448.050 99.900 ;
        RECT 451.950 97.800 454.050 99.900 ;
        RECT 421.950 82.950 424.050 85.050 ;
        RECT 439.950 82.950 442.050 85.050 ;
        RECT 455.400 82.050 456.450 104.400 ;
        RECT 461.400 103.350 462.600 105.600 ;
        RECT 466.950 104.100 469.050 109.050 ;
        RECT 467.400 103.350 468.600 104.100 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 464.400 99.900 465.600 100.650 ;
        RECT 463.950 97.800 466.050 99.900 ;
        RECT 470.400 98.400 471.600 100.650 ;
        RECT 470.400 85.050 471.450 98.400 ;
        RECT 476.400 88.050 477.450 124.950 ;
        RECT 478.950 118.950 481.050 121.050 ;
        RECT 479.400 94.050 480.450 118.950 ;
        RECT 481.950 112.950 484.050 115.050 ;
        RECT 482.400 105.450 483.450 112.950 ;
        RECT 485.400 109.050 486.450 131.400 ;
        RECT 499.950 130.800 502.050 132.900 ;
        RECT 506.400 131.400 507.600 133.650 ;
        RECT 515.400 132.900 516.450 184.950 ;
        RECT 518.400 172.050 519.450 202.950 ;
        RECT 521.400 196.050 522.450 250.950 ;
        RECT 524.400 217.050 525.450 250.950 ;
        RECT 536.400 229.050 537.450 260.100 ;
        RECT 542.400 259.350 543.600 260.100 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 545.400 254.400 546.600 256.650 ;
        RECT 529.950 226.950 532.050 229.050 ;
        RECT 535.950 226.950 538.050 229.050 ;
        RECT 523.950 214.950 526.050 217.050 ;
        RECT 530.400 216.600 531.450 226.950 ;
        RECT 541.950 220.950 544.050 223.050 ;
        RECT 530.400 214.350 531.600 216.600 ;
        RECT 535.950 215.100 538.050 217.200 ;
        RECT 536.400 214.350 537.600 215.100 ;
        RECT 526.950 211.950 529.050 214.050 ;
        RECT 529.950 211.950 532.050 214.050 ;
        RECT 532.950 211.950 535.050 214.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 523.950 208.800 526.050 210.900 ;
        RECT 527.400 209.400 528.600 211.650 ;
        RECT 533.400 209.400 534.600 211.650 ;
        RECT 524.400 199.050 525.450 208.800 ;
        RECT 523.950 196.950 526.050 199.050 ;
        RECT 520.950 193.950 523.050 196.050 ;
        RECT 523.950 189.450 526.050 190.050 ;
        RECT 527.400 189.450 528.450 209.400 ;
        RECT 533.400 199.050 534.450 209.400 ;
        RECT 532.950 196.950 535.050 199.050 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 523.950 188.400 528.450 189.450 ;
        RECT 523.950 187.950 526.050 188.400 ;
        RECT 524.400 183.600 525.450 187.950 ;
        RECT 524.400 181.350 525.600 183.600 ;
        RECT 530.400 183.450 531.450 193.950 ;
        RECT 542.400 187.050 543.450 220.950 ;
        RECT 535.950 184.950 538.050 187.050 ;
        RECT 541.950 184.950 544.050 187.050 ;
        RECT 530.400 182.400 534.450 183.450 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 527.400 177.900 528.600 178.650 ;
        RECT 526.950 175.800 529.050 177.900 ;
        RECT 517.950 169.950 520.050 172.050 ;
        RECT 529.950 169.950 532.050 175.050 ;
        RECT 533.400 166.050 534.450 182.400 ;
        RECT 536.400 172.050 537.450 184.950 ;
        RECT 545.400 183.600 546.450 254.400 ;
        RECT 547.950 250.950 550.050 256.050 ;
        RECT 551.400 250.050 552.450 271.950 ;
        RECT 553.950 262.950 556.050 265.050 ;
        RECT 550.950 247.950 553.050 250.050 ;
        RECT 554.400 247.050 555.450 262.950 ;
        RECT 562.950 261.000 565.050 265.050 ;
        RECT 572.400 262.050 573.450 286.800 ;
        RECT 574.950 277.950 577.050 280.050 ;
        RECT 563.400 259.350 564.600 261.000 ;
        RECT 571.950 259.950 574.050 262.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 565.950 256.950 568.050 259.050 ;
        RECT 560.400 255.900 561.600 256.650 ;
        RECT 559.950 250.950 562.050 255.900 ;
        RECT 566.400 254.400 567.600 256.650 ;
        RECT 566.400 250.050 567.450 254.400 ;
        RECT 571.950 253.950 574.050 258.900 ;
        RECT 575.400 253.050 576.450 277.950 ;
        RECT 578.400 262.050 579.450 287.400 ;
        RECT 590.400 283.050 591.450 287.400 ;
        RECT 595.950 283.950 598.050 286.050 ;
        RECT 589.950 280.950 592.050 283.050 ;
        RECT 580.950 268.950 583.050 271.050 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 581.400 261.600 582.450 268.950 ;
        RECT 581.400 259.350 582.600 261.600 ;
        RECT 586.950 260.100 589.050 265.050 ;
        RECT 587.400 259.350 588.600 260.100 ;
        RECT 592.950 259.950 595.050 262.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 584.400 254.400 585.600 256.650 ;
        RECT 574.950 250.950 577.050 253.050 ;
        RECT 580.950 250.950 583.050 253.050 ;
        RECT 565.950 247.950 568.050 250.050 ;
        RECT 553.950 244.950 556.050 247.050 ;
        RECT 562.950 223.950 565.050 226.050 ;
        RECT 553.950 215.100 556.050 217.200 ;
        RECT 554.400 214.350 555.600 215.100 ;
        RECT 559.950 214.950 562.050 217.050 ;
        RECT 550.950 211.950 553.050 214.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 551.400 210.900 552.600 211.650 ;
        RECT 550.950 208.800 553.050 210.900 ;
        RECT 551.400 202.050 552.450 208.800 ;
        RECT 560.400 204.450 561.450 214.950 ;
        RECT 563.400 207.450 564.450 223.950 ;
        RECT 577.950 220.950 580.050 223.050 ;
        RECT 568.950 215.100 571.050 217.200 ;
        RECT 569.400 214.350 570.600 215.100 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 572.400 210.000 573.600 211.650 ;
        RECT 563.400 206.400 567.450 207.450 ;
        RECT 557.400 203.400 561.450 204.450 ;
        RECT 550.950 199.950 553.050 202.050 ;
        RECT 557.400 193.050 558.450 203.400 ;
        RECT 562.950 202.950 565.050 205.050 ;
        RECT 559.950 199.950 562.050 202.050 ;
        RECT 560.400 196.050 561.450 199.950 ;
        RECT 559.950 193.950 562.050 196.050 ;
        RECT 556.950 190.950 559.050 193.050 ;
        RECT 559.950 184.950 562.050 187.050 ;
        RECT 545.400 181.350 546.600 183.600 ;
        RECT 550.950 182.100 553.050 184.200 ;
        RECT 551.400 181.350 552.600 182.100 ;
        RECT 556.950 181.950 559.050 184.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 542.400 177.900 543.600 178.650 ;
        RECT 541.950 175.800 544.050 177.900 ;
        RECT 548.400 177.000 549.600 178.650 ;
        RECT 547.950 172.950 550.050 177.000 ;
        RECT 535.950 169.950 538.050 172.050 ;
        RECT 532.950 163.950 535.050 166.050 ;
        RECT 553.950 160.950 556.050 163.050 ;
        RECT 538.950 148.950 541.050 151.050 ;
        RECT 523.950 137.100 526.050 139.200 ;
        RECT 529.950 138.000 532.050 142.050 ;
        RECT 524.400 136.350 525.600 137.100 ;
        RECT 530.400 136.350 531.600 138.000 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 526.950 133.950 529.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 521.400 132.900 522.600 133.650 ;
        RECT 514.950 132.450 517.050 132.900 ;
        RECT 512.400 131.400 517.050 132.450 ;
        RECT 506.400 127.050 507.450 131.400 ;
        RECT 505.950 124.950 508.050 127.050 ;
        RECT 512.400 124.050 513.450 131.400 ;
        RECT 514.950 130.800 517.050 131.400 ;
        RECT 520.950 130.800 523.050 132.900 ;
        RECT 527.400 131.400 528.600 133.650 ;
        RECT 511.950 121.950 514.050 124.050 ;
        RECT 499.950 118.950 502.050 121.050 ;
        RECT 490.950 109.950 493.050 112.050 ;
        RECT 484.950 106.950 487.050 109.050 ;
        RECT 491.400 105.600 492.450 109.950 ;
        RECT 485.400 105.450 486.600 105.600 ;
        RECT 482.400 104.400 486.600 105.450 ;
        RECT 485.400 103.350 486.600 104.400 ;
        RECT 491.400 103.350 492.600 105.600 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 488.400 98.400 489.600 100.650 ;
        RECT 494.400 99.450 495.600 100.650 ;
        RECT 494.400 98.400 498.450 99.450 ;
        RECT 478.950 91.950 481.050 94.050 ;
        RECT 488.400 88.050 489.450 98.400 ;
        RECT 493.950 91.950 496.050 94.050 ;
        RECT 475.950 85.950 478.050 88.050 ;
        RECT 487.950 85.950 490.050 88.050 ;
        RECT 469.950 82.950 472.050 85.050 ;
        RECT 427.950 79.050 430.050 82.050 ;
        RECT 454.950 79.950 457.050 82.050 ;
        RECT 424.950 78.000 430.050 79.050 ;
        RECT 424.950 77.400 429.450 78.000 ;
        RECT 424.950 76.950 429.000 77.400 ;
        RECT 433.950 76.950 436.050 79.050 ;
        RECT 412.950 73.950 415.050 76.050 ;
        RECT 427.950 73.950 430.050 76.050 ;
        RECT 406.950 67.950 409.050 70.050 ;
        RECT 391.950 64.950 394.050 67.050 ;
        RECT 382.950 59.100 385.050 61.200 ;
        RECT 392.400 60.600 393.450 64.950 ;
        RECT 383.400 55.050 384.450 59.100 ;
        RECT 392.400 58.350 393.600 60.600 ;
        RECT 397.950 59.100 400.050 61.200 ;
        RECT 403.950 59.100 406.050 61.200 ;
        RECT 413.400 60.600 414.450 73.950 ;
        RECT 398.400 58.350 399.600 59.100 ;
        RECT 388.950 55.950 391.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 382.950 52.950 385.050 55.050 ;
        RECT 389.400 53.400 390.600 55.650 ;
        RECT 395.400 54.900 396.600 55.650 ;
        RECT 404.400 55.050 405.450 59.100 ;
        RECT 413.400 58.350 414.600 60.600 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 419.400 58.350 420.600 59.100 ;
        RECT 428.400 58.050 429.450 73.950 ;
        RECT 434.400 61.050 435.450 76.950 ;
        RECT 442.950 67.950 445.050 70.050 ;
        RECT 454.950 67.950 457.050 70.050 ;
        RECT 433.950 58.950 436.050 61.050 ;
        RECT 436.950 59.100 439.050 61.200 ;
        RECT 443.400 60.600 444.450 67.950 ;
        RECT 448.950 61.200 451.050 64.050 ;
        RECT 437.400 58.350 438.600 59.100 ;
        RECT 443.400 58.350 444.600 60.600 ;
        RECT 448.800 60.000 451.050 61.200 ;
        RECT 448.800 59.100 450.900 60.000 ;
        RECT 451.950 59.100 454.050 61.200 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 389.400 49.050 390.450 53.400 ;
        RECT 394.950 52.800 397.050 54.900 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 388.950 46.950 391.050 49.050 ;
        RECT 395.400 34.050 396.450 52.800 ;
        RECT 404.400 40.050 405.450 52.950 ;
        RECT 403.950 37.950 406.050 40.050 ;
        RECT 407.400 37.050 408.450 55.950 ;
        RECT 416.400 54.900 417.600 55.650 ;
        RECT 415.950 52.800 418.050 54.900 ;
        RECT 422.400 53.400 423.600 55.650 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 419.400 46.050 420.450 49.950 ;
        RECT 422.400 49.050 423.450 53.400 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 421.950 46.950 424.050 49.050 ;
        RECT 418.950 43.950 421.050 46.050 ;
        RECT 422.400 43.050 423.450 46.950 ;
        RECT 421.950 40.950 424.050 43.050 ;
        RECT 425.400 40.050 426.450 52.950 ;
        RECT 427.950 52.800 430.050 54.900 ;
        RECT 433.950 52.950 436.050 55.050 ;
        RECT 440.400 54.900 441.600 55.650 ;
        RECT 418.950 37.950 421.050 40.050 ;
        RECT 424.950 37.950 427.050 40.050 ;
        RECT 406.950 34.950 409.050 37.050 ;
        RECT 394.950 31.950 397.050 34.050 ;
        RECT 385.950 27.000 388.050 31.050 ;
        RECT 386.400 25.350 387.600 27.000 ;
        RECT 391.950 26.100 394.050 28.200 ;
        RECT 400.800 26.100 402.900 28.200 ;
        RECT 403.950 26.100 406.050 28.200 ;
        RECT 412.950 26.100 415.050 28.200 ;
        RECT 419.400 27.600 420.450 37.950 ;
        RECT 392.400 25.350 393.600 26.100 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 394.950 22.950 397.050 25.050 ;
        RECT 389.400 20.400 390.600 22.650 ;
        RECT 395.400 20.400 396.600 22.650 ;
        RECT 401.400 22.050 402.450 26.100 ;
        RECT 368.400 14.400 373.050 16.050 ;
        RECT 369.000 13.950 373.050 14.400 ;
        RECT 379.950 13.950 382.050 16.050 ;
        RECT 352.950 10.950 355.050 13.050 ;
        RECT 389.400 10.050 390.450 20.400 ;
        RECT 295.950 9.450 298.050 10.050 ;
        RECT 301.950 9.450 304.050 10.050 ;
        RECT 295.950 8.400 304.050 9.450 ;
        RECT 295.950 7.950 298.050 8.400 ;
        RECT 301.950 7.950 304.050 8.400 ;
        RECT 328.950 7.950 331.050 10.050 ;
        RECT 334.950 7.950 337.050 10.050 ;
        RECT 346.950 7.950 352.050 10.050 ;
        RECT 355.950 7.950 361.050 10.050 ;
        RECT 388.950 7.950 391.050 10.050 ;
        RECT 395.400 7.050 396.450 20.400 ;
        RECT 400.950 19.950 403.050 22.050 ;
        RECT 404.400 7.050 405.450 26.100 ;
        RECT 413.400 25.350 414.600 26.100 ;
        RECT 419.400 25.350 420.600 27.600 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 415.950 22.950 418.050 25.050 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 410.400 21.900 411.600 22.650 ;
        RECT 409.950 19.800 412.050 21.900 ;
        RECT 416.400 20.400 417.600 22.650 ;
        RECT 416.400 10.050 417.450 20.400 ;
        RECT 428.400 16.050 429.450 52.800 ;
        RECT 434.400 27.600 435.450 52.950 ;
        RECT 439.950 52.800 442.050 54.900 ;
        RECT 446.400 53.400 447.600 55.650 ;
        RECT 452.400 55.050 453.450 59.100 ;
        RECT 446.400 34.050 447.450 53.400 ;
        RECT 451.800 52.950 453.900 55.050 ;
        RECT 455.400 54.900 456.450 67.950 ;
        RECT 475.950 64.950 478.050 67.050 ;
        RECT 466.950 64.050 469.050 64.200 ;
        RECT 469.950 64.050 472.050 64.200 ;
        RECT 466.950 62.100 472.050 64.050 ;
        RECT 468.000 61.950 471.000 62.100 ;
        RECT 460.950 59.100 463.050 61.200 ;
        RECT 461.400 58.350 462.600 59.100 ;
        RECT 466.950 58.950 469.050 61.050 ;
        RECT 467.400 58.350 468.600 58.950 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 464.400 54.900 465.600 55.650 ;
        RECT 454.950 52.800 457.050 54.900 ;
        RECT 463.950 52.800 466.050 54.900 ;
        RECT 470.400 53.400 471.600 55.650 ;
        RECT 476.400 54.900 477.450 64.950 ;
        RECT 478.950 59.100 481.050 61.200 ;
        RECT 487.950 59.100 490.050 61.200 ;
        RECT 494.400 60.600 495.450 91.950 ;
        RECT 497.400 61.050 498.450 98.400 ;
        RECT 466.950 49.950 469.050 52.050 ;
        RECT 463.950 43.950 466.050 46.050 ;
        RECT 445.950 31.950 448.050 34.050 ;
        RECT 434.400 25.350 435.600 27.600 ;
        RECT 439.950 26.100 442.050 28.200 ;
        RECT 448.950 26.100 451.050 28.200 ;
        RECT 457.950 26.100 460.050 28.200 ;
        RECT 464.400 27.600 465.450 43.950 ;
        RECT 467.400 37.050 468.450 49.950 ;
        RECT 466.950 34.950 469.050 37.050 ;
        RECT 470.400 34.050 471.450 53.400 ;
        RECT 475.950 52.800 478.050 54.900 ;
        RECT 476.400 34.050 477.450 52.800 ;
        RECT 479.400 46.050 480.450 59.100 ;
        RECT 488.400 58.350 489.600 59.100 ;
        RECT 494.400 58.350 495.600 60.600 ;
        RECT 496.950 58.950 499.050 61.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 485.400 54.900 486.600 55.650 ;
        RECT 491.400 54.900 492.600 55.650 ;
        RECT 484.950 52.800 487.050 54.900 ;
        RECT 490.950 52.800 493.050 54.900 ;
        RECT 478.950 43.950 481.050 46.050 ;
        RECT 485.400 43.050 486.450 52.800 ;
        RECT 496.950 49.950 499.050 55.050 ;
        RECT 484.950 40.950 487.050 43.050 ;
        RECT 478.950 37.950 481.050 40.050 ;
        RECT 466.950 28.950 469.050 33.900 ;
        RECT 469.950 31.950 472.050 34.050 ;
        RECT 475.950 31.950 478.050 34.050 ;
        RECT 440.400 25.350 441.600 26.100 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 430.950 19.800 433.050 21.900 ;
        RECT 437.400 20.400 438.600 22.650 ;
        RECT 443.400 21.900 444.600 22.650 ;
        RECT 427.950 13.950 430.050 16.050 ;
        RECT 415.950 7.950 418.050 10.050 ;
        RECT 220.950 6.450 223.050 7.050 ;
        RECT 212.400 5.400 223.050 6.450 ;
        RECT 220.950 4.950 223.050 5.400 ;
        RECT 226.950 4.950 229.050 7.050 ;
        RECT 262.950 4.950 265.050 7.050 ;
        RECT 394.950 4.950 397.050 7.050 ;
        RECT 403.950 4.950 406.050 7.050 ;
        RECT 431.400 3.450 432.450 19.800 ;
        RECT 437.400 19.050 438.450 20.400 ;
        RECT 442.950 19.800 445.050 21.900 ;
        RECT 436.950 18.450 439.050 19.050 ;
        RECT 434.400 17.400 439.050 18.450 ;
        RECT 434.400 13.050 435.450 17.400 ;
        RECT 436.950 16.950 439.050 17.400 ;
        RECT 436.950 13.800 439.050 15.900 ;
        RECT 433.950 10.950 436.050 13.050 ;
        RECT 437.400 7.050 438.450 13.800 ;
        RECT 449.400 10.050 450.450 26.100 ;
        RECT 458.400 25.350 459.600 26.100 ;
        RECT 464.400 25.350 465.600 27.600 ;
        RECT 469.800 26.100 471.900 28.200 ;
        RECT 472.950 26.100 475.050 28.200 ;
        RECT 479.400 27.600 480.450 37.950 ;
        RECT 484.950 34.950 487.050 37.050 ;
        RECT 485.400 27.600 486.450 34.950 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 455.400 20.400 456.600 22.650 ;
        RECT 461.400 21.000 462.600 22.650 ;
        RECT 470.400 21.900 471.450 26.100 ;
        RECT 455.400 10.050 456.450 20.400 ;
        RECT 460.950 16.950 463.050 21.000 ;
        RECT 469.950 19.800 472.050 21.900 ;
        RECT 470.400 16.050 471.450 19.800 ;
        RECT 473.400 19.050 474.450 26.100 ;
        RECT 479.400 25.350 480.600 27.600 ;
        RECT 485.400 25.350 486.600 27.600 ;
        RECT 500.400 27.450 501.450 118.950 ;
        RECT 527.400 112.050 528.450 131.400 ;
        RECT 539.400 115.050 540.450 148.950 ;
        RECT 547.950 138.000 550.050 142.050 ;
        RECT 554.400 139.200 555.450 160.950 ;
        RECT 557.400 151.050 558.450 181.950 ;
        RECT 556.950 148.950 559.050 151.050 ;
        RECT 560.400 145.050 561.450 184.950 ;
        RECT 563.400 184.050 564.450 202.950 ;
        RECT 566.400 202.050 567.450 206.400 ;
        RECT 571.950 205.950 574.050 210.000 ;
        RECT 578.400 208.050 579.450 220.950 ;
        RECT 577.950 205.950 580.050 208.050 ;
        RECT 565.950 199.950 568.050 202.050 ;
        RECT 566.400 186.450 567.450 199.950 ;
        RECT 566.400 185.400 570.450 186.450 ;
        RECT 562.950 181.950 565.050 184.050 ;
        RECT 569.400 183.600 570.450 185.400 ;
        RECT 569.400 181.350 570.600 183.600 ;
        RECT 574.950 183.000 577.050 187.050 ;
        RECT 578.400 184.200 579.450 205.950 ;
        RECT 575.400 181.350 576.600 183.000 ;
        RECT 577.950 182.100 580.050 184.200 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 574.950 178.950 577.050 181.050 ;
        RECT 566.400 177.900 567.600 178.650 ;
        RECT 572.400 177.900 573.600 178.650 ;
        RECT 581.400 177.900 582.450 250.950 ;
        RECT 584.400 232.050 585.450 254.400 ;
        RECT 583.950 229.950 586.050 232.050 ;
        RECT 593.400 223.050 594.450 259.950 ;
        RECT 596.400 244.050 597.450 283.950 ;
        RECT 599.400 271.050 600.450 293.100 ;
        RECT 598.950 268.950 601.050 271.050 ;
        RECT 602.400 262.200 603.450 295.950 ;
        RECT 605.400 294.450 606.450 298.950 ;
        RECT 610.800 298.200 612.900 300.300 ;
        RECT 619.800 298.500 621.900 300.600 ;
        RECT 608.400 294.450 609.600 294.600 ;
        RECT 605.400 293.400 609.600 294.450 ;
        RECT 605.400 289.050 606.450 293.400 ;
        RECT 608.400 292.350 609.600 293.400 ;
        RECT 608.100 289.950 610.200 292.050 ;
        RECT 604.950 286.950 607.050 289.050 ;
        RECT 611.100 285.600 612.000 298.200 ;
        RECT 617.400 295.350 618.600 297.600 ;
        RECT 617.100 292.950 619.200 295.050 ;
        RECT 612.900 291.900 615.000 292.200 ;
        RECT 621.000 291.900 621.900 298.500 ;
        RECT 623.400 298.050 624.450 331.950 ;
        RECT 626.400 328.050 627.450 361.950 ;
        RECT 628.950 349.950 631.050 352.050 ;
        RECT 625.950 325.950 628.050 328.050 ;
        RECT 629.400 313.050 630.450 349.950 ;
        RECT 638.400 339.600 639.450 364.800 ;
        RECT 641.400 361.050 642.450 391.950 ;
        RECT 647.400 372.600 648.450 397.950 ;
        RECT 668.400 394.050 669.450 410.400 ;
        RECT 673.950 409.800 676.050 411.900 ;
        RECT 667.950 391.950 670.050 394.050 ;
        RECT 674.400 388.050 675.450 409.800 ;
        RECT 673.950 385.950 676.050 388.050 ;
        RECT 647.400 370.350 648.600 372.600 ;
        RECT 652.950 371.100 655.050 373.200 ;
        RECT 658.950 372.450 661.050 373.200 ;
        RECT 665.400 372.450 666.600 372.600 ;
        RECT 658.950 371.400 666.600 372.450 ;
        RECT 658.950 371.100 661.050 371.400 ;
        RECT 653.400 370.350 654.600 371.100 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 650.400 365.400 651.600 367.650 ;
        RECT 650.400 361.050 651.450 365.400 ;
        RECT 640.950 358.950 643.050 361.050 ;
        RECT 649.950 358.950 652.050 361.050 ;
        RECT 652.950 346.950 655.050 349.050 ;
        RECT 643.950 340.950 646.050 343.050 ;
        RECT 638.400 337.350 639.600 339.600 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 635.400 333.900 636.600 334.650 ;
        RECT 634.950 331.800 637.050 333.900 ;
        RECT 637.950 319.950 640.050 322.050 ;
        RECT 638.400 316.050 639.450 319.950 ;
        RECT 640.950 316.950 643.050 319.050 ;
        RECT 637.950 313.950 640.050 316.050 ;
        RECT 628.950 310.950 631.050 313.050 ;
        RECT 622.950 295.950 625.050 298.050 ;
        RECT 634.950 293.100 637.050 295.200 ;
        RECT 641.400 294.600 642.450 316.950 ;
        RECT 644.400 307.050 645.450 340.950 ;
        RECT 653.400 339.600 654.450 346.950 ;
        RECT 659.400 340.050 660.450 371.100 ;
        RECT 665.400 370.350 666.600 371.400 ;
        RECT 673.950 371.100 676.050 373.200 ;
        RECT 674.400 370.350 675.600 371.100 ;
        RECT 665.100 367.950 667.200 370.050 ;
        RECT 668.400 367.950 670.500 370.050 ;
        RECT 673.800 367.950 675.900 370.050 ;
        RECT 668.400 366.900 669.600 367.650 ;
        RECT 667.950 364.800 670.050 366.900 ;
        RECT 668.400 355.050 669.450 364.800 ;
        RECT 667.950 352.950 670.050 355.050 ;
        RECT 680.400 346.050 681.450 427.950 ;
        RECT 686.400 427.050 687.450 442.800 ;
        RECT 692.400 430.050 693.450 478.950 ;
        RECT 700.950 460.950 703.050 463.050 ;
        RECT 701.400 450.600 702.450 460.950 ;
        RECT 707.400 457.050 708.450 488.400 ;
        RECT 713.400 463.050 714.450 508.950 ;
        RECT 734.400 504.450 735.450 520.950 ;
        RECT 740.400 517.050 741.450 521.400 ;
        RECT 746.400 519.450 747.450 521.400 ;
        RECT 752.400 520.050 753.450 523.950 ;
        RECT 761.400 523.050 762.600 523.650 ;
        RECT 754.950 520.950 757.050 523.050 ;
        RECT 761.400 521.400 766.050 523.050 ;
        RECT 762.000 520.950 766.050 521.400 ;
        RECT 743.400 518.400 747.450 519.450 ;
        RECT 739.950 514.950 742.050 517.050 ;
        RECT 743.400 511.050 744.450 518.400 ;
        RECT 751.950 517.950 754.050 520.050 ;
        RECT 745.950 514.950 748.050 517.050 ;
        RECT 742.950 508.950 745.050 511.050 ;
        RECT 734.400 503.400 738.450 504.450 ;
        RECT 723.000 498.450 727.050 499.050 ;
        RECT 729.000 498.450 733.050 499.050 ;
        RECT 722.400 496.950 727.050 498.450 ;
        RECT 728.400 496.950 733.050 498.450 ;
        RECT 722.400 495.600 723.450 496.950 ;
        RECT 728.400 495.600 729.450 496.950 ;
        RECT 722.400 493.350 723.600 495.600 ;
        RECT 728.400 493.350 729.600 495.600 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 725.400 488.400 726.600 490.650 ;
        RECT 731.400 489.900 732.600 490.650 ;
        RECT 725.400 487.050 726.450 488.400 ;
        RECT 730.950 487.800 733.050 489.900 ;
        RECT 724.950 481.950 727.050 487.050 ;
        RECT 712.950 460.950 715.050 463.050 ;
        RECT 706.950 454.950 709.050 457.050 ;
        RECT 701.400 448.350 702.600 450.600 ;
        RECT 709.950 448.950 712.050 451.050 ;
        RECT 697.950 445.950 700.050 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 698.400 444.900 699.600 445.650 ;
        RECT 697.950 442.800 700.050 444.900 ;
        RECT 704.400 443.400 705.600 445.650 ;
        RECT 710.400 444.900 711.450 448.950 ;
        RECT 704.400 439.050 705.450 443.400 ;
        RECT 709.950 442.800 712.050 444.900 ;
        RECT 703.950 436.950 706.050 439.050 ;
        RECT 713.400 430.050 714.450 460.950 ;
        RECT 718.950 449.100 721.050 451.200 ;
        RECT 726.000 450.600 730.050 451.050 ;
        RECT 719.400 448.350 720.600 449.100 ;
        RECT 725.400 448.950 730.050 450.600 ;
        RECT 725.400 448.350 726.600 448.950 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 722.400 444.900 723.600 445.650 ;
        RECT 721.950 442.800 724.050 444.900 ;
        RECT 727.950 442.950 730.050 445.050 ;
        RECT 728.400 439.050 729.450 442.950 ;
        RECT 731.400 439.050 732.450 487.800 ;
        RECT 737.400 480.450 738.450 503.400 ;
        RECT 739.950 496.950 742.050 502.050 ;
        RECT 746.400 499.050 747.450 514.950 ;
        RECT 755.400 511.050 756.450 520.950 ;
        RECT 767.400 520.050 768.450 527.100 ;
        RECT 770.400 520.050 771.450 562.950 ;
        RECT 785.400 544.050 786.450 595.950 ;
        RECT 788.400 555.450 789.450 643.950 ;
        RECT 814.950 643.800 817.050 645.900 ;
        RECT 811.950 637.950 814.050 640.050 ;
        RECT 793.950 605.100 796.050 607.200 ;
        RECT 799.950 606.000 802.050 610.050 ;
        RECT 794.400 604.350 795.600 605.100 ;
        RECT 800.400 604.350 801.600 606.000 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 802.950 601.950 805.050 604.050 ;
        RECT 797.400 599.400 798.600 601.650 ;
        RECT 803.400 600.900 804.600 601.650 ;
        RECT 812.400 601.050 813.450 637.950 ;
        RECT 824.400 637.050 825.450 709.950 ;
        RECT 847.950 703.950 850.050 706.050 ;
        RECT 832.950 688.950 835.050 691.050 ;
        RECT 844.950 688.950 847.050 691.050 ;
        RECT 833.400 684.600 834.450 688.950 ;
        RECT 833.400 682.350 834.600 684.600 ;
        RECT 838.950 683.100 841.050 685.200 ;
        RECT 839.400 682.350 840.600 683.100 ;
        RECT 829.950 679.950 832.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 830.400 677.400 831.600 679.650 ;
        RECT 836.400 678.900 837.600 679.650 ;
        RECT 845.400 679.050 846.450 688.950 ;
        RECT 830.400 645.450 831.450 677.400 ;
        RECT 835.950 676.800 838.050 678.900 ;
        RECT 844.950 676.950 847.050 679.050 ;
        RECT 848.400 676.050 849.450 703.950 ;
        RECT 853.950 683.100 856.050 685.200 ;
        RECT 860.400 684.600 861.450 721.950 ;
        RECT 863.400 718.050 864.450 733.950 ;
        RECT 866.400 733.050 867.450 742.950 ;
        RECT 865.950 730.950 868.050 733.050 ;
        RECT 875.400 729.600 876.450 751.950 ;
        RECT 884.400 751.050 885.450 755.400 ;
        RECT 886.950 751.950 889.050 754.050 ;
        RECT 883.950 748.950 886.050 751.050 ;
        RECT 880.950 733.950 883.050 736.050 ;
        RECT 881.400 729.600 882.450 733.950 ;
        RECT 875.400 727.350 876.600 729.600 ;
        RECT 881.400 727.350 882.600 729.600 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 877.950 724.950 880.050 727.050 ;
        RECT 880.950 724.950 883.050 727.050 ;
        RECT 872.400 722.400 873.600 724.650 ;
        RECT 878.400 722.400 879.600 724.650 ;
        RECT 862.950 715.950 865.050 718.050 ;
        RECT 872.400 715.050 873.450 722.400 ;
        RECT 871.950 712.950 874.050 715.050 ;
        RECT 878.400 706.050 879.450 722.400 ;
        RECT 877.950 703.950 880.050 706.050 ;
        RECT 877.950 691.950 880.050 694.050 ;
        RECT 854.400 682.350 855.600 683.100 ;
        RECT 860.400 682.350 861.600 684.600 ;
        RECT 865.950 683.100 868.050 685.200 ;
        RECT 871.950 683.100 874.050 685.200 ;
        RECT 878.400 684.600 879.450 691.950 ;
        RECT 887.400 688.050 888.450 751.950 ;
        RECT 893.400 739.050 894.450 790.950 ;
        RECT 896.400 754.050 897.450 794.400 ;
        RECT 917.400 793.050 918.450 800.400 ;
        RECT 916.950 790.950 919.050 793.050 ;
        RECT 926.400 790.050 927.450 806.400 ;
        RECT 929.400 805.350 930.600 806.400 ;
        RECT 929.400 802.950 931.500 805.050 ;
        RECT 934.800 802.950 936.900 805.050 ;
        RECT 919.950 787.950 922.050 790.050 ;
        RECT 925.950 787.950 928.050 790.050 ;
        RECT 916.950 778.950 919.050 781.050 ;
        RECT 907.950 761.100 910.050 763.200 ;
        RECT 908.400 760.350 909.600 761.100 ;
        RECT 901.950 757.950 904.050 760.050 ;
        RECT 904.950 757.950 907.050 760.050 ;
        RECT 907.950 757.950 910.050 760.050 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 905.400 755.400 906.600 757.650 ;
        RECT 911.400 755.400 912.600 757.650 ;
        RECT 895.950 751.950 898.050 754.050 ;
        RECT 905.400 751.050 906.450 755.400 ;
        RECT 904.950 748.950 907.050 751.050 ;
        RECT 892.950 736.950 895.050 739.050 ;
        RECT 893.400 730.200 894.450 736.950 ;
        RECT 907.950 730.950 910.050 733.050 ;
        RECT 892.950 728.100 895.050 730.200 ;
        RECT 898.950 728.100 901.050 730.200 ;
        RECT 893.400 727.350 894.600 728.100 ;
        RECT 899.400 727.350 900.600 728.100 ;
        RECT 892.950 724.950 895.050 727.050 ;
        RECT 895.950 724.950 898.050 727.050 ;
        RECT 898.950 724.950 901.050 727.050 ;
        RECT 901.950 724.950 904.050 727.050 ;
        RECT 896.400 722.400 897.600 724.650 ;
        RECT 902.400 723.900 903.600 724.650 ;
        RECT 908.400 724.050 909.450 730.950 ;
        RECT 911.400 730.050 912.450 755.400 ;
        RECT 917.400 751.050 918.450 778.950 ;
        RECT 920.400 757.050 921.450 787.950 ;
        RECT 925.950 766.950 928.050 769.050 ;
        RECT 926.400 762.600 927.450 766.950 ;
        RECT 926.400 760.350 927.600 762.600 ;
        RECT 934.950 761.100 937.050 763.200 ;
        RECT 925.950 757.950 928.050 760.050 ;
        RECT 928.950 757.950 931.050 760.050 ;
        RECT 919.950 754.950 922.050 757.050 ;
        RECT 929.400 756.900 930.600 757.650 ;
        RECT 928.950 754.800 931.050 756.900 ;
        RECT 935.400 751.050 936.450 761.100 ;
        RECT 916.950 748.950 919.050 751.050 ;
        RECT 925.950 748.950 928.050 751.050 ;
        RECT 934.950 748.950 937.050 751.050 ;
        RECT 919.950 736.950 922.050 739.050 ;
        RECT 910.950 727.950 913.050 730.050 ;
        RECT 913.950 729.000 916.050 733.050 ;
        RECT 920.400 729.600 921.450 736.950 ;
        RECT 914.400 727.350 915.600 729.000 ;
        RECT 920.400 727.350 921.600 729.600 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 916.950 724.950 919.050 727.050 ;
        RECT 919.950 724.950 922.050 727.050 ;
        RECT 889.950 718.950 892.050 721.050 ;
        RECT 886.950 685.950 889.050 688.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 856.950 679.950 859.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 850.950 676.950 853.050 679.050 ;
        RECT 857.400 678.900 858.600 679.650 ;
        RECT 847.950 673.950 850.050 676.050 ;
        RECT 841.950 664.950 844.050 667.050 ;
        RECT 842.400 657.450 843.450 664.950 ;
        RECT 851.400 658.050 852.450 676.950 ;
        RECT 856.950 676.800 859.050 678.900 ;
        RECT 853.950 673.950 856.050 676.050 ;
        RECT 842.400 655.200 843.600 657.450 ;
        RECT 837.900 651.900 840.000 653.700 ;
        RECT 841.800 652.800 843.900 654.900 ;
        RECT 845.100 654.300 847.200 656.400 ;
        RECT 850.950 655.950 853.050 658.050 ;
        RECT 836.400 650.700 845.100 651.900 ;
        RECT 833.100 646.950 835.200 649.050 ;
        RECT 833.400 645.450 834.600 646.650 ;
        RECT 830.400 644.400 834.600 645.450 ;
        RECT 830.400 640.050 831.450 644.400 ;
        RECT 836.400 641.700 837.300 650.700 ;
        RECT 843.000 649.800 845.100 650.700 ;
        RECT 846.000 648.900 846.900 654.300 ;
        RECT 848.400 651.450 849.600 651.600 ;
        RECT 851.400 651.450 852.450 655.950 ;
        RECT 848.400 650.400 852.450 651.450 ;
        RECT 848.400 649.350 849.600 650.400 ;
        RECT 840.000 647.700 846.900 648.900 ;
        RECT 840.000 645.300 840.900 647.700 ;
        RECT 838.800 643.200 840.900 645.300 ;
        RECT 841.800 643.950 843.900 646.050 ;
        RECT 829.950 637.950 832.050 640.050 ;
        RECT 835.500 639.600 837.600 641.700 ;
        RECT 842.400 641.400 843.600 643.650 ;
        RECT 845.700 640.500 846.900 647.700 ;
        RECT 847.800 646.950 849.900 649.050 ;
        RECT 845.100 638.400 847.200 640.500 ;
        RECT 823.950 634.950 826.050 637.050 ;
        RECT 832.950 634.950 835.050 637.050 ;
        RECT 817.950 613.950 820.050 616.050 ;
        RECT 818.400 606.600 819.450 613.950 ;
        RECT 818.400 604.350 819.600 606.600 ;
        RECT 823.950 605.100 826.050 607.200 ;
        RECT 829.950 605.100 832.050 607.200 ;
        RECT 824.400 604.350 825.600 605.100 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 823.950 601.950 826.050 604.050 ;
        RECT 797.400 595.050 798.450 599.400 ;
        RECT 802.950 598.800 805.050 600.900 ;
        RECT 811.950 598.950 814.050 601.050 ;
        RECT 821.400 599.400 822.600 601.650 ;
        RECT 796.950 592.950 799.050 595.050 ;
        RECT 814.950 592.950 817.050 595.050 ;
        RECT 793.950 572.100 796.050 574.200 ;
        RECT 815.400 573.600 816.450 592.950 ;
        RECT 821.400 583.050 822.450 599.400 ;
        RECT 830.400 598.050 831.450 605.100 ;
        RECT 823.950 595.950 826.050 598.050 ;
        RECT 829.950 595.950 832.050 598.050 ;
        RECT 820.950 580.950 823.050 583.050 ;
        RECT 824.400 579.450 825.450 595.950 ;
        RECT 833.400 594.450 834.450 634.950 ;
        RECT 844.950 613.950 847.050 616.050 ;
        RECT 838.950 605.100 841.050 607.200 ;
        RECT 845.400 606.600 846.450 613.950 ;
        RECT 839.400 604.350 840.600 605.100 ;
        RECT 845.400 604.350 846.600 606.600 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 835.950 598.950 838.050 601.050 ;
        RECT 842.400 600.000 843.600 601.650 ;
        RECT 848.400 600.900 849.600 601.650 ;
        RECT 821.400 578.400 825.450 579.450 ;
        RECT 830.400 593.400 834.450 594.450 ;
        RECT 821.400 573.600 822.450 578.400 ;
        RECT 794.400 571.350 795.600 572.100 ;
        RECT 815.400 571.350 816.600 573.600 ;
        RECT 821.400 571.350 822.600 573.600 ;
        RECT 826.950 572.100 829.050 574.200 ;
        RECT 830.400 574.050 831.450 593.400 ;
        RECT 791.100 568.950 793.200 571.050 ;
        RECT 794.400 568.950 796.500 571.050 ;
        RECT 799.800 568.950 801.900 571.050 ;
        RECT 811.950 568.950 814.050 571.050 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 791.400 566.400 792.600 568.650 ;
        RECT 800.400 566.400 801.600 568.650 ;
        RECT 812.400 566.400 813.600 568.650 ;
        RECT 818.400 567.000 819.600 568.650 ;
        RECT 827.400 567.450 828.450 572.100 ;
        RECT 829.950 571.950 832.050 574.050 ;
        RECT 836.400 573.600 837.450 598.950 ;
        RECT 841.950 595.950 844.050 600.000 ;
        RECT 847.950 598.800 850.050 600.900 ;
        RECT 847.950 592.950 850.050 595.050 ;
        RECT 844.950 580.950 847.050 583.050 ;
        RECT 836.400 571.350 837.600 573.600 ;
        RECT 832.950 568.950 835.050 571.050 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 833.400 567.450 834.600 568.650 ;
        RECT 839.400 567.900 840.600 568.650 ;
        RECT 791.400 559.050 792.450 566.400 ;
        RECT 800.400 565.050 801.450 566.400 ;
        RECT 800.400 563.400 805.050 565.050 ;
        RECT 801.000 562.950 805.050 563.400 ;
        RECT 790.950 556.950 793.050 559.050 ;
        RECT 788.400 554.400 792.450 555.450 ;
        RECT 784.950 541.950 787.050 544.050 ;
        RECT 775.500 531.300 777.600 533.400 ;
        RECT 785.100 532.500 787.200 534.600 ;
        RECT 772.950 527.100 775.050 529.200 ;
        RECT 773.400 526.350 774.600 527.100 ;
        RECT 773.100 523.950 775.200 526.050 ;
        RECT 776.400 522.300 777.300 531.300 ;
        RECT 778.800 527.700 780.900 529.800 ;
        RECT 782.400 529.350 783.600 531.600 ;
        RECT 780.000 525.300 780.900 527.700 ;
        RECT 781.800 526.950 783.900 529.050 ;
        RECT 785.700 525.300 786.900 532.500 ;
        RECT 791.400 526.050 792.450 554.400 ;
        RECT 793.950 553.950 796.050 556.050 ;
        RECT 780.000 524.100 786.900 525.300 ;
        RECT 783.000 522.300 785.100 523.200 ;
        RECT 776.400 521.100 785.100 522.300 ;
        RECT 760.950 517.950 763.050 520.050 ;
        RECT 754.950 508.950 757.050 511.050 ;
        RECT 757.950 499.950 760.050 502.050 ;
        RECT 745.950 496.950 748.050 499.050 ;
        RECT 746.400 495.600 747.450 496.950 ;
        RECT 746.400 493.350 747.600 495.600 ;
        RECT 751.950 494.100 754.050 496.200 ;
        RECT 752.400 493.350 753.600 494.100 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 745.950 490.950 748.050 493.050 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 743.400 489.000 744.600 490.650 ;
        RECT 749.400 489.900 750.600 490.650 ;
        RECT 742.950 484.950 745.050 489.000 ;
        RECT 748.950 487.800 751.050 489.900 ;
        RECT 734.400 479.400 738.450 480.450 ;
        RECT 734.400 445.050 735.450 479.400 ;
        RECT 739.950 454.950 742.050 457.050 ;
        RECT 745.950 454.950 748.050 457.050 ;
        RECT 740.400 450.600 741.450 454.950 ;
        RECT 746.400 450.600 747.450 454.950 ;
        RECT 740.400 448.350 741.600 450.600 ;
        RECT 746.400 448.350 747.600 450.600 ;
        RECT 754.950 449.100 757.050 451.200 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 733.950 442.950 736.050 445.050 ;
        RECT 743.400 444.900 744.600 445.650 ;
        RECT 742.950 442.800 745.050 444.900 ;
        RECT 749.400 443.400 750.600 445.650 ;
        RECT 749.400 439.050 750.450 443.400 ;
        RECT 727.800 436.950 729.900 439.050 ;
        RECT 730.950 436.950 733.050 439.050 ;
        RECT 748.950 436.950 751.050 439.050 ;
        RECT 755.400 436.050 756.450 449.100 ;
        RECT 742.950 433.950 745.050 436.050 ;
        RECT 754.950 433.950 757.050 436.050 ;
        RECT 691.950 427.950 694.050 430.050 ;
        RECT 712.950 427.950 715.050 430.050 ;
        RECT 685.950 424.950 688.050 427.050 ;
        RECT 700.950 424.950 703.050 427.050 ;
        RECT 697.950 421.950 700.050 424.050 ;
        RECT 688.950 416.100 691.050 418.200 ;
        RECT 689.400 415.350 690.600 416.100 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 692.400 410.400 693.600 412.650 ;
        RECT 698.400 412.050 699.450 421.950 ;
        RECT 692.400 409.050 693.450 410.400 ;
        RECT 697.950 409.950 700.050 412.050 ;
        RECT 692.400 407.400 697.050 409.050 ;
        RECT 693.000 406.950 697.050 407.400 ;
        RECT 691.950 400.950 694.050 403.050 ;
        RECT 692.400 397.050 693.450 400.950 ;
        RECT 694.950 397.950 697.050 400.050 ;
        RECT 691.950 394.950 694.050 397.050 ;
        RECT 688.950 371.100 691.050 373.200 ;
        RECT 695.400 372.600 696.450 397.950 ;
        RECT 701.400 384.450 702.450 424.950 ;
        RECT 709.950 421.950 712.050 424.050 ;
        RECT 710.400 417.600 711.450 421.950 ;
        RECT 710.400 415.350 711.600 417.600 ;
        RECT 715.950 416.100 718.050 418.200 ;
        RECT 716.400 415.350 717.600 416.100 ;
        RECT 721.950 415.950 724.050 418.050 ;
        RECT 730.950 416.100 733.050 418.200 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 707.400 411.000 708.600 412.650 ;
        RECT 706.950 406.950 709.050 411.000 ;
        RECT 713.400 410.400 714.600 412.650 ;
        RECT 713.400 406.050 714.450 410.400 ;
        RECT 722.400 409.050 723.450 415.950 ;
        RECT 731.400 415.350 732.600 416.100 ;
        RECT 739.950 415.950 742.050 418.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 728.400 410.400 729.600 412.650 ;
        RECT 734.400 411.000 735.600 412.650 ;
        RECT 721.950 406.950 724.050 409.050 ;
        RECT 712.950 403.950 715.050 406.050 ;
        RECT 728.400 391.050 729.450 410.400 ;
        RECT 733.950 408.450 736.050 411.000 ;
        RECT 733.950 407.400 738.450 408.450 ;
        RECT 733.950 406.950 736.050 407.400 ;
        RECT 727.950 388.950 730.050 391.050 ;
        RECT 701.400 383.400 705.450 384.450 ;
        RECT 689.400 370.350 690.600 371.100 ;
        RECT 695.400 370.350 696.600 372.600 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 692.400 365.400 693.600 367.650 ;
        RECT 698.400 365.400 699.600 367.650 ;
        RECT 692.400 361.050 693.450 365.400 ;
        RECT 698.400 361.050 699.450 365.400 ;
        RECT 691.950 358.950 694.050 361.050 ;
        RECT 697.950 358.950 700.050 361.050 ;
        RECT 682.950 352.950 685.050 355.050 ;
        RECT 661.950 343.950 664.050 346.050 ;
        RECT 679.950 343.950 682.050 346.050 ;
        RECT 653.400 337.350 654.600 339.600 ;
        RECT 658.950 337.950 661.050 340.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 652.950 334.950 655.050 337.050 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 650.400 333.900 651.600 334.650 ;
        RECT 656.400 333.900 657.600 334.650 ;
        RECT 649.950 331.800 652.050 333.900 ;
        RECT 655.950 331.800 658.050 333.900 ;
        RECT 662.400 328.050 663.450 343.950 ;
        RECT 670.950 338.100 673.050 340.200 ;
        RECT 679.950 338.100 682.050 340.200 ;
        RECT 671.400 337.350 672.600 338.100 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 664.950 331.800 667.050 333.900 ;
        RECT 668.400 332.400 669.600 334.650 ;
        RECT 674.400 333.900 675.600 334.650 ;
        RECT 649.950 325.950 652.050 328.050 ;
        RECT 661.950 325.950 664.050 328.050 ;
        RECT 643.950 304.950 646.050 307.050 ;
        RECT 650.400 295.200 651.450 325.950 ;
        RECT 655.950 298.950 658.050 301.050 ;
        RECT 635.400 292.350 636.600 293.100 ;
        RECT 641.400 292.350 642.600 294.600 ;
        RECT 649.950 293.100 652.050 295.200 ;
        RECT 656.400 294.600 657.450 298.950 ;
        RECT 665.400 294.600 666.450 331.800 ;
        RECT 668.400 316.050 669.450 332.400 ;
        RECT 673.950 328.950 676.050 333.900 ;
        RECT 680.400 316.050 681.450 338.100 ;
        RECT 683.400 333.900 684.450 352.950 ;
        RECT 697.950 343.950 700.050 346.050 ;
        RECT 691.950 338.100 694.050 340.200 ;
        RECT 698.400 339.600 699.450 343.950 ;
        RECT 692.400 337.350 693.600 338.100 ;
        RECT 698.400 337.350 699.600 339.600 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 697.950 334.950 700.050 337.050 ;
        RECT 682.950 331.800 685.050 333.900 ;
        RECT 689.400 333.000 690.600 334.650 ;
        RECT 695.400 333.900 696.600 334.650 ;
        RECT 688.950 328.950 691.050 333.000 ;
        RECT 694.950 328.950 697.050 333.900 ;
        RECT 689.400 322.050 690.450 328.950 ;
        RECT 688.950 319.950 691.050 322.050 ;
        RECT 704.400 316.050 705.450 383.400 ;
        RECT 721.950 379.950 724.050 382.050 ;
        RECT 712.950 371.100 715.050 373.200 ;
        RECT 722.400 372.600 723.450 379.950 ;
        RECT 713.400 370.350 714.600 371.100 ;
        RECT 722.400 370.350 723.600 372.600 ;
        RECT 713.100 367.950 715.200 370.050 ;
        RECT 718.500 367.950 720.600 370.050 ;
        RECT 721.800 367.950 723.900 370.050 ;
        RECT 719.400 366.900 720.600 367.650 ;
        RECT 728.400 366.900 729.450 388.950 ;
        RECT 737.400 373.200 738.450 407.400 ;
        RECT 740.400 400.050 741.450 415.950 ;
        RECT 743.400 403.050 744.450 433.950 ;
        RECT 758.400 418.200 759.450 499.950 ;
        RECT 761.400 472.050 762.450 517.950 ;
        RECT 763.950 517.800 766.050 519.900 ;
        RECT 766.950 517.950 769.050 520.050 ;
        RECT 769.950 517.950 772.050 520.050 ;
        RECT 777.900 519.300 780.000 521.100 ;
        RECT 781.800 518.100 783.900 520.200 ;
        RECT 786.000 518.700 786.900 524.100 ;
        RECT 787.800 523.950 789.900 526.050 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 788.400 522.450 789.600 523.650 ;
        RECT 788.400 521.400 792.450 522.450 ;
        RECT 764.400 496.050 765.450 517.800 ;
        RECT 782.400 515.550 783.600 517.800 ;
        RECT 785.100 516.600 787.200 518.700 ;
        RECT 782.400 511.050 783.450 515.550 ;
        RECT 791.400 514.050 792.450 521.400 ;
        RECT 790.950 511.950 793.050 514.050 ;
        RECT 781.950 508.950 784.050 511.050 ;
        RECT 794.400 510.450 795.450 553.950 ;
        RECT 812.400 544.050 813.450 566.400 ;
        RECT 817.950 562.950 820.050 567.000 ;
        RECT 827.400 566.400 834.600 567.450 ;
        RECT 811.950 541.950 814.050 544.050 ;
        RECT 830.400 532.050 831.450 566.400 ;
        RECT 838.950 565.800 841.050 567.900 ;
        RECT 832.950 562.950 835.050 565.050 ;
        RECT 829.950 529.950 832.050 532.050 ;
        RECT 805.950 527.100 808.050 529.200 ;
        RECT 820.950 528.450 823.050 529.200 ;
        RECT 833.400 528.600 834.450 562.950 ;
        RECT 839.400 556.050 840.450 565.800 ;
        RECT 845.400 565.050 846.450 580.950 ;
        RECT 844.950 562.950 847.050 565.050 ;
        RECT 848.400 556.050 849.450 592.950 ;
        RECT 850.950 586.950 853.050 592.050 ;
        RECT 854.400 586.050 855.450 673.950 ;
        RECT 866.400 673.050 867.450 683.100 ;
        RECT 872.400 682.350 873.600 683.100 ;
        RECT 878.400 682.350 879.600 684.600 ;
        RECT 871.950 679.950 874.050 682.050 ;
        RECT 874.950 679.950 877.050 682.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 875.400 677.400 876.600 679.650 ;
        RECT 881.400 679.050 882.600 679.650 ;
        RECT 881.400 677.400 886.050 679.050 ;
        RECT 865.950 670.950 868.050 673.050 ;
        RECT 875.400 658.050 876.450 677.400 ;
        RECT 882.000 676.950 886.050 677.400 ;
        RECT 880.950 673.950 883.050 676.050 ;
        RECT 877.950 670.950 880.050 673.050 ;
        RECT 856.950 655.950 859.050 658.050 ;
        RECT 868.950 655.950 871.050 658.050 ;
        RECT 874.950 655.950 877.050 658.050 ;
        RECT 857.400 643.050 858.450 655.950 ;
        RECT 862.950 650.100 865.050 652.200 ;
        RECT 869.400 651.600 870.450 655.950 ;
        RECT 863.400 649.350 864.600 650.100 ;
        RECT 869.400 649.350 870.600 651.600 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 866.400 645.900 867.600 646.650 ;
        RECT 865.950 643.800 868.050 645.900 ;
        RECT 872.400 644.400 873.600 646.650 ;
        RECT 856.950 640.950 859.050 643.050 ;
        RECT 868.950 640.950 871.050 643.050 ;
        RECT 856.950 634.950 859.050 637.050 ;
        RECT 857.400 592.050 858.450 634.950 ;
        RECT 869.400 607.050 870.450 640.950 ;
        RECT 872.400 637.050 873.450 644.400 ;
        RECT 878.400 637.050 879.450 670.950 ;
        RECT 881.400 643.050 882.450 673.950 ;
        RECT 887.400 673.050 888.450 685.950 ;
        RECT 890.400 682.050 891.450 718.950 ;
        RECT 896.400 717.450 897.450 722.400 ;
        RECT 901.950 718.950 904.050 723.900 ;
        RECT 907.950 721.950 910.050 724.050 ;
        RECT 917.400 723.900 918.600 724.650 ;
        RECT 916.950 721.800 919.050 723.900 ;
        RECT 893.400 716.400 897.450 717.450 ;
        RECT 893.400 703.050 894.450 716.400 ;
        RECT 904.950 715.950 907.050 718.050 ;
        RECT 919.950 715.950 922.050 718.050 ;
        RECT 892.950 700.950 895.050 703.050 ;
        RECT 893.400 685.050 894.450 700.950 ;
        RECT 892.950 682.950 895.050 685.050 ;
        RECT 895.950 683.100 898.050 685.200 ;
        RECT 901.950 684.000 904.050 688.050 ;
        RECT 905.400 685.050 906.450 715.950 ;
        RECT 907.950 703.950 910.050 706.050 ;
        RECT 908.400 694.050 909.450 703.950 ;
        RECT 907.950 691.950 910.050 694.050 ;
        RECT 896.400 682.350 897.600 683.100 ;
        RECT 902.400 682.350 903.600 684.000 ;
        RECT 904.950 682.950 907.050 685.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 895.950 679.950 898.050 682.050 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 886.950 670.950 889.050 673.050 ;
        RECT 890.400 667.050 891.450 679.950 ;
        RECT 899.400 678.900 900.600 679.650 ;
        RECT 908.400 679.050 909.450 691.950 ;
        RECT 913.950 683.100 916.050 685.200 ;
        RECT 920.400 684.600 921.450 715.950 ;
        RECT 926.400 703.050 927.450 748.950 ;
        RECT 937.950 742.950 940.050 745.050 ;
        RECT 928.950 728.100 931.050 730.200 ;
        RECT 938.400 729.600 939.450 742.950 ;
        RECT 929.400 706.050 930.450 728.100 ;
        RECT 938.400 727.350 939.600 729.600 ;
        RECT 943.950 728.100 946.050 730.200 ;
        RECT 944.400 727.350 945.600 728.100 ;
        RECT 934.950 724.950 937.050 727.050 ;
        RECT 937.950 724.950 940.050 727.050 ;
        RECT 940.950 724.950 943.050 727.050 ;
        RECT 943.950 724.950 946.050 727.050 ;
        RECT 935.400 723.900 936.600 724.650 ;
        RECT 941.400 723.900 942.600 724.650 ;
        RECT 934.950 721.800 937.050 723.900 ;
        RECT 940.950 721.800 943.050 723.900 ;
        RECT 946.950 721.800 949.050 723.900 ;
        RECT 928.950 703.950 931.050 706.050 ;
        RECT 925.950 700.950 928.050 703.050 ;
        RECT 914.400 682.350 915.600 683.100 ;
        RECT 920.400 682.350 921.600 684.600 ;
        RECT 925.950 683.100 928.050 685.200 ;
        RECT 931.950 683.100 934.050 685.200 ;
        RECT 937.950 683.100 940.050 685.200 ;
        RECT 943.800 683.100 945.900 685.200 ;
        RECT 947.400 685.050 948.450 721.800 ;
        RECT 926.400 682.350 927.600 683.100 ;
        RECT 913.950 679.950 916.050 682.050 ;
        RECT 916.950 679.950 919.050 682.050 ;
        RECT 919.950 679.950 922.050 682.050 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 925.950 679.950 928.050 682.050 ;
        RECT 898.950 676.800 901.050 678.900 ;
        RECT 907.950 676.950 910.050 679.050 ;
        RECT 917.400 677.400 918.600 679.650 ;
        RECT 923.400 678.900 924.600 679.650 ;
        RECT 901.950 673.950 904.050 676.050 ;
        RECT 889.950 664.950 892.050 667.050 ;
        RECT 890.400 651.600 891.450 664.950 ;
        RECT 890.400 649.350 891.600 651.600 ;
        RECT 895.950 650.100 898.050 652.200 ;
        RECT 896.400 649.350 897.600 650.100 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 895.950 646.950 898.050 649.050 ;
        RECT 887.400 644.400 888.600 646.650 ;
        RECT 893.400 644.400 894.600 646.650 ;
        RECT 880.950 640.950 883.050 643.050 ;
        RECT 871.950 634.950 874.050 637.050 ;
        RECT 877.950 634.950 880.050 637.050 ;
        RECT 887.400 631.050 888.450 644.400 ;
        RECT 893.400 643.050 894.450 644.400 ;
        RECT 892.950 640.950 895.050 643.050 ;
        RECT 902.400 642.450 903.450 673.950 ;
        RECT 917.400 673.050 918.450 677.400 ;
        RECT 922.950 676.800 925.050 678.900 ;
        RECT 923.400 675.450 924.450 676.800 ;
        RECT 920.400 674.400 924.450 675.450 ;
        RECT 904.950 670.950 907.050 673.050 ;
        RECT 916.950 670.950 919.050 673.050 ;
        RECT 905.400 645.450 906.450 670.950 ;
        RECT 910.950 650.100 913.050 652.200 ;
        RECT 911.400 649.350 912.600 650.100 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 914.400 645.900 915.600 646.650 ;
        RECT 905.400 644.400 909.450 645.450 ;
        RECT 902.400 641.400 906.450 642.450 ;
        RECT 871.950 628.950 874.050 631.050 ;
        RECT 886.950 628.950 889.050 631.050 ;
        RECT 859.950 606.600 864.000 607.050 ;
        RECT 859.950 604.950 864.600 606.600 ;
        RECT 868.950 604.950 871.050 607.050 ;
        RECT 863.400 604.350 864.600 604.950 ;
        RECT 872.400 604.050 873.450 628.950 ;
        RECT 880.950 605.100 883.050 607.200 ;
        RECT 881.400 604.350 882.600 605.100 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 871.950 601.950 874.050 604.050 ;
        RECT 877.950 601.950 880.050 604.050 ;
        RECT 880.950 601.950 883.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 859.950 598.950 862.050 601.050 ;
        RECT 866.400 600.000 867.600 601.650 ;
        RECT 860.400 594.450 861.450 598.950 ;
        RECT 865.950 595.950 868.050 600.000 ;
        RECT 868.950 598.950 871.050 601.050 ;
        RECT 878.400 600.450 879.600 601.650 ;
        RECT 875.400 599.400 879.600 600.450 ;
        RECT 884.400 599.400 885.600 601.650 ;
        RECT 865.950 594.450 868.050 594.900 ;
        RECT 860.400 593.400 868.050 594.450 ;
        RECT 865.950 592.800 868.050 593.400 ;
        RECT 856.950 589.950 859.050 592.050 ;
        RECT 859.950 589.950 862.050 592.050 ;
        RECT 853.950 583.950 856.050 586.050 ;
        RECT 860.400 583.050 861.450 589.950 ;
        RECT 865.950 589.800 868.050 591.900 ;
        RECT 862.950 586.950 865.050 589.050 ;
        RECT 859.950 580.950 862.050 583.050 ;
        RECT 856.950 572.100 859.050 574.200 ;
        RECT 863.400 573.600 864.450 586.950 ;
        RECT 866.400 574.050 867.450 589.800 ;
        RECT 857.400 571.350 858.600 572.100 ;
        RECT 863.400 571.350 864.600 573.600 ;
        RECT 865.950 571.950 868.050 574.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 854.400 567.900 855.600 568.650 ;
        RECT 853.950 565.800 856.050 567.900 ;
        RECT 860.400 567.000 861.600 568.650 ;
        RECT 859.950 562.950 862.050 567.000 ;
        RECT 869.400 562.050 870.450 598.950 ;
        RECT 875.400 595.050 876.450 599.400 ;
        RECT 874.950 592.950 877.050 595.050 ;
        RECT 884.400 586.050 885.450 599.400 ;
        RECT 889.950 598.800 892.050 600.900 ;
        RECT 883.950 583.950 886.050 586.050 ;
        RECT 877.950 580.950 880.050 583.050 ;
        RECT 878.400 573.600 879.450 580.950 ;
        RECT 890.400 577.050 891.450 598.800 ;
        RECT 893.400 589.050 894.450 640.950 ;
        RECT 895.950 605.100 898.050 607.200 ;
        RECT 901.950 605.100 904.050 607.200 ;
        RECT 905.400 606.600 906.450 641.400 ;
        RECT 908.400 631.050 909.450 644.400 ;
        RECT 913.950 643.800 916.050 645.900 ;
        RECT 920.400 640.050 921.450 674.400 ;
        RECT 932.400 673.050 933.450 683.100 ;
        RECT 938.400 682.350 939.600 683.100 ;
        RECT 944.400 682.350 945.600 683.100 ;
        RECT 946.950 682.950 949.050 685.050 ;
        RECT 937.950 679.950 940.050 682.050 ;
        RECT 940.950 679.950 943.050 682.050 ;
        RECT 943.950 679.950 946.050 682.050 ;
        RECT 941.400 678.900 942.600 679.650 ;
        RECT 940.950 676.800 943.050 678.900 ;
        RECT 931.950 670.950 934.050 673.050 ;
        RECT 940.950 670.950 943.050 673.050 ;
        RECT 925.950 661.950 928.050 664.050 ;
        RECT 926.400 651.600 927.450 661.950 ;
        RECT 926.400 649.350 927.600 651.600 ;
        RECT 931.950 650.100 934.050 652.200 ;
        RECT 932.400 649.350 933.600 650.100 ;
        RECT 925.950 646.950 928.050 649.050 ;
        RECT 928.950 646.950 931.050 649.050 ;
        RECT 931.950 646.950 934.050 649.050 ;
        RECT 934.950 646.950 937.050 649.050 ;
        RECT 929.400 645.000 930.600 646.650 ;
        RECT 928.950 640.950 931.050 645.000 ;
        RECT 935.400 644.400 936.600 646.650 ;
        RECT 935.400 640.050 936.450 644.400 ;
        RECT 937.950 642.450 940.050 643.050 ;
        RECT 941.400 642.450 942.450 670.950 ;
        RECT 937.950 641.400 942.450 642.450 ;
        RECT 937.950 640.950 940.050 641.400 ;
        RECT 919.950 637.950 922.050 640.050 ;
        RECT 934.950 637.950 937.050 640.050 ;
        RECT 907.950 628.950 910.050 631.050 ;
        RECT 892.950 586.950 895.050 589.050 ;
        RECT 896.400 583.050 897.450 605.100 ;
        RECT 902.400 598.050 903.450 605.100 ;
        RECT 905.400 604.350 906.600 606.600 ;
        RECT 913.950 605.100 916.050 607.200 ;
        RECT 914.400 604.350 915.600 605.100 ;
        RECT 905.400 601.950 907.500 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 920.100 601.950 922.200 604.050 ;
        RECT 911.400 600.900 912.600 601.650 ;
        RECT 910.950 598.800 913.050 600.900 ;
        RECT 920.400 599.400 921.600 601.650 ;
        RECT 901.950 595.950 904.050 598.050 ;
        RECT 910.950 595.650 913.050 597.750 ;
        RECT 895.950 580.950 898.050 583.050 ;
        RECT 878.400 571.350 879.600 573.600 ;
        RECT 883.950 573.000 886.050 577.050 ;
        RECT 889.950 574.950 892.050 577.050 ;
        RECT 884.400 571.350 885.600 573.000 ;
        RECT 874.950 568.950 877.050 571.050 ;
        RECT 877.950 568.950 880.050 571.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 871.950 565.950 874.050 568.050 ;
        RECT 881.400 567.900 882.600 568.650 ;
        RECT 859.950 559.800 862.050 561.900 ;
        RECT 868.950 559.950 871.050 562.050 ;
        RECT 872.400 561.450 873.450 565.950 ;
        RECT 880.950 565.800 883.050 567.900 ;
        RECT 890.400 562.050 891.450 574.950 ;
        RECT 892.950 572.100 895.050 574.200 ;
        RECT 898.950 572.100 901.050 574.200 ;
        RECT 904.950 573.000 907.050 577.050 ;
        RECT 872.400 560.400 876.450 561.450 ;
        RECT 838.950 553.950 841.050 556.050 ;
        RECT 847.950 553.950 850.050 556.050 ;
        RECT 844.950 547.950 847.050 550.050 ;
        RECT 835.950 529.950 838.050 532.050 ;
        RECT 824.400 528.450 825.600 528.600 ;
        RECT 820.950 527.400 825.600 528.450 ;
        RECT 820.950 527.100 823.050 527.400 ;
        RECT 806.400 526.350 807.600 527.100 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 808.950 523.950 811.050 526.050 ;
        RECT 803.400 522.900 804.600 523.650 ;
        RECT 802.950 520.800 805.050 522.900 ;
        RECT 809.400 522.000 810.600 523.650 ;
        RECT 808.950 517.950 811.050 522.000 ;
        RECT 802.950 511.950 805.050 514.050 ;
        RECT 791.400 509.400 795.450 510.450 ;
        RECT 769.950 499.950 772.050 502.050 ;
        RECT 781.950 499.950 784.050 502.050 ;
        RECT 763.950 493.950 766.050 496.050 ;
        RECT 770.400 495.600 771.450 499.950 ;
        RECT 770.400 493.350 771.600 495.600 ;
        RECT 775.950 494.100 778.050 496.200 ;
        RECT 776.400 493.350 777.600 494.100 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 772.950 490.950 775.050 493.050 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 767.400 489.900 768.600 490.650 ;
        RECT 766.950 487.800 769.050 489.900 ;
        RECT 773.400 488.400 774.600 490.650 ;
        RECT 760.950 469.950 763.050 472.050 ;
        RECT 767.400 463.050 768.450 487.800 ;
        RECT 773.400 475.050 774.450 488.400 ;
        RECT 778.950 484.950 781.050 487.050 ;
        RECT 772.950 472.950 775.050 475.050 ;
        RECT 760.950 460.950 763.050 463.050 ;
        RECT 766.950 460.950 769.050 463.050 ;
        RECT 761.400 451.050 762.450 460.950 ;
        RECT 766.950 454.950 769.050 457.050 ;
        RECT 760.950 448.950 763.050 451.050 ;
        RECT 767.400 450.600 768.450 454.950 ;
        RECT 767.400 448.350 768.600 450.600 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 766.950 445.950 769.050 448.050 ;
        RECT 760.950 442.950 763.050 445.050 ;
        RECT 764.400 443.400 765.600 445.650 ;
        RECT 761.400 424.050 762.450 442.950 ;
        RECT 764.400 430.050 765.450 443.400 ;
        RECT 763.950 427.950 766.050 430.050 ;
        RECT 760.950 421.950 763.050 424.050 ;
        RECT 748.950 416.100 751.050 418.200 ;
        RECT 757.950 416.100 760.050 418.200 ;
        RECT 761.400 417.450 762.450 421.950 ;
        RECT 764.400 417.450 765.600 417.600 ;
        RECT 761.400 416.400 765.600 417.450 ;
        RECT 749.400 415.350 750.600 416.100 ;
        RECT 764.400 415.350 765.600 416.400 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 763.950 412.950 766.050 415.050 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 752.400 411.000 753.600 412.650 ;
        RECT 751.950 406.950 754.050 411.000 ;
        RECT 757.950 409.950 760.050 412.050 ;
        RECT 767.400 410.400 768.600 412.650 ;
        RECT 773.400 412.050 774.450 472.950 ;
        RECT 775.950 463.950 778.050 466.050 ;
        RECT 742.950 400.950 745.050 403.050 ;
        RECT 739.950 397.950 742.050 400.050 ;
        RECT 754.950 397.950 757.050 400.050 ;
        RECT 742.950 388.950 745.050 391.050 ;
        RECT 736.950 371.100 739.050 373.200 ;
        RECT 743.400 372.600 744.450 388.950 ;
        RECT 737.400 370.350 738.600 371.100 ;
        RECT 743.400 370.350 744.600 372.600 ;
        RECT 748.950 371.100 751.050 373.200 ;
        RECT 749.400 370.350 750.600 371.100 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 739.950 367.950 742.050 370.050 ;
        RECT 742.950 367.950 745.050 370.050 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 740.400 366.900 741.600 367.650 ;
        RECT 718.950 364.800 721.050 366.900 ;
        RECT 727.950 364.800 730.050 366.900 ;
        RECT 739.950 364.800 742.050 366.900 ;
        RECT 746.400 365.400 747.600 367.650 ;
        RECT 746.400 358.050 747.450 365.400 ;
        RECT 755.400 361.050 756.450 397.950 ;
        RECT 754.950 358.950 757.050 361.050 ;
        RECT 745.950 355.950 748.050 358.050 ;
        RECT 746.400 346.050 747.450 355.950 ;
        RECT 748.950 346.950 751.050 349.050 ;
        RECT 755.400 348.450 756.450 358.950 ;
        RECT 752.400 347.400 756.450 348.450 ;
        RECT 733.950 343.950 736.050 346.050 ;
        RECT 745.950 343.950 748.050 346.050 ;
        RECT 715.950 338.100 718.050 340.200 ;
        RECT 721.950 338.100 724.050 340.200 ;
        RECT 734.400 339.600 735.450 343.950 ;
        RECT 749.400 340.050 750.450 346.950 ;
        RECT 716.400 337.350 717.600 338.100 ;
        RECT 722.400 337.350 723.600 338.100 ;
        RECT 734.400 337.350 735.600 339.600 ;
        RECT 742.950 337.950 745.050 340.050 ;
        RECT 748.950 337.950 751.050 340.050 ;
        RECT 752.400 339.600 753.450 347.400 ;
        RECT 758.400 339.600 759.450 409.950 ;
        RECT 767.400 409.050 768.450 410.400 ;
        RECT 772.950 409.950 775.050 412.050 ;
        RECT 776.400 409.050 777.450 463.950 ;
        RECT 779.400 451.050 780.450 484.950 ;
        RECT 782.400 466.050 783.450 499.950 ;
        RECT 791.400 496.200 792.450 509.400 ;
        RECT 790.950 494.100 793.050 496.200 ;
        RECT 796.950 495.000 799.050 499.050 ;
        RECT 791.400 493.350 792.600 494.100 ;
        RECT 797.400 493.350 798.600 495.000 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 790.950 490.950 793.050 493.050 ;
        RECT 793.950 490.950 796.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 788.400 488.400 789.600 490.650 ;
        RECT 794.400 489.000 795.600 490.650 ;
        RECT 781.950 463.950 784.050 466.050 ;
        RECT 788.400 460.050 789.450 488.400 ;
        RECT 793.950 484.950 796.050 489.000 ;
        RECT 790.950 472.950 793.050 475.050 ;
        RECT 787.950 457.950 790.050 460.050 ;
        RECT 778.950 448.950 781.050 451.050 ;
        RECT 784.950 449.100 787.050 451.200 ;
        RECT 791.400 450.600 792.450 472.950 ;
        RECT 803.400 469.050 804.450 511.950 ;
        RECT 821.400 505.050 822.450 527.100 ;
        RECT 824.400 526.350 825.600 527.400 ;
        RECT 833.400 526.350 834.600 528.600 ;
        RECT 824.100 523.950 826.200 526.050 ;
        RECT 829.500 523.950 831.600 526.050 ;
        RECT 832.800 523.950 834.900 526.050 ;
        RECT 830.400 521.400 831.600 523.650 ;
        RECT 830.400 520.050 831.450 521.400 ;
        RECT 829.950 519.450 832.050 520.050 ;
        RECT 829.950 519.000 834.450 519.450 ;
        RECT 829.950 518.400 835.050 519.000 ;
        RECT 829.950 517.950 832.050 518.400 ;
        RECT 832.950 514.950 835.050 518.400 ;
        RECT 820.950 502.950 823.050 505.050 ;
        RECT 823.950 496.950 826.050 499.050 ;
        RECT 832.950 498.450 835.050 499.050 ;
        RECT 836.400 498.450 837.450 529.950 ;
        RECT 845.400 528.600 846.450 547.950 ;
        RECT 845.400 526.350 846.600 528.600 ;
        RECT 850.950 527.100 853.050 529.200 ;
        RECT 851.400 526.350 852.600 527.100 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 850.950 523.950 853.050 526.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 841.950 520.950 844.050 523.050 ;
        RECT 848.400 521.400 849.600 523.650 ;
        RECT 854.400 522.900 855.600 523.650 ;
        RECT 860.400 523.050 861.450 559.800 ;
        RECT 862.950 553.950 865.050 556.050 ;
        RECT 842.400 514.050 843.450 520.950 ;
        RECT 841.950 511.950 844.050 514.050 ;
        RECT 848.400 508.050 849.450 521.400 ;
        RECT 853.950 520.800 856.050 522.900 ;
        RECT 859.950 520.950 862.050 523.050 ;
        RECT 863.400 517.050 864.450 553.950 ;
        RECT 868.950 527.100 871.050 529.200 ;
        RECT 875.400 528.600 876.450 560.400 ;
        RECT 889.950 559.950 892.050 562.050 ;
        RECT 893.400 556.050 894.450 572.100 ;
        RECT 899.400 571.350 900.600 572.100 ;
        RECT 905.400 571.350 906.600 573.000 ;
        RECT 898.950 568.950 901.050 571.050 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 902.400 567.900 903.600 568.650 ;
        RECT 901.950 565.800 904.050 567.900 ;
        RECT 907.950 559.950 910.050 562.050 ;
        RECT 892.950 553.950 895.050 556.050 ;
        RECT 889.950 532.950 892.050 535.050 ;
        RECT 869.400 526.350 870.600 527.100 ;
        RECT 875.400 526.350 876.600 528.600 ;
        RECT 880.950 528.000 883.050 532.050 ;
        RECT 886.950 529.950 889.050 532.050 ;
        RECT 881.400 526.350 882.600 528.000 ;
        RECT 868.950 523.950 871.050 526.050 ;
        RECT 871.950 523.950 874.050 526.050 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 880.950 523.950 883.050 526.050 ;
        RECT 865.950 520.800 868.050 522.900 ;
        RECT 872.400 521.400 873.600 523.650 ;
        RECT 878.400 522.900 879.600 523.650 ;
        RECT 856.950 514.950 859.050 517.050 ;
        RECT 862.950 514.950 865.050 517.050 ;
        RECT 847.950 505.950 850.050 508.050 ;
        RECT 844.950 502.950 847.050 505.050 ;
        RECT 832.950 497.400 837.450 498.450 ;
        RECT 805.950 493.950 808.050 496.050 ;
        RECT 814.950 494.100 817.050 496.200 ;
        RECT 802.950 466.950 805.050 469.050 ;
        RECT 793.950 463.950 796.050 466.050 ;
        RECT 794.400 457.050 795.450 463.950 ;
        RECT 806.400 460.050 807.450 493.950 ;
        RECT 815.400 493.350 816.600 494.100 ;
        RECT 811.950 490.950 814.050 493.050 ;
        RECT 814.950 490.950 817.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 812.400 488.400 813.600 490.650 ;
        RECT 818.400 489.900 819.600 490.650 ;
        RECT 824.400 489.900 825.450 496.950 ;
        RECT 832.950 495.000 835.050 497.400 ;
        RECT 833.400 493.350 834.600 495.000 ;
        RECT 838.950 494.100 841.050 496.200 ;
        RECT 839.400 493.350 840.600 494.100 ;
        RECT 829.950 490.950 832.050 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 812.400 484.050 813.450 488.400 ;
        RECT 817.950 487.800 820.050 489.900 ;
        RECT 823.950 487.800 826.050 489.900 ;
        RECT 830.400 489.000 831.600 490.650 ;
        RECT 811.950 481.950 814.050 484.050 ;
        RECT 820.950 481.950 823.050 487.050 ;
        RECT 829.950 484.950 832.050 489.000 ;
        RECT 836.400 488.400 837.600 490.650 ;
        RECT 836.400 486.450 837.450 488.400 ;
        RECT 841.950 487.950 844.050 490.050 ;
        RECT 836.400 485.400 840.450 486.450 ;
        RECT 817.950 472.950 820.050 475.050 ;
        RECT 796.950 457.950 799.050 460.050 ;
        RECT 805.950 457.950 808.050 460.050 ;
        RECT 793.950 454.950 796.050 457.050 ;
        RECT 785.400 448.350 786.600 449.100 ;
        RECT 791.400 448.350 792.600 450.600 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 787.950 445.950 790.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 778.950 442.950 781.050 445.050 ;
        RECT 782.400 443.400 783.600 445.650 ;
        RECT 788.400 443.400 789.600 445.650 ;
        RECT 779.400 439.050 780.450 442.950 ;
        RECT 778.950 436.950 781.050 439.050 ;
        RECT 782.400 418.200 783.450 443.400 ;
        RECT 788.400 441.450 789.450 443.400 ;
        RECT 793.950 442.950 796.050 445.050 ;
        RECT 788.400 440.400 792.450 441.450 ;
        RECT 787.950 436.950 790.050 439.050 ;
        RECT 781.950 416.100 784.050 418.200 ;
        RECT 788.400 417.600 789.450 436.950 ;
        RECT 791.400 433.050 792.450 440.400 ;
        RECT 790.950 430.950 793.050 433.050 ;
        RECT 782.400 415.350 783.600 416.100 ;
        RECT 788.400 415.350 789.600 417.600 ;
        RECT 794.400 417.450 795.450 442.950 ;
        RECT 797.400 421.050 798.450 457.950 ;
        RECT 805.950 454.800 808.050 456.900 ;
        RECT 799.950 451.950 802.050 454.050 ;
        RECT 796.950 418.950 799.050 421.050 ;
        RECT 794.400 416.400 798.450 417.450 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 784.950 412.950 787.050 415.050 ;
        RECT 787.950 412.950 790.050 415.050 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 785.400 411.000 786.600 412.650 ;
        RECT 791.400 411.900 792.600 412.650 ;
        RECT 767.400 406.950 772.050 409.050 ;
        RECT 775.950 406.950 778.050 409.050 ;
        RECT 784.950 406.950 787.050 411.000 ;
        RECT 790.950 409.800 793.050 411.900 ;
        RECT 767.400 403.050 768.450 406.950 ;
        RECT 766.950 400.950 769.050 403.050 ;
        RECT 769.950 379.950 772.050 382.050 ;
        RECT 787.950 379.950 790.050 382.050 ;
        RECT 763.950 371.100 766.050 373.200 ;
        RECT 770.400 372.600 771.450 379.950 ;
        RECT 781.950 376.950 784.050 379.050 ;
        RECT 764.400 370.350 765.600 371.100 ;
        RECT 770.400 370.350 771.600 372.600 ;
        RECT 778.950 371.100 781.050 373.200 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 769.950 367.950 772.050 370.050 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 760.950 364.950 763.050 367.050 ;
        RECT 767.400 365.400 768.600 367.650 ;
        RECT 773.400 365.400 774.600 367.650 ;
        RECT 779.400 366.450 780.450 371.100 ;
        RECT 776.400 365.400 780.450 366.450 ;
        RECT 761.400 349.050 762.450 364.950 ;
        RECT 767.400 358.050 768.450 365.400 ;
        RECT 766.950 355.950 769.050 358.050 ;
        RECT 760.950 346.950 763.050 349.050 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 713.400 332.400 714.600 334.650 ;
        RECT 719.400 333.000 720.600 334.650 ;
        RECT 737.400 333.900 738.600 334.650 ;
        RECT 713.400 322.050 714.450 332.400 ;
        RECT 718.950 328.950 721.050 333.000 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 743.400 328.050 744.450 337.950 ;
        RECT 752.400 337.350 753.600 339.600 ;
        RECT 758.400 337.350 759.600 339.600 ;
        RECT 766.950 338.100 769.050 340.200 ;
        RECT 773.400 339.450 774.450 365.400 ;
        RECT 776.400 340.200 777.450 365.400 ;
        RECT 782.400 364.050 783.450 376.950 ;
        RECT 788.400 372.600 789.450 379.950 ;
        RECT 797.400 376.050 798.450 416.400 ;
        RECT 800.400 411.450 801.450 451.950 ;
        RECT 806.400 450.600 807.450 454.800 ;
        RECT 806.400 448.350 807.600 450.600 ;
        RECT 811.950 450.000 814.050 454.050 ;
        RECT 818.400 451.050 819.450 472.950 ;
        RECT 812.400 448.350 813.600 450.000 ;
        RECT 817.950 448.950 820.050 451.050 ;
        RECT 805.950 445.950 808.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 809.400 443.400 810.600 445.650 ;
        RECT 815.400 445.050 816.600 445.650 ;
        RECT 815.400 443.400 820.050 445.050 ;
        RECT 809.400 424.050 810.450 443.400 ;
        RECT 816.000 442.950 820.050 443.400 ;
        RECT 821.400 442.050 822.450 481.950 ;
        RECT 826.950 449.100 829.050 451.200 ;
        RECT 832.950 450.000 835.050 454.050 ;
        RECT 839.400 451.050 840.450 485.400 ;
        RECT 842.400 481.050 843.450 487.950 ;
        RECT 841.950 478.950 844.050 481.050 ;
        RECT 827.400 448.350 828.600 449.100 ;
        RECT 833.400 448.350 834.600 450.000 ;
        RECT 838.950 448.950 841.050 451.050 ;
        RECT 841.950 449.100 844.050 451.200 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 829.950 445.950 832.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 830.400 443.400 831.600 445.650 ;
        RECT 836.400 444.000 837.600 445.650 ;
        RECT 842.400 444.450 843.450 449.100 ;
        RECT 814.950 439.950 817.050 442.050 ;
        RECT 820.950 439.950 823.050 442.050 ;
        RECT 808.950 421.950 811.050 424.050 ;
        RECT 805.950 417.000 808.050 421.050 ;
        RECT 806.400 415.350 807.600 417.000 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 809.400 411.900 810.600 412.650 ;
        RECT 815.400 412.050 816.450 439.950 ;
        RECT 830.400 433.050 831.450 443.400 ;
        RECT 835.950 439.950 838.050 444.000 ;
        RECT 839.400 443.400 843.450 444.450 ;
        RECT 839.400 436.050 840.450 443.400 ;
        RECT 845.400 442.050 846.450 502.950 ;
        RECT 857.400 499.050 858.450 514.950 ;
        RECT 859.950 511.950 862.050 514.050 ;
        RECT 850.950 494.100 853.050 496.200 ;
        RECT 856.950 495.000 859.050 499.050 ;
        RECT 860.400 496.050 861.450 511.950 ;
        RECT 851.400 493.350 852.600 494.100 ;
        RECT 857.400 493.350 858.600 495.000 ;
        RECT 859.950 493.950 862.050 496.050 ;
        RECT 850.950 490.950 853.050 493.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 847.950 487.950 850.050 490.050 ;
        RECT 854.400 489.900 855.600 490.650 ;
        RECT 848.400 451.050 849.450 487.950 ;
        RECT 853.950 487.800 856.050 489.900 ;
        RECT 859.950 487.950 862.050 490.050 ;
        RECT 860.400 474.450 861.450 487.950 ;
        RECT 863.400 478.050 864.450 514.950 ;
        RECT 866.400 496.050 867.450 520.800 ;
        RECT 872.400 517.050 873.450 521.400 ;
        RECT 877.950 520.800 880.050 522.900 ;
        RECT 871.950 514.950 874.050 517.050 ;
        RECT 865.950 493.950 868.050 496.050 ;
        RECT 872.400 495.600 873.450 514.950 ;
        RECT 887.400 508.050 888.450 529.950 ;
        RECT 890.400 529.200 891.450 532.950 ;
        RECT 895.950 531.450 900.000 532.050 ;
        RECT 895.950 529.950 900.450 531.450 ;
        RECT 889.950 527.100 892.050 529.200 ;
        RECT 899.400 528.600 900.450 529.950 ;
        RECT 886.950 505.950 889.050 508.050 ;
        RECT 886.950 499.950 889.050 502.050 ;
        RECT 872.400 493.350 873.600 495.600 ;
        RECT 877.950 494.100 880.050 496.200 ;
        RECT 878.400 493.350 879.600 494.100 ;
        RECT 883.950 493.950 886.050 496.050 ;
        RECT 868.950 490.950 871.050 493.050 ;
        RECT 871.950 490.950 874.050 493.050 ;
        RECT 874.950 490.950 877.050 493.050 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 865.950 484.950 868.050 490.050 ;
        RECT 869.400 489.000 870.600 490.650 ;
        RECT 875.400 489.000 876.600 490.650 ;
        RECT 884.400 490.050 885.450 493.950 ;
        RECT 868.950 484.950 871.050 489.000 ;
        RECT 874.950 484.950 877.050 489.000 ;
        RECT 883.950 487.950 886.050 490.050 ;
        RECT 862.950 475.950 865.050 478.050 ;
        RECT 860.400 473.400 864.450 474.450 ;
        RECT 853.950 454.950 856.050 457.050 ;
        RECT 854.400 451.200 855.450 454.950 ;
        RECT 847.950 448.950 850.050 451.050 ;
        RECT 853.950 449.100 856.050 451.200 ;
        RECT 859.950 449.100 862.050 451.200 ;
        RECT 863.400 451.050 864.450 473.400 ;
        RECT 854.400 448.350 855.600 449.100 ;
        RECT 860.400 448.350 861.600 449.100 ;
        RECT 862.950 448.950 865.050 451.050 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 847.950 444.450 850.050 445.050 ;
        RECT 851.400 444.450 852.600 445.650 ;
        RECT 847.950 443.400 852.600 444.450 ;
        RECT 857.400 444.000 858.600 445.650 ;
        RECT 847.950 442.950 850.050 443.400 ;
        RECT 841.950 439.950 844.050 442.050 ;
        RECT 844.950 439.950 847.050 442.050 ;
        RECT 838.950 433.950 841.050 436.050 ;
        RECT 829.950 430.950 832.050 433.050 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 823.950 416.100 826.050 418.200 ;
        RECT 830.400 417.600 831.450 424.950 ;
        RECT 824.400 415.350 825.600 416.100 ;
        RECT 830.400 415.350 831.600 417.600 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 802.950 411.450 805.050 411.900 ;
        RECT 800.400 410.400 805.050 411.450 ;
        RECT 802.950 409.800 805.050 410.400 ;
        RECT 808.950 409.800 811.050 411.900 ;
        RECT 814.950 409.950 817.050 412.050 ;
        RECT 820.950 409.950 823.050 412.050 ;
        RECT 827.400 410.400 828.600 412.650 ;
        RECT 833.400 410.400 834.600 412.650 ;
        RECT 796.950 373.950 799.050 376.050 ;
        RECT 788.400 370.350 789.600 372.600 ;
        RECT 793.950 371.100 796.050 373.200 ;
        RECT 794.400 370.350 795.600 371.100 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 790.950 367.950 793.050 370.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 791.400 365.400 792.600 367.650 ;
        RECT 797.400 366.450 798.600 367.650 ;
        RECT 803.400 366.450 804.450 409.800 ;
        RECT 805.950 388.950 808.050 391.050 ;
        RECT 806.400 373.050 807.450 388.950 ;
        RECT 821.400 382.050 822.450 409.950 ;
        RECT 827.400 408.450 828.450 410.400 ;
        RECT 824.400 407.400 828.450 408.450 ;
        RECT 820.950 379.950 823.050 382.050 ;
        RECT 811.950 376.950 814.050 379.050 ;
        RECT 805.950 370.950 808.050 373.050 ;
        RECT 812.400 372.600 813.450 376.950 ;
        RECT 812.400 370.350 813.600 372.600 ;
        RECT 817.950 371.100 820.050 373.200 ;
        RECT 818.400 370.350 819.600 371.100 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 809.400 366.900 810.600 367.650 ;
        RECT 797.400 365.400 804.450 366.450 ;
        RECT 781.950 361.950 784.050 364.050 ;
        RECT 787.950 358.950 790.050 361.050 ;
        RECT 781.950 343.950 784.050 346.050 ;
        RECT 770.400 338.400 774.450 339.450 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 757.950 334.950 760.050 337.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 755.400 333.900 756.600 334.650 ;
        RECT 761.400 333.900 762.600 334.650 ;
        RECT 754.950 331.800 757.050 333.900 ;
        RECT 760.950 331.800 763.050 333.900 ;
        RECT 767.400 333.450 768.450 338.100 ;
        RECT 764.400 332.400 768.450 333.450 ;
        RECT 755.400 330.300 756.450 331.800 ;
        RECT 760.950 330.300 763.050 330.750 ;
        RECT 755.400 329.250 763.050 330.300 ;
        RECT 760.950 328.650 763.050 329.250 ;
        RECT 764.400 328.050 765.450 332.400 ;
        RECT 770.400 328.050 771.450 338.400 ;
        RECT 775.950 338.100 778.050 340.200 ;
        RECT 782.400 339.600 783.450 343.950 ;
        RECT 788.400 340.050 789.450 358.950 ;
        RECT 791.400 355.050 792.450 365.400 ;
        RECT 808.950 364.800 811.050 366.900 ;
        RECT 815.400 365.400 816.600 367.650 ;
        RECT 793.950 361.950 796.050 364.050 ;
        RECT 790.950 352.950 793.050 355.050 ;
        RECT 790.950 343.950 793.050 346.050 ;
        RECT 776.400 337.350 777.600 338.100 ;
        RECT 782.400 337.350 783.600 339.600 ;
        RECT 787.950 337.950 790.050 340.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 779.400 333.000 780.600 334.650 ;
        RECT 785.400 333.900 786.600 334.650 ;
        RECT 778.950 328.950 781.050 333.000 ;
        RECT 784.950 331.800 787.050 333.900 ;
        RECT 787.950 331.950 790.050 334.050 ;
        RECT 791.400 333.900 792.450 343.950 ;
        RECT 794.400 340.050 795.450 361.950 ;
        RECT 805.950 349.950 808.050 352.050 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 799.950 339.000 802.050 343.050 ;
        RECT 806.400 339.600 807.450 349.950 ;
        RECT 809.400 349.050 810.450 364.800 ;
        RECT 811.950 361.950 814.050 364.050 ;
        RECT 808.950 346.950 811.050 349.050 ;
        RECT 800.400 337.350 801.600 339.000 ;
        RECT 806.400 337.350 807.600 339.600 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 797.400 333.900 798.600 334.650 ;
        RECT 803.400 333.900 804.600 334.650 ;
        RECT 742.950 325.950 745.050 328.050 ;
        RECT 763.950 325.950 766.050 328.050 ;
        RECT 769.950 325.950 772.050 328.050 ;
        RECT 712.950 319.950 715.050 322.050 ;
        RECT 667.950 313.950 670.050 316.050 ;
        RECT 679.950 313.950 682.050 316.050 ;
        RECT 691.950 313.950 694.050 316.050 ;
        RECT 703.950 313.950 706.050 316.050 ;
        RECT 680.400 301.050 681.450 313.950 ;
        RECT 692.400 307.050 693.450 313.950 ;
        RECT 745.950 310.950 748.050 313.050 ;
        RECT 754.950 310.950 757.050 313.050 ;
        RECT 700.950 307.950 703.050 310.050 ;
        RECT 691.950 304.950 694.050 307.050 ;
        RECT 679.950 298.950 682.050 301.050 ;
        RECT 612.900 291.000 621.900 291.900 ;
        RECT 612.900 290.100 615.000 291.000 ;
        RECT 618.000 289.200 620.100 290.100 ;
        RECT 612.900 288.000 620.100 289.200 ;
        RECT 612.900 287.100 615.000 288.000 ;
        RECT 610.500 283.500 612.600 285.600 ;
        RECT 617.100 284.100 619.200 286.200 ;
        RECT 621.000 285.900 621.900 291.000 ;
        RECT 622.800 289.950 624.900 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 623.400 288.450 624.600 289.650 ;
        RECT 623.400 287.400 627.450 288.450 ;
        RECT 638.400 288.000 639.600 289.650 ;
        RECT 620.400 283.800 622.500 285.900 ;
        RECT 617.400 281.550 618.600 283.800 ;
        RECT 626.400 283.050 627.450 287.400 ;
        RECT 637.950 283.950 640.050 288.000 ;
        RECT 617.400 274.050 618.450 281.550 ;
        RECT 625.950 280.950 628.050 283.050 ;
        RECT 643.950 277.950 646.050 280.050 ;
        RECT 616.950 271.950 619.050 274.050 ;
        RECT 616.950 268.800 619.050 270.900 ;
        RECT 601.950 260.100 604.050 262.200 ;
        RECT 607.950 260.100 610.050 262.200 ;
        RECT 602.400 259.350 603.600 260.100 ;
        RECT 608.400 259.350 609.600 260.100 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 605.400 254.400 606.600 256.650 ;
        RECT 611.400 255.000 612.600 256.650 ;
        RECT 595.950 241.950 598.050 244.050 ;
        RECT 595.950 229.950 598.050 232.050 ;
        RECT 592.950 220.950 595.050 223.050 ;
        RECT 589.950 215.100 592.050 217.200 ;
        RECT 590.400 214.350 591.600 215.100 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 587.400 209.400 588.600 211.650 ;
        RECT 587.400 202.050 588.450 209.400 ;
        RECT 586.950 199.950 589.050 202.050 ;
        RECT 583.950 187.950 586.050 190.050 ;
        RECT 592.950 187.950 595.050 190.050 ;
        RECT 584.400 184.050 585.450 187.950 ;
        RECT 583.950 181.950 586.050 184.050 ;
        RECT 586.950 182.100 589.050 187.050 ;
        RECT 593.400 183.600 594.450 187.950 ;
        RECT 596.400 186.450 597.450 229.950 ;
        RECT 605.400 226.050 606.450 254.400 ;
        RECT 610.950 250.950 613.050 255.000 ;
        RECT 617.400 241.050 618.450 268.800 ;
        RECT 634.950 265.950 637.050 268.050 ;
        RECT 635.400 265.200 636.600 265.950 ;
        RECT 622.950 262.950 625.050 265.050 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 620.400 253.050 621.450 259.950 ;
        RECT 623.400 255.450 624.450 262.950 ;
        RECT 630.900 261.900 633.000 263.700 ;
        RECT 634.800 262.800 636.900 264.900 ;
        RECT 638.100 264.300 640.200 266.400 ;
        RECT 629.400 260.700 638.100 261.900 ;
        RECT 626.100 256.950 628.200 259.050 ;
        RECT 626.400 255.450 627.600 256.650 ;
        RECT 623.400 254.400 627.600 255.450 ;
        RECT 619.950 250.950 622.050 253.050 ;
        RECT 629.400 251.700 630.300 260.700 ;
        RECT 636.000 259.800 638.100 260.700 ;
        RECT 639.000 258.900 639.900 264.300 ;
        RECT 641.400 261.450 642.600 261.600 ;
        RECT 644.400 261.450 645.450 277.950 ;
        RECT 646.950 271.950 649.050 274.050 ;
        RECT 641.400 260.400 645.450 261.450 ;
        RECT 641.400 259.350 642.600 260.400 ;
        RECT 633.000 257.700 639.900 258.900 ;
        RECT 633.000 255.300 633.900 257.700 ;
        RECT 631.800 253.200 633.900 255.300 ;
        RECT 634.800 253.950 636.900 256.050 ;
        RECT 628.500 249.600 630.600 251.700 ;
        RECT 635.400 251.400 636.600 253.650 ;
        RECT 638.700 250.500 639.900 257.700 ;
        RECT 640.800 256.950 642.900 259.050 ;
        RECT 643.950 256.950 646.050 259.050 ;
        RECT 638.100 248.400 640.200 250.500 ;
        RECT 616.950 238.950 619.050 241.050 ;
        RECT 625.950 238.950 628.050 241.050 ;
        RECT 619.950 232.950 622.050 235.050 ;
        RECT 610.950 229.950 613.050 232.050 ;
        RECT 604.950 223.950 607.050 226.050 ;
        RECT 598.950 214.950 601.050 217.050 ;
        RECT 604.950 215.100 607.050 217.200 ;
        RECT 611.400 216.600 612.450 229.950 ;
        RECT 599.400 208.050 600.450 214.950 ;
        RECT 605.400 214.350 606.600 215.100 ;
        RECT 611.400 214.350 612.600 216.600 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 608.400 210.000 609.600 211.650 ;
        RECT 598.950 207.450 601.050 208.050 ;
        RECT 598.950 206.400 603.450 207.450 ;
        RECT 598.950 205.950 601.050 206.400 ;
        RECT 598.950 186.450 601.050 190.050 ;
        RECT 596.400 185.400 601.050 186.450 ;
        RECT 587.400 181.350 588.600 182.100 ;
        RECT 593.400 181.350 594.600 183.600 ;
        RECT 598.950 181.950 601.050 185.400 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 565.950 175.800 568.050 177.900 ;
        RECT 571.950 175.800 574.050 177.900 ;
        RECT 580.950 175.800 583.050 177.900 ;
        RECT 583.950 175.950 586.050 178.050 ;
        RECT 590.400 177.900 591.600 178.650 ;
        RECT 596.400 177.900 597.600 178.650 ;
        RECT 602.400 177.900 603.450 206.400 ;
        RECT 604.950 205.950 607.050 208.050 ;
        RECT 607.950 207.450 610.050 210.000 ;
        RECT 614.400 209.400 615.600 211.650 ;
        RECT 607.950 206.400 612.450 207.450 ;
        RECT 607.950 205.950 610.050 206.400 ;
        RECT 605.400 184.050 606.450 205.950 ;
        RECT 604.950 181.950 607.050 184.050 ;
        RECT 611.400 183.600 612.450 206.400 ;
        RECT 614.400 205.050 615.450 209.400 ;
        RECT 613.950 202.950 616.050 205.050 ;
        RECT 620.400 196.050 621.450 232.950 ;
        RECT 622.950 215.100 625.050 217.200 ;
        RECT 626.400 217.050 627.450 238.950 ;
        RECT 644.400 235.050 645.450 256.950 ;
        RECT 647.400 255.900 648.450 271.950 ;
        RECT 650.400 262.050 651.450 293.100 ;
        RECT 656.400 292.350 657.600 294.600 ;
        RECT 665.400 292.350 666.600 294.600 ;
        RECT 682.950 293.100 685.050 295.200 ;
        RECT 683.400 292.350 684.600 293.100 ;
        RECT 656.100 289.950 658.200 292.050 ;
        RECT 659.400 289.950 661.500 292.050 ;
        RECT 664.800 289.950 666.900 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 659.400 287.400 660.600 289.650 ;
        RECT 680.400 288.900 681.600 289.650 ;
        RECT 659.400 280.050 660.450 287.400 ;
        RECT 679.950 286.800 682.050 288.900 ;
        RECT 686.400 288.000 687.600 289.650 ;
        RECT 685.950 283.950 688.050 288.000 ;
        RECT 692.400 286.050 693.450 304.950 ;
        RECT 701.400 304.050 702.450 307.950 ;
        RECT 700.950 301.950 703.050 304.050 ;
        RECT 730.950 301.950 733.050 304.050 ;
        RECT 701.400 294.600 702.450 301.950 ;
        RECT 701.400 292.350 702.600 294.600 ;
        RECT 706.950 294.000 709.050 298.050 ;
        RECT 712.950 295.950 715.050 298.050 ;
        RECT 707.400 292.350 708.600 294.000 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 704.400 287.400 705.600 289.650 ;
        RECT 713.400 288.900 714.450 295.950 ;
        RECT 731.400 294.600 732.450 301.950 ;
        RECT 746.400 294.600 747.450 310.950 ;
        RECT 755.400 298.050 756.450 310.950 ;
        RECT 757.950 304.950 760.050 307.050 ;
        RECT 754.950 295.950 757.050 298.050 ;
        RECT 722.400 294.450 723.600 294.600 ;
        RECT 719.400 293.400 723.600 294.450 ;
        RECT 691.950 283.950 694.050 286.050 ;
        RECT 658.950 277.950 661.050 280.050 ;
        RECT 664.950 262.950 667.050 268.050 ;
        RECT 692.400 265.050 693.450 283.950 ;
        RECT 667.950 262.950 670.050 265.050 ;
        RECT 649.950 259.950 652.050 262.050 ;
        RECT 655.950 260.100 658.050 262.200 ;
        RECT 656.400 259.350 657.600 260.100 ;
        RECT 664.950 259.800 667.050 261.900 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 653.400 255.900 654.600 256.650 ;
        RECT 646.950 253.800 649.050 255.900 ;
        RECT 652.950 253.800 655.050 255.900 ;
        RECT 659.400 255.000 660.600 256.650 ;
        RECT 643.950 232.950 646.050 235.050 ;
        RECT 640.950 223.950 643.050 226.050 ;
        RECT 634.950 219.450 637.050 220.050 ;
        RECT 634.950 219.000 639.450 219.450 ;
        RECT 634.950 218.400 640.050 219.000 ;
        RECT 623.400 205.050 624.450 215.100 ;
        RECT 625.950 214.950 628.050 217.050 ;
        RECT 628.950 215.100 631.050 217.200 ;
        RECT 634.950 216.000 637.050 218.400 ;
        RECT 629.400 214.350 630.600 215.100 ;
        RECT 635.400 214.350 636.600 216.000 ;
        RECT 637.950 214.950 640.050 218.400 ;
        RECT 628.950 211.950 631.050 214.050 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 625.950 205.950 628.050 211.050 ;
        RECT 632.400 210.900 633.600 211.650 ;
        RECT 631.950 208.800 634.050 210.900 ;
        RECT 622.950 202.950 625.050 205.050 ;
        RECT 619.950 193.950 622.050 196.050 ;
        RECT 625.950 187.950 628.050 190.050 ;
        RECT 626.400 184.050 627.450 187.950 ;
        RECT 611.400 181.350 612.600 183.600 ;
        RECT 617.400 183.450 618.600 183.600 ;
        RECT 617.400 182.400 624.450 183.450 ;
        RECT 617.400 181.350 618.600 182.400 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 608.400 177.900 609.600 178.650 ;
        RECT 559.950 142.950 562.050 145.050 ;
        RECT 548.400 136.350 549.600 138.000 ;
        RECT 553.950 137.100 556.050 139.200 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 574.950 137.100 577.050 139.200 ;
        RECT 584.400 139.050 585.450 175.950 ;
        RECT 589.950 175.800 592.050 177.900 ;
        RECT 595.950 175.800 598.050 177.900 ;
        RECT 601.950 175.800 604.050 177.900 ;
        RECT 607.950 175.800 610.050 177.900 ;
        RECT 614.400 177.000 615.600 178.650 ;
        RECT 613.950 172.950 616.050 177.000 ;
        RECT 589.950 148.950 592.050 151.050 ;
        RECT 586.950 142.950 589.050 145.050 ;
        RECT 581.400 138.450 582.600 138.600 ;
        RECT 583.950 138.450 586.050 139.050 ;
        RECT 581.400 137.400 586.050 138.450 ;
        RECT 554.400 136.350 555.600 137.100 ;
        RECT 569.400 136.350 570.600 137.100 ;
        RECT 575.400 136.350 576.600 137.100 ;
        RECT 581.400 136.350 582.600 137.400 ;
        RECT 583.950 136.950 586.050 137.400 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 545.400 132.900 546.600 133.650 ;
        RECT 544.950 130.800 547.050 132.900 ;
        RECT 551.400 131.400 552.600 133.650 ;
        RECT 572.400 131.400 573.600 133.650 ;
        RECT 578.400 132.900 579.600 133.650 ;
        RECT 551.400 127.050 552.450 131.400 ;
        RECT 568.950 127.950 571.050 130.050 ;
        RECT 550.950 124.950 553.050 127.050 ;
        RECT 538.950 112.950 541.050 115.050 ;
        RECT 523.800 111.000 525.900 112.050 ;
        RECT 523.800 109.950 526.050 111.000 ;
        RECT 526.950 109.950 529.050 112.050 ;
        RECT 565.950 109.950 568.050 112.050 ;
        RECT 523.950 108.450 526.050 109.950 ;
        RECT 523.950 108.000 528.450 108.450 ;
        RECT 524.400 107.400 528.450 108.000 ;
        RECT 505.950 104.100 508.050 106.200 ;
        RECT 511.950 104.100 514.050 106.200 ;
        RECT 520.950 104.100 523.050 106.200 ;
        RECT 527.400 105.600 528.450 107.400 ;
        RECT 506.400 103.350 507.600 104.100 ;
        RECT 512.400 103.350 513.600 104.100 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 509.400 99.900 510.600 100.650 ;
        RECT 508.950 97.800 511.050 99.900 ;
        RECT 515.400 98.400 516.600 100.650 ;
        RECT 509.400 79.050 510.450 97.800 ;
        RECT 515.400 94.050 516.450 98.400 ;
        RECT 521.400 96.450 522.450 104.100 ;
        RECT 527.400 103.350 528.600 105.600 ;
        RECT 532.950 104.100 535.050 106.200 ;
        RECT 533.400 103.350 534.600 104.100 ;
        RECT 544.950 103.950 547.050 106.050 ;
        RECT 550.950 104.100 553.050 106.200 ;
        RECT 556.950 105.000 559.050 109.050 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 530.400 99.900 531.600 100.650 ;
        RECT 529.950 97.800 532.050 99.900 ;
        RECT 536.400 98.400 537.600 100.650 ;
        RECT 521.400 95.400 525.450 96.450 ;
        RECT 514.950 91.950 517.050 94.050 ;
        RECT 520.950 82.950 523.050 85.050 ;
        RECT 508.950 76.950 511.050 79.050 ;
        RECT 508.950 59.100 511.050 61.200 ;
        RECT 514.950 59.100 517.050 61.200 ;
        RECT 509.400 58.350 510.600 59.100 ;
        RECT 515.400 58.350 516.600 59.100 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 506.400 53.400 507.600 55.650 ;
        RECT 512.400 54.900 513.600 55.650 ;
        RECT 521.400 55.050 522.450 82.950 ;
        RECT 524.400 76.050 525.450 95.400 ;
        RECT 530.400 93.450 531.450 97.800 ;
        RECT 530.400 92.400 534.450 93.450 ;
        RECT 529.950 88.950 532.050 91.050 ;
        RECT 523.950 73.950 526.050 76.050 ;
        RECT 506.400 43.050 507.450 53.400 ;
        RECT 511.950 52.800 514.050 54.900 ;
        RECT 520.950 52.950 523.050 55.050 ;
        RECT 524.400 52.050 525.450 73.950 ;
        RECT 530.400 61.200 531.450 88.950 ;
        RECT 533.400 76.050 534.450 92.400 ;
        RECT 536.400 91.050 537.450 98.400 ;
        RECT 535.950 88.950 538.050 91.050 ;
        RECT 545.400 84.450 546.450 103.950 ;
        RECT 551.400 103.350 552.600 104.100 ;
        RECT 557.400 103.350 558.600 105.000 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 554.400 99.900 555.600 100.650 ;
        RECT 560.400 99.900 561.600 100.650 ;
        RECT 566.400 99.900 567.450 109.950 ;
        RECT 569.400 99.900 570.450 127.950 ;
        RECT 572.400 109.050 573.450 131.400 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 583.950 130.950 586.050 133.050 ;
        RECT 587.400 132.900 588.450 142.950 ;
        RECT 584.400 124.050 585.450 130.950 ;
        RECT 586.950 130.800 589.050 132.900 ;
        RECT 583.950 121.950 586.050 124.050 ;
        RECT 571.950 106.950 574.050 109.050 ;
        RECT 577.950 105.000 580.050 109.050 ;
        RECT 590.400 106.200 591.450 148.950 ;
        RECT 595.950 142.950 598.050 145.050 ;
        RECT 596.400 138.600 597.450 142.950 ;
        RECT 623.400 142.050 624.450 182.400 ;
        RECT 625.950 181.950 628.050 184.050 ;
        RECT 628.950 183.000 631.050 187.050 ;
        RECT 634.950 183.000 637.050 187.050 ;
        RECT 641.400 184.050 642.450 223.950 ;
        RECT 647.400 220.050 648.450 253.800 ;
        RECT 658.950 250.950 661.050 255.000 ;
        RECT 665.400 226.050 666.450 259.800 ;
        RECT 668.400 253.050 669.450 262.950 ;
        RECT 673.950 260.100 676.050 265.050 ;
        RECT 679.950 261.000 682.050 265.050 ;
        RECT 685.950 262.950 688.050 265.050 ;
        RECT 691.950 262.950 694.050 265.050 ;
        RECT 674.400 259.350 675.600 260.100 ;
        RECT 680.400 259.350 681.600 261.000 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 670.950 253.950 673.050 256.050 ;
        RECT 677.400 255.000 678.600 256.650 ;
        RECT 667.950 250.950 670.050 253.050 ;
        RECT 664.950 223.950 667.050 226.050 ;
        RECT 646.950 217.950 649.050 220.050 ;
        RECT 649.950 215.100 652.050 217.200 ;
        RECT 650.400 214.350 651.600 215.100 ;
        RECT 658.950 214.950 661.050 217.050 ;
        RECT 664.950 215.100 667.050 217.200 ;
        RECT 671.400 216.600 672.450 253.950 ;
        RECT 676.950 250.950 679.050 255.000 ;
        RECT 686.400 253.050 687.450 262.950 ;
        RECT 704.400 262.200 705.450 287.400 ;
        RECT 712.950 286.800 715.050 288.900 ;
        RECT 719.400 277.050 720.450 293.400 ;
        RECT 722.400 292.350 723.600 293.400 ;
        RECT 731.400 294.450 732.600 294.600 ;
        RECT 731.400 293.400 735.450 294.450 ;
        RECT 731.400 292.350 732.600 293.400 ;
        RECT 722.100 289.950 724.200 292.050 ;
        RECT 725.400 289.950 727.500 292.050 ;
        RECT 730.800 289.950 732.900 292.050 ;
        RECT 725.400 288.900 726.600 289.650 ;
        RECT 724.950 286.800 727.050 288.900 ;
        RECT 718.950 274.950 721.050 277.050 ;
        RECT 718.950 268.950 721.050 271.050 ;
        RECT 706.950 262.950 709.050 265.050 ;
        RECT 694.950 260.100 697.050 262.200 ;
        RECT 703.950 260.100 706.050 262.200 ;
        RECT 695.400 259.350 696.600 260.100 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 692.400 255.000 693.600 256.650 ;
        RECT 698.400 255.900 699.600 256.650 ;
        RECT 685.950 250.950 688.050 253.050 ;
        RECT 691.950 250.950 694.050 255.000 ;
        RECT 697.950 253.800 700.050 255.900 ;
        RECT 676.950 241.950 679.050 244.050 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 649.950 211.950 652.050 214.050 ;
        RECT 652.950 211.950 655.050 214.050 ;
        RECT 643.950 205.950 646.050 210.900 ;
        RECT 647.400 209.400 648.600 211.650 ;
        RECT 653.400 210.900 654.600 211.650 ;
        RECT 647.400 205.050 648.450 209.400 ;
        RECT 652.950 208.800 655.050 210.900 ;
        RECT 646.950 202.950 649.050 205.050 ;
        RECT 659.400 199.050 660.450 214.950 ;
        RECT 665.400 214.350 666.600 215.100 ;
        RECT 671.400 214.350 672.600 216.600 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 670.950 211.950 673.050 214.050 ;
        RECT 668.400 210.900 669.600 211.650 ;
        RECT 667.950 208.800 670.050 210.900 ;
        RECT 661.950 199.950 664.050 202.050 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 658.950 196.950 661.050 199.050 ;
        RECT 643.950 184.950 646.050 187.050 ;
        RECT 629.400 181.350 630.600 183.000 ;
        RECT 635.400 181.350 636.600 183.000 ;
        RECT 640.950 181.950 643.050 184.050 ;
        RECT 628.950 178.950 631.050 181.050 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 632.400 177.900 633.600 178.650 ;
        RECT 638.400 177.900 639.600 178.650 ;
        RECT 631.950 175.800 634.050 177.900 ;
        RECT 637.950 175.800 640.050 177.900 ;
        RECT 644.400 151.050 645.450 184.950 ;
        RECT 647.400 169.050 648.450 196.950 ;
        RECT 652.950 190.950 655.050 193.050 ;
        RECT 653.400 183.600 654.450 190.950 ;
        RECT 653.400 181.350 654.600 183.600 ;
        RECT 659.400 183.450 660.600 183.600 ;
        RECT 662.400 183.450 663.450 199.950 ;
        RECT 677.400 187.050 678.450 241.950 ;
        RECT 682.950 223.950 685.050 226.050 ;
        RECT 679.950 215.100 682.050 217.200 ;
        RECT 683.400 217.050 684.450 223.950 ;
        RECT 704.400 220.050 705.450 260.100 ;
        RECT 680.400 211.050 681.450 215.100 ;
        RECT 682.950 214.950 685.050 217.050 ;
        RECT 685.950 215.100 688.050 217.200 ;
        RECT 691.950 216.000 694.050 220.050 ;
        RECT 686.400 214.350 687.600 215.100 ;
        RECT 692.400 214.350 693.600 216.000 ;
        RECT 697.950 214.950 700.050 220.050 ;
        RECT 703.950 217.950 706.050 220.050 ;
        RECT 700.950 214.950 703.050 217.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 694.950 211.950 697.050 214.050 ;
        RECT 679.950 208.950 682.050 211.050 ;
        RECT 689.400 210.000 690.600 211.650 ;
        RECT 688.950 205.950 691.050 210.000 ;
        RECT 695.400 209.400 696.600 211.650 ;
        RECT 685.950 199.950 688.050 202.050 ;
        RECT 670.950 184.950 673.050 187.050 ;
        RECT 676.950 184.950 679.050 187.050 ;
        RECT 659.400 182.400 663.450 183.450 ;
        RECT 659.400 181.350 660.600 182.400 ;
        RECT 667.950 182.100 670.050 184.200 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 656.400 177.900 657.600 178.650 ;
        RECT 668.400 178.050 669.450 182.100 ;
        RECT 655.950 175.800 658.050 177.900 ;
        RECT 667.950 175.950 670.050 178.050 ;
        RECT 646.950 166.950 649.050 169.050 ;
        RECT 671.400 151.050 672.450 184.950 ;
        RECT 679.950 182.100 682.050 184.200 ;
        RECT 680.400 181.350 681.600 182.100 ;
        RECT 674.100 178.950 676.200 181.050 ;
        RECT 679.500 178.950 681.600 181.050 ;
        RECT 682.800 178.950 684.900 181.050 ;
        RECT 674.400 176.400 675.600 178.650 ;
        RECT 683.400 177.900 684.600 178.650 ;
        RECT 674.400 163.050 675.450 176.400 ;
        RECT 682.950 175.800 685.050 177.900 ;
        RECT 683.400 169.050 684.450 175.800 ;
        RECT 682.950 166.950 685.050 169.050 ;
        RECT 673.950 160.950 676.050 163.050 ;
        RECT 686.400 157.050 687.450 199.950 ;
        RECT 695.400 193.050 696.450 209.400 ;
        RECT 701.400 202.050 702.450 214.950 ;
        RECT 704.400 210.900 705.450 217.950 ;
        RECT 707.400 217.050 708.450 262.950 ;
        RECT 712.950 260.100 715.050 262.200 ;
        RECT 719.400 261.600 720.450 268.950 ;
        RECT 725.400 265.050 726.450 286.800 ;
        RECT 727.950 274.950 730.050 277.050 ;
        RECT 724.950 262.950 727.050 265.050 ;
        RECT 713.400 259.350 714.600 260.100 ;
        RECT 719.400 259.350 720.600 261.600 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 716.400 255.000 717.600 256.650 ;
        RECT 722.400 256.050 723.600 256.650 ;
        RECT 715.950 250.950 718.050 255.000 ;
        RECT 722.400 254.400 727.050 256.050 ;
        RECT 723.000 253.950 727.050 254.400 ;
        RECT 725.400 250.050 726.450 253.950 ;
        RECT 724.950 247.950 727.050 250.050 ;
        RECT 709.950 223.950 712.050 226.050 ;
        RECT 706.950 214.950 709.050 217.050 ;
        RECT 710.400 216.600 711.450 223.950 ;
        RECT 725.400 220.050 726.450 247.950 ;
        RECT 710.400 214.350 711.600 216.600 ;
        RECT 715.950 216.000 718.050 220.050 ;
        RECT 724.950 217.950 727.050 220.050 ;
        RECT 728.400 217.200 729.450 274.950 ;
        RECT 734.400 265.050 735.450 293.400 ;
        RECT 746.400 292.350 747.600 294.600 ;
        RECT 751.950 293.100 754.050 295.200 ;
        RECT 752.400 292.350 753.600 293.100 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 748.950 289.950 751.050 292.050 ;
        RECT 751.950 289.950 754.050 292.050 ;
        RECT 749.400 288.900 750.600 289.650 ;
        RECT 758.400 289.050 759.450 304.950 ;
        RECT 760.950 298.950 763.050 301.050 ;
        RECT 748.950 286.800 751.050 288.900 ;
        RECT 757.950 286.950 760.050 289.050 ;
        RECT 751.950 268.950 754.050 271.050 ;
        RECT 733.950 262.950 736.050 265.050 ;
        RECT 736.950 261.000 739.050 265.050 ;
        RECT 737.400 259.350 738.600 261.000 ;
        RECT 742.950 260.100 745.050 262.200 ;
        RECT 743.400 259.350 744.600 260.100 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 736.950 256.950 739.050 259.050 ;
        RECT 739.950 256.950 742.050 259.050 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 745.950 256.950 748.050 259.050 ;
        RECT 734.400 255.900 735.600 256.650 ;
        RECT 733.950 253.800 736.050 255.900 ;
        RECT 740.400 254.400 741.600 256.650 ;
        RECT 746.400 254.400 747.600 256.650 ;
        RECT 740.400 220.050 741.450 254.400 ;
        RECT 746.400 241.050 747.450 254.400 ;
        RECT 752.400 253.050 753.450 268.950 ;
        RECT 761.400 265.050 762.450 298.950 ;
        RECT 766.800 298.200 768.900 300.300 ;
        RECT 775.800 298.500 777.900 300.600 ;
        RECT 763.950 293.100 766.050 295.200 ;
        RECT 764.400 292.350 765.600 293.100 ;
        RECT 764.100 289.950 766.200 292.050 ;
        RECT 767.100 285.600 768.000 298.200 ;
        RECT 773.400 295.350 774.600 297.600 ;
        RECT 773.100 292.950 775.200 295.050 ;
        RECT 768.900 291.900 771.000 292.200 ;
        RECT 777.000 291.900 777.900 298.500 ;
        RECT 781.950 293.100 784.050 295.200 ;
        RECT 788.400 294.450 789.450 331.950 ;
        RECT 790.950 331.800 793.050 333.900 ;
        RECT 796.950 331.800 799.050 333.900 ;
        RECT 802.950 331.800 805.050 333.900 ;
        RECT 808.950 333.450 811.050 333.900 ;
        RECT 812.400 333.450 813.450 361.950 ;
        RECT 815.400 355.050 816.450 365.400 ;
        RECT 817.950 358.950 820.050 361.050 ;
        RECT 814.950 352.950 817.050 355.050 ;
        RECT 818.400 349.050 819.450 358.950 ;
        RECT 824.400 352.050 825.450 407.400 ;
        RECT 833.400 406.050 834.450 410.400 ;
        RECT 832.950 403.950 835.050 406.050 ;
        RECT 839.400 397.050 840.450 433.950 ;
        RECT 842.400 427.050 843.450 439.950 ;
        RECT 841.950 424.950 844.050 427.050 ;
        RECT 848.400 417.600 849.450 442.950 ;
        RECT 856.950 439.950 859.050 444.000 ;
        RECT 862.950 442.950 865.050 445.050 ;
        RECT 856.950 424.950 859.050 427.050 ;
        RECT 848.400 415.350 849.600 417.600 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 845.400 411.450 846.600 412.650 ;
        RECT 851.400 411.900 852.600 412.650 ;
        RECT 842.400 410.400 846.600 411.450 ;
        RECT 842.400 400.050 843.450 410.400 ;
        RECT 850.950 409.800 853.050 411.900 ;
        RECT 844.950 403.950 847.050 406.050 ;
        RECT 841.950 397.950 844.050 400.050 ;
        RECT 838.950 394.950 841.050 397.050 ;
        RECT 832.950 376.950 835.050 379.050 ;
        RECT 833.400 372.600 834.450 376.950 ;
        RECT 833.400 370.350 834.600 372.600 ;
        RECT 838.950 372.000 841.050 376.050 ;
        RECT 842.400 373.050 843.450 397.950 ;
        RECT 839.400 370.350 840.600 372.000 ;
        RECT 841.950 370.950 844.050 373.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 835.950 367.950 838.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 830.400 365.400 831.600 367.650 ;
        RECT 836.400 365.400 837.600 367.650 ;
        RECT 830.400 361.050 831.450 365.400 ;
        RECT 829.950 358.950 832.050 361.050 ;
        RECT 836.400 360.450 837.450 365.400 ;
        RECT 841.950 364.950 844.050 367.050 ;
        RECT 836.400 359.400 840.450 360.450 ;
        RECT 835.950 355.950 838.050 358.050 ;
        RECT 823.950 349.950 826.050 352.050 ;
        RECT 817.950 346.950 820.050 349.050 ;
        RECT 821.400 347.400 828.450 348.450 ;
        RECT 821.400 343.050 822.450 347.400 ;
        RECT 823.950 343.950 826.050 346.050 ;
        RECT 814.950 340.950 817.050 343.050 ;
        RECT 820.950 340.950 823.050 343.050 ;
        RECT 808.950 332.400 813.450 333.450 ;
        RECT 808.950 328.950 811.050 332.400 ;
        RECT 805.950 310.950 808.050 313.050 ;
        RECT 790.950 304.950 793.050 307.050 ;
        RECT 785.400 293.400 789.450 294.450 ;
        RECT 791.400 294.600 792.450 304.950 ;
        RECT 768.900 291.000 777.900 291.900 ;
        RECT 768.900 290.100 771.000 291.000 ;
        RECT 774.000 289.200 776.100 290.100 ;
        RECT 768.900 288.000 776.100 289.200 ;
        RECT 768.900 287.100 771.000 288.000 ;
        RECT 766.500 283.500 768.600 285.600 ;
        RECT 773.100 284.100 775.200 286.200 ;
        RECT 777.000 285.900 777.900 291.000 ;
        RECT 778.800 289.950 780.900 292.050 ;
        RECT 779.400 288.900 780.600 289.650 ;
        RECT 778.950 286.800 781.050 288.900 ;
        RECT 776.400 283.800 778.500 285.900 ;
        RECT 773.400 282.000 774.600 283.800 ;
        RECT 772.950 277.950 775.050 282.000 ;
        RECT 782.400 280.050 783.450 293.100 ;
        RECT 781.950 277.950 784.050 280.050 ;
        RECT 785.400 268.050 786.450 293.400 ;
        RECT 791.400 292.350 792.600 294.600 ;
        RECT 796.950 293.100 799.050 295.200 ;
        RECT 797.400 292.350 798.600 293.100 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 794.400 287.400 795.600 289.650 ;
        RECT 800.400 288.900 801.600 289.650 ;
        RECT 794.400 277.050 795.450 287.400 ;
        RECT 799.950 286.800 802.050 288.900 ;
        RECT 802.950 286.950 805.050 289.050 ;
        RECT 800.400 283.050 801.450 286.800 ;
        RECT 799.950 280.950 802.050 283.050 ;
        RECT 793.950 274.950 796.050 277.050 ;
        RECT 784.950 265.950 787.050 268.050 ;
        RECT 793.950 265.950 796.050 268.050 ;
        RECT 760.950 262.950 763.050 265.050 ;
        RECT 772.950 262.950 775.050 265.050 ;
        RECT 761.400 261.600 762.450 262.950 ;
        RECT 761.400 259.350 762.600 261.600 ;
        RECT 766.950 260.100 769.050 262.200 ;
        RECT 767.400 259.350 768.600 260.100 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 758.400 254.400 759.600 256.650 ;
        RECT 764.400 255.000 765.600 256.650 ;
        RECT 751.950 250.950 754.050 253.050 ;
        RECT 745.950 238.950 748.050 241.050 ;
        RECT 716.400 214.350 717.600 216.000 ;
        RECT 727.950 215.100 730.050 217.200 ;
        RECT 730.950 216.000 733.050 220.050 ;
        RECT 739.950 217.950 742.050 220.050 ;
        RECT 731.400 214.350 732.600 216.000 ;
        RECT 736.950 215.100 739.050 217.200 ;
        RECT 737.400 214.350 738.600 215.100 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 715.950 211.950 718.050 214.050 ;
        RECT 718.950 211.950 721.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 713.400 210.900 714.600 211.650 ;
        RECT 703.950 208.800 706.050 210.900 ;
        RECT 712.950 208.800 715.050 210.900 ;
        RECT 719.400 209.400 720.600 211.650 ;
        RECT 734.400 209.400 735.600 211.650 ;
        RECT 740.400 209.400 741.600 211.650 ;
        RECT 746.400 210.900 747.450 238.950 ;
        RECT 758.400 238.050 759.450 254.400 ;
        RECT 763.950 250.950 766.050 255.000 ;
        RECT 764.400 244.050 765.450 250.950 ;
        RECT 763.950 241.950 766.050 244.050 ;
        RECT 757.950 235.950 760.050 238.050 ;
        RECT 773.400 226.050 774.450 262.950 ;
        RECT 781.950 261.000 784.050 265.050 ;
        RECT 782.400 259.350 783.600 261.000 ;
        RECT 787.950 260.100 790.050 262.200 ;
        RECT 788.400 259.350 789.600 260.100 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 779.400 254.400 780.600 256.650 ;
        RECT 785.400 254.400 786.600 256.650 ;
        RECT 779.400 238.050 780.450 254.400 ;
        RECT 785.400 244.050 786.450 254.400 ;
        RECT 784.950 241.950 787.050 244.050 ;
        RECT 778.950 235.950 781.050 238.050 ;
        RECT 772.950 223.950 775.050 226.050 ;
        RECT 748.950 217.950 751.050 220.050 ;
        RECT 700.950 199.950 703.050 202.050 ;
        RECT 694.950 190.950 697.050 193.050 ;
        RECT 691.950 187.950 694.050 190.050 ;
        RECT 688.950 184.950 691.050 187.050 ;
        RECT 689.400 172.050 690.450 184.950 ;
        RECT 692.400 178.050 693.450 187.950 ;
        RECT 697.950 183.000 700.050 187.050 ;
        RECT 701.400 186.450 702.450 199.950 ;
        RECT 719.400 196.050 720.450 209.400 ;
        RECT 734.400 208.050 735.450 209.400 ;
        RECT 734.400 206.400 739.050 208.050 ;
        RECT 735.000 205.950 739.050 206.400 ;
        RECT 712.950 193.950 715.050 196.050 ;
        RECT 718.950 193.950 721.050 196.050 ;
        RECT 701.400 185.400 705.450 186.450 ;
        RECT 704.400 183.600 705.450 185.400 ;
        RECT 698.400 181.350 699.600 183.000 ;
        RECT 704.400 181.350 705.600 183.600 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 691.950 175.950 694.050 178.050 ;
        RECT 701.400 176.400 702.600 178.650 ;
        RECT 688.950 169.950 691.050 172.050 ;
        RECT 694.950 169.950 697.050 172.050 ;
        RECT 685.950 154.950 688.050 157.050 ;
        RECT 625.950 148.950 628.050 151.050 ;
        RECT 643.950 148.950 646.050 151.050 ;
        RECT 670.950 148.950 673.050 151.050 ;
        RECT 596.400 136.350 597.600 138.600 ;
        RECT 601.950 138.000 604.050 142.050 ;
        RECT 622.950 139.950 625.050 142.050 ;
        RECT 602.400 136.350 603.600 138.000 ;
        RECT 613.950 137.100 616.050 139.200 ;
        RECT 619.950 137.100 622.050 139.200 ;
        RECT 626.400 138.600 627.450 148.950 ;
        RECT 637.950 139.950 640.050 142.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 592.950 130.950 595.050 133.050 ;
        RECT 599.400 132.900 600.600 133.650 ;
        RECT 593.400 112.050 594.450 130.950 ;
        RECT 598.950 130.800 601.050 132.900 ;
        RECT 605.400 131.400 606.600 133.650 ;
        RECT 595.950 112.950 598.050 115.050 ;
        RECT 592.950 109.950 595.050 112.050 ;
        RECT 596.400 108.450 597.450 112.950 ;
        RECT 593.400 107.400 597.450 108.450 ;
        RECT 605.400 108.450 606.450 131.400 ;
        RECT 614.400 127.050 615.450 137.100 ;
        RECT 620.400 136.350 621.600 137.100 ;
        RECT 626.400 136.350 627.600 138.600 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 623.400 132.900 624.600 133.650 ;
        RECT 622.950 130.800 625.050 132.900 ;
        RECT 629.400 131.400 630.600 133.650 ;
        RECT 638.400 132.900 639.450 139.950 ;
        RECT 644.400 138.600 645.450 148.950 ;
        RECT 644.400 136.350 645.600 138.600 ;
        RECT 649.950 137.100 652.050 139.200 ;
        RECT 658.950 137.100 661.050 139.200 ;
        RECT 667.950 137.100 670.050 139.200 ;
        RECT 673.950 137.100 676.050 139.200 ;
        RECT 686.400 138.450 687.450 154.950 ;
        RECT 688.950 145.950 691.050 148.050 ;
        RECT 683.400 137.400 687.450 138.450 ;
        RECT 689.400 138.600 690.450 145.950 ;
        RECT 695.400 139.200 696.450 169.950 ;
        RECT 701.400 160.050 702.450 176.400 ;
        RECT 700.950 157.950 703.050 160.050 ;
        RECT 713.400 151.050 714.450 193.950 ;
        RECT 740.400 190.050 741.450 209.400 ;
        RECT 745.950 208.800 748.050 210.900 ;
        RECT 749.400 199.050 750.450 217.950 ;
        RECT 754.950 215.100 757.050 217.200 ;
        RECT 760.950 216.000 763.050 220.050 ;
        RECT 772.950 217.950 775.050 220.050 ;
        RECT 755.400 214.350 756.600 215.100 ;
        RECT 761.400 214.350 762.600 216.000 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 758.400 210.900 759.600 211.650 ;
        RECT 757.950 208.800 760.050 210.900 ;
        RECT 764.400 209.400 765.600 211.650 ;
        RECT 764.400 205.050 765.450 209.400 ;
        RECT 763.950 202.950 766.050 205.050 ;
        RECT 748.950 196.950 751.050 199.050 ;
        RECT 754.950 190.950 757.050 193.050 ;
        RECT 718.950 187.950 721.050 190.050 ;
        RECT 739.950 187.950 742.050 190.050 ;
        RECT 719.400 184.200 720.450 187.950 ;
        RECT 718.950 182.100 721.050 184.200 ;
        RECT 724.950 183.000 727.050 187.050 ;
        RECT 741.000 186.450 745.050 187.050 ;
        RECT 740.400 184.950 745.050 186.450 ;
        RECT 748.950 184.950 751.050 187.050 ;
        RECT 751.950 184.950 754.050 187.050 ;
        RECT 719.400 181.350 720.600 182.100 ;
        RECT 725.400 181.350 726.600 183.000 ;
        RECT 730.950 181.950 733.050 184.050 ;
        RECT 740.400 183.600 741.450 184.950 ;
        RECT 718.950 178.950 721.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 722.400 176.400 723.600 178.650 ;
        RECT 731.400 177.900 732.450 181.950 ;
        RECT 740.400 181.350 741.600 183.600 ;
        RECT 736.950 178.950 739.050 181.050 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 737.400 177.900 738.600 178.650 ;
        RECT 743.400 177.900 744.600 178.650 ;
        RECT 722.400 175.050 723.450 176.400 ;
        RECT 730.950 175.800 733.050 177.900 ;
        RECT 736.950 175.800 739.050 177.900 ;
        RECT 742.950 175.800 745.050 177.900 ;
        RECT 745.950 175.950 748.050 178.050 ;
        RECT 749.400 177.900 750.450 184.950 ;
        RECT 752.400 178.050 753.450 184.950 ;
        RECT 755.400 178.050 756.450 190.950 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 763.950 182.100 766.050 184.200 ;
        RECT 764.400 181.350 765.600 182.100 ;
        RECT 758.100 178.950 760.200 181.050 ;
        RECT 763.500 178.950 765.600 181.050 ;
        RECT 766.800 178.950 768.900 181.050 ;
        RECT 722.400 173.400 727.050 175.050 ;
        RECT 723.000 172.950 727.050 173.400 ;
        RECT 731.400 172.050 732.450 175.800 ;
        RECT 730.950 169.950 733.050 172.050 ;
        RECT 736.950 171.450 739.050 174.750 ;
        RECT 742.950 171.450 745.050 172.050 ;
        RECT 736.950 171.000 745.050 171.450 ;
        RECT 737.400 170.400 745.050 171.000 ;
        RECT 742.950 169.950 745.050 170.400 ;
        RECT 742.950 157.950 745.050 160.050 ;
        RECT 703.950 148.950 706.050 151.050 ;
        RECT 712.950 148.950 715.050 151.050 ;
        RECT 650.400 136.350 651.600 137.100 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 647.400 132.900 648.600 133.650 ;
        RECT 629.400 130.050 630.450 131.400 ;
        RECT 637.950 130.800 640.050 132.900 ;
        RECT 646.950 130.800 649.050 132.900 ;
        RECT 653.400 131.400 654.600 133.650 ;
        RECT 629.400 128.400 634.050 130.050 ;
        RECT 630.000 127.950 634.050 128.400 ;
        RECT 613.950 124.950 616.050 127.050 ;
        RECT 628.950 124.950 631.050 127.050 ;
        RECT 610.950 112.950 613.050 115.050 ;
        RECT 605.400 107.400 609.450 108.450 ;
        RECT 578.400 103.350 579.600 105.000 ;
        RECT 583.950 104.100 586.050 106.200 ;
        RECT 589.950 104.100 592.050 106.200 ;
        RECT 584.400 103.350 585.600 104.100 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 575.400 99.900 576.600 100.650 ;
        RECT 553.950 97.800 556.050 99.900 ;
        RECT 559.950 97.800 562.050 99.900 ;
        RECT 565.800 99.000 567.900 99.900 ;
        RECT 565.800 97.800 568.050 99.000 ;
        RECT 568.950 97.800 571.050 99.900 ;
        RECT 574.950 97.800 577.050 99.900 ;
        RECT 581.400 99.000 582.600 100.650 ;
        RECT 565.950 94.950 568.050 97.800 ;
        RECT 580.950 94.950 583.050 99.000 ;
        RECT 586.950 97.950 589.050 100.050 ;
        RECT 593.400 99.450 594.450 107.400 ;
        RECT 601.950 104.100 604.050 106.200 ;
        RECT 602.400 103.350 603.600 104.100 ;
        RECT 596.100 100.950 598.200 103.050 ;
        RECT 601.500 100.950 603.600 103.050 ;
        RECT 604.800 100.950 606.900 103.050 ;
        RECT 596.400 99.450 597.600 100.650 ;
        RECT 593.400 98.400 597.600 99.450 ;
        RECT 605.400 98.400 606.600 100.650 ;
        RECT 550.950 91.950 553.050 94.050 ;
        RECT 545.400 83.400 549.450 84.450 ;
        RECT 544.950 79.950 547.050 82.050 ;
        RECT 532.950 73.950 535.050 76.050 ;
        RECT 535.950 64.950 538.050 67.050 ;
        RECT 529.950 59.100 532.050 61.200 ;
        RECT 536.400 60.600 537.450 64.950 ;
        RECT 530.400 58.350 531.600 59.100 ;
        RECT 536.400 58.350 537.600 60.600 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 526.950 52.950 529.050 55.050 ;
        RECT 533.400 54.000 534.600 55.650 ;
        RECT 539.400 55.050 540.600 55.650 ;
        RECT 545.400 55.050 546.450 79.950 ;
        RECT 523.950 49.950 526.050 52.050 ;
        RECT 505.950 40.950 508.050 43.050 ;
        RECT 517.950 40.950 520.050 43.050 ;
        RECT 518.400 37.050 519.450 40.950 ;
        RECT 517.950 34.950 520.050 37.050 ;
        RECT 497.400 26.400 501.450 27.450 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 482.400 21.900 483.600 22.650 ;
        RECT 488.400 21.900 489.600 22.650 ;
        RECT 497.400 21.900 498.450 26.400 ;
        RECT 505.950 26.100 508.050 28.200 ;
        RECT 511.950 26.100 514.050 28.200 ;
        RECT 506.400 25.350 507.600 26.100 ;
        RECT 512.400 25.350 513.600 26.100 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 487.950 19.800 490.050 21.900 ;
        RECT 472.950 16.950 475.050 19.050 ;
        RECT 496.950 16.950 499.050 21.900 ;
        RECT 503.400 21.000 504.600 22.650 ;
        RECT 509.400 21.000 510.600 22.650 ;
        RECT 502.950 16.950 505.050 21.000 ;
        RECT 508.950 16.950 511.050 21.000 ;
        RECT 518.400 19.050 519.450 34.950 ;
        RECT 527.400 34.050 528.450 52.950 ;
        RECT 532.950 49.950 535.050 54.000 ;
        RECT 539.400 53.400 544.050 55.050 ;
        RECT 540.000 52.950 544.050 53.400 ;
        RECT 544.950 52.950 547.050 55.050 ;
        RECT 548.400 49.050 549.450 83.400 ;
        RECT 551.400 79.050 552.450 91.950 ;
        RECT 587.400 88.050 588.450 97.950 ;
        RECT 605.400 97.050 606.450 98.400 ;
        RECT 604.950 94.950 607.050 97.050 ;
        RECT 556.950 85.950 559.050 88.050 ;
        RECT 586.950 85.950 589.050 88.050 ;
        RECT 550.950 76.950 553.050 79.050 ;
        RECT 550.950 70.950 553.050 73.050 ;
        RECT 551.400 61.050 552.450 70.950 ;
        RECT 557.400 64.050 558.450 85.950 ;
        RECT 592.950 79.950 595.050 82.050 ;
        RECT 565.950 76.950 568.050 79.050 ;
        RECT 556.950 61.950 559.050 64.050 ;
        RECT 550.950 58.950 553.050 61.050 ;
        RECT 553.950 59.100 556.050 61.200 ;
        RECT 562.950 59.100 565.050 61.200 ;
        RECT 554.400 58.350 555.600 59.100 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 557.400 55.050 558.600 55.650 ;
        RECT 557.400 53.400 562.050 55.050 ;
        RECT 558.000 52.950 562.050 53.400 ;
        RECT 547.950 46.950 550.050 49.050 ;
        RECT 559.950 43.950 562.050 46.050 ;
        RECT 560.400 40.050 561.450 43.950 ;
        RECT 563.400 43.050 564.450 59.100 ;
        RECT 566.400 55.050 567.450 76.950 ;
        RECT 580.950 73.950 583.050 76.050 ;
        RECT 574.950 59.100 577.050 61.200 ;
        RECT 581.400 60.600 582.450 73.950 ;
        RECT 589.950 67.950 592.050 70.050 ;
        RECT 575.400 58.350 576.600 59.100 ;
        RECT 581.400 58.350 582.600 60.600 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 580.950 55.950 583.050 58.050 ;
        RECT 565.950 52.800 568.050 55.050 ;
        RECT 572.400 54.900 573.600 55.650 ;
        RECT 578.400 54.900 579.600 55.650 ;
        RECT 590.400 55.050 591.450 67.950 ;
        RECT 593.400 61.200 594.450 79.950 ;
        RECT 605.400 76.050 606.450 94.950 ;
        RECT 608.400 88.050 609.450 107.400 ;
        RECT 611.400 94.050 612.450 112.950 ;
        RECT 619.950 104.100 622.050 106.200 ;
        RECT 620.400 103.350 621.600 104.100 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 617.400 99.900 618.600 100.650 ;
        RECT 616.950 97.800 619.050 99.900 ;
        RECT 623.400 98.400 624.600 100.650 ;
        RECT 623.400 94.050 624.450 98.400 ;
        RECT 629.400 97.050 630.450 124.950 ;
        RECT 637.950 118.950 640.050 121.050 ;
        RECT 638.400 105.600 639.450 118.950 ;
        RECT 643.950 109.950 646.050 112.050 ;
        RECT 644.400 105.600 645.450 109.950 ;
        RECT 649.950 108.450 652.050 109.050 ;
        RECT 653.400 108.450 654.450 131.400 ;
        RECT 655.950 127.950 658.050 133.050 ;
        RECT 659.400 127.050 660.450 137.100 ;
        RECT 668.400 136.350 669.600 137.100 ;
        RECT 674.400 136.350 675.600 137.100 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 658.950 124.950 661.050 127.050 ;
        RECT 662.400 115.050 663.450 133.950 ;
        RECT 671.400 131.400 672.600 133.650 ;
        RECT 677.400 131.400 678.600 133.650 ;
        RECT 683.400 132.900 684.450 137.400 ;
        RECT 689.400 136.350 690.600 138.600 ;
        RECT 694.950 137.100 697.050 139.200 ;
        RECT 695.400 136.350 696.600 137.100 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 667.950 124.950 670.050 130.050 ;
        RECT 671.400 129.450 672.450 131.400 ;
        RECT 671.400 128.400 675.450 129.450 ;
        RECT 661.950 112.950 664.050 115.050 ;
        RECT 667.950 112.950 670.050 115.050 ;
        RECT 655.950 109.950 658.050 112.050 ;
        RECT 649.950 107.400 654.450 108.450 ;
        RECT 649.950 106.950 652.050 107.400 ;
        RECT 638.400 103.350 639.600 105.600 ;
        RECT 644.400 103.350 645.600 105.600 ;
        RECT 650.400 103.050 651.450 106.950 ;
        RECT 656.400 105.450 657.450 109.950 ;
        RECT 653.400 104.400 657.450 105.450 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 635.400 100.050 636.600 100.650 ;
        RECT 631.950 98.400 636.600 100.050 ;
        RECT 641.400 99.900 642.600 100.650 ;
        RECT 631.950 97.950 636.450 98.400 ;
        RECT 628.950 94.950 631.050 97.050 ;
        RECT 635.400 96.300 636.450 97.950 ;
        RECT 640.950 97.800 643.050 99.900 ;
        RECT 646.950 97.950 649.050 100.050 ;
        RECT 640.950 96.300 643.050 96.750 ;
        RECT 635.400 95.250 643.050 96.300 ;
        RECT 640.950 94.650 643.050 95.250 ;
        RECT 610.950 91.950 613.050 94.050 ;
        RECT 622.950 91.950 625.050 94.050 ;
        RECT 607.950 85.950 610.050 88.050 ;
        RECT 598.950 73.950 601.050 76.050 ;
        RECT 604.950 73.950 607.050 76.050 ;
        RECT 592.950 59.100 595.050 61.200 ;
        RECT 599.400 60.600 600.450 73.950 ;
        RECT 599.400 58.350 600.600 60.600 ;
        RECT 604.950 60.000 607.050 64.050 ;
        RECT 608.400 60.450 609.450 85.950 ;
        RECT 610.950 76.950 613.050 79.050 ;
        RECT 611.400 64.050 612.450 76.950 ;
        RECT 619.950 70.950 622.050 73.050 ;
        RECT 640.950 70.950 643.050 73.050 ;
        RECT 610.950 61.950 613.050 64.050 ;
        RECT 620.400 61.200 621.450 70.950 ;
        RECT 605.400 58.350 606.600 60.000 ;
        RECT 608.400 59.400 612.450 60.450 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 604.950 55.950 607.050 58.050 ;
        RECT 571.950 52.800 574.050 54.900 ;
        RECT 577.950 52.800 580.050 54.900 ;
        RECT 589.950 52.950 592.050 55.050 ;
        RECT 596.400 53.400 597.600 55.650 ;
        RECT 602.400 54.900 603.600 55.650 ;
        RECT 611.400 54.900 612.450 59.400 ;
        RECT 619.950 59.100 622.050 61.200 ;
        RECT 625.950 60.000 628.050 64.050 ;
        RECT 631.950 61.950 634.050 64.050 ;
        RECT 620.400 58.350 621.600 59.100 ;
        RECT 626.400 58.350 627.600 60.000 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 596.400 46.050 597.450 53.400 ;
        RECT 601.950 52.800 604.050 54.900 ;
        RECT 610.950 52.800 613.050 54.900 ;
        RECT 617.400 53.400 618.600 55.650 ;
        RECT 623.400 53.400 624.600 55.650 ;
        RECT 632.400 54.900 633.450 61.950 ;
        RECT 641.400 60.600 642.450 70.950 ;
        RECT 647.400 64.050 648.450 97.950 ;
        RECT 653.400 97.050 654.450 104.400 ;
        RECT 661.950 104.100 664.050 106.200 ;
        RECT 668.400 105.600 669.450 112.950 ;
        RECT 662.400 103.350 663.600 104.100 ;
        RECT 668.400 103.350 669.600 105.600 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 659.400 98.400 660.600 100.650 ;
        RECT 665.400 99.900 666.600 100.650 ;
        RECT 652.950 94.950 655.050 97.050 ;
        RECT 659.400 94.050 660.450 98.400 ;
        RECT 664.950 97.800 667.050 99.900 ;
        RECT 670.950 97.950 673.050 100.050 ;
        RECT 658.950 91.950 661.050 94.050 ;
        RECT 671.400 67.050 672.450 97.950 ;
        RECT 674.400 88.050 675.450 128.400 ;
        RECT 677.400 124.050 678.450 131.400 ;
        RECT 682.950 130.800 685.050 132.900 ;
        RECT 692.400 131.400 693.600 133.650 ;
        RECT 698.400 132.900 699.600 133.650 ;
        RECT 688.950 124.950 691.050 127.050 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 676.950 112.950 679.050 115.050 ;
        RECT 673.950 85.950 676.050 88.050 ;
        RECT 649.950 66.450 652.050 67.050 ;
        RECT 649.950 65.400 654.450 66.450 ;
        RECT 649.950 64.950 652.050 65.400 ;
        RECT 646.950 61.950 649.050 64.050 ;
        RECT 641.400 58.350 642.600 60.600 ;
        RECT 647.400 60.450 648.600 60.600 ;
        RECT 650.400 60.450 651.450 64.950 ;
        RECT 647.400 59.400 651.450 60.450 ;
        RECT 647.400 58.350 648.600 59.400 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 565.950 43.950 571.050 46.050 ;
        RECT 595.950 43.950 598.050 46.050 ;
        RECT 562.950 40.950 565.050 43.050 ;
        RECT 617.400 40.050 618.450 53.400 ;
        RECT 623.400 49.050 624.450 53.400 ;
        RECT 631.950 52.800 634.050 54.900 ;
        RECT 638.400 53.400 639.600 55.650 ;
        RECT 644.400 54.900 645.600 55.650 ;
        RECT 622.950 46.950 625.050 49.050 ;
        RECT 559.950 37.950 562.050 40.050 ;
        RECT 574.950 37.950 577.050 40.050 ;
        RECT 586.950 37.950 589.050 40.050 ;
        RECT 598.950 37.950 601.050 40.050 ;
        RECT 607.950 37.950 610.050 40.050 ;
        RECT 616.950 37.950 619.050 40.050 ;
        RECT 562.800 34.950 564.900 37.050 ;
        RECT 565.950 34.950 568.050 37.050 ;
        RECT 526.950 31.950 529.050 34.050 ;
        RECT 520.950 25.950 523.050 28.050 ;
        RECT 526.950 26.100 529.050 28.200 ;
        RECT 532.950 27.000 535.050 31.050 ;
        RECT 517.950 16.950 520.050 19.050 ;
        RECT 521.400 16.050 522.450 25.950 ;
        RECT 527.400 25.350 528.600 26.100 ;
        RECT 533.400 25.350 534.600 27.000 ;
        RECT 541.950 25.950 544.050 28.050 ;
        RECT 547.950 26.100 550.050 28.200 ;
        RECT 553.950 27.000 556.050 31.050 ;
        RECT 563.400 28.200 564.450 34.950 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 530.400 21.900 531.600 22.650 ;
        RECT 536.400 21.900 537.600 22.650 ;
        RECT 529.950 16.950 532.050 21.900 ;
        RECT 535.950 19.800 538.050 21.900 ;
        RECT 457.950 13.950 460.050 16.050 ;
        RECT 469.950 13.950 472.050 16.050 ;
        RECT 490.950 13.950 496.050 16.050 ;
        RECT 504.000 15.900 507.000 16.050 ;
        RECT 502.950 13.950 508.050 15.900 ;
        RECT 520.950 13.950 523.050 16.050 ;
        RECT 448.950 7.950 451.050 10.050 ;
        RECT 454.950 7.950 457.050 10.050 ;
        RECT 458.400 7.050 459.450 13.950 ;
        RECT 502.950 13.800 505.050 13.950 ;
        RECT 505.950 13.800 508.050 13.950 ;
        RECT 433.950 5.400 438.450 7.050 ;
        RECT 433.950 4.950 438.000 5.400 ;
        RECT 457.950 4.950 460.050 7.050 ;
        RECT 505.950 6.450 508.050 7.050 ;
        RECT 511.950 6.450 514.050 7.050 ;
        RECT 505.950 5.400 514.050 6.450 ;
        RECT 505.950 4.950 508.050 5.400 ;
        RECT 511.950 4.950 514.050 5.400 ;
        RECT 542.400 4.050 543.450 25.950 ;
        RECT 548.400 25.350 549.600 26.100 ;
        RECT 554.400 25.350 555.600 27.000 ;
        RECT 562.950 26.100 565.050 28.200 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 551.400 21.000 552.600 22.650 ;
        RECT 550.950 16.950 553.050 21.000 ;
        RECT 557.400 20.400 558.600 22.650 ;
        RECT 566.400 21.900 567.450 34.950 ;
        RECT 575.400 27.600 576.450 37.950 ;
        RECT 575.400 25.350 576.600 27.600 ;
        RECT 580.950 26.100 583.050 28.200 ;
        RECT 581.400 25.350 582.600 26.100 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 572.400 21.900 573.600 22.650 ;
        RECT 578.400 21.900 579.600 22.650 ;
        RECT 557.400 16.050 558.450 20.400 ;
        RECT 565.950 19.800 568.050 21.900 ;
        RECT 571.950 19.800 574.050 21.900 ;
        RECT 577.950 19.800 580.050 21.900 ;
        RECT 556.950 13.950 559.050 16.050 ;
        RECT 587.400 7.050 588.450 37.950 ;
        RECT 589.950 31.950 592.050 34.050 ;
        RECT 590.400 19.050 591.450 31.950 ;
        RECT 599.400 27.600 600.450 37.950 ;
        RECT 599.400 25.350 600.600 27.600 ;
        RECT 604.950 26.100 607.050 28.200 ;
        RECT 608.400 28.050 609.450 37.950 ;
        RECT 617.400 31.050 618.450 37.950 ;
        RECT 628.950 31.950 631.050 34.050 ;
        RECT 610.950 28.950 613.050 31.050 ;
        RECT 616.950 28.950 619.050 31.050 ;
        RECT 605.400 25.350 606.600 26.100 ;
        RECT 607.950 25.950 610.050 28.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 596.400 21.000 597.600 22.650 ;
        RECT 602.400 21.900 603.600 22.650 ;
        RECT 611.400 21.900 612.450 28.950 ;
        RECT 613.950 25.950 616.050 28.050 ;
        RECT 622.950 26.100 625.050 28.200 ;
        RECT 629.400 27.600 630.450 31.950 ;
        RECT 638.400 31.050 639.450 53.400 ;
        RECT 643.950 52.800 646.050 54.900 ;
        RECT 653.400 49.050 654.450 65.400 ;
        RECT 670.950 64.950 673.050 67.050 ;
        RECT 658.950 59.100 661.050 61.200 ;
        RECT 664.950 59.100 667.050 61.200 ;
        RECT 659.400 58.350 660.600 59.100 ;
        RECT 665.400 58.350 666.600 59.100 ;
        RECT 670.950 58.950 673.050 61.050 ;
        RECT 673.950 59.100 676.050 61.200 ;
        RECT 677.400 61.050 678.450 112.950 ;
        RECT 689.400 106.200 690.450 124.950 ;
        RECT 692.400 108.450 693.450 131.400 ;
        RECT 697.950 130.800 700.050 132.900 ;
        RECT 697.950 109.950 700.050 112.050 ;
        RECT 692.400 108.000 696.450 108.450 ;
        RECT 692.400 107.400 697.050 108.000 ;
        RECT 682.950 104.100 685.050 106.200 ;
        RECT 688.950 104.100 691.050 106.200 ;
        RECT 683.400 103.350 684.600 104.100 ;
        RECT 689.400 103.350 690.600 104.100 ;
        RECT 694.950 103.950 697.050 107.400 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 686.400 98.400 687.600 100.650 ;
        RECT 692.400 99.900 693.600 100.650 ;
        RECT 686.400 88.050 687.450 98.400 ;
        RECT 691.950 97.800 694.050 99.900 ;
        RECT 694.950 97.950 697.050 100.050 ;
        RECT 698.400 99.900 699.450 109.950 ;
        RECT 704.400 105.450 705.450 148.950 ;
        RECT 706.950 145.950 709.050 148.050 ;
        RECT 727.950 145.950 730.050 148.050 ;
        RECT 707.400 121.050 708.450 145.950 ;
        RECT 715.950 137.100 718.050 139.200 ;
        RECT 721.950 137.100 724.050 139.200 ;
        RECT 716.400 136.350 717.600 137.100 ;
        RECT 722.400 136.350 723.600 137.100 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 713.400 132.900 714.600 133.650 ;
        RECT 712.950 130.800 715.050 132.900 ;
        RECT 719.400 131.400 720.600 133.650 ;
        RECT 712.950 124.950 715.050 127.050 ;
        RECT 706.950 118.950 709.050 121.050 ;
        RECT 706.950 109.950 709.050 112.050 ;
        RECT 701.400 104.400 705.450 105.450 ;
        RECT 707.400 105.600 708.450 109.950 ;
        RECT 713.400 105.600 714.450 124.950 ;
        RECT 685.950 85.950 688.050 88.050 ;
        RECT 682.950 64.950 685.050 67.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 662.400 53.400 663.600 55.650 ;
        RECT 652.950 46.950 655.050 49.050 ;
        RECT 640.950 37.950 643.050 40.050 ;
        RECT 629.400 27.450 630.600 27.600 ;
        RECT 631.950 27.450 634.050 31.050 ;
        RECT 637.950 28.950 640.050 31.050 ;
        RECT 629.400 27.000 634.050 27.450 ;
        RECT 629.400 26.400 633.450 27.000 ;
        RECT 589.950 13.950 592.050 19.050 ;
        RECT 595.950 16.950 598.050 21.000 ;
        RECT 601.950 19.800 604.050 21.900 ;
        RECT 610.950 19.800 613.050 21.900 ;
        RECT 614.400 10.050 615.450 25.950 ;
        RECT 623.400 25.350 624.600 26.100 ;
        RECT 629.400 25.350 630.600 26.400 ;
        RECT 634.950 25.950 637.050 28.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 620.400 21.000 621.600 22.650 ;
        RECT 626.400 21.900 627.600 22.650 ;
        RECT 619.950 16.950 622.050 21.000 ;
        RECT 625.950 19.800 628.050 21.900 ;
        RECT 635.400 16.050 636.450 25.950 ;
        RECT 638.400 21.900 639.450 28.950 ;
        RECT 641.400 28.050 642.450 37.950 ;
        RECT 662.400 34.050 663.450 53.400 ;
        RECT 646.950 31.950 649.050 34.050 ;
        RECT 661.950 31.950 664.050 34.050 ;
        RECT 640.950 25.950 643.050 28.050 ;
        RECT 647.400 27.600 648.450 31.950 ;
        RECT 671.400 31.050 672.450 58.950 ;
        RECT 674.400 46.050 675.450 59.100 ;
        RECT 676.950 58.950 679.050 61.050 ;
        RECT 683.400 60.600 684.450 64.950 ;
        RECT 683.400 58.350 684.600 60.600 ;
        RECT 688.950 59.100 691.050 61.200 ;
        RECT 689.400 58.350 690.600 59.100 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 680.400 54.900 681.600 55.650 ;
        RECT 686.400 54.900 687.600 55.650 ;
        RECT 695.400 54.900 696.450 97.950 ;
        RECT 697.950 97.800 700.050 99.900 ;
        RECT 701.400 88.050 702.450 104.400 ;
        RECT 707.400 103.350 708.600 105.600 ;
        RECT 713.400 103.350 714.600 105.600 ;
        RECT 719.400 105.450 720.450 131.400 ;
        RECT 728.400 127.050 729.450 145.950 ;
        RECT 736.950 137.100 739.050 139.200 ;
        RECT 737.400 136.350 738.600 137.100 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 734.400 131.400 735.600 133.650 ;
        RECT 734.400 127.050 735.450 131.400 ;
        RECT 739.950 130.950 742.050 133.050 ;
        RECT 727.950 124.950 730.050 127.050 ;
        RECT 733.950 124.950 736.050 127.050 ;
        RECT 734.400 121.050 735.450 124.950 ;
        RECT 740.400 121.050 741.450 130.950 ;
        RECT 733.950 118.950 736.050 121.050 ;
        RECT 739.950 118.950 742.050 121.050 ;
        RECT 743.400 118.050 744.450 157.950 ;
        RECT 746.400 157.050 747.450 175.950 ;
        RECT 748.800 175.800 750.900 177.900 ;
        RECT 751.950 175.950 754.050 178.050 ;
        RECT 754.950 175.950 757.050 178.050 ;
        RECT 758.400 177.000 759.600 178.650 ;
        RECT 767.400 177.900 768.600 178.650 ;
        RECT 751.950 169.950 754.050 174.900 ;
        RECT 757.950 172.950 760.050 177.000 ;
        RECT 766.950 175.800 769.050 177.900 ;
        RECT 763.950 172.950 766.050 175.050 ;
        RECT 756.000 171.900 759.000 172.050 ;
        RECT 754.950 169.950 760.050 171.900 ;
        RECT 754.950 169.800 757.050 169.950 ;
        RECT 757.950 169.800 760.050 169.950 ;
        RECT 751.950 160.950 754.050 163.050 ;
        RECT 745.950 154.950 748.050 157.050 ;
        RECT 752.400 138.600 753.450 160.950 ;
        RECT 764.400 160.050 765.450 172.950 ;
        RECT 763.950 157.950 766.050 160.050 ;
        RECT 752.400 136.350 753.600 138.600 ;
        RECT 757.950 137.100 760.050 139.200 ;
        RECT 758.400 136.350 759.600 137.100 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 749.400 131.400 750.600 133.650 ;
        RECT 755.400 132.900 756.600 133.650 ;
        RECT 764.400 132.900 765.450 157.950 ;
        RECT 770.400 154.050 771.450 187.950 ;
        RECT 769.950 151.950 772.050 154.050 ;
        RECT 773.400 148.050 774.450 217.950 ;
        RECT 779.400 217.200 780.450 235.950 ;
        RECT 794.400 228.450 795.450 265.950 ;
        RECT 803.400 261.600 804.450 286.950 ;
        RECT 806.400 277.050 807.450 310.950 ;
        RECT 809.400 289.050 810.450 328.950 ;
        RECT 815.400 328.050 816.450 340.950 ;
        RECT 824.400 340.200 825.450 343.950 ;
        RECT 827.400 343.050 828.450 347.400 ;
        RECT 829.950 343.950 832.050 346.050 ;
        RECT 826.950 340.950 829.050 343.050 ;
        RECT 823.950 338.100 826.050 340.200 ;
        RECT 830.400 339.600 831.450 343.950 ;
        RECT 824.400 337.350 825.600 338.100 ;
        RECT 830.400 337.350 831.600 339.600 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 821.400 332.400 822.600 334.650 ;
        RECT 827.400 333.000 828.600 334.650 ;
        RECT 821.400 328.050 822.450 332.400 ;
        RECT 826.950 328.950 829.050 333.000 ;
        RECT 814.950 325.950 817.050 328.050 ;
        RECT 820.950 325.950 823.050 328.050 ;
        RECT 836.400 327.450 837.450 355.950 ;
        RECT 839.400 352.050 840.450 359.400 ;
        RECT 838.950 349.950 841.050 352.050 ;
        RECT 842.400 339.450 843.450 364.950 ;
        RECT 845.400 364.050 846.450 403.950 ;
        RECT 857.400 403.050 858.450 424.950 ;
        RECT 859.950 421.950 862.050 424.050 ;
        RECT 860.400 406.050 861.450 421.950 ;
        RECT 863.400 418.200 864.450 442.950 ;
        RECT 866.400 433.050 867.450 484.950 ;
        RECT 871.950 466.950 874.050 469.050 ;
        RECT 868.950 451.950 871.050 454.050 ;
        RECT 865.950 430.950 868.050 433.050 ;
        RECT 869.400 424.050 870.450 451.950 ;
        RECT 872.400 451.050 873.450 466.950 ;
        RECT 887.400 463.050 888.450 499.950 ;
        RECT 890.400 496.050 891.450 527.100 ;
        RECT 899.400 526.350 900.600 528.600 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 896.400 521.400 897.600 523.650 ;
        RECT 902.400 521.400 903.600 523.650 ;
        RECT 896.400 514.050 897.450 521.400 ;
        RECT 895.950 511.950 898.050 514.050 ;
        RECT 902.400 511.050 903.450 521.400 ;
        RECT 901.950 508.950 904.050 511.050 ;
        RECT 895.950 505.950 898.050 508.050 ;
        RECT 889.950 493.950 892.050 496.050 ;
        RECT 896.400 495.600 897.450 505.950 ;
        RECT 908.400 502.050 909.450 559.950 ;
        RECT 907.950 499.950 910.050 502.050 ;
        RECT 903.000 495.600 907.050 496.050 ;
        RECT 896.400 493.350 897.600 495.600 ;
        RECT 902.400 493.950 907.050 495.600 ;
        RECT 907.950 493.950 910.050 496.050 ;
        RECT 902.400 493.350 903.600 493.950 ;
        RECT 892.950 490.950 895.050 493.050 ;
        RECT 895.950 490.950 898.050 493.050 ;
        RECT 898.950 490.950 901.050 493.050 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 893.400 490.050 894.600 490.650 ;
        RECT 889.950 488.400 894.600 490.050 ;
        RECT 899.400 488.400 900.600 490.650 ;
        RECT 889.950 487.950 894.000 488.400 ;
        RECT 889.950 484.800 892.050 486.900 ;
        RECT 886.950 460.950 889.050 463.050 ;
        RECT 880.950 457.950 883.050 460.050 ;
        RECT 871.950 448.950 874.050 451.050 ;
        RECT 874.950 450.000 877.050 454.050 ;
        RECT 881.400 450.600 882.450 457.950 ;
        RECT 875.400 448.350 876.600 450.000 ;
        RECT 881.400 448.350 882.600 450.600 ;
        RECT 874.950 445.950 877.050 448.050 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 871.950 442.950 874.050 445.050 ;
        RECT 878.400 443.400 879.600 445.650 ;
        RECT 884.400 444.900 885.600 445.650 ;
        RECT 890.400 445.050 891.450 484.800 ;
        RECT 892.950 472.950 895.050 475.050 ;
        RECT 893.400 451.050 894.450 472.950 ;
        RECT 899.400 454.050 900.450 488.400 ;
        RECT 908.400 487.050 909.450 493.950 ;
        RECT 911.400 489.450 912.450 595.650 ;
        RECT 916.950 580.950 919.050 583.050 ;
        RECT 913.950 577.950 916.050 580.050 ;
        RECT 914.400 574.050 915.450 577.950 ;
        RECT 913.950 571.950 916.050 574.050 ;
        RECT 917.400 573.600 918.450 580.950 ;
        RECT 920.400 580.050 921.450 599.400 ;
        RECT 935.400 598.050 936.450 637.950 ;
        RECT 934.950 595.950 937.050 598.050 ;
        RECT 919.950 577.950 922.050 580.050 ;
        RECT 931.950 577.950 934.050 580.050 ;
        RECT 917.400 571.350 918.600 573.600 ;
        RECT 922.950 572.100 925.050 577.050 ;
        RECT 923.400 571.350 924.600 572.100 ;
        RECT 916.950 568.950 919.050 571.050 ;
        RECT 919.950 568.950 922.050 571.050 ;
        RECT 922.950 568.950 925.050 571.050 ;
        RECT 925.950 568.950 928.050 571.050 ;
        RECT 920.400 567.900 921.600 568.650 ;
        RECT 919.950 565.800 922.050 567.900 ;
        RECT 926.400 567.450 927.600 568.650 ;
        RECT 926.400 566.400 930.450 567.450 ;
        RECT 920.400 564.450 921.450 565.800 ;
        RECT 917.400 563.400 921.450 564.450 ;
        RECT 917.400 528.600 918.450 563.400 ;
        RECT 929.400 556.050 930.450 566.400 ;
        RECT 928.950 553.950 931.050 556.050 ;
        RECT 925.950 547.950 928.050 550.050 ;
        RECT 917.400 526.350 918.600 528.600 ;
        RECT 916.950 523.950 919.050 526.050 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 913.950 520.950 916.050 523.050 ;
        RECT 920.400 522.000 921.600 523.650 ;
        RECT 926.400 523.050 927.450 547.950 ;
        RECT 914.400 511.050 915.450 520.950 ;
        RECT 919.950 517.950 922.050 522.000 ;
        RECT 925.950 520.950 928.050 523.050 ;
        RECT 925.950 517.800 928.050 519.900 ;
        RECT 919.950 511.950 922.050 514.050 ;
        RECT 913.950 508.950 916.050 511.050 ;
        RECT 914.400 496.050 915.450 508.950 ;
        RECT 913.950 493.950 916.050 496.050 ;
        RECT 920.400 495.600 921.450 511.950 ;
        RECT 926.400 496.050 927.450 517.800 ;
        RECT 920.400 493.350 921.600 495.600 ;
        RECT 925.950 493.950 928.050 496.050 ;
        RECT 916.950 490.950 919.050 493.050 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 922.950 490.950 925.050 493.050 ;
        RECT 911.400 488.400 915.450 489.450 ;
        RECT 901.950 484.950 904.050 487.050 ;
        RECT 907.950 484.950 910.050 487.050 ;
        RECT 902.400 460.050 903.450 484.950 ;
        RECT 904.950 475.950 907.050 478.050 ;
        RECT 901.950 457.950 904.050 460.050 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 898.950 450.000 901.050 454.050 ;
        RECT 905.400 450.600 906.450 475.950 ;
        RECT 910.950 469.950 913.050 472.050 ;
        RECT 907.950 460.950 910.050 463.050 ;
        RECT 908.400 451.050 909.450 460.950 ;
        RECT 899.400 448.350 900.600 450.000 ;
        RECT 905.400 448.350 906.600 450.600 ;
        RECT 907.950 448.950 910.050 451.050 ;
        RECT 895.950 445.950 898.050 448.050 ;
        RECT 898.950 445.950 901.050 448.050 ;
        RECT 901.950 445.950 904.050 448.050 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 872.400 427.050 873.450 442.950 ;
        RECT 874.950 433.950 877.050 436.050 ;
        RECT 871.950 424.950 874.050 427.050 ;
        RECT 868.950 421.950 871.050 424.050 ;
        RECT 875.400 421.050 876.450 433.950 ;
        RECT 874.950 418.950 877.050 421.050 ;
        RECT 862.950 416.100 865.050 418.200 ;
        RECT 871.950 416.100 874.050 418.200 ;
        RECT 863.400 411.900 864.450 416.100 ;
        RECT 872.400 415.350 873.600 416.100 ;
        RECT 866.100 412.950 868.200 415.050 ;
        RECT 871.500 412.950 873.600 415.050 ;
        RECT 874.800 412.950 876.900 415.050 ;
        RECT 862.950 409.800 865.050 411.900 ;
        RECT 866.400 410.400 867.600 412.650 ;
        RECT 875.400 411.900 876.600 412.650 ;
        RECT 859.950 403.950 862.050 406.050 ;
        RECT 856.950 400.950 859.050 403.050 ;
        RECT 853.950 379.950 856.050 382.050 ;
        RECT 847.950 373.950 850.050 376.050 ;
        RECT 844.950 361.950 847.050 364.050 ;
        RECT 845.400 346.050 846.450 361.950 ;
        RECT 848.400 358.050 849.450 373.950 ;
        RECT 854.400 372.600 855.450 379.950 ;
        RECT 854.400 370.350 855.600 372.600 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 857.400 366.450 858.600 367.650 ;
        RECT 859.950 366.450 862.050 367.050 ;
        RECT 857.400 365.400 862.050 366.450 ;
        RECT 859.950 364.950 862.050 365.400 ;
        RECT 853.950 358.950 856.050 361.050 ;
        RECT 847.950 355.950 850.050 358.050 ;
        RECT 844.950 343.950 847.050 346.050 ;
        RECT 846.000 342.900 849.000 343.050 ;
        RECT 844.950 342.450 849.000 342.900 ;
        RECT 844.950 340.950 849.450 342.450 ;
        RECT 844.950 340.800 847.050 340.950 ;
        RECT 839.400 338.400 843.450 339.450 ;
        RECT 848.400 339.600 849.450 340.950 ;
        RECT 854.400 339.600 855.450 358.950 ;
        RECT 839.400 333.450 840.450 338.400 ;
        RECT 848.400 337.350 849.600 339.600 ;
        RECT 854.400 337.350 855.600 339.600 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 845.400 333.900 846.600 334.650 ;
        RECT 839.400 332.400 843.450 333.450 ;
        RECT 838.950 327.450 841.050 328.050 ;
        RECT 836.400 326.400 841.050 327.450 ;
        RECT 838.950 325.950 841.050 326.400 ;
        RECT 817.800 298.200 819.900 300.300 ;
        RECT 826.800 298.500 828.900 300.600 ;
        RECT 814.950 294.450 817.050 295.200 ;
        RECT 812.400 293.400 817.050 294.450 ;
        RECT 808.950 286.950 811.050 289.050 ;
        RECT 812.400 280.050 813.450 293.400 ;
        RECT 814.950 293.100 817.050 293.400 ;
        RECT 815.400 292.350 816.600 293.100 ;
        RECT 815.100 289.950 817.200 292.050 ;
        RECT 818.100 285.600 819.000 298.200 ;
        RECT 824.400 295.350 825.600 297.600 ;
        RECT 824.100 292.950 826.200 295.050 ;
        RECT 819.900 291.900 822.000 292.200 ;
        RECT 828.000 291.900 828.900 298.500 ;
        RECT 819.900 291.000 828.900 291.900 ;
        RECT 819.900 290.100 822.000 291.000 ;
        RECT 825.000 289.200 827.100 290.100 ;
        RECT 819.900 288.000 827.100 289.200 ;
        RECT 819.900 287.100 822.000 288.000 ;
        RECT 817.500 283.500 819.600 285.600 ;
        RECT 824.100 284.100 826.200 286.200 ;
        RECT 828.000 285.900 828.900 291.000 ;
        RECT 829.800 289.950 831.900 292.050 ;
        RECT 830.400 288.900 831.600 289.650 ;
        RECT 829.950 286.800 832.050 288.900 ;
        RECT 827.400 283.800 829.500 285.900 ;
        RECT 824.400 281.550 825.600 283.800 ;
        RECT 811.950 277.950 814.050 280.050 ;
        RECT 805.950 274.950 808.050 277.050 ;
        RECT 824.400 265.050 825.450 281.550 ;
        RECT 839.400 280.050 840.450 325.950 ;
        RECT 838.950 277.950 841.050 280.050 ;
        RECT 803.400 259.350 804.600 261.600 ;
        RECT 808.950 261.000 811.050 265.050 ;
        RECT 817.950 262.950 820.050 265.050 ;
        RECT 823.950 262.950 826.050 265.050 ;
        RECT 809.400 259.350 810.600 261.000 ;
        RECT 811.950 259.950 817.050 262.050 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 800.400 255.900 801.600 256.650 ;
        RECT 806.400 255.900 807.600 256.650 ;
        RECT 818.400 255.900 819.450 262.950 ;
        RECT 820.950 261.600 825.000 262.050 ;
        RECT 820.950 259.950 825.600 261.600 ;
        RECT 829.950 260.100 832.050 262.200 ;
        RECT 824.400 259.350 825.600 259.950 ;
        RECT 830.400 259.350 831.600 260.100 ;
        RECT 838.950 259.950 841.050 262.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 799.950 253.800 802.050 255.900 ;
        RECT 805.950 253.800 808.050 255.900 ;
        RECT 817.950 253.800 820.050 255.900 ;
        RECT 827.400 254.400 828.600 256.650 ;
        RECT 833.400 255.900 834.600 256.650 ;
        RECT 832.950 255.450 835.050 255.900 ;
        RECT 832.950 254.400 837.450 255.450 ;
        RECT 791.400 227.400 795.450 228.450 ;
        RECT 784.950 223.950 787.050 226.050 ;
        RECT 778.950 215.100 781.050 217.200 ;
        RECT 785.400 216.600 786.450 223.950 ;
        RECT 779.400 214.350 780.600 215.100 ;
        RECT 785.400 214.350 786.600 216.600 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 782.400 209.400 783.600 211.650 ;
        RECT 782.400 196.050 783.450 209.400 ;
        RECT 781.950 193.950 784.050 196.050 ;
        RECT 784.950 187.950 787.050 190.050 ;
        RECT 778.950 182.100 781.050 184.200 ;
        RECT 785.400 183.600 786.450 187.950 ;
        RECT 791.400 184.050 792.450 227.400 ;
        RECT 793.950 223.950 796.050 226.050 ;
        RECT 794.400 210.900 795.450 223.950 ;
        RECT 800.400 223.050 801.450 253.800 ;
        RECT 827.400 252.450 828.450 254.400 ;
        RECT 832.950 253.800 835.050 254.400 ;
        RECT 824.400 251.400 828.450 252.450 ;
        RECT 824.400 238.050 825.450 251.400 ;
        RECT 832.950 250.650 835.050 252.750 ;
        RECT 823.950 235.950 826.050 238.050 ;
        RECT 799.950 220.950 802.050 223.050 ;
        RECT 799.950 215.100 802.050 217.200 ;
        RECT 805.950 215.100 808.050 217.200 ;
        RECT 814.950 215.100 817.050 217.200 ;
        RECT 824.400 216.600 825.450 235.950 ;
        RECT 800.400 214.350 801.600 215.100 ;
        RECT 806.400 214.350 807.600 215.100 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 803.400 210.900 804.600 211.650 ;
        RECT 793.950 208.800 796.050 210.900 ;
        RECT 802.950 208.800 805.050 210.900 ;
        RECT 809.400 209.400 810.600 211.650 ;
        RECT 809.400 204.450 810.450 209.400 ;
        RECT 815.400 205.050 816.450 215.100 ;
        RECT 824.400 214.350 825.600 216.600 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 826.950 211.950 829.050 214.050 ;
        RECT 821.400 209.400 822.600 211.650 ;
        RECT 827.400 209.400 828.600 211.650 ;
        RECT 833.400 211.050 834.450 250.650 ;
        RECT 817.950 205.950 820.050 208.050 ;
        RECT 809.400 203.400 813.450 204.450 ;
        RECT 808.950 199.950 811.050 202.050 ;
        RECT 779.400 181.350 780.600 182.100 ;
        RECT 785.400 181.350 786.600 183.600 ;
        RECT 790.950 181.950 793.050 184.050 ;
        RECT 796.950 182.100 799.050 184.200 ;
        RECT 802.950 182.100 805.050 184.200 ;
        RECT 809.400 183.600 810.450 199.950 ;
        RECT 812.400 187.050 813.450 203.400 ;
        RECT 814.950 202.950 817.050 205.050 ;
        RECT 818.400 199.050 819.450 205.950 ;
        RECT 821.400 205.050 822.450 209.400 ;
        RECT 820.950 204.450 823.050 205.050 ;
        RECT 820.950 203.400 825.450 204.450 ;
        RECT 820.950 202.950 823.050 203.400 ;
        RECT 817.950 196.950 820.050 199.050 ;
        RECT 820.950 187.950 823.050 190.050 ;
        RECT 811.950 184.950 814.050 187.050 ;
        RECT 817.950 184.950 820.050 187.050 ;
        RECT 778.950 178.950 781.050 181.050 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 782.400 177.900 783.600 178.650 ;
        RECT 781.950 175.800 784.050 177.900 ;
        RECT 788.400 176.400 789.600 178.650 ;
        RECT 788.400 166.050 789.450 176.400 ;
        RECT 794.400 172.050 795.450 178.950 ;
        RECT 793.950 169.950 796.050 172.050 ;
        RECT 797.400 166.050 798.450 182.100 ;
        RECT 803.400 181.350 804.600 182.100 ;
        RECT 809.400 181.350 810.600 183.600 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 799.950 172.950 802.050 178.050 ;
        RECT 806.400 176.400 807.600 178.650 ;
        RECT 812.400 176.400 813.600 178.650 ;
        RECT 806.400 172.050 807.450 176.400 ;
        RECT 805.950 169.950 808.050 172.050 ;
        RECT 775.950 163.950 778.050 166.050 ;
        RECT 787.950 163.950 790.050 166.050 ;
        RECT 796.950 163.950 799.050 166.050 ;
        RECT 772.950 145.950 775.050 148.050 ;
        RECT 769.950 137.100 772.050 139.200 ;
        RECT 776.400 139.050 777.450 163.950 ;
        RECT 805.950 160.950 808.050 163.050 ;
        RECT 802.950 154.950 805.050 157.050 ;
        RECT 799.950 151.950 802.050 154.050 ;
        RECT 787.950 148.950 790.050 151.050 ;
        RECT 781.950 145.950 784.050 148.050 ;
        RECT 770.400 136.350 771.600 137.100 ;
        RECT 775.950 136.950 778.050 139.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 773.400 132.900 774.600 133.650 ;
        RECT 749.400 129.450 750.450 131.400 ;
        RECT 754.950 130.800 757.050 132.900 ;
        RECT 763.950 130.800 766.050 132.900 ;
        RECT 772.950 130.800 775.050 132.900 ;
        RECT 749.400 128.400 753.450 129.450 ;
        RECT 748.950 124.950 751.050 127.050 ;
        RECT 742.950 115.950 745.050 118.050 ;
        RECT 730.950 112.950 733.050 115.050 ;
        RECT 731.400 105.600 732.450 112.950 ;
        RECT 719.400 104.400 723.450 105.450 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 703.950 97.950 706.050 100.050 ;
        RECT 710.400 99.900 711.600 100.650 ;
        RECT 704.400 94.050 705.450 97.950 ;
        RECT 709.950 97.800 712.050 99.900 ;
        RECT 716.400 98.400 717.600 100.650 ;
        RECT 722.400 99.900 723.450 104.400 ;
        RECT 731.400 103.350 732.600 105.600 ;
        RECT 736.950 105.000 739.050 109.050 ;
        RECT 745.950 106.950 748.050 109.050 ;
        RECT 737.400 103.350 738.600 105.000 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 734.400 99.900 735.600 100.650 ;
        RECT 716.400 94.050 717.450 98.400 ;
        RECT 721.950 97.800 724.050 99.900 ;
        RECT 733.950 97.800 736.050 99.900 ;
        RECT 740.400 98.400 741.600 100.650 ;
        RECT 703.950 91.950 706.050 94.050 ;
        RECT 715.950 91.950 718.050 94.050 ;
        RECT 721.950 91.950 724.050 94.050 ;
        RECT 700.950 85.950 703.050 88.050 ;
        RECT 701.400 61.200 702.450 85.950 ;
        RECT 704.400 79.050 705.450 91.950 ;
        RECT 703.950 76.950 706.050 79.050 ;
        RECT 718.950 76.950 721.050 79.050 ;
        RECT 706.950 64.950 709.050 67.050 ;
        RECT 700.950 59.100 703.050 61.200 ;
        RECT 707.400 60.600 708.450 64.950 ;
        RECT 707.400 58.350 708.600 60.600 ;
        RECT 712.950 59.100 715.050 61.200 ;
        RECT 713.400 58.350 714.600 59.100 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 679.950 52.800 682.050 54.900 ;
        RECT 685.950 52.800 688.050 54.900 ;
        RECT 694.950 52.800 697.050 54.900 ;
        RECT 704.400 53.400 705.600 55.650 ;
        RECT 710.400 54.900 711.600 55.650 ;
        RECT 704.400 49.050 705.450 53.400 ;
        RECT 709.950 52.800 712.050 54.900 ;
        RECT 679.950 46.950 682.050 49.050 ;
        RECT 703.800 46.950 705.900 49.050 ;
        RECT 706.950 46.950 709.050 49.050 ;
        RECT 673.950 43.950 676.050 46.050 ;
        RECT 649.950 28.950 655.050 31.050 ;
        RECT 670.950 28.950 673.050 31.050 ;
        RECT 676.950 28.950 679.050 31.050 ;
        RECT 647.400 25.350 648.600 27.600 ;
        RECT 653.400 27.450 654.600 27.600 ;
        RECT 653.400 26.400 660.450 27.450 ;
        RECT 653.400 25.350 654.600 26.400 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 644.400 21.900 645.600 22.650 ;
        RECT 650.400 21.900 651.600 22.650 ;
        RECT 637.950 19.800 640.050 21.900 ;
        RECT 643.950 19.800 646.050 21.900 ;
        RECT 649.950 19.800 652.050 21.900 ;
        RECT 659.400 16.050 660.450 26.400 ;
        RECT 667.950 26.100 670.050 28.200 ;
        RECT 668.400 25.350 669.600 26.100 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 665.400 20.400 666.600 22.650 ;
        RECT 671.400 21.900 672.600 22.650 ;
        RECT 665.400 18.450 666.450 20.400 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 665.400 17.400 669.450 18.450 ;
        RECT 634.950 13.950 637.050 16.050 ;
        RECT 658.950 13.950 661.050 16.050 ;
        RECT 661.950 13.950 667.050 16.050 ;
        RECT 668.400 13.050 669.450 17.400 ;
        RECT 677.400 13.050 678.450 28.950 ;
        RECT 680.400 21.900 681.450 46.950 ;
        RECT 700.800 45.000 702.900 46.050 ;
        RECT 700.800 43.950 703.050 45.000 ;
        RECT 688.950 40.950 691.050 43.050 ;
        RECT 700.950 42.450 703.050 43.950 ;
        RECT 707.400 42.450 708.450 46.950 ;
        RECT 700.950 42.000 708.450 42.450 ;
        RECT 701.400 41.400 708.450 42.000 ;
        RECT 689.400 27.600 690.450 40.950 ;
        RECT 719.400 34.050 720.450 76.950 ;
        RECT 722.400 54.900 723.450 91.950 ;
        RECT 734.400 63.450 735.450 97.800 ;
        RECT 740.400 88.050 741.450 98.400 ;
        RECT 746.400 94.050 747.450 106.950 ;
        RECT 749.400 106.050 750.450 124.950 ;
        RECT 752.400 115.050 753.450 128.400 ;
        RECT 760.950 118.950 763.050 121.050 ;
        RECT 751.950 112.950 754.050 115.050 ;
        RECT 748.950 103.950 751.050 106.050 ;
        RECT 754.950 104.100 757.050 106.200 ;
        RECT 761.400 106.050 762.450 118.950 ;
        RECT 763.950 115.950 766.050 118.050 ;
        RECT 755.400 103.350 756.600 104.100 ;
        RECT 760.950 103.950 763.050 106.050 ;
        RECT 751.950 100.950 754.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 752.400 99.900 753.600 100.650 ;
        RECT 758.400 99.900 759.600 100.650 ;
        RECT 764.400 99.900 765.450 115.950 ;
        RECT 766.950 103.950 769.050 106.050 ;
        RECT 775.950 104.100 778.050 106.200 ;
        RECT 782.400 106.050 783.450 145.950 ;
        RECT 784.950 142.950 787.050 148.050 ;
        RECT 785.400 139.050 786.450 142.950 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 788.400 138.600 789.450 148.950 ;
        RECT 788.400 136.350 789.600 138.600 ;
        RECT 793.950 137.100 796.050 139.200 ;
        RECT 800.400 139.050 801.450 151.950 ;
        RECT 794.400 136.350 795.600 137.100 ;
        RECT 799.950 136.950 802.050 139.050 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 791.400 131.400 792.600 133.650 ;
        RECT 797.400 131.400 798.600 133.650 ;
        RECT 785.400 106.200 786.450 130.950 ;
        RECT 791.400 112.050 792.450 131.400 ;
        RECT 797.400 118.050 798.450 131.400 ;
        RECT 799.950 130.950 802.050 133.050 ;
        RECT 800.400 124.050 801.450 130.950 ;
        RECT 799.950 121.950 802.050 124.050 ;
        RECT 796.950 115.950 799.050 118.050 ;
        RECT 790.950 109.950 793.050 112.050 ;
        RECT 803.400 109.050 804.450 154.950 ;
        RECT 806.400 145.050 807.450 160.950 ;
        RECT 812.400 160.050 813.450 176.400 ;
        RECT 814.950 175.950 817.050 178.050 ;
        RECT 811.950 157.950 814.050 160.050 ;
        RECT 815.400 154.050 816.450 175.950 ;
        RECT 818.400 172.050 819.450 184.950 ;
        RECT 817.950 169.950 820.050 172.050 ;
        RECT 821.400 154.050 822.450 187.950 ;
        RECT 824.400 184.050 825.450 203.400 ;
        RECT 827.400 196.050 828.450 209.400 ;
        RECT 832.950 208.950 835.050 211.050 ;
        RECT 826.950 193.950 829.050 196.050 ;
        RECT 827.400 187.050 828.450 193.950 ;
        RECT 829.950 190.950 832.050 193.050 ;
        RECT 826.950 184.950 829.050 187.050 ;
        RECT 823.950 181.950 826.050 184.050 ;
        RECT 830.400 183.600 831.450 190.950 ;
        RECT 836.400 184.050 837.450 254.400 ;
        RECT 839.400 247.050 840.450 259.950 ;
        RECT 842.400 253.050 843.450 332.400 ;
        RECT 844.950 331.800 847.050 333.900 ;
        RECT 851.400 332.400 852.600 334.650 ;
        RECT 851.400 328.050 852.450 332.400 ;
        RECT 850.950 325.950 853.050 328.050 ;
        RECT 860.400 313.050 861.450 364.950 ;
        RECT 863.400 333.450 864.450 409.800 ;
        RECT 866.400 400.050 867.450 410.400 ;
        RECT 874.950 409.800 877.050 411.900 ;
        RECT 878.400 406.050 879.450 443.400 ;
        RECT 883.950 442.800 886.050 444.900 ;
        RECT 889.950 442.950 892.050 445.050 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 896.400 443.400 897.600 445.650 ;
        RECT 902.400 444.900 903.600 445.650 ;
        RECT 880.950 439.950 883.050 442.050 ;
        RECT 881.400 412.050 882.450 439.950 ;
        RECT 883.950 433.950 886.050 436.050 ;
        RECT 880.950 409.950 883.050 412.050 ;
        RECT 884.400 411.450 885.450 433.950 ;
        RECT 893.400 417.600 894.450 442.950 ;
        RECT 896.400 421.050 897.450 443.400 ;
        RECT 901.950 442.800 904.050 444.900 ;
        RECT 911.400 427.050 912.450 469.950 ;
        RECT 914.400 469.050 915.450 488.400 ;
        RECT 917.400 488.400 918.600 490.650 ;
        RECT 923.400 488.400 924.600 490.650 ;
        RECT 917.400 484.050 918.450 488.400 ;
        RECT 919.950 484.950 922.050 487.050 ;
        RECT 916.950 481.950 919.050 484.050 ;
        RECT 916.950 475.950 919.050 478.050 ;
        RECT 917.400 472.050 918.450 475.950 ;
        RECT 916.950 469.950 919.050 472.050 ;
        RECT 913.950 466.950 916.050 469.050 ;
        RECT 917.400 454.050 918.450 469.950 ;
        RECT 920.400 454.050 921.450 484.950 ;
        RECT 923.400 481.050 924.450 488.400 ;
        RECT 925.950 487.950 928.050 490.050 ;
        RECT 922.950 478.950 925.050 481.050 ;
        RECT 916.950 451.950 919.050 454.050 ;
        RECT 919.950 450.000 922.050 454.050 ;
        RECT 926.400 453.450 927.450 487.950 ;
        RECT 929.400 475.050 930.450 553.950 ;
        RECT 932.400 550.050 933.450 577.950 ;
        RECT 934.800 572.100 936.900 574.200 ;
        RECT 938.400 574.050 939.450 640.950 ;
        RECT 943.950 577.950 946.050 580.050 ;
        RECT 935.400 568.050 936.450 572.100 ;
        RECT 937.950 571.950 940.050 574.050 ;
        RECT 944.400 573.600 945.450 577.950 ;
        RECT 944.400 571.350 945.600 573.600 ;
        RECT 940.950 568.950 943.050 571.050 ;
        RECT 943.950 568.950 946.050 571.050 ;
        RECT 934.950 565.950 937.050 568.050 ;
        RECT 941.400 567.900 942.600 568.650 ;
        RECT 940.950 565.800 943.050 567.900 ;
        RECT 946.950 565.950 949.050 568.050 ;
        RECT 931.950 547.950 934.050 550.050 ;
        RECT 934.950 532.950 937.050 535.050 ;
        RECT 935.400 528.600 936.450 532.950 ;
        RECT 935.400 526.350 936.600 528.600 ;
        RECT 940.950 527.100 943.050 529.200 ;
        RECT 941.400 526.350 942.600 527.100 ;
        RECT 934.950 523.950 937.050 526.050 ;
        RECT 937.950 523.950 940.050 526.050 ;
        RECT 940.950 523.950 943.050 526.050 ;
        RECT 938.400 521.400 939.600 523.650 ;
        RECT 938.400 499.050 939.450 521.400 ;
        RECT 943.950 520.950 946.050 523.050 ;
        RECT 940.950 516.450 943.050 517.050 ;
        RECT 944.400 516.450 945.450 520.950 ;
        RECT 940.950 515.400 945.450 516.450 ;
        RECT 940.950 514.950 943.050 515.400 ;
        RECT 931.950 496.950 934.050 499.050 ;
        RECT 937.950 496.950 940.050 499.050 ;
        RECT 932.400 490.050 933.450 496.950 ;
        RECT 941.400 495.600 942.450 514.950 ;
        RECT 947.400 508.050 948.450 565.950 ;
        RECT 946.950 505.950 949.050 508.050 ;
        RECT 941.400 493.350 942.600 495.600 ;
        RECT 937.950 490.950 940.050 493.050 ;
        RECT 940.950 490.950 943.050 493.050 ;
        RECT 943.950 490.950 946.050 493.050 ;
        RECT 931.950 487.950 934.050 490.050 ;
        RECT 938.400 489.900 939.600 490.650 ;
        RECT 931.950 484.800 934.050 486.900 ;
        RECT 937.950 484.950 940.050 489.900 ;
        RECT 944.400 488.400 945.600 490.650 ;
        RECT 928.950 472.950 931.050 475.050 ;
        RECT 926.400 453.000 930.450 453.450 ;
        RECT 926.400 452.400 931.050 453.000 ;
        RECT 920.400 448.350 921.600 450.000 ;
        RECT 925.950 449.100 928.050 451.200 ;
        RECT 926.400 448.350 927.600 449.100 ;
        RECT 928.950 448.950 931.050 452.400 ;
        RECT 916.950 445.950 919.050 448.050 ;
        RECT 919.950 445.950 922.050 448.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 925.950 445.950 928.050 448.050 ;
        RECT 917.400 444.900 918.600 445.650 ;
        RECT 923.400 444.900 924.600 445.650 ;
        RECT 916.950 442.800 919.050 444.900 ;
        RECT 922.950 442.800 925.050 444.900 ;
        RECT 932.400 444.450 933.450 484.800 ;
        RECT 944.400 481.050 945.450 488.400 ;
        RECT 943.950 478.950 946.050 481.050 ;
        RECT 937.950 469.950 940.050 472.050 ;
        RECT 934.950 448.950 937.050 454.050 ;
        RECT 938.400 450.600 939.450 469.950 ;
        RECT 946.950 466.950 949.050 469.050 ;
        RECT 938.400 448.350 939.600 450.600 ;
        RECT 937.950 445.950 940.050 448.050 ;
        RECT 940.950 445.950 943.050 448.050 ;
        RECT 929.400 443.400 933.450 444.450 ;
        RECT 941.400 443.400 942.600 445.650 ;
        RECT 919.950 439.950 922.050 442.050 ;
        RECT 910.950 424.950 913.050 427.050 ;
        RECT 895.950 418.950 898.050 421.050 ;
        RECT 893.400 415.350 894.600 417.600 ;
        RECT 904.950 416.100 907.050 418.200 ;
        RECT 913.950 416.100 916.050 418.200 ;
        RECT 920.400 417.600 921.450 439.950 ;
        RECT 925.950 436.950 928.050 439.050 ;
        RECT 922.950 424.950 925.050 427.050 ;
        RECT 923.400 418.050 924.450 424.950 ;
        RECT 889.950 412.950 892.050 415.050 ;
        RECT 892.950 412.950 895.050 415.050 ;
        RECT 895.950 412.950 898.050 415.050 ;
        RECT 890.400 411.900 891.600 412.650 ;
        RECT 884.400 410.400 888.450 411.450 ;
        RECT 877.950 403.950 880.050 406.050 ;
        RECT 865.950 397.950 868.050 400.050 ;
        RECT 865.950 371.100 868.050 373.200 ;
        RECT 868.950 372.600 873.000 373.050 ;
        RECT 866.400 361.050 867.450 371.100 ;
        RECT 868.950 370.950 873.600 372.600 ;
        RECT 877.950 372.000 880.050 376.050 ;
        RECT 872.400 370.350 873.600 370.950 ;
        RECT 878.400 370.350 879.600 372.000 ;
        RECT 871.950 367.950 874.050 370.050 ;
        RECT 874.950 367.950 877.050 370.050 ;
        RECT 877.950 367.950 880.050 370.050 ;
        RECT 880.950 367.950 883.050 370.050 ;
        RECT 875.400 366.000 876.600 367.650 ;
        RECT 881.400 366.000 882.600 367.650 ;
        RECT 874.950 361.950 877.050 366.000 ;
        RECT 880.950 361.950 883.050 366.000 ;
        RECT 887.400 361.050 888.450 410.400 ;
        RECT 889.950 409.800 892.050 411.900 ;
        RECT 896.400 410.400 897.600 412.650 ;
        RECT 896.400 409.050 897.450 410.400 ;
        RECT 905.400 409.050 906.450 416.100 ;
        RECT 914.400 415.350 915.600 416.100 ;
        RECT 920.400 415.350 921.600 417.600 ;
        RECT 922.950 415.950 925.050 418.050 ;
        RECT 910.950 412.950 913.050 415.050 ;
        RECT 913.950 412.950 916.050 415.050 ;
        RECT 916.950 412.950 919.050 415.050 ;
        RECT 919.950 412.950 922.050 415.050 ;
        RECT 911.400 412.050 912.600 412.650 ;
        RECT 907.950 410.400 912.600 412.050 ;
        RECT 917.400 411.900 918.600 412.650 ;
        RECT 907.950 409.950 912.000 410.400 ;
        RECT 916.950 409.800 919.050 411.900 ;
        RECT 922.950 409.950 925.050 412.050 ;
        RECT 895.950 408.450 898.050 409.050 ;
        RECT 893.400 407.400 898.050 408.450 ;
        RECT 889.950 373.950 892.050 376.050 ;
        RECT 865.950 358.950 868.050 361.050 ;
        RECT 877.950 358.950 880.050 361.050 ;
        RECT 886.950 358.950 889.050 361.050 ;
        RECT 871.950 338.100 874.050 340.200 ;
        RECT 878.400 339.600 879.450 358.950 ;
        RECT 890.400 352.050 891.450 373.950 ;
        RECT 893.400 373.050 894.450 407.400 ;
        RECT 895.950 406.950 898.050 407.400 ;
        RECT 904.950 406.950 907.050 409.050 ;
        RECT 910.950 403.950 913.050 406.050 ;
        RECT 907.950 400.950 910.050 403.050 ;
        RECT 895.950 379.950 898.050 382.050 ;
        RECT 892.950 370.950 895.050 373.050 ;
        RECT 896.400 372.600 897.450 379.950 ;
        RECT 896.400 370.350 897.600 372.600 ;
        RECT 901.950 371.100 904.050 373.200 ;
        RECT 908.400 373.050 909.450 400.950 ;
        RECT 902.400 370.350 903.600 371.100 ;
        RECT 907.950 370.950 910.050 373.050 ;
        RECT 895.950 367.950 898.050 370.050 ;
        RECT 898.950 367.950 901.050 370.050 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 892.950 364.950 895.050 367.050 ;
        RECT 899.400 365.400 900.600 367.650 ;
        RECT 905.400 365.400 906.600 367.650 ;
        RECT 889.950 349.950 892.050 352.050 ;
        RECT 893.400 346.050 894.450 364.950 ;
        RECT 899.400 355.050 900.450 365.400 ;
        RECT 905.400 358.050 906.450 365.400 ;
        RECT 911.400 364.050 912.450 403.950 ;
        RECT 923.400 379.050 924.450 409.950 ;
        RECT 926.400 409.050 927.450 436.950 ;
        RECT 925.950 406.950 928.050 409.050 ;
        RECT 929.400 405.450 930.450 443.400 ;
        RECT 931.950 439.950 934.050 442.050 ;
        RECT 937.950 439.950 940.050 442.050 ;
        RECT 932.400 418.050 933.450 439.950 ;
        RECT 938.400 418.200 939.450 439.950 ;
        RECT 941.400 436.050 942.450 443.400 ;
        RECT 947.400 439.050 948.450 466.950 ;
        RECT 946.950 436.950 949.050 439.050 ;
        RECT 940.950 433.950 943.050 436.050 ;
        RECT 931.950 415.950 934.050 418.050 ;
        RECT 937.950 416.100 940.050 418.200 ;
        RECT 938.400 415.350 939.600 416.100 ;
        RECT 946.950 415.950 949.050 418.050 ;
        RECT 934.950 412.950 937.050 415.050 ;
        RECT 937.950 412.950 940.050 415.050 ;
        RECT 940.950 412.950 943.050 415.050 ;
        RECT 935.400 410.400 936.600 412.650 ;
        RECT 941.400 410.400 942.600 412.650 ;
        RECT 935.400 408.450 936.450 410.400 ;
        RECT 935.400 407.400 939.450 408.450 ;
        RECT 931.950 405.450 934.050 406.050 ;
        RECT 929.400 404.400 934.050 405.450 ;
        RECT 931.950 403.950 934.050 404.400 ;
        RECT 922.950 376.950 925.050 379.050 ;
        RECT 913.950 373.950 916.050 376.050 ;
        RECT 910.950 361.950 913.050 364.050 ;
        RECT 904.950 355.950 907.050 358.050 ;
        RECT 898.950 352.950 901.050 355.050 ;
        RECT 886.950 343.950 889.050 346.050 ;
        RECT 892.950 343.950 895.050 346.050 ;
        RECT 872.400 337.350 873.600 338.100 ;
        RECT 878.400 337.350 879.600 339.600 ;
        RECT 883.950 337.950 886.050 340.050 ;
        RECT 868.950 334.950 871.050 337.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 869.400 333.450 870.600 334.650 ;
        RECT 863.400 332.400 870.600 333.450 ;
        RECT 875.400 332.400 876.600 334.650 ;
        RECT 859.950 310.950 862.050 313.050 ;
        RECT 847.800 298.500 849.900 300.600 ;
        RECT 845.100 289.950 847.200 292.050 ;
        RECT 848.100 291.300 849.300 298.500 ;
        RECT 851.400 295.350 852.600 297.600 ;
        RECT 857.400 297.300 859.500 299.400 ;
        RECT 851.100 292.950 853.200 295.050 ;
        RECT 854.100 293.700 856.200 295.800 ;
        RECT 854.100 291.300 855.000 293.700 ;
        RECT 848.100 290.100 855.000 291.300 ;
        RECT 845.400 288.900 846.600 289.650 ;
        RECT 844.950 286.800 847.050 288.900 ;
        RECT 848.100 284.700 849.000 290.100 ;
        RECT 849.900 288.300 852.000 289.200 ;
        RECT 857.700 288.300 858.600 297.300 ;
        RECT 859.950 293.100 862.050 295.200 ;
        RECT 860.400 292.350 861.600 293.100 ;
        RECT 859.800 289.950 861.900 292.050 ;
        RECT 849.900 287.100 858.600 288.300 ;
        RECT 847.800 282.600 849.900 284.700 ;
        RECT 851.100 284.100 853.200 286.200 ;
        RECT 855.000 285.300 857.100 287.100 ;
        RECT 851.400 281.550 852.600 283.800 ;
        RECT 847.950 277.950 850.050 280.050 ;
        RECT 848.400 261.600 849.450 277.950 ;
        RECT 851.400 265.050 852.450 281.550 ;
        RECT 850.950 262.950 853.050 265.050 ;
        RECT 848.400 259.350 849.600 261.600 ;
        RECT 853.950 261.000 856.050 265.050 ;
        RECT 862.950 262.950 865.050 265.050 ;
        RECT 854.400 259.350 855.600 261.000 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 856.950 256.950 859.050 259.050 ;
        RECT 851.400 254.400 852.600 256.650 ;
        RECT 857.400 256.050 858.600 256.650 ;
        RECT 857.400 254.400 862.050 256.050 ;
        RECT 841.950 250.950 844.050 253.050 ;
        RECT 847.950 247.950 850.050 250.050 ;
        RECT 838.950 244.950 841.050 247.050 ;
        RECT 841.950 220.950 844.050 223.050 ;
        RECT 842.400 216.600 843.450 220.950 ;
        RECT 848.400 217.200 849.450 247.950 ;
        RECT 851.400 238.050 852.450 254.400 ;
        RECT 858.000 253.950 862.050 254.400 ;
        RECT 856.950 250.950 859.050 253.050 ;
        RECT 850.950 235.950 853.050 238.050 ;
        RECT 842.400 214.350 843.600 216.600 ;
        RECT 847.950 215.100 850.050 217.200 ;
        RECT 848.400 214.350 849.600 215.100 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 850.950 211.950 853.050 214.050 ;
        RECT 838.950 208.950 841.050 211.050 ;
        RECT 845.400 210.900 846.600 211.650 ;
        RECT 830.400 181.350 831.600 183.600 ;
        RECT 835.950 181.950 838.050 184.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 827.400 177.900 828.600 178.650 ;
        RECT 833.400 177.900 834.600 178.650 ;
        RECT 826.950 175.800 829.050 177.900 ;
        RECT 832.950 175.800 835.050 177.900 ;
        RECT 835.950 175.950 838.050 178.050 ;
        RECT 839.400 177.450 840.450 208.950 ;
        RECT 844.950 208.800 847.050 210.900 ;
        RECT 851.400 209.400 852.600 211.650 ;
        RECT 844.950 202.950 847.050 205.050 ;
        RECT 841.950 181.950 844.050 187.050 ;
        RECT 845.400 183.600 846.450 202.950 ;
        RECT 851.400 196.050 852.450 209.400 ;
        RECT 850.950 193.950 853.050 196.050 ;
        RECT 857.400 192.450 858.450 250.950 ;
        RECT 860.400 250.050 861.450 253.950 ;
        RECT 859.950 247.950 862.050 250.050 ;
        RECT 863.400 246.450 864.450 262.950 ;
        RECT 866.400 253.050 867.450 332.400 ;
        RECT 875.400 315.450 876.450 332.400 ;
        RECT 884.400 331.050 885.450 337.950 ;
        RECT 883.950 328.950 886.050 331.050 ;
        RECT 887.400 319.050 888.450 343.950 ;
        RECT 892.950 338.100 895.050 340.200 ;
        RECT 898.950 338.100 901.050 340.200 ;
        RECT 907.950 338.100 910.050 340.200 ;
        RECT 911.400 340.050 912.450 361.950 ;
        RECT 914.400 358.050 915.450 373.950 ;
        RECT 922.950 372.000 925.050 375.900 ;
        RECT 928.950 372.000 931.050 376.050 ;
        RECT 932.400 373.050 933.450 403.950 ;
        RECT 934.950 373.950 937.050 376.050 ;
        RECT 923.400 370.350 924.600 372.000 ;
        RECT 929.400 370.350 930.600 372.000 ;
        RECT 931.950 370.950 934.050 373.050 ;
        RECT 919.950 367.950 922.050 370.050 ;
        RECT 922.950 367.950 925.050 370.050 ;
        RECT 925.950 367.950 928.050 370.050 ;
        RECT 928.950 367.950 931.050 370.050 ;
        RECT 916.950 364.950 919.050 367.050 ;
        RECT 920.400 366.900 921.600 367.650 ;
        RECT 913.950 355.950 916.050 358.050 ;
        RECT 914.400 343.050 915.450 355.950 ;
        RECT 913.950 340.950 916.050 343.050 ;
        RECT 893.400 337.350 894.600 338.100 ;
        RECT 899.400 337.350 900.600 338.100 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 896.400 332.400 897.600 334.650 ;
        RECT 902.400 333.450 903.600 334.650 ;
        RECT 904.950 333.450 907.050 334.050 ;
        RECT 902.400 332.400 907.050 333.450 ;
        RECT 886.950 316.950 889.050 319.050 ;
        RECT 872.400 314.400 876.450 315.450 ;
        RECT 868.950 304.950 871.050 307.050 ;
        RECT 869.400 280.050 870.450 304.950 ;
        RECT 872.400 295.050 873.450 314.400 ;
        RECT 896.400 298.050 897.450 332.400 ;
        RECT 904.950 331.950 907.050 332.400 ;
        RECT 898.950 328.950 904.050 331.050 ;
        RECT 898.950 316.950 901.050 319.050 ;
        RECT 871.950 292.950 874.050 295.050 ;
        RECT 877.950 294.000 880.050 298.050 ;
        RECT 889.950 295.950 892.050 298.050 ;
        RECT 895.950 295.950 898.050 298.050 ;
        RECT 878.400 292.350 879.600 294.000 ;
        RECT 883.950 293.100 886.050 295.200 ;
        RECT 884.400 292.350 885.600 293.100 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 877.950 289.950 880.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 875.400 288.900 876.600 289.650 ;
        RECT 874.950 283.950 877.050 288.900 ;
        RECT 881.400 287.400 882.600 289.650 ;
        RECT 890.400 288.450 891.450 295.950 ;
        RECT 899.400 294.600 900.450 316.950 ;
        RECT 905.400 295.050 906.450 331.950 ;
        RECT 899.400 292.350 900.600 294.600 ;
        RECT 904.950 292.950 907.050 295.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 898.950 289.950 901.050 292.050 ;
        RECT 901.950 289.950 904.050 292.050 ;
        RECT 890.400 287.400 894.450 288.450 ;
        RECT 896.400 288.000 897.600 289.650 ;
        RECT 881.400 285.450 882.450 287.400 ;
        RECT 881.400 284.400 885.450 285.450 ;
        RECT 868.950 277.950 871.050 280.050 ;
        RECT 880.950 277.950 883.050 280.050 ;
        RECT 874.950 260.100 877.050 262.200 ;
        RECT 881.400 261.600 882.450 277.950 ;
        RECT 884.400 271.050 885.450 284.400 ;
        RECT 889.950 277.950 892.050 280.050 ;
        RECT 883.950 268.950 886.050 271.050 ;
        RECT 875.400 259.350 876.600 260.100 ;
        RECT 881.400 259.350 882.600 261.600 ;
        RECT 886.950 260.100 889.050 262.200 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 880.950 256.950 883.050 259.050 ;
        RECT 872.400 254.400 873.600 256.650 ;
        RECT 878.400 254.400 879.600 256.650 ;
        RECT 865.950 250.950 868.050 253.050 ;
        RECT 872.400 247.050 873.450 254.400 ;
        RECT 878.400 252.450 879.450 254.400 ;
        RECT 875.400 251.400 879.450 252.450 ;
        RECT 860.400 245.400 864.450 246.450 ;
        RECT 860.400 217.050 861.450 245.400 ;
        RECT 871.950 244.950 874.050 247.050 ;
        RECT 875.400 243.450 876.450 251.400 ;
        RECT 880.950 250.950 883.050 253.050 ;
        RECT 877.950 247.950 880.050 250.050 ;
        RECT 872.400 243.000 876.450 243.450 ;
        RECT 872.400 242.400 877.050 243.000 ;
        RECT 868.950 220.950 871.050 223.050 ;
        RECT 859.950 214.950 862.050 217.050 ;
        RECT 862.950 215.100 865.050 217.200 ;
        RECT 869.400 216.600 870.450 220.950 ;
        RECT 872.400 220.050 873.450 242.400 ;
        RECT 874.950 238.950 877.050 242.400 ;
        RECT 874.950 232.950 877.050 235.050 ;
        RECT 871.950 217.950 874.050 220.050 ;
        RECT 875.400 217.050 876.450 232.950 ;
        RECT 863.400 214.350 864.600 215.100 ;
        RECT 869.400 214.350 870.600 216.600 ;
        RECT 874.950 214.950 877.050 217.050 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 859.950 205.950 862.050 211.050 ;
        RECT 866.400 210.900 867.600 211.650 ;
        RECT 872.400 210.900 873.600 211.650 ;
        RECT 878.400 211.050 879.450 247.950 ;
        RECT 865.950 208.800 868.050 210.900 ;
        RECT 871.950 208.800 874.050 210.900 ;
        RECT 874.950 208.950 877.050 211.050 ;
        RECT 877.950 208.950 880.050 211.050 ;
        RECT 881.400 210.450 882.450 250.950 ;
        RECT 887.400 250.050 888.450 260.100 ;
        RECT 883.950 247.950 886.050 250.050 ;
        RECT 886.950 247.950 889.050 250.050 ;
        RECT 884.400 235.050 885.450 247.950 ;
        RECT 886.950 244.800 889.050 246.900 ;
        RECT 883.950 232.950 886.050 235.050 ;
        RECT 883.950 226.950 886.050 229.050 ;
        RECT 884.400 217.050 885.450 226.950 ;
        RECT 883.950 214.950 886.050 217.050 ;
        RECT 887.400 216.600 888.450 244.800 ;
        RECT 890.400 220.050 891.450 277.950 ;
        RECT 893.400 262.050 894.450 287.400 ;
        RECT 895.950 283.950 898.050 288.000 ;
        RECT 902.400 287.400 903.600 289.650 ;
        RECT 902.400 280.050 903.450 287.400 ;
        RECT 904.950 286.950 907.050 289.050 ;
        RECT 901.950 277.950 904.050 280.050 ;
        RECT 905.400 265.050 906.450 286.950 ;
        RECT 908.400 271.050 909.450 338.100 ;
        RECT 910.950 337.950 913.050 340.050 ;
        RECT 917.400 339.600 918.450 364.950 ;
        RECT 919.950 364.800 922.050 366.900 ;
        RECT 926.400 366.000 927.600 367.650 ;
        RECT 925.950 364.050 928.050 366.000 ;
        RECT 925.800 363.000 928.050 364.050 ;
        RECT 925.800 361.950 927.900 363.000 ;
        RECT 928.950 361.950 931.050 364.050 ;
        RECT 925.950 340.950 928.050 343.050 ;
        RECT 917.400 337.350 918.600 339.600 ;
        RECT 913.950 334.950 916.050 337.050 ;
        RECT 916.950 334.950 919.050 337.050 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 910.950 331.950 913.050 334.050 ;
        RECT 914.400 333.000 915.600 334.650 ;
        RECT 911.400 310.050 912.450 331.950 ;
        RECT 913.950 328.950 916.050 333.000 ;
        RECT 920.400 332.400 921.600 334.650 ;
        RECT 916.950 328.950 919.050 331.050 ;
        RECT 913.950 310.950 916.050 313.050 ;
        RECT 910.950 307.950 913.050 310.050 ;
        RECT 910.950 298.950 913.050 301.050 ;
        RECT 911.400 295.050 912.450 298.950 ;
        RECT 914.400 298.050 915.450 310.950 ;
        RECT 917.400 301.050 918.450 328.950 ;
        RECT 916.950 298.950 919.050 301.050 ;
        RECT 920.400 298.200 921.450 332.400 ;
        RECT 922.950 328.950 925.050 334.050 ;
        RECT 922.950 304.950 925.050 307.050 ;
        RECT 910.950 292.950 913.050 295.050 ;
        RECT 913.950 294.000 916.050 298.050 ;
        RECT 919.950 296.100 922.050 298.200 ;
        RECT 923.400 298.050 924.450 304.950 ;
        RECT 922.950 295.950 925.050 298.050 ;
        RECT 926.400 295.200 927.450 340.950 ;
        RECT 914.400 292.350 915.600 294.000 ;
        RECT 919.950 292.950 922.050 295.050 ;
        RECT 925.950 293.100 928.050 295.200 ;
        RECT 920.400 292.350 921.600 292.950 ;
        RECT 913.950 289.950 916.050 292.050 ;
        RECT 916.950 289.950 919.050 292.050 ;
        RECT 919.950 289.950 922.050 292.050 ;
        RECT 922.950 289.950 925.050 292.050 ;
        RECT 910.950 286.950 913.050 289.050 ;
        RECT 917.400 288.900 918.600 289.650 ;
        RECT 923.400 288.900 924.600 289.650 ;
        RECT 907.950 268.950 910.050 271.050 ;
        RECT 904.950 262.950 907.050 265.050 ;
        RECT 892.950 259.950 895.050 262.050 ;
        RECT 898.950 260.100 901.050 262.200 ;
        RECT 905.400 261.600 906.450 262.950 ;
        RECT 911.400 262.050 912.450 286.950 ;
        RECT 916.950 286.800 919.050 288.900 ;
        RECT 922.950 286.800 925.050 288.900 ;
        RECT 925.950 286.950 928.050 289.050 ;
        RECT 916.950 277.950 919.050 280.050 ;
        RECT 913.950 262.950 916.050 265.050 ;
        RECT 899.400 259.350 900.600 260.100 ;
        RECT 905.400 259.350 906.600 261.600 ;
        RECT 910.950 259.950 913.050 262.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 901.950 256.950 904.050 259.050 ;
        RECT 904.950 256.950 907.050 259.050 ;
        RECT 910.950 256.800 913.050 258.900 ;
        RECT 892.950 253.950 895.050 256.050 ;
        RECT 896.400 254.400 897.600 256.650 ;
        RECT 902.400 254.400 903.600 256.650 ;
        RECT 893.400 247.050 894.450 253.950 ;
        RECT 896.400 250.050 897.450 254.400 ;
        RECT 902.400 252.450 903.450 254.400 ;
        RECT 907.950 253.950 910.050 256.050 ;
        RECT 899.400 251.400 903.450 252.450 ;
        RECT 895.950 247.950 898.050 250.050 ;
        RECT 892.950 244.950 895.050 247.050 ;
        RECT 899.400 241.050 900.450 251.400 ;
        RECT 901.950 249.450 906.000 250.050 ;
        RECT 901.950 247.950 906.450 249.450 ;
        RECT 901.950 244.800 904.050 246.900 ;
        RECT 898.950 238.950 901.050 241.050 ;
        RECT 902.400 234.450 903.450 244.800 ;
        RECT 905.400 238.050 906.450 247.950 ;
        RECT 904.950 235.950 907.050 238.050 ;
        RECT 902.400 233.400 906.450 234.450 ;
        RECT 897.000 231.450 901.050 232.050 ;
        RECT 896.400 231.000 901.050 231.450 ;
        RECT 895.950 229.950 901.050 231.000 ;
        RECT 895.950 226.950 898.050 229.950 ;
        RECT 898.950 223.950 901.050 226.050 ;
        RECT 889.950 217.950 892.050 220.050 ;
        RECT 887.400 214.350 888.600 216.600 ;
        RECT 892.950 215.100 895.050 217.200 ;
        RECT 899.400 217.050 900.450 223.950 ;
        RECT 901.950 217.950 904.050 220.050 ;
        RECT 893.400 214.350 894.600 215.100 ;
        RECT 898.950 214.950 901.050 217.050 ;
        RECT 886.950 211.950 889.050 214.050 ;
        RECT 889.950 211.950 892.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 895.950 211.950 898.050 214.050 ;
        RECT 881.400 209.400 885.450 210.450 ;
        RECT 862.950 199.950 865.050 202.050 ;
        RECT 857.400 191.400 861.450 192.450 ;
        RECT 850.950 187.950 853.050 190.050 ;
        RECT 851.400 183.600 852.450 187.950 ;
        RECT 845.400 181.350 846.600 183.600 ;
        RECT 851.400 181.350 852.600 183.600 ;
        RECT 844.950 178.950 847.050 181.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 839.400 176.400 843.450 177.450 ;
        RECT 833.400 169.050 834.450 175.800 ;
        RECT 836.400 172.050 837.450 175.950 ;
        RECT 835.950 169.950 838.050 172.050 ;
        RECT 832.950 166.950 835.050 169.050 ;
        RECT 814.950 151.950 817.050 154.050 ;
        RECT 820.950 151.950 823.050 154.050 ;
        RECT 826.950 151.950 829.050 154.050 ;
        RECT 829.950 151.950 832.050 154.050 ;
        RECT 808.950 148.950 811.050 151.050 ;
        RECT 805.950 142.950 808.050 145.050 ;
        RECT 809.400 138.600 810.450 148.950 ;
        RECT 814.950 145.950 817.050 148.050 ;
        RECT 815.400 138.600 816.450 145.950 ;
        RECT 823.950 139.950 826.050 142.050 ;
        RECT 809.400 136.350 810.600 138.600 ;
        RECT 815.400 136.350 816.600 138.600 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 812.400 132.900 813.600 133.650 ;
        RECT 818.400 132.900 819.600 133.650 ;
        RECT 824.400 133.050 825.450 139.950 ;
        RECT 811.950 130.800 814.050 132.900 ;
        RECT 817.950 130.800 820.050 132.900 ;
        RECT 823.950 130.950 826.050 133.050 ;
        RECT 812.400 124.050 813.450 130.800 ;
        RECT 820.950 124.950 823.050 127.050 ;
        RECT 805.950 121.950 808.050 124.050 ;
        RECT 811.950 121.950 814.050 124.050 ;
        RECT 806.400 112.050 807.450 121.950 ;
        RECT 808.950 115.950 811.050 118.050 ;
        RECT 805.950 109.950 808.050 112.050 ;
        RECT 802.950 106.950 805.050 109.050 ;
        RECT 751.950 97.800 754.050 99.900 ;
        RECT 757.950 97.800 760.050 99.900 ;
        RECT 763.950 97.800 766.050 99.900 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 764.400 88.050 765.450 97.800 ;
        RECT 767.400 94.050 768.450 103.950 ;
        RECT 776.400 103.350 777.600 104.100 ;
        RECT 781.950 103.950 784.050 106.050 ;
        RECT 784.950 104.100 787.050 106.200 ;
        RECT 787.950 103.950 790.050 106.050 ;
        RECT 793.950 104.100 796.050 106.200 ;
        RECT 799.950 104.100 802.050 106.200 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 773.400 100.050 774.600 100.650 ;
        RECT 769.950 98.400 774.600 100.050 ;
        RECT 779.400 98.400 780.600 100.650 ;
        RECT 769.950 97.950 774.000 98.400 ;
        RECT 769.950 94.800 772.050 96.900 ;
        RECT 766.950 91.950 769.050 94.050 ;
        RECT 739.950 87.450 742.050 88.050 ;
        RECT 739.950 86.400 744.450 87.450 ;
        RECT 739.950 85.950 742.050 86.400 ;
        RECT 731.400 62.400 735.450 63.450 ;
        RECT 731.400 60.600 732.450 62.400 ;
        RECT 731.400 58.350 732.600 60.600 ;
        RECT 736.950 59.100 739.050 61.200 ;
        RECT 737.400 58.350 738.600 59.100 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 721.950 52.800 724.050 54.900 ;
        RECT 728.400 53.400 729.600 55.650 ;
        RECT 734.400 54.900 735.600 55.650 ;
        RECT 743.400 54.900 744.450 86.400 ;
        RECT 763.950 85.950 766.050 88.050 ;
        RECT 770.400 67.050 771.450 94.800 ;
        RECT 779.400 88.050 780.450 98.400 ;
        RECT 788.400 88.050 789.450 103.950 ;
        RECT 794.400 103.350 795.600 104.100 ;
        RECT 800.400 103.350 801.600 104.100 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 797.400 99.900 798.600 100.650 ;
        RECT 796.950 97.800 799.050 99.900 ;
        RECT 803.400 98.400 804.600 100.650 ;
        RECT 778.950 85.950 781.050 88.050 ;
        RECT 787.950 85.950 790.050 88.050 ;
        RECT 797.400 85.050 798.450 97.800 ;
        RECT 799.950 94.950 802.050 97.050 ;
        RECT 796.950 82.950 799.050 85.050 ;
        RECT 769.950 64.950 772.050 67.050 ;
        RECT 748.950 59.100 751.050 61.200 ;
        RECT 757.950 59.100 760.050 61.200 ;
        RECT 763.950 59.100 766.050 61.200 ;
        RECT 770.400 60.600 771.450 64.950 ;
        RECT 749.400 58.350 750.600 59.100 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 752.400 54.900 753.600 55.650 ;
        RECT 728.400 49.050 729.450 53.400 ;
        RECT 733.950 52.800 736.050 54.900 ;
        RECT 742.950 52.800 745.050 54.900 ;
        RECT 751.950 52.800 754.050 54.900 ;
        RECT 727.950 46.950 730.050 49.050 ;
        RECT 758.400 46.050 759.450 59.100 ;
        RECT 764.400 58.350 765.600 59.100 ;
        RECT 770.400 58.350 771.600 60.600 ;
        RECT 784.950 59.100 787.050 61.200 ;
        RECT 790.950 60.000 793.050 64.050 ;
        RECT 785.400 58.350 786.600 59.100 ;
        RECT 791.400 58.350 792.600 60.000 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 769.950 55.950 772.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 767.400 53.400 768.600 55.650 ;
        RECT 782.400 53.400 783.600 55.650 ;
        RECT 788.400 54.900 789.600 55.650 ;
        RECT 800.400 54.900 801.450 94.950 ;
        RECT 803.400 88.050 804.450 98.400 ;
        RECT 802.950 85.950 805.050 88.050 ;
        RECT 809.400 63.450 810.450 115.950 ;
        RECT 821.400 109.050 822.450 124.950 ;
        RECT 811.950 106.950 814.050 109.050 ;
        RECT 812.400 64.050 813.450 106.950 ;
        RECT 820.950 105.000 823.050 109.050 ;
        RECT 827.400 106.200 828.450 151.950 ;
        RECT 830.400 139.050 831.450 151.950 ;
        RECT 832.950 148.950 835.050 151.050 ;
        RECT 829.950 136.950 832.050 139.050 ;
        RECT 833.400 138.600 834.450 148.950 ;
        RECT 838.950 145.950 841.050 148.050 ;
        RECT 839.400 138.600 840.450 145.950 ;
        RECT 842.400 145.050 843.450 176.400 ;
        RECT 848.400 176.400 849.600 178.650 ;
        RECT 854.400 177.450 855.600 178.650 ;
        RECT 854.400 176.400 858.450 177.450 ;
        RECT 848.400 157.050 849.450 176.400 ;
        RECT 853.950 172.950 856.050 175.050 ;
        RECT 847.950 154.950 850.050 157.050 ;
        RECT 841.950 142.950 844.050 145.050 ;
        RECT 847.950 142.950 850.050 145.050 ;
        RECT 833.400 136.350 834.600 138.600 ;
        RECT 839.400 136.350 840.600 138.600 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 836.400 131.400 837.600 133.650 ;
        RECT 842.400 133.050 843.600 133.650 ;
        RECT 842.400 131.400 847.050 133.050 ;
        RECT 836.400 124.050 837.450 131.400 ;
        RECT 843.000 130.950 847.050 131.400 ;
        RECT 841.950 127.950 844.050 130.050 ;
        RECT 835.950 121.950 838.050 124.050 ;
        RECT 832.950 115.950 835.050 118.050 ;
        RECT 829.950 112.950 832.050 115.050 ;
        RECT 821.400 103.350 822.600 105.000 ;
        RECT 826.950 104.100 829.050 106.200 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 818.400 99.900 819.600 100.650 ;
        RECT 817.950 97.800 820.050 99.900 ;
        RECT 824.400 99.450 825.600 100.650 ;
        RECT 830.400 99.900 831.450 112.950 ;
        RECT 833.400 106.050 834.450 115.950 ;
        RECT 842.400 112.050 843.450 127.950 ;
        RECT 844.950 121.950 847.050 124.050 ;
        RECT 841.950 109.950 844.050 112.050 ;
        RECT 832.950 103.950 835.050 106.050 ;
        RECT 838.950 104.100 841.050 106.200 ;
        RECT 845.400 105.600 846.450 121.950 ;
        RECT 848.400 118.050 849.450 142.950 ;
        RECT 850.950 139.950 853.050 142.050 ;
        RECT 847.950 115.950 850.050 118.050 ;
        RECT 851.400 106.050 852.450 139.950 ;
        RECT 854.400 139.050 855.450 172.950 ;
        RECT 857.400 169.050 858.450 176.400 ;
        RECT 860.400 175.050 861.450 191.400 ;
        RECT 859.950 172.950 862.050 175.050 ;
        RECT 856.950 166.950 859.050 169.050 ;
        RECT 863.400 163.050 864.450 199.950 ;
        RECT 866.400 193.050 867.450 208.800 ;
        RECT 872.400 193.050 873.450 208.800 ;
        RECT 875.400 199.050 876.450 208.950 ;
        RECT 877.950 199.950 880.050 205.050 ;
        RECT 874.950 196.950 877.050 199.050 ;
        RECT 865.950 190.950 868.050 193.050 ;
        RECT 871.950 190.950 874.050 193.050 ;
        RECT 874.950 187.950 877.050 190.050 ;
        RECT 865.950 183.600 870.000 184.050 ;
        RECT 875.400 183.600 876.450 187.950 ;
        RECT 865.950 181.950 870.600 183.600 ;
        RECT 869.400 181.350 870.600 181.950 ;
        RECT 875.400 181.350 876.600 183.600 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 865.950 175.950 868.050 178.050 ;
        RECT 872.400 177.900 873.600 178.650 ;
        RECT 878.400 177.900 879.600 178.650 ;
        RECT 866.400 169.050 867.450 175.950 ;
        RECT 871.950 175.800 874.050 177.900 ;
        RECT 877.950 175.800 880.050 177.900 ;
        RECT 884.400 175.050 885.450 209.400 ;
        RECT 890.400 209.400 891.600 211.650 ;
        RECT 896.400 209.400 897.600 211.650 ;
        RECT 886.950 205.950 889.050 208.050 ;
        RECT 887.400 184.050 888.450 205.950 ;
        RECT 890.400 193.050 891.450 209.400 ;
        RECT 892.950 205.950 895.050 208.050 ;
        RECT 889.950 190.950 892.050 193.050 ;
        RECT 893.400 190.050 894.450 205.950 ;
        RECT 896.400 205.050 897.450 209.400 ;
        RECT 895.950 202.950 898.050 205.050 ;
        RECT 895.950 196.950 898.050 199.050 ;
        RECT 892.950 187.950 895.050 190.050 ;
        RECT 896.400 186.450 897.450 196.950 ;
        RECT 898.950 193.950 901.050 196.050 ;
        RECT 893.400 185.400 897.450 186.450 ;
        RECT 886.950 181.950 889.050 184.050 ;
        RECT 893.400 183.600 894.450 185.400 ;
        RECT 899.400 184.200 900.450 193.950 ;
        RECT 893.400 181.350 894.600 183.600 ;
        RECT 898.950 182.100 901.050 184.200 ;
        RECT 902.400 183.450 903.450 217.950 ;
        RECT 905.400 217.050 906.450 233.400 ;
        RECT 908.400 226.050 909.450 253.950 ;
        RECT 911.400 250.050 912.450 256.800 ;
        RECT 910.950 247.950 913.050 250.050 ;
        RECT 910.950 235.950 913.050 238.050 ;
        RECT 907.950 223.950 910.050 226.050 ;
        RECT 904.950 214.950 907.050 217.050 ;
        RECT 911.400 216.600 912.450 235.950 ;
        RECT 914.400 220.050 915.450 262.950 ;
        RECT 917.400 262.050 918.450 277.950 ;
        RECT 926.400 274.050 927.450 286.950 ;
        RECT 929.400 280.050 930.450 361.950 ;
        RECT 935.400 351.450 936.450 373.950 ;
        RECT 938.400 361.050 939.450 407.400 ;
        RECT 941.400 406.050 942.450 410.400 ;
        RECT 943.950 406.950 946.050 409.050 ;
        RECT 940.950 403.950 943.050 406.050 ;
        RECT 940.950 376.950 943.050 379.050 ;
        RECT 937.950 358.950 940.050 361.050 ;
        RECT 932.400 350.400 936.450 351.450 ;
        RECT 932.400 340.050 933.450 350.400 ;
        RECT 941.400 343.050 942.450 376.950 ;
        RECT 944.400 364.050 945.450 406.950 ;
        RECT 943.950 361.950 946.050 364.050 ;
        RECT 943.950 358.800 946.050 360.900 ;
        RECT 940.950 340.950 943.050 343.050 ;
        RECT 931.950 337.950 934.050 340.050 ;
        RECT 937.950 338.100 940.050 340.200 ;
        RECT 944.400 339.600 945.450 358.800 ;
        RECT 947.400 340.050 948.450 415.950 ;
        RECT 938.400 337.350 939.600 338.100 ;
        RECT 944.400 337.350 945.600 339.600 ;
        RECT 946.950 337.950 949.050 340.050 ;
        RECT 934.950 334.950 937.050 337.050 ;
        RECT 937.950 334.950 940.050 337.050 ;
        RECT 940.950 334.950 943.050 337.050 ;
        RECT 943.950 334.950 946.050 337.050 ;
        RECT 935.400 332.400 936.600 334.650 ;
        RECT 941.400 332.400 942.600 334.650 ;
        RECT 935.400 313.050 936.450 332.400 ;
        RECT 937.950 328.950 940.050 331.050 ;
        RECT 941.400 330.450 942.450 332.400 ;
        RECT 946.950 331.950 949.050 334.050 ;
        RECT 941.400 329.400 945.450 330.450 ;
        RECT 934.950 310.950 937.050 313.050 ;
        RECT 938.400 298.050 939.450 328.950 ;
        RECT 940.950 307.950 943.050 310.050 ;
        RECT 937.950 295.950 940.050 298.050 ;
        RECT 934.950 293.100 937.050 295.200 ;
        RECT 941.400 294.600 942.450 307.950 ;
        RECT 944.400 295.050 945.450 329.400 ;
        RECT 935.400 292.350 936.600 293.100 ;
        RECT 941.400 292.350 942.600 294.600 ;
        RECT 943.950 292.950 946.050 295.050 ;
        RECT 934.950 289.950 937.050 292.050 ;
        RECT 937.950 289.950 940.050 292.050 ;
        RECT 940.950 289.950 943.050 292.050 ;
        RECT 938.400 288.900 939.600 289.650 ;
        RECT 931.950 286.800 934.050 288.900 ;
        RECT 937.950 286.800 940.050 288.900 ;
        RECT 928.950 277.950 931.050 280.050 ;
        RECT 925.950 271.950 928.050 274.050 ;
        RECT 919.950 268.950 922.050 271.050 ;
        RECT 916.950 259.950 919.050 262.050 ;
        RECT 920.400 261.600 921.450 268.950 ;
        RECT 920.400 259.350 921.600 261.600 ;
        RECT 925.950 260.100 928.050 262.200 ;
        RECT 932.400 262.050 933.450 286.800 ;
        RECT 943.950 283.950 946.050 286.050 ;
        RECT 934.950 271.950 937.050 274.050 ;
        RECT 926.400 259.350 927.600 260.100 ;
        RECT 931.950 259.950 934.050 262.050 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 922.950 256.950 925.050 259.050 ;
        RECT 925.950 256.950 928.050 259.050 ;
        RECT 928.950 256.950 931.050 259.050 ;
        RECT 916.950 250.950 919.050 256.050 ;
        RECT 923.400 254.400 924.600 256.650 ;
        RECT 929.400 255.900 930.600 256.650 ;
        RECT 916.950 229.950 919.050 232.050 ;
        RECT 913.950 217.950 916.050 220.050 ;
        RECT 917.400 216.600 918.450 229.950 ;
        RECT 923.400 223.050 924.450 254.400 ;
        RECT 928.950 253.800 931.050 255.900 ;
        RECT 931.950 253.950 934.050 256.050 ;
        RECT 925.950 250.950 928.050 253.050 ;
        RECT 922.950 220.950 925.050 223.050 ;
        RECT 922.950 217.800 925.050 219.900 ;
        RECT 911.400 214.350 912.600 216.600 ;
        RECT 917.400 214.350 918.600 216.600 ;
        RECT 907.950 211.950 910.050 214.050 ;
        RECT 910.950 211.950 913.050 214.050 ;
        RECT 913.950 211.950 916.050 214.050 ;
        RECT 916.950 211.950 919.050 214.050 ;
        RECT 904.950 208.950 907.050 211.050 ;
        RECT 908.400 210.900 909.600 211.650 ;
        RECT 914.400 210.900 915.600 211.650 ;
        RECT 923.400 210.900 924.450 217.800 ;
        RECT 905.400 187.050 906.450 208.950 ;
        RECT 907.950 208.800 910.050 210.900 ;
        RECT 913.950 208.800 916.050 210.900 ;
        RECT 922.950 208.800 925.050 210.900 ;
        RECT 918.000 207.600 922.050 208.050 ;
        RECT 917.400 205.950 922.050 207.600 ;
        RECT 907.950 202.950 910.050 205.050 ;
        RECT 908.400 199.050 909.450 202.950 ;
        RECT 917.400 199.050 918.450 205.950 ;
        RECT 919.950 202.800 922.050 204.900 ;
        RECT 908.400 197.400 913.050 199.050 ;
        RECT 909.000 196.950 913.050 197.400 ;
        RECT 916.950 196.950 919.050 199.050 ;
        RECT 917.400 193.050 918.450 196.950 ;
        RECT 916.950 190.950 919.050 193.050 ;
        RECT 920.400 189.450 921.450 202.800 ;
        RECT 923.400 202.050 924.450 208.800 ;
        RECT 922.950 199.950 925.050 202.050 ;
        RECT 926.400 198.450 927.450 250.950 ;
        RECT 928.950 247.950 931.050 250.050 ;
        RECT 929.400 217.050 930.450 247.950 ;
        RECT 928.950 214.950 931.050 217.050 ;
        RECT 932.400 216.600 933.450 253.950 ;
        RECT 935.400 247.050 936.450 271.950 ;
        RECT 937.950 265.950 940.050 268.050 ;
        RECT 938.400 262.050 939.450 265.950 ;
        RECT 944.400 265.050 945.450 283.950 ;
        RECT 947.400 268.050 948.450 331.950 ;
        RECT 946.950 265.950 949.050 268.050 ;
        RECT 943.950 262.950 946.050 265.050 ;
        RECT 937.950 259.950 940.050 262.050 ;
        RECT 945.000 261.600 949.050 262.050 ;
        RECT 944.400 259.950 949.050 261.600 ;
        RECT 944.400 259.350 945.600 259.950 ;
        RECT 940.950 256.950 943.050 259.050 ;
        RECT 943.950 256.950 946.050 259.050 ;
        RECT 937.950 253.950 940.050 256.050 ;
        RECT 941.400 255.900 942.600 256.650 ;
        RECT 934.950 244.950 937.050 247.050 ;
        RECT 934.950 235.950 937.050 238.050 ;
        RECT 935.400 219.450 936.450 235.950 ;
        RECT 938.400 223.050 939.450 253.950 ;
        RECT 940.950 253.800 943.050 255.900 ;
        RECT 946.950 253.950 949.050 256.050 ;
        RECT 943.950 247.950 946.050 250.050 ;
        RECT 944.400 232.050 945.450 247.950 ;
        RECT 943.950 229.950 946.050 232.050 ;
        RECT 937.950 220.950 940.050 223.050 ;
        RECT 943.950 220.950 946.050 223.050 ;
        RECT 935.400 218.400 939.450 219.450 ;
        RECT 938.400 216.600 939.450 218.400 ;
        RECT 944.400 217.050 945.450 220.950 ;
        RECT 932.400 214.350 933.600 216.600 ;
        RECT 938.400 214.350 939.600 216.600 ;
        RECT 943.950 214.950 946.050 217.050 ;
        RECT 931.950 211.950 934.050 214.050 ;
        RECT 934.950 211.950 937.050 214.050 ;
        RECT 937.950 211.950 940.050 214.050 ;
        RECT 940.950 211.950 943.050 214.050 ;
        RECT 928.950 208.950 931.050 211.050 ;
        RECT 935.400 209.400 936.600 211.650 ;
        RECT 941.400 209.400 942.600 211.650 ;
        RECT 929.400 205.050 930.450 208.950 ;
        RECT 928.950 202.950 931.050 205.050 ;
        RECT 935.400 202.050 936.450 209.400 ;
        RECT 937.950 202.950 940.050 205.050 ;
        RECT 934.950 199.950 937.050 202.050 ;
        RECT 917.400 188.400 921.450 189.450 ;
        RECT 923.400 197.400 927.450 198.450 ;
        RECT 904.950 184.950 907.050 187.050 ;
        RECT 902.400 182.400 906.450 183.450 ;
        RECT 899.400 181.350 900.600 182.100 ;
        RECT 889.950 178.950 892.050 181.050 ;
        RECT 892.950 178.950 895.050 181.050 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 886.950 175.950 889.050 178.050 ;
        RECT 890.400 176.400 891.600 178.650 ;
        RECT 896.400 176.400 897.600 178.650 ;
        RECT 871.950 172.650 874.050 174.750 ;
        RECT 883.950 172.950 886.050 175.050 ;
        RECT 865.950 166.950 868.050 169.050 ;
        RECT 862.950 160.950 865.050 163.050 ;
        RECT 853.950 136.950 856.050 139.050 ;
        RECT 859.950 138.000 862.050 142.050 ;
        RECT 865.950 138.000 868.050 142.050 ;
        RECT 860.400 136.350 861.600 138.000 ;
        RECT 866.400 136.350 867.600 138.000 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 853.950 130.950 856.050 133.050 ;
        RECT 857.400 131.400 858.600 133.650 ;
        RECT 863.400 132.000 864.600 133.650 ;
        RECT 839.400 103.350 840.600 104.100 ;
        RECT 845.400 103.350 846.600 105.600 ;
        RECT 850.950 103.950 853.050 106.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 829.950 99.450 832.050 99.900 ;
        RECT 824.400 98.400 832.050 99.450 ;
        RECT 829.950 97.800 832.050 98.400 ;
        RECT 820.950 94.950 823.050 97.050 ;
        RECT 832.950 94.950 835.050 100.050 ;
        RECT 836.400 99.900 837.600 100.650 ;
        RECT 835.950 97.800 838.050 99.900 ;
        RECT 842.400 98.400 843.600 100.650 ;
        RECT 848.400 99.000 849.600 100.650 ;
        RECT 806.400 62.400 810.450 63.450 ;
        RECT 806.400 61.200 807.450 62.400 ;
        RECT 811.950 61.950 814.050 64.050 ;
        RECT 805.950 59.100 808.050 61.200 ;
        RECT 812.400 60.600 813.450 61.950 ;
        RECT 806.400 58.350 807.600 59.100 ;
        RECT 812.400 58.350 813.600 60.600 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 811.950 55.950 814.050 58.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 767.400 49.050 768.450 53.400 ;
        RECT 766.950 46.950 769.050 49.050 ;
        RECT 757.800 43.950 759.900 46.050 ;
        RECT 760.950 43.950 763.050 46.050 ;
        RECT 721.950 37.950 724.050 40.050 ;
        RECT 694.950 31.950 697.050 34.050 ;
        RECT 706.950 31.950 709.050 34.050 ;
        RECT 718.950 31.950 721.050 34.050 ;
        RECT 695.400 27.600 696.450 31.950 ;
        RECT 707.400 27.600 708.450 31.950 ;
        RECT 689.400 25.350 690.600 27.600 ;
        RECT 695.400 25.350 696.600 27.600 ;
        RECT 707.400 25.350 708.600 27.600 ;
        RECT 712.950 26.100 715.050 28.200 ;
        RECT 713.400 25.350 714.600 26.100 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 715.950 22.950 718.050 25.050 ;
        RECT 686.400 21.900 687.600 22.650 ;
        RECT 679.950 19.800 682.050 21.900 ;
        RECT 685.950 19.800 688.050 21.900 ;
        RECT 692.400 20.400 693.600 22.650 ;
        RECT 710.400 20.400 711.600 22.650 ;
        RECT 716.400 21.000 717.600 22.650 ;
        RECT 686.400 16.050 687.450 19.800 ;
        RECT 692.400 16.050 693.450 20.400 ;
        RECT 710.400 16.050 711.450 20.400 ;
        RECT 715.950 16.950 718.050 21.000 ;
        RECT 722.400 16.050 723.450 37.950 ;
        RECT 736.950 34.950 739.050 37.050 ;
        RECT 754.950 34.950 757.050 37.050 ;
        RECT 724.950 25.950 727.050 28.050 ;
        RECT 730.950 26.100 733.050 28.200 ;
        RECT 737.400 27.600 738.450 34.950 ;
        RECT 755.400 27.600 756.450 34.950 ;
        RECT 761.400 27.600 762.450 43.950 ;
        RECT 775.950 34.950 778.050 37.050 ;
        RECT 685.950 13.950 688.050 16.050 ;
        RECT 691.950 13.950 694.050 16.050 ;
        RECT 709.950 13.950 712.050 16.050 ;
        RECT 721.950 13.950 724.050 16.050 ;
        RECT 667.950 10.950 670.050 13.050 ;
        RECT 676.950 10.950 679.050 13.050 ;
        RECT 613.950 7.950 616.050 10.050 ;
        RECT 725.400 7.050 726.450 25.950 ;
        RECT 731.400 25.350 732.600 26.100 ;
        RECT 737.400 25.350 738.600 27.600 ;
        RECT 755.400 25.350 756.600 27.600 ;
        RECT 761.400 25.350 762.600 27.600 ;
        RECT 766.950 25.950 769.050 28.050 ;
        RECT 776.400 27.600 777.450 34.950 ;
        RECT 782.400 31.050 783.450 53.400 ;
        RECT 787.950 52.800 790.050 54.900 ;
        RECT 799.950 54.450 802.050 54.900 ;
        RECT 797.400 54.000 802.050 54.450 ;
        RECT 809.400 54.000 810.600 55.650 ;
        RECT 796.950 53.400 802.050 54.000 ;
        RECT 796.950 49.950 799.050 53.400 ;
        RECT 799.950 52.800 802.050 53.400 ;
        RECT 805.950 49.950 808.050 52.050 ;
        RECT 808.950 49.950 811.050 54.000 ;
        RECT 815.400 53.400 816.600 55.650 ;
        RECT 821.400 55.050 822.450 94.950 ;
        RECT 842.400 79.050 843.450 98.400 ;
        RECT 847.950 94.950 850.050 99.000 ;
        RECT 854.400 97.050 855.450 130.950 ;
        RECT 857.400 127.050 858.450 131.400 ;
        RECT 862.950 127.950 865.050 132.000 ;
        RECT 872.400 129.450 873.450 172.650 ;
        RECT 874.950 157.950 877.050 160.050 ;
        RECT 875.400 132.450 876.450 157.950 ;
        RECT 883.950 154.950 886.050 157.050 ;
        RECT 877.950 142.950 880.050 145.050 ;
        RECT 878.400 139.050 879.450 142.950 ;
        RECT 877.950 136.950 880.050 139.050 ;
        RECT 884.400 138.600 885.450 154.950 ;
        RECT 887.400 145.050 888.450 175.950 ;
        RECT 890.400 175.050 891.450 176.400 ;
        RECT 889.950 172.950 892.050 175.050 ;
        RECT 886.950 142.950 889.050 145.050 ;
        RECT 890.400 144.450 891.450 172.950 ;
        RECT 896.400 169.050 897.450 176.400 ;
        RECT 905.400 175.050 906.450 182.400 ;
        RECT 910.950 182.100 913.050 184.200 ;
        RECT 917.400 183.600 918.450 188.400 ;
        RECT 923.400 184.050 924.450 197.400 ;
        RECT 931.950 190.950 934.050 193.050 ;
        RECT 925.800 187.950 927.900 190.050 ;
        RECT 928.950 187.950 931.050 190.050 ;
        RECT 911.400 181.350 912.600 182.100 ;
        RECT 917.400 181.350 918.600 183.600 ;
        RECT 922.950 181.950 925.050 184.050 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 913.950 178.950 916.050 181.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 907.950 175.950 910.050 178.050 ;
        RECT 914.400 176.400 915.600 178.650 ;
        RECT 920.400 176.400 921.600 178.650 ;
        RECT 904.950 172.950 907.050 175.050 ;
        RECT 895.950 166.950 898.050 169.050 ;
        RECT 898.950 151.950 901.050 154.050 ;
        RECT 890.400 143.400 894.450 144.450 ;
        RECT 884.400 136.350 885.600 138.600 ;
        RECT 889.950 137.100 892.050 139.200 ;
        RECT 893.400 139.050 894.450 143.400 ;
        RECT 890.400 136.350 891.600 137.100 ;
        RECT 892.950 136.950 895.050 139.050 ;
        RECT 895.950 137.100 898.050 139.200 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 881.400 132.450 882.600 133.650 ;
        RECT 875.400 131.400 882.600 132.450 ;
        RECT 887.400 131.400 888.600 133.650 ;
        RECT 872.400 128.400 876.450 129.450 ;
        RECT 856.950 124.950 859.050 127.050 ;
        RECT 856.950 103.950 859.050 106.050 ;
        RECT 868.950 104.100 871.050 106.200 ;
        RECT 857.400 97.050 858.450 103.950 ;
        RECT 869.400 103.350 870.600 104.100 ;
        RECT 859.950 99.450 862.050 103.050 ;
        RECT 863.100 100.950 865.200 103.050 ;
        RECT 868.500 100.950 870.600 103.050 ;
        RECT 871.800 100.950 873.900 103.050 ;
        RECT 863.400 99.450 864.600 100.650 ;
        RECT 872.400 99.900 873.600 100.650 ;
        RECT 859.950 99.000 864.600 99.450 ;
        RECT 860.400 98.400 864.600 99.000 ;
        RECT 871.950 97.800 874.050 99.900 ;
        RECT 853.950 94.950 856.050 97.050 ;
        RECT 856.950 94.950 859.050 97.050 ;
        RECT 865.950 94.950 868.050 97.050 ;
        RECT 875.400 96.450 876.450 128.400 ;
        RECT 878.400 115.050 879.450 131.400 ;
        RECT 887.400 124.050 888.450 131.400 ;
        RECT 892.950 130.950 895.050 133.050 ;
        RECT 880.950 121.950 883.050 124.050 ;
        RECT 886.950 121.950 889.050 124.050 ;
        RECT 877.950 112.950 880.050 115.050 ;
        RECT 881.400 106.050 882.450 121.950 ;
        RECT 893.400 121.050 894.450 130.950 ;
        RECT 896.400 130.050 897.450 137.100 ;
        RECT 895.950 127.950 898.050 130.050 ;
        RECT 895.950 124.800 898.050 126.900 ;
        RECT 892.950 118.950 895.050 121.050 ;
        RECT 896.400 117.450 897.450 124.800 ;
        RECT 899.400 124.050 900.450 151.950 ;
        RECT 908.400 151.050 909.450 175.950 ;
        RECT 910.950 172.950 913.050 175.050 ;
        RECT 907.950 148.950 910.050 151.050 ;
        RECT 904.950 137.100 907.050 139.200 ;
        RECT 911.400 138.600 912.450 172.950 ;
        RECT 914.400 169.050 915.450 176.400 ;
        RECT 913.950 166.950 916.050 169.050 ;
        RECT 920.400 145.050 921.450 176.400 ;
        RECT 922.950 175.950 925.050 178.050 ;
        RECT 919.950 142.950 922.050 145.050 ;
        RECT 905.400 136.350 906.600 137.100 ;
        RECT 911.400 136.350 912.600 138.600 ;
        RECT 916.950 138.000 919.050 142.050 ;
        RECT 917.400 136.350 918.600 138.000 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 913.950 133.950 916.050 136.050 ;
        RECT 916.950 133.950 919.050 136.050 ;
        RECT 908.400 132.900 909.600 133.650 ;
        RECT 914.400 132.900 915.600 133.650 ;
        RECT 901.950 130.800 904.050 132.900 ;
        RECT 907.950 130.800 910.050 132.900 ;
        RECT 913.950 130.800 916.050 132.900 ;
        RECT 898.950 121.950 901.050 124.050 ;
        RECT 893.400 116.400 897.450 117.450 ;
        RECT 883.950 106.950 886.050 112.050 ;
        RECT 886.950 109.050 889.050 109.200 ;
        RECT 886.950 107.100 892.050 109.050 ;
        RECT 888.000 106.950 892.050 107.100 ;
        RECT 880.950 105.450 883.050 106.050 ;
        RECT 872.400 95.400 876.450 96.450 ;
        RECT 878.400 104.400 883.050 105.450 ;
        RECT 841.950 76.950 844.050 79.050 ;
        RECT 826.950 73.950 829.050 76.050 ;
        RECT 827.400 60.600 828.450 73.950 ;
        RECT 853.950 70.950 856.050 73.050 ;
        RECT 827.400 58.350 828.600 60.600 ;
        RECT 832.950 59.100 835.050 61.200 ;
        RECT 844.950 59.100 847.050 61.200 ;
        RECT 854.400 60.600 855.450 70.950 ;
        RECT 857.400 64.050 858.450 94.950 ;
        RECT 862.950 67.950 865.050 70.050 ;
        RECT 856.950 61.950 859.050 64.050 ;
        RECT 833.400 58.350 834.600 59.100 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 835.950 55.950 838.050 58.050 ;
        RECT 781.950 28.950 784.050 31.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 734.400 21.900 735.600 22.650 ;
        RECT 740.400 21.900 741.600 22.650 ;
        RECT 752.400 21.900 753.600 22.650 ;
        RECT 733.950 19.800 736.050 21.900 ;
        RECT 739.950 19.800 742.050 21.900 ;
        RECT 751.950 19.800 754.050 21.900 ;
        RECT 758.400 21.000 759.600 22.650 ;
        RECT 757.950 16.950 760.050 21.000 ;
        RECT 767.400 13.050 768.450 25.950 ;
        RECT 776.400 25.350 777.600 27.600 ;
        RECT 782.400 27.450 783.600 27.600 ;
        RECT 782.400 26.400 789.450 27.450 ;
        RECT 782.400 25.350 783.600 26.400 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 778.950 22.950 781.050 25.050 ;
        RECT 781.950 22.950 784.050 25.050 ;
        RECT 773.400 21.900 774.600 22.650 ;
        RECT 772.950 19.800 775.050 21.900 ;
        RECT 779.400 21.000 780.600 22.650 ;
        RECT 778.950 16.950 781.050 21.000 ;
        RECT 788.400 19.050 789.450 26.400 ;
        RECT 790.950 26.100 793.050 28.200 ;
        RECT 799.950 26.100 802.050 28.200 ;
        RECT 806.400 27.600 807.450 49.950 ;
        RECT 811.950 43.950 814.050 46.050 ;
        RECT 787.950 16.950 790.050 19.050 ;
        RECT 766.950 10.950 769.050 13.050 ;
        RECT 791.400 7.050 792.450 26.100 ;
        RECT 800.400 25.350 801.600 26.100 ;
        RECT 806.400 25.350 807.600 27.600 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 799.950 22.950 802.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 797.400 21.900 798.600 22.650 ;
        RECT 796.950 19.800 799.050 21.900 ;
        RECT 803.400 21.000 804.600 22.650 ;
        RECT 797.400 13.050 798.450 19.800 ;
        RECT 799.950 15.450 802.050 19.050 ;
        RECT 802.950 16.950 805.050 21.000 ;
        RECT 808.950 15.450 811.050 16.050 ;
        RECT 799.950 15.000 811.050 15.450 ;
        RECT 800.400 14.400 811.050 15.000 ;
        RECT 808.950 13.950 811.050 14.400 ;
        RECT 796.950 10.950 799.050 13.050 ;
        RECT 812.400 10.050 813.450 43.950 ;
        RECT 815.400 40.050 816.450 53.400 ;
        RECT 820.950 52.950 823.050 55.050 ;
        RECT 830.400 54.900 831.600 55.650 ;
        RECT 829.950 52.800 832.050 54.900 ;
        RECT 836.400 53.400 837.600 55.650 ;
        RECT 829.950 43.950 832.050 46.050 ;
        RECT 814.950 37.950 817.050 40.050 ;
        RECT 823.950 26.100 826.050 28.200 ;
        RECT 830.400 27.600 831.450 43.950 ;
        RECT 836.400 40.050 837.450 53.400 ;
        RECT 845.400 46.050 846.450 59.100 ;
        RECT 854.400 58.350 855.600 60.600 ;
        RECT 859.950 59.100 862.050 61.200 ;
        RECT 863.400 61.050 864.450 67.950 ;
        RECT 860.400 58.350 861.600 59.100 ;
        RECT 862.950 58.950 865.050 61.050 ;
        RECT 866.400 58.050 867.450 94.950 ;
        RECT 868.950 61.950 871.050 64.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 853.950 55.950 856.050 58.050 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 859.950 55.950 862.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 851.400 54.900 852.600 55.650 ;
        RECT 857.400 54.900 858.600 55.650 ;
        RECT 864.000 54.900 867.000 55.050 ;
        RECT 850.950 52.800 853.050 54.900 ;
        RECT 856.950 52.800 859.050 54.900 ;
        RECT 862.950 52.950 868.050 54.900 ;
        RECT 862.950 52.800 865.050 52.950 ;
        RECT 865.950 52.800 868.050 52.950 ;
        RECT 869.400 49.050 870.450 61.950 ;
        RECT 872.400 61.050 873.450 95.400 ;
        RECT 878.400 64.200 879.450 104.400 ;
        RECT 880.950 103.950 883.050 104.400 ;
        RECT 886.950 103.950 889.050 106.050 ;
        RECT 893.400 105.600 894.450 116.400 ;
        RECT 887.400 103.350 888.600 103.950 ;
        RECT 893.400 103.350 894.600 105.600 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 889.950 100.950 892.050 103.050 ;
        RECT 892.950 100.950 895.050 103.050 ;
        RECT 884.400 99.900 885.600 100.650 ;
        RECT 883.950 97.800 886.050 99.900 ;
        RECT 890.400 98.400 891.600 100.650 ;
        RECT 884.400 66.450 885.450 97.800 ;
        RECT 890.400 94.050 891.450 98.400 ;
        RECT 889.950 91.950 892.050 94.050 ;
        RECT 889.950 73.950 892.050 76.050 ;
        RECT 884.400 65.400 888.450 66.450 ;
        RECT 877.950 62.100 880.050 64.200 ;
        RECT 871.950 58.950 874.050 61.050 ;
        RECT 877.950 58.950 880.050 61.050 ;
        RECT 883.950 60.000 886.050 64.050 ;
        RECT 887.400 61.050 888.450 65.400 ;
        RECT 878.400 58.350 879.600 58.950 ;
        RECT 884.400 58.350 885.600 60.000 ;
        RECT 886.950 58.950 889.050 61.050 ;
        RECT 874.950 55.950 877.050 58.050 ;
        RECT 877.950 55.950 880.050 58.050 ;
        RECT 880.950 55.950 883.050 58.050 ;
        RECT 883.950 55.950 886.050 58.050 ;
        RECT 871.950 52.950 874.050 55.050 ;
        RECT 875.400 53.400 876.600 55.650 ;
        RECT 881.400 53.400 882.600 55.650 ;
        RECT 847.950 46.950 850.050 49.050 ;
        RECT 868.950 46.950 871.050 49.050 ;
        RECT 844.950 43.950 847.050 46.050 ;
        RECT 835.950 37.950 838.050 40.050 ;
        RECT 848.400 27.600 849.450 46.950 ;
        RECT 850.950 43.950 853.050 46.050 ;
        RECT 872.400 45.450 873.450 52.950 ;
        RECT 869.400 44.400 873.450 45.450 ;
        RECT 851.400 40.050 852.450 43.950 ;
        RECT 850.950 37.950 853.050 40.050 ;
        RECT 869.400 27.600 870.450 44.400 ;
        RECT 875.400 37.050 876.450 53.400 ;
        RECT 881.400 49.050 882.450 53.400 ;
        RECT 880.950 46.950 883.050 49.050 ;
        RECT 874.950 34.950 877.050 37.050 ;
        RECT 890.400 30.450 891.450 73.950 ;
        RECT 902.400 70.050 903.450 130.800 ;
        RECT 923.400 130.050 924.450 175.950 ;
        RECT 926.400 172.050 927.450 187.950 ;
        RECT 925.950 169.950 928.050 172.050 ;
        RECT 925.950 139.950 928.050 142.050 ;
        RECT 904.950 127.950 907.050 130.050 ;
        RECT 922.950 127.950 925.050 130.050 ;
        RECT 901.950 67.950 904.050 70.050 ;
        RECT 902.400 64.050 903.450 67.950 ;
        RECT 901.950 61.950 904.050 64.050 ;
        RECT 898.950 59.100 901.050 61.200 ;
        RECT 905.400 60.600 906.450 127.950 ;
        RECT 926.400 127.050 927.450 139.950 ;
        RECT 929.400 139.050 930.450 187.950 ;
        RECT 932.400 184.050 933.450 190.950 ;
        RECT 938.400 186.450 939.450 202.950 ;
        RECT 941.400 193.050 942.450 209.400 ;
        RECT 943.950 208.950 946.050 211.050 ;
        RECT 940.950 190.950 943.050 193.050 ;
        RECT 944.400 190.050 945.450 208.950 ;
        RECT 943.950 187.950 946.050 190.050 ;
        RECT 938.400 185.400 942.450 186.450 ;
        RECT 931.950 181.950 934.050 184.050 ;
        RECT 934.950 182.100 937.050 184.200 ;
        RECT 941.400 183.600 942.450 185.400 ;
        RECT 947.400 184.050 948.450 253.950 ;
        RECT 935.400 181.350 936.600 182.100 ;
        RECT 941.400 181.350 942.600 183.600 ;
        RECT 946.950 181.950 949.050 184.050 ;
        RECT 934.950 178.950 937.050 181.050 ;
        RECT 937.950 178.950 940.050 181.050 ;
        RECT 940.950 178.950 943.050 181.050 ;
        RECT 943.950 178.950 946.050 181.050 ;
        RECT 931.950 175.950 934.050 178.050 ;
        RECT 938.400 176.400 939.600 178.650 ;
        RECT 944.400 176.400 945.600 178.650 ;
        RECT 932.400 139.200 933.450 175.950 ;
        RECT 934.950 172.950 937.050 175.050 ;
        RECT 935.400 142.050 936.450 172.950 ;
        RECT 938.400 172.050 939.450 176.400 ;
        RECT 937.950 169.950 940.050 172.050 ;
        RECT 944.400 163.050 945.450 176.400 ;
        RECT 946.950 172.950 949.050 175.050 ;
        RECT 943.950 160.950 946.050 163.050 ;
        RECT 937.950 151.950 940.050 154.050 ;
        RECT 947.400 153.450 948.450 172.950 ;
        RECT 944.400 152.400 948.450 153.450 ;
        RECT 934.950 139.950 937.050 142.050 ;
        RECT 928.950 136.950 931.050 139.050 ;
        RECT 931.950 137.100 934.050 139.200 ;
        RECT 938.400 138.600 939.450 151.950 ;
        RECT 944.400 139.050 945.450 152.400 ;
        RECT 946.950 148.950 949.050 151.050 ;
        RECT 932.400 136.350 933.600 137.100 ;
        RECT 938.400 136.350 939.600 138.600 ;
        RECT 943.950 136.950 946.050 139.050 ;
        RECT 931.950 133.950 934.050 136.050 ;
        RECT 934.950 133.950 937.050 136.050 ;
        RECT 937.950 133.950 940.050 136.050 ;
        RECT 940.950 133.950 943.050 136.050 ;
        RECT 928.950 130.950 931.050 133.050 ;
        RECT 935.400 131.400 936.600 133.650 ;
        RECT 941.400 132.900 942.600 133.650 ;
        RECT 947.400 133.050 948.450 148.950 ;
        RECT 925.950 124.950 928.050 127.050 ;
        RECT 919.950 115.950 922.050 118.050 ;
        RECT 910.950 112.950 913.050 115.050 ;
        RECT 911.400 105.600 912.450 112.950 ;
        RECT 920.400 105.600 921.450 115.950 ;
        RECT 911.400 103.350 912.600 105.600 ;
        RECT 920.400 103.350 921.600 105.600 ;
        RECT 910.800 100.950 912.900 103.050 ;
        RECT 916.950 100.950 919.050 103.050 ;
        RECT 919.950 100.950 922.050 103.050 ;
        RECT 925.500 100.950 927.600 103.050 ;
        RECT 917.400 98.400 918.600 100.650 ;
        RECT 926.400 98.400 927.600 100.650 ;
        RECT 917.400 88.050 918.450 98.400 ;
        RECT 926.400 94.050 927.450 98.400 ;
        RECT 925.950 91.950 928.050 94.050 ;
        RECT 916.950 85.950 919.050 88.050 ;
        RECT 929.400 76.050 930.450 130.950 ;
        RECT 931.950 127.950 934.050 130.050 ;
        RECT 928.950 73.950 931.050 76.050 ;
        RECT 905.400 60.450 906.600 60.600 ;
        RECT 907.950 60.450 910.050 64.050 ;
        RECT 910.950 61.950 913.050 64.050 ;
        RECT 905.400 60.000 910.050 60.450 ;
        RECT 905.400 59.400 909.450 60.000 ;
        RECT 899.400 58.350 900.600 59.100 ;
        RECT 905.400 58.350 906.600 59.400 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 898.950 55.950 901.050 58.050 ;
        RECT 901.950 55.950 904.050 58.050 ;
        RECT 904.950 55.950 907.050 58.050 ;
        RECT 896.400 53.400 897.600 55.650 ;
        RECT 902.400 53.400 903.600 55.650 ;
        RECT 911.400 55.050 912.450 61.950 ;
        RECT 919.950 60.000 922.050 64.050 ;
        RECT 920.400 58.350 921.600 60.000 ;
        RECT 925.950 59.100 928.050 61.200 ;
        RECT 926.400 58.350 927.600 59.100 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 919.950 55.950 922.050 58.050 ;
        RECT 922.950 55.950 925.050 58.050 ;
        RECT 925.950 55.950 928.050 58.050 ;
        RECT 896.400 46.050 897.450 53.400 ;
        RECT 895.950 43.950 898.050 46.050 ;
        RECT 902.400 43.050 903.450 53.400 ;
        RECT 910.950 52.950 913.050 55.050 ;
        RECT 917.400 54.900 918.600 55.650 ;
        RECT 916.950 52.800 919.050 54.900 ;
        RECT 923.400 53.400 924.600 55.650 ;
        RECT 904.950 49.950 907.050 52.050 ;
        RECT 901.950 40.950 904.050 43.050 ;
        RECT 887.400 29.400 891.450 30.450 ;
        RECT 887.400 27.600 888.450 29.400 ;
        RECT 824.400 25.350 825.600 26.100 ;
        RECT 830.400 25.350 831.600 27.600 ;
        RECT 848.400 25.350 849.600 27.600 ;
        RECT 863.400 27.450 864.600 27.600 ;
        RECT 857.400 26.400 864.600 27.450 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 829.950 22.950 832.050 25.050 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 817.950 16.950 820.050 22.050 ;
        RECT 821.400 21.000 822.600 22.650 ;
        RECT 827.400 21.000 828.600 22.650 ;
        RECT 820.950 16.950 823.050 21.000 ;
        RECT 826.950 16.950 829.050 21.000 ;
        RECT 839.400 16.050 840.450 22.950 ;
        RECT 845.400 21.000 846.600 22.650 ;
        RECT 844.950 16.950 847.050 21.000 ;
        RECT 857.400 19.050 858.450 26.400 ;
        RECT 863.400 25.350 864.600 26.400 ;
        RECT 869.400 25.350 870.600 27.600 ;
        RECT 887.400 25.350 888.600 27.600 ;
        RECT 892.950 27.000 895.050 31.050 ;
        RECT 893.400 25.350 894.600 27.000 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 868.950 22.950 871.050 25.050 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 895.950 22.950 898.050 25.050 ;
        RECT 866.400 21.900 867.600 22.650 ;
        RECT 865.950 19.800 868.050 21.900 ;
        RECT 872.400 20.400 873.600 22.650 ;
        RECT 890.400 20.400 891.600 22.650 ;
        RECT 896.400 20.400 897.600 22.650 ;
        RECT 905.400 21.900 906.450 49.950 ;
        RECT 919.950 46.950 922.050 49.050 ;
        RECT 913.950 40.950 916.050 43.050 ;
        RECT 914.400 27.600 915.450 40.950 ;
        RECT 920.400 27.600 921.450 46.950 ;
        RECT 923.400 43.050 924.450 53.400 ;
        RECT 922.950 40.950 925.050 43.050 ;
        RECT 932.400 34.050 933.450 127.950 ;
        RECT 935.400 127.050 936.450 131.400 ;
        RECT 940.950 130.800 943.050 132.900 ;
        RECT 946.950 130.950 949.050 133.050 ;
        RECT 943.950 127.950 946.050 130.050 ;
        RECT 934.950 124.950 937.050 127.050 ;
        RECT 937.950 121.950 940.050 124.050 ;
        RECT 934.950 61.950 937.050 64.050 ;
        RECT 931.950 31.950 934.050 34.050 ;
        RECT 935.400 28.200 936.450 61.950 ;
        RECT 938.400 49.050 939.450 121.950 ;
        RECT 940.950 106.950 943.050 109.050 ;
        RECT 937.950 46.950 940.050 49.050 ;
        RECT 914.400 25.350 915.600 27.600 ;
        RECT 920.400 25.350 921.600 27.600 ;
        RECT 925.950 26.100 928.050 28.200 ;
        RECT 934.950 26.100 937.050 28.200 ;
        RECT 910.950 22.950 913.050 25.050 ;
        RECT 913.950 22.950 916.050 25.050 ;
        RECT 916.950 22.950 919.050 25.050 ;
        RECT 919.950 22.950 922.050 25.050 ;
        RECT 911.400 21.900 912.600 22.650 ;
        RECT 917.400 21.900 918.600 22.650 ;
        RECT 856.950 16.950 859.050 19.050 ;
        RECT 825.000 15.900 828.000 16.050 ;
        RECT 823.950 13.950 829.050 15.900 ;
        RECT 838.950 13.950 841.050 16.050 ;
        RECT 823.950 13.800 826.050 13.950 ;
        RECT 826.950 13.800 829.050 13.950 ;
        RECT 872.400 10.050 873.450 20.400 ;
        RECT 811.950 7.950 814.050 10.050 ;
        RECT 871.950 7.950 874.050 10.050 ;
        RECT 890.400 7.050 891.450 20.400 ;
        RECT 896.400 16.050 897.450 20.400 ;
        RECT 904.950 19.800 907.050 21.900 ;
        RECT 910.950 19.800 913.050 21.900 ;
        RECT 916.950 19.800 919.050 21.900 ;
        RECT 895.950 13.950 898.050 16.050 ;
        RECT 926.400 10.050 927.450 26.100 ;
        RECT 935.400 25.350 936.600 26.100 ;
        RECT 931.950 22.950 934.050 25.050 ;
        RECT 934.950 22.950 937.050 25.050 ;
        RECT 932.400 21.900 933.600 22.650 ;
        RECT 931.950 19.800 934.050 21.900 ;
        RECT 925.950 7.950 928.050 10.050 ;
        RECT 941.400 7.050 942.450 106.950 ;
        RECT 944.400 16.050 945.450 127.950 ;
        RECT 943.950 13.950 946.050 16.050 ;
        RECT 586.950 4.950 589.050 7.050 ;
        RECT 724.950 4.950 727.050 7.050 ;
        RECT 790.950 4.950 793.050 7.050 ;
        RECT 889.950 4.950 892.050 7.050 ;
        RECT 940.950 4.950 943.050 7.050 ;
        RECT 436.950 3.450 439.050 4.050 ;
        RECT 431.400 2.400 439.050 3.450 ;
        RECT 436.950 1.950 439.050 2.400 ;
        RECT 508.950 3.450 511.050 4.050 ;
        RECT 514.950 3.450 517.050 4.050 ;
        RECT 508.950 2.400 517.050 3.450 ;
        RECT 508.950 1.950 511.050 2.400 ;
        RECT 514.950 1.950 517.050 2.400 ;
        RECT 541.950 1.950 544.050 4.050 ;
      LAYER metal3 ;
        RECT 244.950 933.600 247.050 934.050 ;
        RECT 274.950 933.600 277.050 934.050 ;
        RECT 244.950 932.400 277.050 933.600 ;
        RECT 244.950 931.950 247.050 932.400 ;
        RECT 274.950 931.950 277.050 932.400 ;
        RECT 220.950 930.600 223.050 931.050 ;
        RECT 256.950 930.600 259.050 931.050 ;
        RECT 220.950 929.400 259.050 930.600 ;
        RECT 220.950 928.950 223.050 929.400 ;
        RECT 256.950 928.950 259.050 929.400 ;
        RECT 352.950 930.600 355.050 931.050 ;
        RECT 442.950 930.600 445.050 931.050 ;
        RECT 352.950 929.400 445.050 930.600 ;
        RECT 352.950 928.950 355.050 929.400 ;
        RECT 442.950 928.950 445.050 929.400 ;
        RECT 16.950 927.600 19.050 928.050 ;
        RECT 106.950 927.600 109.050 928.050 ;
        RECT 16.950 926.400 109.050 927.600 ;
        RECT 16.950 925.950 19.050 926.400 ;
        RECT 106.950 925.950 109.050 926.400 ;
        RECT 286.950 927.600 289.050 928.050 ;
        RECT 658.950 927.600 661.050 928.050 ;
        RECT 286.950 926.400 661.050 927.600 ;
        RECT 286.950 925.950 289.050 926.400 ;
        RECT 658.950 925.950 661.050 926.400 ;
        RECT 55.950 924.600 58.050 925.050 ;
        RECT 97.950 924.600 100.050 925.050 ;
        RECT 55.950 923.400 100.050 924.600 ;
        RECT 55.950 922.950 58.050 923.400 ;
        RECT 97.950 922.950 100.050 923.400 ;
        RECT 121.950 924.600 124.050 925.050 ;
        RECT 184.950 924.600 187.050 925.050 ;
        RECT 250.950 924.600 253.050 925.050 ;
        RECT 121.950 923.400 253.050 924.600 ;
        RECT 121.950 922.950 124.050 923.400 ;
        RECT 184.950 922.950 187.050 923.400 ;
        RECT 250.950 922.950 253.050 923.400 ;
        RECT 754.950 924.600 757.050 924.900 ;
        RECT 793.950 924.600 796.050 925.050 ;
        RECT 754.950 923.400 796.050 924.600 ;
        RECT 754.950 922.800 757.050 923.400 ;
        RECT 793.950 922.950 796.050 923.400 ;
        RECT 898.950 924.600 901.050 925.050 ;
        RECT 922.950 924.600 925.050 925.050 ;
        RECT 898.950 923.400 925.050 924.600 ;
        RECT 898.950 922.950 901.050 923.400 ;
        RECT 922.950 922.950 925.050 923.400 ;
        RECT 100.950 921.600 103.050 922.050 ;
        RECT 112.950 921.600 115.050 922.050 ;
        RECT 100.950 920.400 115.050 921.600 ;
        RECT 100.950 919.950 103.050 920.400 ;
        RECT 112.950 919.950 115.050 920.400 ;
        RECT 202.950 921.600 205.050 922.050 ;
        RECT 214.950 921.600 217.050 922.050 ;
        RECT 202.950 920.400 217.050 921.600 ;
        RECT 202.950 919.950 205.050 920.400 ;
        RECT 214.950 919.950 217.050 920.400 ;
        RECT 406.950 921.750 409.050 922.200 ;
        RECT 412.950 921.750 415.050 922.200 ;
        RECT 406.950 920.550 415.050 921.750 ;
        RECT 406.950 920.100 409.050 920.550 ;
        RECT 412.950 920.100 415.050 920.550 ;
        RECT 496.950 921.600 499.050 922.200 ;
        RECT 505.950 921.600 508.050 922.200 ;
        RECT 580.950 921.600 583.050 922.050 ;
        RECT 595.950 921.600 598.050 922.200 ;
        RECT 496.950 920.400 598.050 921.600 ;
        RECT 496.950 920.100 499.050 920.400 ;
        RECT 505.950 920.100 508.050 920.400 ;
        RECT 52.950 918.750 55.050 919.200 ;
        RECT 61.950 918.750 64.050 919.200 ;
        RECT 52.950 917.550 64.050 918.750 ;
        RECT 52.950 917.100 55.050 917.550 ;
        RECT 61.950 917.100 64.050 917.550 ;
        RECT 67.950 918.750 70.050 919.200 ;
        RECT 76.950 918.750 79.050 919.200 ;
        RECT 67.950 917.550 79.050 918.750 ;
        RECT 67.950 917.100 70.050 917.550 ;
        RECT 76.950 917.100 79.050 917.550 ;
        RECT 82.950 917.100 85.050 919.200 ;
        RECT 106.950 918.600 109.050 919.200 ;
        RECT 86.400 917.400 109.050 918.600 ;
        RECT 53.400 915.600 54.600 917.100 ;
        RECT 83.400 915.600 84.600 917.100 ;
        RECT 53.400 914.400 84.600 915.600 ;
        RECT 86.400 912.900 87.600 917.400 ;
        RECT 106.950 917.100 109.050 917.400 ;
        RECT 136.950 918.750 139.050 919.200 ;
        RECT 142.950 918.750 145.050 919.200 ;
        RECT 136.950 917.550 145.050 918.750 ;
        RECT 136.950 917.100 139.050 917.550 ;
        RECT 142.950 917.100 145.050 917.550 ;
        RECT 148.950 918.600 151.050 919.200 ;
        RECT 157.950 918.750 160.050 919.200 ;
        RECT 163.950 918.750 166.050 919.200 ;
        RECT 157.950 918.600 166.050 918.750 ;
        RECT 148.950 917.550 166.050 918.600 ;
        RECT 148.950 917.400 160.050 917.550 ;
        RECT 148.950 917.100 151.050 917.400 ;
        RECT 157.950 917.100 160.050 917.400 ;
        RECT 163.950 917.100 166.050 917.550 ;
        RECT 169.950 917.100 172.050 919.200 ;
        RECT 190.950 917.100 193.050 919.200 ;
        RECT 208.950 918.600 211.050 919.200 ;
        RECT 226.950 918.600 229.050 919.200 ;
        RECT 208.950 917.400 229.050 918.600 ;
        RECT 208.950 917.100 211.050 917.400 ;
        RECT 226.950 917.100 229.050 917.400 ;
        RECT 232.950 918.750 235.050 919.200 ;
        RECT 241.950 918.750 244.050 919.200 ;
        RECT 232.950 917.550 244.050 918.750 ;
        RECT 280.950 918.600 283.050 919.200 ;
        RECT 232.950 917.100 235.050 917.550 ;
        RECT 241.950 917.100 244.050 917.550 ;
        RECT 275.400 917.400 283.050 918.600 ;
        RECT 97.950 915.600 100.050 916.050 ;
        RECT 121.950 915.600 124.050 916.050 ;
        RECT 97.950 914.400 124.050 915.600 ;
        RECT 137.400 915.600 138.600 917.100 ;
        RECT 170.400 915.600 171.600 917.100 ;
        RECT 137.400 914.400 171.600 915.600 ;
        RECT 97.950 913.950 100.050 914.400 ;
        RECT 121.950 913.950 124.050 914.400 ;
        RECT 85.950 910.800 88.050 912.900 ;
        RECT 139.950 912.450 142.050 912.900 ;
        RECT 145.950 912.450 148.050 912.900 ;
        RECT 139.950 911.250 148.050 912.450 ;
        RECT 139.950 910.800 142.050 911.250 ;
        RECT 145.950 910.800 148.050 911.250 ;
        RECT 166.950 912.600 169.050 912.900 ;
        RECT 191.400 912.600 192.600 917.100 ;
        RECT 166.950 911.400 192.600 912.600 ;
        RECT 193.950 912.450 196.050 912.900 ;
        RECT 205.950 912.450 208.050 912.900 ;
        RECT 166.950 910.800 169.050 911.400 ;
        RECT 193.950 911.250 208.050 912.450 ;
        RECT 193.950 910.800 196.050 911.250 ;
        RECT 205.950 910.800 208.050 911.250 ;
        RECT 211.950 912.600 214.050 912.900 ;
        RECT 220.950 912.600 223.050 913.050 ;
        RECT 211.950 911.400 223.050 912.600 ;
        RECT 211.950 910.800 214.050 911.400 ;
        RECT 220.950 910.950 223.050 911.400 ;
        RECT 259.950 912.600 262.050 912.900 ;
        RECT 275.400 912.600 276.600 917.400 ;
        RECT 280.950 917.100 283.050 917.400 ;
        RECT 340.950 918.600 343.050 919.200 ;
        RECT 340.950 918.000 351.600 918.600 ;
        RECT 340.950 917.400 352.050 918.000 ;
        RECT 340.950 917.100 343.050 917.400 ;
        RECT 349.950 913.950 352.050 917.400 ;
        RECT 382.950 914.100 385.050 916.200 ;
        RECT 448.950 915.750 451.050 916.200 ;
        RECT 472.950 915.750 475.050 916.200 ;
        RECT 497.400 916.050 498.600 920.100 ;
        RECT 580.950 919.950 583.050 920.400 ;
        RECT 595.950 920.100 598.050 920.400 ;
        RECT 865.950 921.600 868.050 922.050 ;
        RECT 889.950 921.600 892.050 922.050 ;
        RECT 913.950 921.600 916.050 922.050 ;
        RECT 937.950 921.600 940.050 922.050 ;
        RECT 865.950 920.400 940.050 921.600 ;
        RECT 865.950 919.950 868.050 920.400 ;
        RECT 889.950 919.950 892.050 920.400 ;
        RECT 913.950 919.950 916.050 920.400 ;
        RECT 937.950 919.950 940.050 920.400 ;
        RECT 673.950 918.600 676.050 919.200 ;
        RECT 694.950 918.600 697.050 919.050 ;
        RECT 673.950 917.400 697.050 918.600 ;
        RECT 673.950 917.100 676.050 917.400 ;
        RECT 694.950 916.950 697.050 917.400 ;
        RECT 802.950 918.750 805.050 919.200 ;
        RECT 808.950 918.750 811.050 919.200 ;
        RECT 802.950 917.550 811.050 918.750 ;
        RECT 802.950 917.100 805.050 917.550 ;
        RECT 808.950 917.100 811.050 917.550 ;
        RECT 820.950 918.750 823.050 919.200 ;
        RECT 832.950 918.750 835.050 919.200 ;
        RECT 820.950 917.550 835.050 918.750 ;
        RECT 838.950 918.600 841.050 919.200 ;
        RECT 820.950 917.100 823.050 917.550 ;
        RECT 832.950 917.100 835.050 917.550 ;
        RECT 836.400 917.400 841.050 918.600 ;
        RECT 448.950 914.550 475.050 915.750 ;
        RECT 448.950 914.100 451.050 914.550 ;
        RECT 472.950 914.100 475.050 914.550 ;
        RECT 493.950 914.400 498.600 916.050 ;
        RECT 529.950 915.600 532.050 916.200 ;
        RECT 500.400 914.400 532.050 915.600 ;
        RECT 259.950 911.400 276.600 912.600 ;
        RECT 277.950 912.450 280.050 912.900 ;
        RECT 286.950 912.450 289.050 912.900 ;
        RECT 259.950 910.800 262.050 911.400 ;
        RECT 277.950 911.250 289.050 912.450 ;
        RECT 277.950 910.800 280.050 911.250 ;
        RECT 286.950 910.800 289.050 911.250 ;
        RECT 322.950 912.600 325.050 912.900 ;
        RECT 337.950 912.600 340.050 912.900 ;
        RECT 346.950 912.600 349.050 913.050 ;
        RECT 322.950 911.400 349.050 912.600 ;
        RECT 383.400 912.600 384.600 914.100 ;
        RECT 493.950 913.950 498.000 914.400 ;
        RECT 397.950 912.600 400.050 913.050 ;
        RECT 383.400 911.400 400.050 912.600 ;
        RECT 322.950 910.800 325.050 911.400 ;
        RECT 337.950 910.800 340.050 911.400 ;
        RECT 346.950 910.950 349.050 911.400 ;
        RECT 397.950 910.950 400.050 911.400 ;
        RECT 490.950 912.600 493.050 913.050 ;
        RECT 500.400 912.600 501.600 914.400 ;
        RECT 529.950 914.100 532.050 914.400 ;
        RECT 574.950 915.750 577.050 916.200 ;
        RECT 619.950 915.750 622.050 916.200 ;
        RECT 574.950 914.550 622.050 915.750 ;
        RECT 574.950 914.100 577.050 914.550 ;
        RECT 619.950 914.100 622.050 914.550 ;
        RECT 697.950 915.450 700.050 915.900 ;
        RECT 718.950 915.450 721.050 915.900 ;
        RECT 697.950 914.250 721.050 915.450 ;
        RECT 697.950 913.800 700.050 914.250 ;
        RECT 718.950 913.800 721.050 914.250 ;
        RECT 836.400 913.050 837.600 917.400 ;
        RECT 838.950 917.100 841.050 917.400 ;
        RECT 490.950 911.400 501.600 912.600 ;
        RECT 556.950 912.600 559.050 913.050 ;
        RECT 643.950 912.600 646.050 913.050 ;
        RECT 556.950 911.400 646.050 912.600 ;
        RECT 490.950 910.950 493.050 911.400 ;
        RECT 556.950 910.950 559.050 911.400 ;
        RECT 643.950 910.950 646.050 911.400 ;
        RECT 658.950 912.600 661.050 913.050 ;
        RECT 670.950 912.600 673.050 912.900 ;
        RECT 658.950 911.400 673.050 912.600 ;
        RECT 658.950 910.950 661.050 911.400 ;
        RECT 670.950 910.800 673.050 911.400 ;
        RECT 808.950 912.600 811.050 913.050 ;
        RECT 817.950 912.600 820.050 912.900 ;
        RECT 808.950 911.400 820.050 912.600 ;
        RECT 808.950 910.950 811.050 911.400 ;
        RECT 817.950 910.800 820.050 911.400 ;
        RECT 835.950 910.950 838.050 913.050 ;
        RECT 883.950 912.450 886.050 912.900 ;
        RECT 889.950 912.450 892.050 912.900 ;
        RECT 883.950 911.250 892.050 912.450 ;
        RECT 883.950 910.800 886.050 911.250 ;
        RECT 889.950 910.800 892.050 911.250 ;
        RECT 88.950 909.600 91.050 910.050 ;
        RECT 136.950 909.600 139.050 910.050 ;
        RECT 88.950 908.400 139.050 909.600 ;
        RECT 88.950 907.950 91.050 908.400 ;
        RECT 136.950 907.950 139.050 908.400 ;
        RECT 187.950 909.600 190.050 910.050 ;
        RECT 241.950 909.600 244.050 910.050 ;
        RECT 187.950 908.400 244.050 909.600 ;
        RECT 187.950 907.950 190.050 908.400 ;
        RECT 241.950 907.950 244.050 908.400 ;
        RECT 565.950 909.600 568.050 910.050 ;
        RECT 583.950 909.600 586.050 910.050 ;
        RECT 565.950 908.400 586.050 909.600 ;
        RECT 565.950 907.950 568.050 908.400 ;
        RECT 583.950 907.950 586.050 908.400 ;
        RECT 655.950 909.600 658.050 910.050 ;
        RECT 706.950 909.600 709.050 910.050 ;
        RECT 655.950 908.400 709.050 909.600 ;
        RECT 655.950 907.950 658.050 908.400 ;
        RECT 706.950 907.950 709.050 908.400 ;
        RECT 40.950 906.600 43.050 907.050 ;
        RECT 55.950 906.600 58.050 907.050 ;
        RECT 40.950 905.400 58.050 906.600 ;
        RECT 40.950 904.950 43.050 905.400 ;
        RECT 55.950 904.950 58.050 905.400 ;
        RECT 109.950 906.600 112.050 907.050 ;
        RECT 130.950 906.600 133.050 907.050 ;
        RECT 109.950 905.400 133.050 906.600 ;
        RECT 109.950 904.950 112.050 905.400 ;
        RECT 130.950 904.950 133.050 905.400 ;
        RECT 139.950 906.600 142.050 906.900 ;
        RECT 157.950 906.600 160.050 907.050 ;
        RECT 901.800 906.600 903.900 907.050 ;
        RECT 139.950 905.400 160.050 906.600 ;
        RECT 139.950 904.800 142.050 905.400 ;
        RECT 157.950 904.950 160.050 905.400 ;
        RECT 857.400 905.400 903.900 906.600 ;
        RECT 52.950 903.600 55.050 904.050 ;
        RECT 67.800 903.600 69.900 904.050 ;
        RECT 52.950 902.400 69.900 903.600 ;
        RECT 52.950 901.950 55.050 902.400 ;
        RECT 67.800 901.950 69.900 902.400 ;
        RECT 70.950 903.600 73.050 904.050 ;
        RECT 88.950 903.600 91.050 904.050 ;
        RECT 70.950 902.400 91.050 903.600 ;
        RECT 70.950 901.950 73.050 902.400 ;
        RECT 88.950 901.950 91.050 902.400 ;
        RECT 151.950 903.600 154.050 904.050 ;
        RECT 202.950 903.600 205.050 904.050 ;
        RECT 229.950 903.600 232.050 904.050 ;
        RECT 151.950 902.400 232.050 903.600 ;
        RECT 151.950 901.950 154.050 902.400 ;
        RECT 202.950 901.950 205.050 902.400 ;
        RECT 229.950 901.950 232.050 902.400 ;
        RECT 241.950 903.600 244.050 904.050 ;
        RECT 298.950 903.600 301.050 904.050 ;
        RECT 406.950 903.600 409.050 904.050 ;
        RECT 427.950 903.600 430.050 904.050 ;
        RECT 241.950 902.400 301.050 903.600 ;
        RECT 368.400 903.000 430.050 903.600 ;
        RECT 241.950 901.950 244.050 902.400 ;
        RECT 298.950 901.950 301.050 902.400 ;
        RECT 367.950 902.400 430.050 903.000 ;
        RECT 94.950 900.600 97.050 901.050 ;
        RECT 100.950 900.600 103.050 901.050 ;
        RECT 106.950 900.600 109.050 901.050 ;
        RECT 94.950 899.400 109.050 900.600 ;
        RECT 94.950 898.950 97.050 899.400 ;
        RECT 100.950 898.950 103.050 899.400 ;
        RECT 106.950 898.950 109.050 899.400 ;
        RECT 139.950 900.600 142.050 901.050 ;
        RECT 199.950 900.600 202.050 901.050 ;
        RECT 139.950 899.400 202.050 900.600 ;
        RECT 139.950 898.950 142.050 899.400 ;
        RECT 199.950 898.950 202.050 899.400 ;
        RECT 205.950 900.600 208.050 901.050 ;
        RECT 238.950 900.600 241.050 901.050 ;
        RECT 205.950 899.400 241.050 900.600 ;
        RECT 205.950 898.950 208.050 899.400 ;
        RECT 238.950 898.950 241.050 899.400 ;
        RECT 367.950 898.950 370.050 902.400 ;
        RECT 406.950 901.950 409.050 902.400 ;
        RECT 427.950 901.950 430.050 902.400 ;
        RECT 511.950 903.600 514.050 904.050 ;
        RECT 565.950 903.600 568.050 904.050 ;
        RECT 511.950 902.400 568.050 903.600 ;
        RECT 511.950 901.950 514.050 902.400 ;
        RECT 565.950 901.950 568.050 902.400 ;
        RECT 718.950 903.600 721.050 904.050 ;
        RECT 857.400 903.600 858.600 905.400 ;
        RECT 901.800 904.950 903.900 905.400 ;
        RECT 904.950 906.600 907.050 907.050 ;
        RECT 919.950 906.600 922.050 907.050 ;
        RECT 904.950 905.400 922.050 906.600 ;
        RECT 904.950 904.950 907.050 905.400 ;
        RECT 919.950 904.950 922.050 905.400 ;
        RECT 718.950 902.400 858.600 903.600 ;
        RECT 877.950 903.600 880.050 904.050 ;
        RECT 895.950 903.600 898.050 904.050 ;
        RECT 877.950 902.400 898.050 903.600 ;
        RECT 718.950 901.950 721.050 902.400 ;
        RECT 877.950 901.950 880.050 902.400 ;
        RECT 895.950 901.950 898.050 902.400 ;
        RECT 412.950 900.600 415.050 901.050 ;
        RECT 454.950 900.600 457.050 901.050 ;
        RECT 493.950 900.600 496.050 901.050 ;
        RECT 412.950 899.400 496.050 900.600 ;
        RECT 412.950 898.950 415.050 899.400 ;
        RECT 454.950 898.950 457.050 899.400 ;
        RECT 493.950 898.950 496.050 899.400 ;
        RECT 598.950 900.600 601.050 901.050 ;
        RECT 655.950 900.600 658.050 901.050 ;
        RECT 598.950 899.400 658.050 900.600 ;
        RECT 598.950 898.950 601.050 899.400 ;
        RECT 655.950 898.950 658.050 899.400 ;
        RECT 700.950 900.600 703.050 901.050 ;
        RECT 724.950 900.600 727.050 901.050 ;
        RECT 700.950 899.400 727.050 900.600 ;
        RECT 700.950 898.950 703.050 899.400 ;
        RECT 724.950 898.950 727.050 899.400 ;
        RECT 802.950 900.600 805.050 901.050 ;
        RECT 820.800 900.600 822.900 901.050 ;
        RECT 802.950 899.400 822.900 900.600 ;
        RECT 802.950 898.950 805.050 899.400 ;
        RECT 820.800 898.950 822.900 899.400 ;
        RECT 823.950 900.600 826.050 901.050 ;
        RECT 838.950 900.600 841.050 901.050 ;
        RECT 823.950 899.400 841.050 900.600 ;
        RECT 823.950 898.950 826.050 899.400 ;
        RECT 838.950 898.950 841.050 899.400 ;
        RECT 844.950 900.600 847.050 901.050 ;
        RECT 862.950 900.600 865.050 901.050 ;
        RECT 844.950 899.400 865.050 900.600 ;
        RECT 844.950 898.950 847.050 899.400 ;
        RECT 862.950 898.950 865.050 899.400 ;
        RECT 127.950 897.600 130.050 898.050 ;
        RECT 133.950 897.600 136.050 898.050 ;
        RECT 127.950 896.400 136.050 897.600 ;
        RECT 127.950 895.950 130.050 896.400 ;
        RECT 133.950 895.950 136.050 896.400 ;
        RECT 388.950 897.600 391.050 898.050 ;
        RECT 424.950 897.600 427.050 898.050 ;
        RECT 436.950 897.600 439.050 898.050 ;
        RECT 388.950 896.400 439.050 897.600 ;
        RECT 388.950 895.950 391.050 896.400 ;
        RECT 424.950 895.950 427.050 896.400 ;
        RECT 436.950 895.950 439.050 896.400 ;
        RECT 481.950 897.600 484.050 898.050 ;
        RECT 490.950 897.600 493.050 898.050 ;
        RECT 481.950 896.400 493.050 897.600 ;
        RECT 481.950 895.950 484.050 896.400 ;
        RECT 490.950 895.950 493.050 896.400 ;
        RECT 616.950 897.600 619.050 898.050 ;
        RECT 727.950 897.600 730.050 898.050 ;
        RECT 616.950 896.400 730.050 897.600 ;
        RECT 616.950 895.950 619.050 896.400 ;
        RECT 727.950 895.950 730.050 896.400 ;
        RECT 91.950 894.600 94.050 895.050 ;
        RECT 148.950 894.600 151.050 895.050 ;
        RECT 91.950 893.400 151.050 894.600 ;
        RECT 91.950 892.950 94.050 893.400 ;
        RECT 148.950 892.950 151.050 893.400 ;
        RECT 196.950 894.600 199.050 895.050 ;
        RECT 217.950 894.600 220.050 895.050 ;
        RECT 196.950 893.400 220.050 894.600 ;
        RECT 196.950 892.950 199.050 893.400 ;
        RECT 217.950 892.950 220.050 893.400 ;
        RECT 223.950 894.600 226.050 895.050 ;
        RECT 256.950 894.600 259.050 895.050 ;
        RECT 223.950 893.400 259.050 894.600 ;
        RECT 223.950 892.950 226.050 893.400 ;
        RECT 256.950 892.950 259.050 893.400 ;
        RECT 262.950 894.600 265.050 895.050 ;
        RECT 295.950 894.600 298.050 895.050 ;
        RECT 262.950 893.400 298.050 894.600 ;
        RECT 262.950 892.950 265.050 893.400 ;
        RECT 295.950 892.950 298.050 893.400 ;
        RECT 499.950 894.600 502.050 895.050 ;
        RECT 517.950 894.600 520.050 895.050 ;
        RECT 499.950 893.400 520.050 894.600 ;
        RECT 499.950 892.950 502.050 893.400 ;
        RECT 517.950 892.950 520.050 893.400 ;
        RECT 733.950 894.600 736.050 895.050 ;
        RECT 745.950 894.600 748.050 895.050 ;
        RECT 835.950 894.600 838.050 895.050 ;
        RECT 733.950 893.400 838.050 894.600 ;
        RECT 733.950 892.950 736.050 893.400 ;
        RECT 745.950 892.950 748.050 893.400 ;
        RECT 835.950 892.950 838.050 893.400 ;
        RECT 13.950 891.600 16.050 892.050 ;
        RECT 64.950 891.600 67.050 892.050 ;
        RECT 13.950 890.400 67.050 891.600 ;
        RECT 13.950 889.950 16.050 890.400 ;
        RECT 64.950 889.950 67.050 890.400 ;
        RECT 85.950 891.600 88.050 892.050 ;
        RECT 166.950 891.600 169.050 892.050 ;
        RECT 85.950 890.400 169.050 891.600 ;
        RECT 85.950 889.950 88.050 890.400 ;
        RECT 166.950 889.950 169.050 890.400 ;
        RECT 220.950 891.600 223.050 892.050 ;
        RECT 229.950 891.600 232.050 892.050 ;
        RECT 259.950 891.600 262.050 892.050 ;
        RECT 220.950 890.400 262.050 891.600 ;
        RECT 220.950 889.950 223.050 890.400 ;
        RECT 229.950 889.950 232.050 890.400 ;
        RECT 259.950 889.950 262.050 890.400 ;
        RECT 307.950 891.600 310.050 892.050 ;
        RECT 337.950 891.600 340.050 892.050 ;
        RECT 448.950 891.600 451.050 892.050 ;
        RECT 307.950 890.400 340.050 891.600 ;
        RECT 307.950 889.950 310.050 890.400 ;
        RECT 337.950 889.950 340.050 890.400 ;
        RECT 410.400 890.400 451.050 891.600 ;
        RECT 154.950 888.600 157.050 889.050 ;
        RECT 125.400 887.400 157.050 888.600 ;
        RECT 19.950 884.100 22.050 886.200 ;
        RECT 25.950 885.750 28.050 886.200 ;
        RECT 37.950 885.750 40.050 886.200 ;
        RECT 25.950 884.550 40.050 885.750 ;
        RECT 25.950 884.100 28.050 884.550 ;
        RECT 37.950 884.100 40.050 884.550 ;
        RECT 55.950 884.100 58.050 886.200 ;
        RECT 100.950 884.100 103.050 886.200 ;
        RECT 115.950 885.600 118.050 886.200 ;
        RECT 125.400 886.050 126.600 887.400 ;
        RECT 154.950 886.950 157.050 887.400 ;
        RECT 160.950 886.950 163.050 889.050 ;
        RECT 379.950 888.600 382.050 889.050 ;
        RECT 410.400 888.600 411.600 890.400 ;
        RECT 448.950 889.950 451.050 890.400 ;
        RECT 463.950 891.600 466.050 892.050 ;
        RECT 496.950 891.600 499.050 892.050 ;
        RECT 463.950 890.400 499.050 891.600 ;
        RECT 463.950 889.950 466.050 890.400 ;
        RECT 496.950 889.950 499.050 890.400 ;
        RECT 580.950 891.600 583.050 892.050 ;
        RECT 589.950 891.600 592.050 892.050 ;
        RECT 580.950 890.400 592.050 891.600 ;
        RECT 580.950 889.950 583.050 890.400 ;
        RECT 589.950 889.950 592.050 890.400 ;
        RECT 685.950 891.600 688.050 892.050 ;
        RECT 709.950 891.600 712.050 892.050 ;
        RECT 685.950 890.400 712.050 891.600 ;
        RECT 685.950 889.950 688.050 890.400 ;
        RECT 709.950 889.950 712.050 890.400 ;
        RECT 760.950 891.600 763.050 892.050 ;
        RECT 775.950 891.600 778.050 892.050 ;
        RECT 787.950 891.600 790.050 892.050 ;
        RECT 760.950 890.400 790.050 891.600 ;
        RECT 760.950 889.950 763.050 890.400 ;
        RECT 775.950 889.950 778.050 890.400 ;
        RECT 787.950 889.950 790.050 890.400 ;
        RECT 826.950 891.600 829.050 892.050 ;
        RECT 871.950 891.600 874.050 892.050 ;
        RECT 892.950 891.600 895.050 892.050 ;
        RECT 826.950 890.400 895.050 891.600 ;
        RECT 826.950 889.950 829.050 890.400 ;
        RECT 871.950 889.950 874.050 890.400 ;
        RECT 892.950 889.950 895.050 890.400 ;
        RECT 379.950 887.400 411.600 888.600 ;
        RECT 535.950 888.600 538.050 889.050 ;
        RECT 556.950 888.600 559.050 889.050 ;
        RECT 607.950 888.600 610.050 889.050 ;
        RECT 535.950 887.400 610.050 888.600 ;
        RECT 379.950 886.950 382.050 887.400 ;
        RECT 535.950 886.950 538.050 887.400 ;
        RECT 556.950 886.950 559.050 887.400 ;
        RECT 607.950 886.950 610.050 887.400 ;
        RECT 844.950 888.600 847.050 889.200 ;
        RECT 886.950 888.600 889.050 889.050 ;
        RECT 844.950 887.400 889.050 888.600 ;
        RECT 844.950 887.100 847.050 887.400 ;
        RECT 886.950 886.950 889.050 887.400 ;
        RECT 901.950 888.600 904.050 889.050 ;
        RECT 913.950 888.600 916.050 889.050 ;
        RECT 901.950 887.400 916.050 888.600 ;
        RECT 901.950 886.950 904.050 887.400 ;
        RECT 913.950 886.950 916.050 887.400 ;
        RECT 124.950 885.600 127.050 886.050 ;
        RECT 115.950 884.400 127.050 885.600 ;
        RECT 115.950 884.100 118.050 884.400 ;
        RECT 20.400 880.050 21.600 884.100 ;
        RECT 56.400 880.050 57.600 884.100 ;
        RECT 101.400 880.050 102.600 884.100 ;
        RECT 124.950 883.950 127.050 884.400 ;
        RECT 157.950 884.100 160.050 886.200 ;
        RECT 20.400 878.400 25.050 880.050 ;
        RECT 21.000 877.950 25.050 878.400 ;
        RECT 34.950 879.450 37.050 879.900 ;
        RECT 46.950 879.450 49.050 879.900 ;
        RECT 34.950 878.250 49.050 879.450 ;
        RECT 34.950 877.800 37.050 878.250 ;
        RECT 46.950 877.800 49.050 878.250 ;
        RECT 52.950 878.400 57.600 880.050 ;
        RECT 58.950 879.600 61.050 879.900 ;
        RECT 79.950 879.600 82.050 879.900 ;
        RECT 85.950 879.600 88.050 880.050 ;
        RECT 58.950 878.400 88.050 879.600 ;
        RECT 101.400 878.400 106.050 880.050 ;
        RECT 52.950 877.950 57.000 878.400 ;
        RECT 58.950 877.800 61.050 878.400 ;
        RECT 79.950 877.800 82.050 878.400 ;
        RECT 85.950 877.950 88.050 878.400 ;
        RECT 102.000 877.950 106.050 878.400 ;
        RECT 130.950 879.600 133.050 879.900 ;
        RECT 148.950 879.600 151.050 879.900 ;
        RECT 130.950 879.450 151.050 879.600 ;
        RECT 154.950 879.450 157.050 879.900 ;
        RECT 130.950 878.400 157.050 879.450 ;
        RECT 130.950 877.800 133.050 878.400 ;
        RECT 148.950 878.250 157.050 878.400 ;
        RECT 148.950 877.800 151.050 878.250 ;
        RECT 154.950 877.800 157.050 878.250 ;
        RECT 158.400 877.050 159.600 884.100 ;
        RECT 161.400 879.900 162.600 886.950 ;
        RECT 175.950 885.600 178.050 886.200 ;
        RECT 187.950 885.600 190.050 886.050 ;
        RECT 205.950 885.600 208.050 886.050 ;
        RECT 175.950 884.400 208.050 885.600 ;
        RECT 175.950 884.100 178.050 884.400 ;
        RECT 187.950 883.950 190.050 884.400 ;
        RECT 205.950 883.950 208.050 884.400 ;
        RECT 214.950 884.100 217.050 886.200 ;
        RECT 259.950 885.600 262.050 886.200 ;
        RECT 277.950 885.600 280.050 886.200 ;
        RECT 259.950 884.400 280.050 885.600 ;
        RECT 259.950 884.100 262.050 884.400 ;
        RECT 277.950 884.100 280.050 884.400 ;
        RECT 310.950 885.750 313.050 886.200 ;
        RECT 316.950 885.750 319.050 886.200 ;
        RECT 310.950 884.550 319.050 885.750 ;
        RECT 310.950 884.100 313.050 884.550 ;
        RECT 316.950 884.100 319.050 884.550 ;
        RECT 322.950 884.100 325.050 886.200 ;
        RECT 343.950 885.600 346.050 886.200 ;
        RECT 361.950 885.750 364.050 886.200 ;
        RECT 376.950 885.750 379.050 886.200 ;
        RECT 343.950 884.400 360.600 885.600 ;
        RECT 343.950 884.100 346.050 884.400 ;
        RECT 160.950 877.800 163.050 879.900 ;
        RECT 166.950 879.450 169.050 879.900 ;
        RECT 178.950 879.450 181.050 879.900 ;
        RECT 166.950 878.250 181.050 879.450 ;
        RECT 166.950 877.800 169.050 878.250 ;
        RECT 178.950 877.800 181.050 878.250 ;
        RECT 187.950 879.450 190.050 879.900 ;
        RECT 193.950 879.450 196.050 879.900 ;
        RECT 187.950 878.250 196.050 879.450 ;
        RECT 187.950 877.800 190.050 878.250 ;
        RECT 193.950 877.800 196.050 878.250 ;
        RECT 199.950 879.600 202.050 879.900 ;
        RECT 215.400 879.600 216.600 884.100 ;
        RECT 199.950 878.400 216.600 879.600 ;
        RECT 229.950 879.450 232.050 879.900 ;
        RECT 235.950 879.450 238.050 879.900 ;
        RECT 199.950 877.800 202.050 878.400 ;
        RECT 229.950 878.250 238.050 879.450 ;
        RECT 229.950 877.800 232.050 878.250 ;
        RECT 235.950 877.800 238.050 878.250 ;
        RECT 298.950 879.600 301.050 879.900 ;
        RECT 310.950 879.600 313.050 880.050 ;
        RECT 298.950 878.400 313.050 879.600 ;
        RECT 323.400 879.600 324.600 884.100 ;
        RECT 359.400 879.900 360.600 884.400 ;
        RECT 361.950 884.550 379.050 885.750 ;
        RECT 361.950 884.100 364.050 884.550 ;
        RECT 376.950 884.100 379.050 884.550 ;
        RECT 412.950 885.750 415.050 886.200 ;
        RECT 421.950 885.750 424.050 886.200 ;
        RECT 412.950 884.550 424.050 885.750 ;
        RECT 412.950 884.100 415.050 884.550 ;
        RECT 421.950 884.100 424.050 884.550 ;
        RECT 427.950 885.600 430.050 886.050 ;
        RECT 469.950 885.750 472.050 886.200 ;
        RECT 475.950 885.750 478.050 886.200 ;
        RECT 469.950 885.600 478.050 885.750 ;
        RECT 427.950 884.550 478.050 885.600 ;
        RECT 427.950 884.400 472.050 884.550 ;
        RECT 427.950 883.950 430.050 884.400 ;
        RECT 469.950 884.100 472.050 884.400 ;
        RECT 475.950 884.100 478.050 884.550 ;
        RECT 496.950 885.750 499.050 886.200 ;
        RECT 505.950 885.750 508.050 886.200 ;
        RECT 496.950 884.550 508.050 885.750 ;
        RECT 496.950 884.100 499.050 884.550 ;
        RECT 505.950 884.100 508.050 884.550 ;
        RECT 511.950 883.950 514.050 886.050 ;
        RECT 523.950 885.600 526.050 886.200 ;
        RECT 535.950 885.600 538.050 886.200 ;
        RECT 523.950 884.400 538.050 885.600 ;
        RECT 523.950 884.100 526.050 884.400 ;
        RECT 535.950 884.100 538.050 884.400 ;
        RECT 541.950 885.750 544.050 886.200 ;
        RECT 547.950 885.750 550.050 886.200 ;
        RECT 541.950 884.550 550.050 885.750 ;
        RECT 541.950 884.100 544.050 884.550 ;
        RECT 547.950 884.100 550.050 884.550 ;
        RECT 580.950 885.600 583.050 886.200 ;
        RECT 586.950 885.600 589.050 886.050 ;
        RECT 580.950 884.400 589.050 885.600 ;
        RECT 580.950 884.100 583.050 884.400 ;
        RECT 586.950 883.950 589.050 884.400 ;
        RECT 622.950 885.750 625.050 886.200 ;
        RECT 697.950 885.750 700.050 886.200 ;
        RECT 622.950 884.550 700.050 885.750 ;
        RECT 622.950 884.100 625.050 884.550 ;
        RECT 697.950 884.100 700.050 884.550 ;
        RECT 742.950 885.600 745.050 886.050 ;
        RECT 754.950 885.600 757.050 886.200 ;
        RECT 742.950 884.400 757.050 885.600 ;
        RECT 742.950 883.950 745.050 884.400 ;
        RECT 754.950 884.100 757.050 884.400 ;
        RECT 781.950 885.600 784.050 886.200 ;
        RECT 805.950 885.750 808.050 886.200 ;
        RECT 814.950 885.750 817.050 886.200 ;
        RECT 781.950 884.400 804.600 885.600 ;
        RECT 781.950 884.100 784.050 884.400 ;
        RECT 334.950 879.600 337.050 879.900 ;
        RECT 323.400 878.400 337.050 879.600 ;
        RECT 298.950 877.800 301.050 878.400 ;
        RECT 310.950 877.950 313.050 878.400 ;
        RECT 334.950 877.800 337.050 878.400 ;
        RECT 340.950 879.450 343.050 879.900 ;
        RECT 352.950 879.450 355.050 879.900 ;
        RECT 340.950 878.250 355.050 879.450 ;
        RECT 340.950 877.800 343.050 878.250 ;
        RECT 352.950 877.800 355.050 878.250 ;
        RECT 358.950 877.800 361.050 879.900 ;
        RECT 364.950 879.600 367.050 879.900 ;
        RECT 379.950 879.600 382.050 880.050 ;
        RECT 364.950 878.400 382.050 879.600 ;
        RECT 364.950 877.800 367.050 878.400 ;
        RECT 379.950 877.950 382.050 878.400 ;
        RECT 484.950 879.450 487.050 879.900 ;
        RECT 493.950 879.450 496.050 879.900 ;
        RECT 484.950 878.250 496.050 879.450 ;
        RECT 512.400 879.600 513.600 883.950 ;
        RECT 628.950 881.100 631.050 883.200 ;
        RECT 664.950 882.600 667.050 882.900 ;
        RECT 685.950 882.600 688.050 883.050 ;
        RECT 664.950 881.400 688.050 882.600 ;
        RECT 514.950 879.600 517.050 879.900 ;
        RECT 512.400 878.400 517.050 879.600 ;
        RECT 484.950 877.800 487.050 878.250 ;
        RECT 493.950 877.800 496.050 878.250 ;
        RECT 514.950 877.800 517.050 878.400 ;
        RECT 520.950 879.600 523.050 879.900 ;
        RECT 547.950 879.600 550.050 880.050 ;
        RECT 520.950 878.400 550.050 879.600 ;
        RECT 520.950 877.800 523.050 878.400 ;
        RECT 547.950 877.950 550.050 878.400 ;
        RECT 586.950 879.450 589.050 879.900 ;
        RECT 595.950 879.450 598.050 879.900 ;
        RECT 586.950 878.250 598.050 879.450 ;
        RECT 586.950 877.800 589.050 878.250 ;
        RECT 595.950 877.800 598.050 878.250 ;
        RECT 607.950 879.450 610.050 879.900 ;
        RECT 619.950 879.600 622.050 879.900 ;
        RECT 629.400 879.600 630.600 881.100 ;
        RECT 664.950 880.800 667.050 881.400 ;
        RECT 685.950 880.950 688.050 881.400 ;
        RECT 691.950 880.950 694.050 883.050 ;
        RECT 803.400 882.600 804.600 884.400 ;
        RECT 805.950 884.550 817.050 885.750 ;
        RECT 829.950 885.600 832.050 886.050 ;
        RECT 805.950 884.100 808.050 884.550 ;
        RECT 814.950 884.100 817.050 884.550 ;
        RECT 818.400 884.400 832.050 885.600 ;
        RECT 803.400 882.000 813.600 882.600 ;
        RECT 803.400 881.400 814.050 882.000 ;
        RECT 619.950 879.450 630.600 879.600 ;
        RECT 607.950 878.400 630.600 879.450 ;
        RECT 607.950 878.250 622.050 878.400 ;
        RECT 607.950 877.800 610.050 878.250 ;
        RECT 619.950 877.800 622.050 878.250 ;
        RECT 124.950 876.600 127.050 877.050 ;
        RECT 136.950 876.600 139.050 877.050 ;
        RECT 124.950 875.400 139.050 876.600 ;
        RECT 124.950 874.950 127.050 875.400 ;
        RECT 136.950 874.950 139.050 875.400 ;
        RECT 157.950 874.950 160.050 877.050 ;
        RECT 205.950 876.600 208.050 877.050 ;
        RECT 217.950 876.600 220.050 877.050 ;
        RECT 205.950 875.400 220.050 876.600 ;
        RECT 205.950 874.950 208.050 875.400 ;
        RECT 217.950 874.950 220.050 875.400 ;
        RECT 370.950 876.600 373.050 877.050 ;
        RECT 385.950 876.600 388.050 877.050 ;
        RECT 370.950 875.400 388.050 876.600 ;
        RECT 370.950 874.950 373.050 875.400 ;
        RECT 385.950 874.950 388.050 875.400 ;
        RECT 397.950 876.600 400.050 877.050 ;
        RECT 409.950 876.600 412.050 877.050 ;
        RECT 397.950 875.400 412.050 876.600 ;
        RECT 397.950 874.950 400.050 875.400 ;
        RECT 409.950 874.950 412.050 875.400 ;
        RECT 433.950 876.600 436.050 877.050 ;
        RECT 466.950 876.600 469.050 877.050 ;
        RECT 433.950 875.400 469.050 876.600 ;
        RECT 433.950 874.950 436.050 875.400 ;
        RECT 466.950 874.950 469.050 875.400 ;
        RECT 502.950 876.600 505.050 877.050 ;
        RECT 679.950 876.600 682.050 877.050 ;
        RECT 502.950 875.400 682.050 876.600 ;
        RECT 502.950 874.950 505.050 875.400 ;
        RECT 679.950 874.950 682.050 875.400 ;
        RECT 685.950 876.600 688.050 877.050 ;
        RECT 692.400 876.600 693.600 880.950 ;
        RECT 712.950 879.450 715.050 879.900 ;
        RECT 718.950 879.450 721.050 879.900 ;
        RECT 712.950 878.250 721.050 879.450 ;
        RECT 712.950 877.800 715.050 878.250 ;
        RECT 718.950 877.800 721.050 878.250 ;
        RECT 745.950 879.450 748.050 879.900 ;
        RECT 772.950 879.450 775.050 879.900 ;
        RECT 745.950 878.250 775.050 879.450 ;
        RECT 745.950 877.800 748.050 878.250 ;
        RECT 772.950 877.800 775.050 878.250 ;
        RECT 787.950 879.600 790.050 880.050 ;
        RECT 796.950 879.600 799.050 879.900 ;
        RECT 787.950 878.400 799.050 879.600 ;
        RECT 787.950 877.950 790.050 878.400 ;
        RECT 796.950 877.800 799.050 878.400 ;
        RECT 811.950 877.950 814.050 881.400 ;
        RECT 818.400 879.900 819.600 884.400 ;
        RECT 829.950 883.950 832.050 884.400 ;
        RECT 835.950 885.600 838.050 886.050 ;
        RECT 841.950 885.600 844.050 886.050 ;
        RECT 835.950 884.400 844.050 885.600 ;
        RECT 835.950 883.950 838.050 884.400 ;
        RECT 841.950 883.950 844.050 884.400 ;
        RECT 853.950 885.750 856.050 886.200 ;
        RECT 862.950 885.750 865.050 886.200 ;
        RECT 853.950 884.550 865.050 885.750 ;
        RECT 853.950 884.100 856.050 884.550 ;
        RECT 862.950 884.100 865.050 884.550 ;
        RECT 886.950 884.100 889.050 886.200 ;
        RECT 922.950 885.600 925.050 886.050 ;
        RECT 928.950 885.600 931.050 886.200 ;
        RECT 922.950 884.400 931.050 885.600 ;
        RECT 887.400 882.600 888.600 884.100 ;
        RECT 922.950 883.950 925.050 884.400 ;
        RECT 928.950 884.100 931.050 884.400 ;
        RECT 887.400 881.400 891.600 882.600 ;
        RECT 817.950 877.800 820.050 879.900 ;
        RECT 844.950 879.600 847.050 879.900 ;
        RECT 877.950 879.600 880.050 880.050 ;
        RECT 883.950 879.600 886.050 879.900 ;
        RECT 844.950 878.400 886.050 879.600 ;
        RECT 890.400 879.600 891.600 881.400 ;
        RECT 913.950 879.600 916.050 879.900 ;
        RECT 890.400 878.400 916.050 879.600 ;
        RECT 844.950 877.800 847.050 878.400 ;
        RECT 877.950 877.950 880.050 878.400 ;
        RECT 883.950 877.800 886.050 878.400 ;
        RECT 913.950 877.800 916.050 878.400 ;
        RECT 685.950 875.400 693.600 876.600 ;
        RECT 685.950 874.950 688.050 875.400 ;
        RECT 40.950 873.600 43.050 874.050 ;
        RECT 64.950 873.600 67.050 874.050 ;
        RECT 40.950 872.400 67.050 873.600 ;
        RECT 40.950 871.950 43.050 872.400 ;
        RECT 64.950 871.950 67.050 872.400 ;
        RECT 73.950 873.600 76.050 874.050 ;
        RECT 109.950 873.600 112.050 874.050 ;
        RECT 73.950 872.400 112.050 873.600 ;
        RECT 73.950 871.950 76.050 872.400 ;
        RECT 109.950 871.950 112.050 872.400 ;
        RECT 154.950 873.600 157.050 874.050 ;
        RECT 172.950 873.600 175.050 874.050 ;
        RECT 154.950 872.400 175.050 873.600 ;
        RECT 154.950 871.950 157.050 872.400 ;
        RECT 172.950 871.950 175.050 872.400 ;
        RECT 220.950 873.600 223.050 874.050 ;
        RECT 256.950 873.600 259.050 874.050 ;
        RECT 289.950 873.600 292.050 874.050 ;
        RECT 337.950 873.600 340.050 874.050 ;
        RECT 220.950 872.400 340.050 873.600 ;
        RECT 220.950 871.950 223.050 872.400 ;
        RECT 256.950 871.950 259.050 872.400 ;
        RECT 289.950 871.950 292.050 872.400 ;
        RECT 337.950 871.950 340.050 872.400 ;
        RECT 349.950 873.600 352.050 874.050 ;
        RECT 403.950 873.600 406.050 874.050 ;
        RECT 349.950 872.400 406.050 873.600 ;
        RECT 349.950 871.950 352.050 872.400 ;
        RECT 403.950 871.950 406.050 872.400 ;
        RECT 469.950 873.600 472.050 874.050 ;
        RECT 496.950 873.600 499.050 874.050 ;
        RECT 469.950 872.400 499.050 873.600 ;
        RECT 469.950 871.950 472.050 872.400 ;
        RECT 496.950 871.950 499.050 872.400 ;
        RECT 547.950 873.600 550.050 874.050 ;
        RECT 601.950 873.600 604.050 874.050 ;
        RECT 613.950 873.600 616.050 874.050 ;
        RECT 547.950 872.400 616.050 873.600 ;
        RECT 680.400 873.600 681.600 874.950 ;
        RECT 784.950 873.600 787.050 874.050 ;
        RECT 841.950 873.600 844.050 874.050 ;
        RECT 680.400 872.400 844.050 873.600 ;
        RECT 547.950 871.950 550.050 872.400 ;
        RECT 601.950 871.950 604.050 872.400 ;
        RECT 613.950 871.950 616.050 872.400 ;
        RECT 784.950 871.950 787.050 872.400 ;
        RECT 841.950 871.950 844.050 872.400 ;
        RECT 868.950 873.600 871.050 874.050 ;
        RECT 889.950 873.600 892.050 874.050 ;
        RECT 868.950 872.400 892.050 873.600 ;
        RECT 868.950 871.950 871.050 872.400 ;
        RECT 889.950 871.950 892.050 872.400 ;
        RECT 22.950 870.600 25.050 871.050 ;
        RECT 52.950 870.600 55.050 871.050 ;
        RECT 22.950 869.400 55.050 870.600 ;
        RECT 65.400 870.600 66.600 871.950 ;
        RECT 118.950 870.600 121.050 871.050 ;
        RECT 65.400 869.400 121.050 870.600 ;
        RECT 22.950 868.950 25.050 869.400 ;
        RECT 52.950 868.950 55.050 869.400 ;
        RECT 118.950 868.950 121.050 869.400 ;
        RECT 409.950 870.600 412.050 871.050 ;
        RECT 460.950 870.600 463.050 871.050 ;
        RECT 409.950 869.400 463.050 870.600 ;
        RECT 409.950 868.950 412.050 869.400 ;
        RECT 460.950 868.950 463.050 869.400 ;
        RECT 538.950 870.600 541.050 871.050 ;
        RECT 577.950 870.600 580.050 871.050 ;
        RECT 538.950 869.400 580.050 870.600 ;
        RECT 538.950 868.950 541.050 869.400 ;
        RECT 577.950 868.950 580.050 869.400 ;
        RECT 682.950 870.600 685.050 871.050 ;
        RECT 694.950 870.600 697.050 871.050 ;
        RECT 682.950 869.400 697.050 870.600 ;
        RECT 682.950 868.950 685.050 869.400 ;
        RECT 694.950 868.950 697.050 869.400 ;
        RECT 706.950 870.600 709.050 871.050 ;
        RECT 730.950 870.600 733.050 871.050 ;
        RECT 706.950 869.400 733.050 870.600 ;
        RECT 706.950 868.950 709.050 869.400 ;
        RECT 730.950 868.950 733.050 869.400 ;
        RECT 751.950 870.600 754.050 871.050 ;
        RECT 796.950 870.600 799.050 871.050 ;
        RECT 751.950 869.400 799.050 870.600 ;
        RECT 751.950 868.950 754.050 869.400 ;
        RECT 796.950 868.950 799.050 869.400 ;
        RECT 811.950 870.600 814.050 871.050 ;
        RECT 853.950 870.600 856.050 871.050 ;
        RECT 811.950 869.400 856.050 870.600 ;
        RECT 811.950 868.950 814.050 869.400 ;
        RECT 853.950 868.950 856.050 869.400 ;
        RECT 43.950 867.600 46.050 868.050 ;
        RECT 73.950 867.600 76.050 868.050 ;
        RECT 43.950 866.400 76.050 867.600 ;
        RECT 43.950 865.950 46.050 866.400 ;
        RECT 73.950 865.950 76.050 866.400 ;
        RECT 157.950 867.600 160.050 868.050 ;
        RECT 220.950 867.600 223.050 868.050 ;
        RECT 157.950 866.400 223.050 867.600 ;
        RECT 157.950 865.950 160.050 866.400 ;
        RECT 220.950 865.950 223.050 866.400 ;
        RECT 334.950 867.600 337.050 868.050 ;
        RECT 373.950 867.600 376.050 868.050 ;
        RECT 469.950 867.600 472.050 868.050 ;
        RECT 757.950 867.600 760.050 868.050 ;
        RECT 808.950 867.600 811.050 868.050 ;
        RECT 334.950 866.400 811.050 867.600 ;
        RECT 334.950 865.950 337.050 866.400 ;
        RECT 373.950 865.950 376.050 866.400 ;
        RECT 469.950 865.950 472.050 866.400 ;
        RECT 757.950 865.950 760.050 866.400 ;
        RECT 808.950 865.950 811.050 866.400 ;
        RECT 337.950 864.600 340.050 865.050 ;
        RECT 409.950 864.600 412.050 865.050 ;
        RECT 337.950 863.400 412.050 864.600 ;
        RECT 337.950 862.950 340.050 863.400 ;
        RECT 409.950 862.950 412.050 863.400 ;
        RECT 433.950 864.600 436.050 865.050 ;
        RECT 463.950 864.600 466.050 865.050 ;
        RECT 433.950 863.400 466.050 864.600 ;
        RECT 433.950 862.950 436.050 863.400 ;
        RECT 463.950 862.950 466.050 863.400 ;
        RECT 694.950 864.600 697.050 865.050 ;
        RECT 805.950 864.600 808.050 865.050 ;
        RECT 835.950 864.600 838.050 865.050 ;
        RECT 694.950 863.400 838.050 864.600 ;
        RECT 694.950 862.950 697.050 863.400 ;
        RECT 805.950 862.950 808.050 863.400 ;
        RECT 835.950 862.950 838.050 863.400 ;
        RECT 97.950 861.600 100.050 862.050 ;
        RECT 154.950 861.600 157.050 862.050 ;
        RECT 97.950 860.400 157.050 861.600 ;
        RECT 97.950 859.950 100.050 860.400 ;
        RECT 154.950 859.950 157.050 860.400 ;
        RECT 430.950 861.600 433.050 862.050 ;
        RECT 478.950 861.600 481.050 862.050 ;
        RECT 430.950 860.400 481.050 861.600 ;
        RECT 430.950 859.950 433.050 860.400 ;
        RECT 478.950 859.950 481.050 860.400 ;
        RECT 547.950 861.600 550.050 862.050 ;
        RECT 637.950 861.600 640.050 862.050 ;
        RECT 547.950 860.400 640.050 861.600 ;
        RECT 547.950 859.950 550.050 860.400 ;
        RECT 637.950 859.950 640.050 860.400 ;
        RECT 643.950 861.600 646.050 862.050 ;
        RECT 673.950 861.600 676.050 862.050 ;
        RECT 643.950 860.400 676.050 861.600 ;
        RECT 643.950 859.950 646.050 860.400 ;
        RECT 673.950 859.950 676.050 860.400 ;
        RECT 58.950 858.600 61.050 859.050 ;
        RECT 67.950 858.600 70.050 859.050 ;
        RECT 91.950 858.600 94.050 859.050 ;
        RECT 58.950 857.400 94.050 858.600 ;
        RECT 58.950 856.950 61.050 857.400 ;
        RECT 67.950 856.950 70.050 857.400 ;
        RECT 91.950 856.950 94.050 857.400 ;
        RECT 367.950 858.600 370.050 859.050 ;
        RECT 427.950 858.600 430.050 859.050 ;
        RECT 784.950 858.600 787.050 859.050 ;
        RECT 823.950 858.600 826.050 859.050 ;
        RECT 874.950 858.600 877.050 859.050 ;
        RECT 367.950 857.400 430.050 858.600 ;
        RECT 367.950 856.950 370.050 857.400 ;
        RECT 427.950 856.950 430.050 857.400 ;
        RECT 533.400 857.400 687.600 858.600 ;
        RECT 463.950 855.600 466.050 856.050 ;
        RECT 533.400 855.600 534.600 857.400 ;
        RECT 463.950 854.400 534.600 855.600 ;
        RECT 553.950 855.600 556.050 856.050 ;
        RECT 613.950 855.600 616.050 856.050 ;
        RECT 553.950 854.400 616.050 855.600 ;
        RECT 686.400 855.600 687.600 857.400 ;
        RECT 784.950 857.400 877.050 858.600 ;
        RECT 784.950 856.950 787.050 857.400 ;
        RECT 823.950 856.950 826.050 857.400 ;
        RECT 874.950 856.950 877.050 857.400 ;
        RECT 718.950 855.600 721.050 856.050 ;
        RECT 686.400 854.400 721.050 855.600 ;
        RECT 463.950 853.950 466.050 854.400 ;
        RECT 553.950 853.950 556.050 854.400 ;
        RECT 613.950 853.950 616.050 854.400 ;
        RECT 718.950 853.950 721.050 854.400 ;
        RECT 751.950 855.600 754.050 856.050 ;
        RECT 772.950 855.600 775.050 856.050 ;
        RECT 751.950 854.400 885.600 855.600 ;
        RECT 751.950 853.950 754.050 854.400 ;
        RECT 772.950 853.950 775.050 854.400 ;
        RECT 884.400 853.050 885.600 854.400 ;
        RECT 52.950 852.600 55.050 853.050 ;
        RECT 73.950 852.600 76.050 853.050 ;
        RECT 103.950 852.600 106.050 853.050 ;
        RECT 52.950 851.400 106.050 852.600 ;
        RECT 52.950 850.950 55.050 851.400 ;
        RECT 73.950 850.950 76.050 851.400 ;
        RECT 103.950 850.950 106.050 851.400 ;
        RECT 199.950 852.600 202.050 853.050 ;
        RECT 439.950 852.600 442.050 853.050 ;
        RECT 199.950 851.400 442.050 852.600 ;
        RECT 199.950 850.950 202.050 851.400 ;
        RECT 439.950 850.950 442.050 851.400 ;
        RECT 637.950 852.600 640.050 853.050 ;
        RECT 694.950 852.600 697.050 853.050 ;
        RECT 637.950 851.400 697.050 852.600 ;
        RECT 637.950 850.950 640.050 851.400 ;
        RECT 694.950 850.950 697.050 851.400 ;
        RECT 760.950 852.600 763.050 853.050 ;
        RECT 784.950 852.600 787.050 853.050 ;
        RECT 760.950 851.400 787.050 852.600 ;
        RECT 760.950 850.950 763.050 851.400 ;
        RECT 784.950 850.950 787.050 851.400 ;
        RECT 817.950 852.600 820.050 853.050 ;
        RECT 850.950 852.600 853.050 853.050 ;
        RECT 817.950 851.400 853.050 852.600 ;
        RECT 817.950 850.950 820.050 851.400 ;
        RECT 850.950 850.950 853.050 851.400 ;
        RECT 883.950 852.600 886.050 853.050 ;
        RECT 922.950 852.600 925.050 853.050 ;
        RECT 883.950 851.400 925.050 852.600 ;
        RECT 883.950 850.950 886.050 851.400 ;
        RECT 922.950 850.950 925.050 851.400 ;
        RECT 394.950 849.600 397.050 850.050 ;
        RECT 406.950 849.600 409.050 850.050 ;
        RECT 394.950 848.400 409.050 849.600 ;
        RECT 394.950 847.950 397.050 848.400 ;
        RECT 406.950 847.950 409.050 848.400 ;
        RECT 589.950 849.600 592.050 850.050 ;
        RECT 628.950 849.600 631.050 850.050 ;
        RECT 589.950 848.400 631.050 849.600 ;
        RECT 589.950 847.950 592.050 848.400 ;
        RECT 628.950 847.950 631.050 848.400 ;
        RECT 634.950 849.600 637.050 850.050 ;
        RECT 700.950 849.600 703.050 850.050 ;
        RECT 724.950 849.600 727.050 850.050 ;
        RECT 634.950 848.400 727.050 849.600 ;
        RECT 634.950 847.950 637.050 848.400 ;
        RECT 700.950 847.950 703.050 848.400 ;
        RECT 724.950 847.950 727.050 848.400 ;
        RECT 787.950 849.600 790.050 850.050 ;
        RECT 832.950 849.600 835.050 850.050 ;
        RECT 862.950 849.600 865.050 850.050 ;
        RECT 904.950 849.600 907.050 850.050 ;
        RECT 787.950 848.400 907.050 849.600 ;
        RECT 787.950 847.950 790.050 848.400 ;
        RECT 832.950 847.950 835.050 848.400 ;
        RECT 862.950 847.950 865.050 848.400 ;
        RECT 904.950 847.950 907.050 848.400 ;
        RECT 64.950 846.600 67.050 847.050 ;
        RECT 88.950 846.600 91.050 847.050 ;
        RECT 196.950 846.600 199.050 847.050 ;
        RECT 64.950 845.400 91.050 846.600 ;
        RECT 64.950 844.950 67.050 845.400 ;
        RECT 88.950 844.950 91.050 845.400 ;
        RECT 107.400 845.400 199.050 846.600 ;
        RECT 16.950 840.750 19.050 841.200 ;
        RECT 28.950 840.750 31.050 841.200 ;
        RECT 16.950 839.550 31.050 840.750 ;
        RECT 16.950 839.100 19.050 839.550 ;
        RECT 28.950 839.100 31.050 839.550 ;
        RECT 40.950 839.100 43.050 841.200 ;
        RECT 19.950 834.600 22.050 834.900 ;
        RECT 41.400 834.600 42.600 839.100 ;
        RECT 46.950 838.950 49.050 841.050 ;
        RECT 76.950 840.750 79.050 841.200 ;
        RECT 82.950 840.750 85.050 841.200 ;
        RECT 76.950 839.550 85.050 840.750 ;
        RECT 76.950 839.100 79.050 839.550 ;
        RECT 82.950 839.100 85.050 839.550 ;
        RECT 88.950 840.750 91.050 841.200 ;
        RECT 97.950 840.750 100.050 841.200 ;
        RECT 88.950 839.550 100.050 840.750 ;
        RECT 88.950 839.100 91.050 839.550 ;
        RECT 97.950 839.100 100.050 839.550 ;
        RECT 47.400 835.050 48.600 838.950 ;
        RECT 72.000 837.600 76.050 838.050 ;
        RECT 71.400 835.950 76.050 837.600 ;
        RECT 19.950 833.400 42.600 834.600 ;
        RECT 19.950 832.800 22.050 833.400 ;
        RECT 46.950 832.950 49.050 835.050 ;
        RECT 61.950 834.600 64.050 834.900 ;
        RECT 71.400 834.600 72.600 835.950 ;
        RECT 107.400 834.900 108.600 845.400 ;
        RECT 196.950 844.950 199.050 845.400 ;
        RECT 214.950 846.600 217.050 847.050 ;
        RECT 271.950 846.600 274.050 847.050 ;
        RECT 214.950 845.400 274.050 846.600 ;
        RECT 214.950 844.950 217.050 845.400 ;
        RECT 271.950 844.950 274.050 845.400 ;
        RECT 280.950 846.600 283.050 847.050 ;
        RECT 295.950 846.600 298.050 847.050 ;
        RECT 280.950 845.400 298.050 846.600 ;
        RECT 280.950 844.950 283.050 845.400 ;
        RECT 295.950 844.950 298.050 845.400 ;
        RECT 319.950 846.600 322.050 847.050 ;
        RECT 334.950 846.600 337.050 847.050 ;
        RECT 319.950 845.400 337.050 846.600 ;
        RECT 319.950 844.950 322.050 845.400 ;
        RECT 334.950 844.950 337.050 845.400 ;
        RECT 445.950 846.600 448.050 847.050 ;
        RECT 487.950 846.600 490.050 847.050 ;
        RECT 445.950 845.400 490.050 846.600 ;
        RECT 445.950 844.950 448.050 845.400 ;
        RECT 487.950 844.950 490.050 845.400 ;
        RECT 577.950 846.600 580.050 847.050 ;
        RECT 694.950 846.600 697.050 847.050 ;
        RECT 778.950 846.600 781.050 847.050 ;
        RECT 577.950 845.400 697.050 846.600 ;
        RECT 577.950 844.950 580.050 845.400 ;
        RECT 694.950 844.950 697.050 845.400 ;
        RECT 740.400 845.400 781.050 846.600 ;
        RECT 397.950 843.600 400.050 844.050 ;
        RECT 433.950 843.600 436.050 844.050 ;
        RECT 397.950 842.400 436.050 843.600 ;
        RECT 397.950 841.950 400.050 842.400 ;
        RECT 433.950 841.950 436.050 842.400 ;
        RECT 685.950 841.950 688.050 844.050 ;
        RECT 718.950 843.600 721.050 844.050 ;
        RECT 740.400 843.600 741.600 845.400 ;
        RECT 778.950 844.950 781.050 845.400 ;
        RECT 718.950 842.400 741.600 843.600 ;
        RECT 832.950 843.600 835.050 844.050 ;
        RECT 841.950 843.600 844.050 844.200 ;
        RECT 832.950 842.400 844.050 843.600 ;
        RECT 718.950 841.950 721.050 842.400 ;
        RECT 832.950 841.950 835.050 842.400 ;
        RECT 841.950 842.100 844.050 842.400 ;
        RECT 895.950 843.600 898.050 844.050 ;
        RECT 904.950 843.600 907.050 844.050 ;
        RECT 895.950 842.400 907.050 843.600 ;
        RECT 895.950 841.950 898.050 842.400 ;
        RECT 904.950 841.950 907.050 842.400 ;
        RECT 109.950 839.100 112.050 841.200 ;
        RECT 115.950 840.750 118.050 841.200 ;
        RECT 121.950 840.750 124.050 841.200 ;
        RECT 115.950 839.550 124.050 840.750 ;
        RECT 115.950 839.100 118.050 839.550 ;
        RECT 121.950 839.100 124.050 839.550 ;
        RECT 127.950 839.100 130.050 841.200 ;
        RECT 148.950 840.600 151.050 841.200 ;
        RECT 157.950 840.600 160.050 841.050 ;
        RECT 148.950 839.400 160.050 840.600 ;
        RECT 148.950 839.100 151.050 839.400 ;
        RECT 110.400 837.600 111.600 839.100 ;
        RECT 128.400 837.600 129.600 839.100 ;
        RECT 157.950 838.950 160.050 839.400 ;
        RECT 190.950 840.600 193.050 841.200 ;
        RECT 208.950 840.600 211.050 841.200 ;
        RECT 190.950 839.400 211.050 840.600 ;
        RECT 190.950 839.100 193.050 839.400 ;
        RECT 208.950 839.100 211.050 839.400 ;
        RECT 232.950 840.600 235.050 841.200 ;
        RECT 244.950 840.600 247.050 841.050 ;
        RECT 232.950 839.400 247.050 840.600 ;
        RECT 232.950 839.100 235.050 839.400 ;
        RECT 244.950 838.950 247.050 839.400 ;
        RECT 262.950 840.750 265.050 841.200 ;
        RECT 271.950 840.750 274.050 841.200 ;
        RECT 262.950 839.550 274.050 840.750 ;
        RECT 262.950 839.100 265.050 839.550 ;
        RECT 271.950 839.100 274.050 839.550 ;
        RECT 280.950 840.600 283.050 841.200 ;
        RECT 292.950 840.600 295.050 841.050 ;
        RECT 319.950 840.600 322.050 841.200 ;
        RECT 280.950 839.400 288.600 840.600 ;
        RECT 280.950 839.100 283.050 839.400 ;
        RECT 287.400 837.600 288.600 839.400 ;
        RECT 292.950 839.400 322.050 840.600 ;
        RECT 292.950 838.950 295.050 839.400 ;
        RECT 319.950 839.100 322.050 839.400 ;
        RECT 325.800 839.100 327.900 841.200 ;
        RECT 343.950 840.600 346.050 841.200 ;
        RECT 355.950 840.750 358.050 841.200 ;
        RECT 361.950 840.750 364.050 841.200 ;
        RECT 343.950 839.400 354.600 840.600 ;
        RECT 343.950 839.100 346.050 839.400 ;
        RECT 110.400 836.400 114.600 837.600 ;
        RECT 128.400 836.400 180.600 837.600 ;
        RECT 287.400 836.400 303.600 837.600 ;
        RECT 61.950 833.400 72.600 834.600 ;
        RECT 61.950 832.800 64.050 833.400 ;
        RECT 106.950 832.800 109.050 834.900 ;
        RECT 113.400 834.600 114.600 836.400 ;
        RECT 179.400 835.050 180.600 836.400 ;
        RECT 124.950 834.600 127.050 834.900 ;
        RECT 113.400 833.400 127.050 834.600 ;
        RECT 124.950 832.800 127.050 833.400 ;
        RECT 178.950 834.600 181.050 835.050 ;
        RECT 302.400 834.900 303.600 836.400 ;
        RECT 205.950 834.600 208.050 834.900 ;
        RECT 178.950 833.400 208.050 834.600 ;
        RECT 178.950 832.950 181.050 833.400 ;
        RECT 205.950 832.800 208.050 833.400 ;
        RECT 211.950 834.450 214.050 834.900 ;
        RECT 244.950 834.450 247.050 834.900 ;
        RECT 211.950 833.250 247.050 834.450 ;
        RECT 211.950 832.800 214.050 833.250 ;
        RECT 244.950 832.800 247.050 833.250 ;
        RECT 301.950 832.800 304.050 834.900 ;
        RECT 22.950 831.600 25.050 832.050 ;
        RECT 31.950 831.600 34.050 832.050 ;
        RECT 22.950 830.400 34.050 831.600 ;
        RECT 22.950 829.950 25.050 830.400 ;
        RECT 31.950 829.950 34.050 830.400 ;
        RECT 43.950 831.600 46.050 832.050 ;
        RECT 52.950 831.600 55.050 832.050 ;
        RECT 85.950 831.600 88.050 832.050 ;
        RECT 43.950 830.400 88.050 831.600 ;
        RECT 43.950 829.950 46.050 830.400 ;
        RECT 52.950 829.950 55.050 830.400 ;
        RECT 85.950 829.950 88.050 830.400 ;
        RECT 283.950 831.600 286.050 832.050 ;
        RECT 295.950 831.600 298.050 832.050 ;
        RECT 283.950 830.400 298.050 831.600 ;
        RECT 326.400 831.600 327.600 839.100 ;
        RECT 353.400 837.600 354.600 839.400 ;
        RECT 355.950 839.550 364.050 840.750 ;
        RECT 355.950 839.100 358.050 839.550 ;
        RECT 361.950 839.100 364.050 839.550 ;
        RECT 373.950 840.600 376.050 841.050 ;
        RECT 385.950 840.600 388.050 841.200 ;
        RECT 373.950 839.400 381.600 840.600 ;
        RECT 373.950 838.950 376.050 839.400 ;
        RECT 380.400 837.600 381.600 839.400 ;
        RECT 385.950 839.400 432.600 840.600 ;
        RECT 385.950 839.100 388.050 839.400 ;
        RECT 394.950 837.600 397.050 838.050 ;
        RECT 431.400 837.600 432.600 839.400 ;
        RECT 436.950 839.100 439.050 841.200 ;
        RECT 454.950 840.750 457.050 841.200 ;
        RECT 478.950 840.750 481.050 841.200 ;
        RECT 454.950 839.550 481.050 840.750 ;
        RECT 454.950 839.100 457.050 839.550 ;
        RECT 478.950 839.100 481.050 839.550 ;
        RECT 529.950 840.600 532.050 841.200 ;
        RECT 535.800 840.600 537.900 841.050 ;
        RECT 529.950 839.400 537.900 840.600 ;
        RECT 529.950 839.100 532.050 839.400 ;
        RECT 353.400 836.400 378.600 837.600 ;
        RECT 380.400 836.400 387.600 837.600 ;
        RECT 349.950 834.600 352.050 835.050 ;
        RECT 355.950 834.600 358.050 835.050 ;
        RECT 349.950 833.400 358.050 834.600 ;
        RECT 377.400 834.600 378.600 836.400 ;
        RECT 382.950 834.600 385.050 834.900 ;
        RECT 377.400 833.400 385.050 834.600 ;
        RECT 386.400 834.600 387.600 836.400 ;
        RECT 394.950 836.400 429.600 837.600 ;
        RECT 431.400 836.400 435.600 837.600 ;
        RECT 394.950 835.950 397.050 836.400 ;
        RECT 428.400 834.900 429.600 836.400 ;
        RECT 434.400 834.900 435.600 836.400 ;
        RECT 437.400 835.050 438.600 839.100 ;
        RECT 535.800 838.950 537.900 839.400 ;
        RECT 538.950 840.600 541.050 841.050 ;
        RECT 547.950 840.600 550.050 841.200 ;
        RECT 538.950 839.400 550.050 840.600 ;
        RECT 538.950 838.950 541.050 839.400 ;
        RECT 547.950 839.100 550.050 839.400 ;
        RECT 568.950 840.600 571.050 841.200 ;
        RECT 583.950 840.600 586.050 841.200 ;
        RECT 568.950 839.400 586.050 840.600 ;
        RECT 568.950 839.100 571.050 839.400 ;
        RECT 583.950 839.100 586.050 839.400 ;
        RECT 610.950 840.600 613.050 841.050 ;
        RECT 619.950 840.600 622.050 841.200 ;
        RECT 610.950 839.400 622.050 840.600 ;
        RECT 610.950 838.950 613.050 839.400 ;
        RECT 619.950 839.100 622.050 839.400 ;
        RECT 637.950 840.600 640.050 841.050 ;
        RECT 652.950 840.600 655.050 841.050 ;
        RECT 637.950 839.400 655.050 840.600 ;
        RECT 637.950 838.950 640.050 839.400 ;
        RECT 652.950 838.950 655.050 839.400 ;
        RECT 686.400 838.050 687.600 841.950 ;
        RECT 697.950 840.750 700.050 841.200 ;
        RECT 712.950 840.750 715.050 841.200 ;
        RECT 697.950 839.550 715.050 840.750 ;
        RECT 697.950 839.100 700.050 839.550 ;
        RECT 712.950 839.100 715.050 839.550 ;
        RECT 739.950 840.750 742.050 841.200 ;
        RECT 766.950 840.750 769.050 841.200 ;
        RECT 739.950 839.550 769.050 840.750 ;
        RECT 739.950 839.100 742.050 839.550 ;
        RECT 766.950 839.100 769.050 839.550 ;
        RECT 871.950 840.600 874.050 841.050 ;
        RECT 889.950 840.750 892.050 841.200 ;
        RECT 901.950 840.750 904.050 841.200 ;
        RECT 889.950 840.600 904.050 840.750 ;
        RECT 871.950 839.550 904.050 840.600 ;
        RECT 871.950 839.400 892.050 839.550 ;
        RECT 871.950 838.950 874.050 839.400 ;
        RECT 889.950 839.100 892.050 839.400 ;
        RECT 901.950 839.100 904.050 839.550 ;
        RECT 685.950 835.950 688.050 838.050 ;
        RECT 691.950 837.600 694.050 838.050 ;
        RECT 736.950 837.600 739.050 838.050 ;
        RECT 691.950 836.400 739.050 837.600 ;
        RECT 691.950 835.950 694.050 836.400 ;
        RECT 736.950 835.950 739.050 836.400 ;
        RECT 409.950 834.600 412.050 834.900 ;
        RECT 386.400 833.400 412.050 834.600 ;
        RECT 349.950 832.950 352.050 833.400 ;
        RECT 355.950 832.950 358.050 833.400 ;
        RECT 382.950 832.800 385.050 833.400 ;
        RECT 409.950 832.800 412.050 833.400 ;
        RECT 427.950 832.800 430.050 834.900 ;
        RECT 433.950 832.800 436.050 834.900 ;
        RECT 437.400 833.400 442.050 835.050 ;
        RECT 438.000 832.950 442.050 833.400 ;
        RECT 445.950 834.450 448.050 834.900 ;
        RECT 451.950 834.450 454.050 834.900 ;
        RECT 445.950 833.250 454.050 834.450 ;
        RECT 445.950 832.800 448.050 833.250 ;
        RECT 451.950 832.800 454.050 833.250 ;
        RECT 463.950 834.450 466.050 834.900 ;
        RECT 472.950 834.450 475.050 834.900 ;
        RECT 463.950 833.250 475.050 834.450 ;
        RECT 463.950 832.800 466.050 833.250 ;
        RECT 472.950 832.800 475.050 833.250 ;
        RECT 478.950 834.600 481.050 835.050 ;
        RECT 526.950 834.600 529.050 834.900 ;
        RECT 478.950 833.400 529.050 834.600 ;
        RECT 478.950 832.950 481.050 833.400 ;
        RECT 526.950 832.800 529.050 833.400 ;
        RECT 541.950 834.600 544.050 834.900 ;
        RECT 565.950 834.600 568.050 834.900 ;
        RECT 541.950 833.400 568.050 834.600 ;
        RECT 541.950 832.800 544.050 833.400 ;
        RECT 565.950 832.800 568.050 833.400 ;
        RECT 709.950 834.600 712.050 834.900 ;
        RECT 748.950 834.600 751.050 834.900 ;
        RECT 709.950 833.400 751.050 834.600 ;
        RECT 709.950 832.800 712.050 833.400 ;
        RECT 748.950 832.800 751.050 833.400 ;
        RECT 775.950 834.600 778.050 834.900 ;
        RECT 787.950 834.600 790.050 835.050 ;
        RECT 775.950 833.400 790.050 834.600 ;
        RECT 775.950 832.800 778.050 833.400 ;
        RECT 787.950 832.950 790.050 833.400 ;
        RECT 850.950 834.450 853.050 834.900 ;
        RECT 859.950 834.450 862.050 834.900 ;
        RECT 850.950 833.250 862.050 834.450 ;
        RECT 850.950 832.800 853.050 833.250 ;
        RECT 859.950 832.800 862.050 833.250 ;
        RECT 865.950 834.450 868.050 834.900 ;
        RECT 871.800 834.450 873.900 834.900 ;
        RECT 865.950 833.250 873.900 834.450 ;
        RECT 865.950 832.800 868.050 833.250 ;
        RECT 871.800 832.800 873.900 833.250 ;
        RECT 874.950 834.450 877.050 834.900 ;
        RECT 907.950 834.450 910.050 834.900 ;
        RECT 874.950 833.250 910.050 834.450 ;
        RECT 874.950 832.800 877.050 833.250 ;
        RECT 907.950 832.800 910.050 833.250 ;
        RECT 337.950 831.600 340.050 832.050 ;
        RECT 326.400 830.400 340.050 831.600 ;
        RECT 283.950 829.950 286.050 830.400 ;
        RECT 295.950 829.950 298.050 830.400 ;
        RECT 337.950 829.950 340.050 830.400 ;
        RECT 370.950 831.600 373.050 832.050 ;
        RECT 376.950 831.600 379.050 832.050 ;
        RECT 370.950 830.400 379.050 831.600 ;
        RECT 370.950 829.950 373.050 830.400 ;
        RECT 376.950 829.950 379.050 830.400 ;
        RECT 475.950 831.600 478.050 832.050 ;
        RECT 490.950 831.600 493.050 832.050 ;
        RECT 475.950 830.400 493.050 831.600 ;
        RECT 475.950 829.950 478.050 830.400 ;
        RECT 490.950 829.950 493.050 830.400 ;
        RECT 586.950 831.600 589.050 832.050 ;
        RECT 604.950 831.600 607.050 832.050 ;
        RECT 622.950 831.600 625.050 832.050 ;
        RECT 691.950 831.600 694.050 832.050 ;
        RECT 586.950 830.400 694.050 831.600 ;
        RECT 586.950 829.950 589.050 830.400 ;
        RECT 604.950 829.950 607.050 830.400 ;
        RECT 622.950 829.950 625.050 830.400 ;
        RECT 691.950 829.950 694.050 830.400 ;
        RECT 13.950 828.600 16.050 829.050 ;
        RECT 28.950 828.600 31.050 828.900 ;
        RECT 13.950 827.400 31.050 828.600 ;
        RECT 13.950 826.950 16.050 827.400 ;
        RECT 28.950 826.800 31.050 827.400 ;
        RECT 67.950 828.600 70.050 829.050 ;
        RECT 79.950 828.600 82.050 829.050 ;
        RECT 67.950 827.400 82.050 828.600 ;
        RECT 67.950 826.950 70.050 827.400 ;
        RECT 79.950 826.950 82.050 827.400 ;
        RECT 118.950 828.600 121.050 829.050 ;
        RECT 130.950 828.600 133.050 829.050 ;
        RECT 145.950 828.600 148.050 829.050 ;
        RECT 118.950 827.400 148.050 828.600 ;
        RECT 118.950 826.950 121.050 827.400 ;
        RECT 130.950 826.950 133.050 827.400 ;
        RECT 145.950 826.950 148.050 827.400 ;
        RECT 166.950 828.600 169.050 829.050 ;
        RECT 199.950 828.600 202.050 829.050 ;
        RECT 166.950 827.400 202.050 828.600 ;
        RECT 166.950 826.950 169.050 827.400 ;
        RECT 199.950 826.950 202.050 827.400 ;
        RECT 253.950 828.600 256.050 829.050 ;
        RECT 265.950 828.600 268.050 829.050 ;
        RECT 253.950 827.400 268.050 828.600 ;
        RECT 253.950 826.950 256.050 827.400 ;
        RECT 265.950 826.950 268.050 827.400 ;
        RECT 277.950 828.600 280.050 829.050 ;
        RECT 292.950 828.600 295.050 829.050 ;
        RECT 277.950 827.400 295.050 828.600 ;
        RECT 277.950 826.950 280.050 827.400 ;
        RECT 292.950 826.950 295.050 827.400 ;
        RECT 307.950 828.600 310.050 829.050 ;
        RECT 340.950 828.600 343.050 829.050 ;
        RECT 307.950 827.400 343.050 828.600 ;
        RECT 307.950 826.950 310.050 827.400 ;
        RECT 340.950 826.950 343.050 827.400 ;
        RECT 397.950 828.600 400.050 828.900 ;
        RECT 409.950 828.600 412.050 829.050 ;
        RECT 397.950 827.400 412.050 828.600 ;
        RECT 397.950 826.800 400.050 827.400 ;
        RECT 409.950 826.950 412.050 827.400 ;
        RECT 457.950 828.600 460.050 829.050 ;
        RECT 508.950 828.600 511.050 829.050 ;
        RECT 457.950 827.400 511.050 828.600 ;
        RECT 457.950 826.950 460.050 827.400 ;
        RECT 508.950 826.950 511.050 827.400 ;
        RECT 727.950 828.600 730.050 829.050 ;
        RECT 760.950 828.600 763.050 829.050 ;
        RECT 727.950 827.400 763.050 828.600 ;
        RECT 727.950 826.950 730.050 827.400 ;
        RECT 760.950 826.950 763.050 827.400 ;
        RECT 769.950 828.600 772.050 829.050 ;
        RECT 880.950 828.600 883.050 829.050 ;
        RECT 769.950 827.400 883.050 828.600 ;
        RECT 769.950 826.950 772.050 827.400 ;
        RECT 880.950 826.950 883.050 827.400 ;
        RECT 37.950 825.600 40.050 826.050 ;
        RECT 46.950 825.600 49.050 826.050 ;
        RECT 37.950 824.400 49.050 825.600 ;
        RECT 37.950 823.950 40.050 824.400 ;
        RECT 46.950 823.950 49.050 824.400 ;
        RECT 454.950 825.600 457.050 826.050 ;
        RECT 487.950 825.600 490.050 826.050 ;
        RECT 454.950 824.400 490.050 825.600 ;
        RECT 454.950 823.950 457.050 824.400 ;
        RECT 487.950 823.950 490.050 824.400 ;
        RECT 565.950 825.600 568.050 826.050 ;
        RECT 571.950 825.600 574.050 826.050 ;
        RECT 565.950 824.400 574.050 825.600 ;
        RECT 565.950 823.950 568.050 824.400 ;
        RECT 571.950 823.950 574.050 824.400 ;
        RECT 610.950 825.600 613.050 826.050 ;
        RECT 736.950 825.600 739.050 826.050 ;
        RECT 781.950 825.600 784.050 826.050 ;
        RECT 610.950 824.400 657.600 825.600 ;
        RECT 610.950 823.950 613.050 824.400 ;
        RECT 656.400 823.050 657.600 824.400 ;
        RECT 736.950 824.400 784.050 825.600 ;
        RECT 736.950 823.950 739.050 824.400 ;
        RECT 781.950 823.950 784.050 824.400 ;
        RECT 82.950 822.600 85.050 823.050 ;
        RECT 97.950 822.600 100.050 823.050 ;
        RECT 82.950 821.400 100.050 822.600 ;
        RECT 82.950 820.950 85.050 821.400 ;
        RECT 97.950 820.950 100.050 821.400 ;
        RECT 322.950 822.600 325.050 823.050 ;
        RECT 340.950 822.600 343.050 823.050 ;
        RECT 322.950 821.400 343.050 822.600 ;
        RECT 322.950 820.950 325.050 821.400 ;
        RECT 340.950 820.950 343.050 821.400 ;
        RECT 352.950 822.600 355.050 823.050 ;
        RECT 445.950 822.600 448.050 823.050 ;
        RECT 352.950 821.400 448.050 822.600 ;
        RECT 352.950 820.950 355.050 821.400 ;
        RECT 445.950 820.950 448.050 821.400 ;
        RECT 451.950 822.600 454.050 823.050 ;
        RECT 460.950 822.600 463.050 823.050 ;
        RECT 451.950 821.400 463.050 822.600 ;
        RECT 451.950 820.950 454.050 821.400 ;
        RECT 460.950 820.950 463.050 821.400 ;
        RECT 490.950 822.600 493.050 823.050 ;
        RECT 529.950 822.600 532.050 823.050 ;
        RECT 490.950 821.400 532.050 822.600 ;
        RECT 490.950 820.950 493.050 821.400 ;
        RECT 529.950 820.950 532.050 821.400 ;
        RECT 535.950 822.600 538.050 823.050 ;
        RECT 628.950 822.600 631.050 823.050 ;
        RECT 535.950 821.400 631.050 822.600 ;
        RECT 656.400 821.400 661.050 823.050 ;
        RECT 535.950 820.950 538.050 821.400 ;
        RECT 628.950 820.950 631.050 821.400 ;
        RECT 657.000 820.950 661.050 821.400 ;
        RECT 673.950 822.600 676.050 823.050 ;
        RECT 679.950 822.600 682.050 823.050 ;
        RECT 712.950 822.600 715.050 823.050 ;
        RECT 673.950 821.400 715.050 822.600 ;
        RECT 673.950 820.950 676.050 821.400 ;
        RECT 679.950 820.950 682.050 821.400 ;
        RECT 712.950 820.950 715.050 821.400 ;
        RECT 796.950 822.600 799.050 823.050 ;
        RECT 886.950 822.600 889.050 823.050 ;
        RECT 796.950 821.400 889.050 822.600 ;
        RECT 796.950 820.950 799.050 821.400 ;
        RECT 886.950 820.950 889.050 821.400 ;
        RECT 70.950 819.600 73.050 820.050 ;
        RECT 112.950 819.600 115.050 820.050 ;
        RECT 70.950 818.400 115.050 819.600 ;
        RECT 70.950 817.950 73.050 818.400 ;
        RECT 112.950 817.950 115.050 818.400 ;
        RECT 334.950 819.600 337.050 820.050 ;
        RECT 373.950 819.600 376.050 820.050 ;
        RECT 334.950 818.400 376.050 819.600 ;
        RECT 334.950 817.950 337.050 818.400 ;
        RECT 373.950 817.950 376.050 818.400 ;
        RECT 379.950 819.600 382.050 820.050 ;
        RECT 457.950 819.600 460.050 820.050 ;
        RECT 379.950 818.400 460.050 819.600 ;
        RECT 379.950 817.950 382.050 818.400 ;
        RECT 457.950 817.950 460.050 818.400 ;
        RECT 463.950 819.600 466.050 820.050 ;
        RECT 475.950 819.600 478.050 820.050 ;
        RECT 463.950 818.400 478.050 819.600 ;
        RECT 463.950 817.950 466.050 818.400 ;
        RECT 475.950 817.950 478.050 818.400 ;
        RECT 487.950 819.600 490.050 820.050 ;
        RECT 535.950 819.600 538.050 819.900 ;
        RECT 487.950 818.400 538.050 819.600 ;
        RECT 487.950 817.950 490.050 818.400 ;
        RECT 535.950 817.800 538.050 818.400 ;
        RECT 724.950 819.600 727.050 820.050 ;
        RECT 745.950 819.600 748.050 820.050 ;
        RECT 775.950 819.600 778.050 820.050 ;
        RECT 790.950 819.600 793.050 820.050 ;
        RECT 724.950 818.400 795.600 819.600 ;
        RECT 724.950 817.950 727.050 818.400 ;
        RECT 745.950 817.950 748.050 818.400 ;
        RECT 775.950 817.950 778.050 818.400 ;
        RECT 790.950 817.950 793.050 818.400 ;
        RECT 16.950 816.600 19.050 817.050 ;
        RECT 22.950 816.600 25.050 817.050 ;
        RECT 16.950 815.400 25.050 816.600 ;
        RECT 16.950 814.950 19.050 815.400 ;
        RECT 22.950 814.950 25.050 815.400 ;
        RECT 175.950 816.600 178.050 817.050 ;
        RECT 235.950 816.600 238.050 817.050 ;
        RECT 175.950 815.400 238.050 816.600 ;
        RECT 175.950 814.950 178.050 815.400 ;
        RECT 235.950 814.950 238.050 815.400 ;
        RECT 271.950 816.600 274.050 817.050 ;
        RECT 334.950 816.600 337.050 816.900 ;
        RECT 271.950 815.400 337.050 816.600 ;
        RECT 271.950 814.950 274.050 815.400 ;
        RECT 334.950 814.800 337.050 815.400 ;
        RECT 406.950 816.600 409.050 817.050 ;
        RECT 556.950 816.600 559.050 817.050 ;
        RECT 406.950 815.400 559.050 816.600 ;
        RECT 406.950 814.950 409.050 815.400 ;
        RECT 556.950 814.950 559.050 815.400 ;
        RECT 658.950 816.600 661.050 817.050 ;
        RECT 769.950 816.600 772.050 817.050 ;
        RECT 658.950 815.400 772.050 816.600 ;
        RECT 794.400 816.600 795.600 818.400 ;
        RECT 886.950 816.600 889.050 817.050 ;
        RECT 794.400 815.400 889.050 816.600 ;
        RECT 658.950 814.950 661.050 815.400 ;
        RECT 769.950 814.950 772.050 815.400 ;
        RECT 886.950 814.950 889.050 815.400 ;
        RECT 46.950 813.600 49.050 814.050 ;
        RECT 55.950 813.600 58.050 814.050 ;
        RECT 46.950 812.400 58.050 813.600 ;
        RECT 46.950 811.950 49.050 812.400 ;
        RECT 55.950 811.950 58.050 812.400 ;
        RECT 94.950 813.600 97.050 814.050 ;
        RECT 115.950 813.600 118.050 814.050 ;
        RECT 127.950 813.600 130.050 814.050 ;
        RECT 94.950 812.400 130.050 813.600 ;
        RECT 94.950 811.950 97.050 812.400 ;
        RECT 115.950 811.950 118.050 812.400 ;
        RECT 127.950 811.950 130.050 812.400 ;
        RECT 157.950 813.600 160.050 814.050 ;
        RECT 166.950 813.600 169.050 814.050 ;
        RECT 157.950 812.400 169.050 813.600 ;
        RECT 157.950 811.950 160.050 812.400 ;
        RECT 166.950 811.950 169.050 812.400 ;
        RECT 322.950 813.600 325.050 814.050 ;
        RECT 397.950 813.600 400.050 814.050 ;
        RECT 322.950 812.400 400.050 813.600 ;
        RECT 322.950 811.950 325.050 812.400 ;
        RECT 397.950 811.950 400.050 812.400 ;
        RECT 445.950 813.600 448.050 814.050 ;
        RECT 502.950 813.600 505.050 814.050 ;
        RECT 445.950 812.400 505.050 813.600 ;
        RECT 445.950 811.950 448.050 812.400 ;
        RECT 502.950 811.950 505.050 812.400 ;
        RECT 514.950 813.600 517.050 814.050 ;
        RECT 547.950 813.600 550.050 814.050 ;
        RECT 514.950 812.400 550.050 813.600 ;
        RECT 514.950 811.950 517.050 812.400 ;
        RECT 547.950 811.950 550.050 812.400 ;
        RECT 613.950 813.600 616.050 814.050 ;
        RECT 649.950 813.600 652.050 814.050 ;
        RECT 613.950 812.400 652.050 813.600 ;
        RECT 613.950 811.950 616.050 812.400 ;
        RECT 649.950 811.950 652.050 812.400 ;
        RECT 661.950 813.600 664.050 814.050 ;
        RECT 673.950 813.600 676.050 814.050 ;
        RECT 709.950 813.600 712.050 814.050 ;
        RECT 661.950 812.400 712.050 813.600 ;
        RECT 661.950 811.950 664.050 812.400 ;
        RECT 673.950 811.950 676.050 812.400 ;
        RECT 709.950 811.950 712.050 812.400 ;
        RECT 895.950 813.600 898.050 814.050 ;
        RECT 925.950 813.600 928.050 814.050 ;
        RECT 895.950 812.400 928.050 813.600 ;
        RECT 895.950 811.950 898.050 812.400 ;
        RECT 925.950 811.950 928.050 812.400 ;
        RECT 40.950 810.600 43.050 811.050 ;
        RECT 88.950 810.600 91.050 811.050 ;
        RECT 136.950 810.600 139.050 811.050 ;
        RECT 178.950 810.600 181.050 811.050 ;
        RECT 184.950 810.600 187.050 811.050 ;
        RECT 40.950 809.400 187.050 810.600 ;
        RECT 40.950 808.950 43.050 809.400 ;
        RECT 88.950 808.950 91.050 809.400 ;
        RECT 136.950 808.950 139.050 809.400 ;
        RECT 178.950 808.950 181.050 809.400 ;
        RECT 184.950 808.950 187.050 809.400 ;
        RECT 334.950 810.600 337.050 811.050 ;
        RECT 394.950 810.600 397.050 811.050 ;
        RECT 334.950 809.400 397.050 810.600 ;
        RECT 334.950 808.950 337.050 809.400 ;
        RECT 394.950 808.950 397.050 809.400 ;
        RECT 439.950 808.950 442.050 811.050 ;
        RECT 460.950 810.600 463.050 811.050 ;
        RECT 505.950 810.600 508.050 811.050 ;
        RECT 583.950 810.600 586.050 811.050 ;
        RECT 460.950 809.400 483.600 810.600 ;
        RECT 460.950 808.950 463.050 809.400 ;
        RECT 1.950 807.750 4.050 808.200 ;
        RECT 22.950 807.750 25.050 808.200 ;
        RECT 1.950 807.600 25.050 807.750 ;
        RECT 40.950 807.600 43.050 808.200 ;
        RECT 1.950 806.550 43.050 807.600 ;
        RECT 1.950 806.100 4.050 806.550 ;
        RECT 22.950 806.400 43.050 806.550 ;
        RECT 22.950 806.100 25.050 806.400 ;
        RECT 40.950 806.100 43.050 806.400 ;
        RECT 58.950 807.750 61.050 808.200 ;
        RECT 76.950 807.750 79.050 808.200 ;
        RECT 58.950 806.550 79.050 807.750 ;
        RECT 58.950 806.100 61.050 806.550 ;
        RECT 76.950 806.100 79.050 806.550 ;
        RECT 106.950 807.750 109.050 808.200 ;
        RECT 112.950 807.750 115.050 808.200 ;
        RECT 106.950 806.550 115.050 807.750 ;
        RECT 106.950 806.100 109.050 806.550 ;
        RECT 112.950 806.100 115.050 806.550 ;
        RECT 145.950 807.750 148.050 808.200 ;
        RECT 160.950 807.750 163.050 808.200 ;
        RECT 145.950 806.550 163.050 807.750 ;
        RECT 145.950 806.100 148.050 806.550 ;
        RECT 160.950 806.100 163.050 806.550 ;
        RECT 190.950 807.600 193.050 808.200 ;
        RECT 199.950 807.750 202.050 808.200 ;
        RECT 205.950 807.750 208.050 808.200 ;
        RECT 190.950 806.400 198.600 807.600 ;
        RECT 190.950 806.100 193.050 806.400 ;
        RECT 197.400 804.600 198.600 806.400 ;
        RECT 199.950 806.550 208.050 807.750 ;
        RECT 199.950 806.100 202.050 806.550 ;
        RECT 205.950 806.100 208.050 806.550 ;
        RECT 211.950 807.600 214.050 808.200 ;
        RECT 229.950 807.600 232.050 808.200 ;
        RECT 211.950 806.400 232.050 807.600 ;
        RECT 211.950 806.100 214.050 806.400 ;
        RECT 229.950 806.100 232.050 806.400 ;
        RECT 244.950 807.750 247.050 808.200 ;
        RECT 250.950 807.750 253.050 808.200 ;
        RECT 244.950 806.550 253.050 807.750 ;
        RECT 244.950 806.100 247.050 806.550 ;
        RECT 250.950 806.100 253.050 806.550 ;
        RECT 277.950 807.600 280.050 808.200 ;
        RECT 313.950 807.600 316.050 808.200 ;
        RECT 277.950 806.400 316.050 807.600 ;
        RECT 277.950 806.100 280.050 806.400 ;
        RECT 313.950 806.100 316.050 806.400 ;
        RECT 337.950 807.600 340.050 808.050 ;
        RECT 355.950 807.750 358.050 808.200 ;
        RECT 361.950 807.750 364.050 808.200 ;
        RECT 355.950 807.600 364.050 807.750 ;
        RECT 403.950 807.600 406.050 808.050 ;
        RECT 337.950 806.550 364.050 807.600 ;
        RECT 337.950 806.400 358.050 806.550 ;
        RECT 337.950 805.950 340.050 806.400 ;
        RECT 355.950 806.100 358.050 806.400 ;
        RECT 361.950 806.100 364.050 806.550 ;
        RECT 395.400 806.400 406.050 807.600 ;
        RECT 197.400 803.400 207.600 804.600 ;
        RECT 28.950 801.450 31.050 801.900 ;
        RECT 37.950 801.450 40.050 801.900 ;
        RECT 28.950 800.250 40.050 801.450 ;
        RECT 28.950 799.800 31.050 800.250 ;
        RECT 37.950 799.800 40.050 800.250 ;
        RECT 55.950 801.450 58.050 801.900 ;
        RECT 61.950 801.450 64.050 801.900 ;
        RECT 55.950 800.250 64.050 801.450 ;
        RECT 55.950 799.800 58.050 800.250 ;
        RECT 61.950 799.800 64.050 800.250 ;
        RECT 121.950 801.450 124.050 801.900 ;
        RECT 127.950 801.450 130.050 801.900 ;
        RECT 121.950 800.250 130.050 801.450 ;
        RECT 121.950 799.800 124.050 800.250 ;
        RECT 127.950 799.800 130.050 800.250 ;
        RECT 151.950 801.600 154.050 802.050 ;
        RECT 163.950 801.600 166.050 801.900 ;
        RECT 151.950 800.400 166.050 801.600 ;
        RECT 151.950 799.950 154.050 800.400 ;
        RECT 163.950 799.800 166.050 800.400 ;
        RECT 169.950 801.450 172.050 801.900 ;
        RECT 175.950 801.450 178.050 801.900 ;
        RECT 169.950 800.250 178.050 801.450 ;
        RECT 169.950 799.800 172.050 800.250 ;
        RECT 175.950 799.800 178.050 800.250 ;
        RECT 193.950 801.600 196.050 801.900 ;
        RECT 199.950 801.600 202.050 802.050 ;
        RECT 193.950 800.400 202.050 801.600 ;
        RECT 206.400 801.600 207.600 803.400 ;
        RECT 215.400 803.400 228.600 804.600 ;
        RECT 215.400 801.900 216.600 803.400 ;
        RECT 214.950 801.600 217.050 801.900 ;
        RECT 206.400 800.400 217.050 801.600 ;
        RECT 227.400 801.600 228.600 803.400 ;
        RECT 238.950 801.600 241.050 801.900 ;
        RECT 227.400 800.400 241.050 801.600 ;
        RECT 193.950 799.800 196.050 800.400 ;
        RECT 199.950 799.950 202.050 800.400 ;
        RECT 214.950 799.800 217.050 800.400 ;
        RECT 238.950 799.800 241.050 800.400 ;
        RECT 253.950 801.600 256.050 801.900 ;
        RECT 268.950 801.600 271.050 801.900 ;
        RECT 253.950 800.400 271.050 801.600 ;
        RECT 253.950 799.800 256.050 800.400 ;
        RECT 268.950 799.800 271.050 800.400 ;
        RECT 340.950 801.450 343.050 801.900 ;
        RECT 346.950 801.450 349.050 801.900 ;
        RECT 340.950 800.250 349.050 801.450 ;
        RECT 340.950 799.800 343.050 800.250 ;
        RECT 346.950 799.800 349.050 800.250 ;
        RECT 382.950 801.600 385.050 802.050 ;
        RECT 395.400 801.600 396.600 806.400 ;
        RECT 403.950 805.950 406.050 806.400 ;
        RECT 415.950 807.600 418.050 808.200 ;
        RECT 430.950 807.600 433.050 808.050 ;
        RECT 415.950 806.400 433.050 807.600 ;
        RECT 415.950 806.100 418.050 806.400 ;
        RECT 430.950 805.950 433.050 806.400 ;
        RECT 382.950 800.400 396.600 801.600 ;
        RECT 382.950 799.950 385.050 800.400 ;
        RECT 13.950 798.600 16.050 799.050 ;
        RECT 29.400 798.600 30.600 799.800 ;
        RECT 440.400 799.050 441.600 808.950 ;
        RECT 445.950 804.750 448.050 805.200 ;
        RECT 460.950 804.750 463.050 805.200 ;
        RECT 482.400 804.900 483.600 809.400 ;
        RECT 505.950 809.400 586.050 810.600 ;
        RECT 505.950 808.950 508.050 809.400 ;
        RECT 583.950 808.950 586.050 809.400 ;
        RECT 733.950 810.600 736.050 811.050 ;
        RECT 757.950 810.600 760.050 811.050 ;
        RECT 766.950 810.600 769.050 811.050 ;
        RECT 733.950 809.400 769.050 810.600 ;
        RECT 733.950 808.950 736.050 809.400 ;
        RECT 757.950 808.950 760.050 809.400 ;
        RECT 766.950 808.950 769.050 809.400 ;
        RECT 517.950 807.600 520.050 808.050 ;
        RECT 577.950 807.600 580.050 808.050 ;
        RECT 517.950 806.400 580.050 807.600 ;
        RECT 517.950 805.950 520.050 806.400 ;
        RECT 577.950 805.950 580.050 806.400 ;
        RECT 583.950 807.600 586.050 808.200 ;
        RECT 592.950 807.600 595.050 808.050 ;
        RECT 583.950 806.400 595.050 807.600 ;
        RECT 583.950 806.100 586.050 806.400 ;
        RECT 592.950 805.950 595.050 806.400 ;
        RECT 607.950 807.750 610.050 808.200 ;
        RECT 613.950 807.750 616.050 808.200 ;
        RECT 607.950 806.550 616.050 807.750 ;
        RECT 607.950 806.100 610.050 806.550 ;
        RECT 613.950 806.100 616.050 806.550 ;
        RECT 643.950 807.600 646.050 808.050 ;
        RECT 655.950 807.600 658.050 808.050 ;
        RECT 643.950 806.400 658.050 807.600 ;
        RECT 643.950 805.950 646.050 806.400 ;
        RECT 655.950 805.950 658.050 806.400 ;
        RECT 667.950 806.100 670.050 808.200 ;
        RECT 709.950 807.750 712.050 808.200 ;
        RECT 721.950 807.750 724.050 808.050 ;
        RECT 730.950 807.750 733.050 808.200 ;
        RECT 709.950 806.550 733.050 807.750 ;
        RECT 709.950 806.100 712.050 806.550 ;
        RECT 445.950 803.550 463.050 804.750 ;
        RECT 445.950 803.100 448.050 803.550 ;
        RECT 460.950 803.100 463.050 803.550 ;
        RECT 481.950 802.800 484.050 804.900 ;
        RECT 502.950 801.600 505.050 805.050 ;
        RECT 508.950 804.600 511.050 805.050 ;
        RECT 595.950 804.600 598.050 805.050 ;
        RECT 508.950 803.400 598.050 804.600 ;
        RECT 508.950 802.950 511.050 803.400 ;
        RECT 595.950 802.950 598.050 803.400 ;
        RECT 511.950 801.600 514.050 802.050 ;
        RECT 502.950 801.000 514.050 801.600 ;
        RECT 503.400 800.400 514.050 801.000 ;
        RECT 511.950 799.950 514.050 800.400 ;
        RECT 526.950 801.600 529.050 801.900 ;
        RECT 538.950 801.600 541.050 802.050 ;
        RECT 526.950 801.450 541.050 801.600 ;
        RECT 550.950 801.450 553.050 801.900 ;
        RECT 526.950 800.400 553.050 801.450 ;
        RECT 526.950 799.800 529.050 800.400 ;
        RECT 538.950 800.250 553.050 800.400 ;
        RECT 538.950 799.950 541.050 800.250 ;
        RECT 550.950 799.800 553.050 800.250 ;
        RECT 556.950 801.450 559.050 801.900 ;
        RECT 562.950 801.450 565.050 801.900 ;
        RECT 556.950 800.250 565.050 801.450 ;
        RECT 556.950 799.800 559.050 800.250 ;
        RECT 562.950 799.800 565.050 800.250 ;
        RECT 568.950 801.600 571.050 801.900 ;
        RECT 574.800 801.600 576.900 802.050 ;
        RECT 568.950 800.400 576.900 801.600 ;
        RECT 568.950 799.800 571.050 800.400 ;
        RECT 574.800 799.950 576.900 800.400 ;
        RECT 577.950 801.600 580.050 802.050 ;
        RECT 589.950 801.600 592.050 801.900 ;
        RECT 577.950 800.400 592.050 801.600 ;
        RECT 577.950 799.950 580.050 800.400 ;
        RECT 589.950 799.800 592.050 800.400 ;
        RECT 652.950 801.450 655.050 801.900 ;
        RECT 658.800 801.450 660.900 801.900 ;
        RECT 652.950 800.250 660.900 801.450 ;
        RECT 652.950 799.800 655.050 800.250 ;
        RECT 658.800 799.800 660.900 800.250 ;
        RECT 661.950 801.600 664.050 802.050 ;
        RECT 668.400 801.600 669.600 806.100 ;
        RECT 721.950 805.950 724.050 806.550 ;
        RECT 730.950 806.100 733.050 806.550 ;
        RECT 898.950 807.750 901.050 808.200 ;
        RECT 913.950 807.750 916.050 808.200 ;
        RECT 898.950 806.550 916.050 807.750 ;
        RECT 898.950 806.100 901.050 806.550 ;
        RECT 913.950 806.100 916.050 806.550 ;
        RECT 661.950 800.400 669.600 801.600 ;
        RECT 676.950 801.600 679.050 801.900 ;
        RECT 688.950 801.600 691.050 801.900 ;
        RECT 832.950 801.600 835.050 805.050 ;
        RECT 859.950 804.450 862.050 804.900 ;
        RECT 880.950 804.450 883.050 804.900 ;
        RECT 859.950 803.250 883.050 804.450 ;
        RECT 859.950 802.800 862.050 803.250 ;
        RECT 880.950 802.800 883.050 803.250 ;
        RECT 676.950 800.400 691.050 801.600 ;
        RECT 661.950 799.950 664.050 800.400 ;
        RECT 676.950 799.800 679.050 800.400 ;
        RECT 688.950 799.800 691.050 800.400 ;
        RECT 827.400 800.400 837.600 801.600 ;
        RECT 13.950 797.400 30.600 798.600 ;
        RECT 46.950 798.600 49.050 799.050 ;
        RECT 52.950 798.600 55.050 799.050 ;
        RECT 46.950 797.400 55.050 798.600 ;
        RECT 13.950 796.950 16.050 797.400 ;
        RECT 46.950 796.950 49.050 797.400 ;
        RECT 52.950 796.950 55.050 797.400 ;
        RECT 97.950 798.600 100.050 799.050 ;
        RECT 106.950 798.600 109.050 799.050 ;
        RECT 112.950 798.600 115.050 799.050 ;
        RECT 157.950 798.600 160.050 799.050 ;
        RECT 97.950 797.400 160.050 798.600 ;
        RECT 97.950 796.950 100.050 797.400 ;
        RECT 106.950 796.950 109.050 797.400 ;
        RECT 112.950 796.950 115.050 797.400 ;
        RECT 157.950 796.950 160.050 797.400 ;
        RECT 379.950 798.600 382.050 799.050 ;
        RECT 406.950 798.600 409.050 799.050 ;
        RECT 379.950 797.400 409.050 798.600 ;
        RECT 379.950 796.950 382.050 797.400 ;
        RECT 406.950 796.950 409.050 797.400 ;
        RECT 439.950 796.950 442.050 799.050 ;
        RECT 481.950 798.600 484.050 799.050 ;
        RECT 496.950 798.600 499.050 799.050 ;
        RECT 481.950 797.400 499.050 798.600 ;
        RECT 481.950 796.950 484.050 797.400 ;
        RECT 496.950 796.950 499.050 797.400 ;
        RECT 505.950 798.450 508.050 798.900 ;
        RECT 517.950 798.450 520.050 798.900 ;
        RECT 505.950 797.250 520.050 798.450 ;
        RECT 505.950 796.800 508.050 797.250 ;
        RECT 517.950 796.800 520.050 797.250 ;
        RECT 625.950 798.600 628.050 799.050 ;
        RECT 646.950 798.600 649.050 799.050 ;
        RECT 679.950 798.600 682.050 799.050 ;
        RECT 697.950 798.600 700.050 799.050 ;
        RECT 625.950 797.400 700.050 798.600 ;
        RECT 625.950 796.950 628.050 797.400 ;
        RECT 646.950 796.950 649.050 797.400 ;
        RECT 679.950 796.950 682.050 797.400 ;
        RECT 697.950 796.950 700.050 797.400 ;
        RECT 703.950 798.600 706.050 799.050 ;
        RECT 712.950 798.600 715.050 799.050 ;
        RECT 827.400 798.900 828.600 800.400 ;
        RECT 836.400 798.900 837.600 800.400 ;
        RECT 703.950 797.400 715.050 798.600 ;
        RECT 703.950 796.950 706.050 797.400 ;
        RECT 712.950 796.950 715.050 797.400 ;
        RECT 826.950 796.800 829.050 798.900 ;
        RECT 835.950 796.800 838.050 798.900 ;
        RECT 115.950 795.600 118.050 796.050 ;
        RECT 133.950 795.600 136.050 796.050 ;
        RECT 115.950 794.400 136.050 795.600 ;
        RECT 115.950 793.950 118.050 794.400 ;
        RECT 133.950 793.950 136.050 794.400 ;
        RECT 229.950 795.600 232.050 796.050 ;
        RECT 322.950 795.600 325.050 796.050 ;
        RECT 229.950 794.400 325.050 795.600 ;
        RECT 229.950 793.950 232.050 794.400 ;
        RECT 322.950 793.950 325.050 794.400 ;
        RECT 367.950 795.600 370.050 796.050 ;
        RECT 430.950 795.600 433.050 796.050 ;
        RECT 523.800 795.600 525.900 796.050 ;
        RECT 367.950 794.400 525.900 795.600 ;
        RECT 367.950 793.950 370.050 794.400 ;
        RECT 430.950 793.950 433.050 794.400 ;
        RECT 523.800 793.950 525.900 794.400 ;
        RECT 526.950 795.600 529.050 796.050 ;
        RECT 535.950 795.600 538.050 796.050 ;
        RECT 526.950 794.400 538.050 795.600 ;
        RECT 526.950 793.950 529.050 794.400 ;
        RECT 535.950 793.950 538.050 794.400 ;
        RECT 547.950 795.600 550.050 796.050 ;
        RECT 610.950 795.600 613.050 796.050 ;
        RECT 547.950 794.400 613.050 795.600 ;
        RECT 547.950 793.950 550.050 794.400 ;
        RECT 610.950 793.950 613.050 794.400 ;
        RECT 637.950 795.600 640.050 796.050 ;
        RECT 670.950 795.600 673.050 796.050 ;
        RECT 637.950 794.400 673.050 795.600 ;
        RECT 637.950 793.950 640.050 794.400 ;
        RECT 670.950 793.950 673.050 794.400 ;
        RECT 34.950 792.600 37.050 793.050 ;
        RECT 43.950 792.600 46.050 793.050 ;
        RECT 58.950 792.600 61.050 793.050 ;
        RECT 34.950 791.400 61.050 792.600 ;
        RECT 34.950 790.950 37.050 791.400 ;
        RECT 43.950 790.950 46.050 791.400 ;
        RECT 58.950 790.950 61.050 791.400 ;
        RECT 82.950 792.600 85.050 793.050 ;
        RECT 91.950 792.600 94.050 793.050 ;
        RECT 82.950 791.400 94.050 792.600 ;
        RECT 82.950 790.950 85.050 791.400 ;
        RECT 91.950 790.950 94.050 791.400 ;
        RECT 157.950 792.600 160.050 793.050 ;
        RECT 187.950 792.600 190.050 793.050 ;
        RECT 208.950 792.600 211.050 793.050 ;
        RECT 157.950 791.400 211.050 792.600 ;
        RECT 157.950 790.950 160.050 791.400 ;
        RECT 187.950 790.950 190.050 791.400 ;
        RECT 208.950 790.950 211.050 791.400 ;
        RECT 262.950 792.600 265.050 793.050 ;
        RECT 457.950 792.600 460.050 793.050 ;
        RECT 505.950 792.600 508.050 793.050 ;
        RECT 262.950 791.400 357.600 792.600 ;
        RECT 262.950 790.950 265.050 791.400 ;
        RECT 94.950 789.600 97.050 790.050 ;
        RECT 109.950 789.600 112.050 790.050 ;
        RECT 94.950 788.400 112.050 789.600 ;
        RECT 94.950 787.950 97.050 788.400 ;
        RECT 109.950 787.950 112.050 788.400 ;
        RECT 250.950 789.600 253.050 790.050 ;
        RECT 352.950 789.600 355.050 790.050 ;
        RECT 250.950 788.400 355.050 789.600 ;
        RECT 356.400 789.600 357.600 791.400 ;
        RECT 457.950 791.400 508.050 792.600 ;
        RECT 524.400 792.600 525.600 793.950 ;
        RECT 580.950 792.600 583.050 793.050 ;
        RECT 697.950 792.600 700.050 793.050 ;
        RECT 736.950 792.600 739.050 793.050 ;
        RECT 524.400 791.400 739.050 792.600 ;
        RECT 457.950 790.950 460.050 791.400 ;
        RECT 505.950 790.950 508.050 791.400 ;
        RECT 580.950 790.950 583.050 791.400 ;
        RECT 697.950 790.950 700.050 791.400 ;
        RECT 736.950 790.950 739.050 791.400 ;
        RECT 892.950 792.600 895.050 793.050 ;
        RECT 916.950 792.600 919.050 793.050 ;
        RECT 892.950 791.400 919.050 792.600 ;
        RECT 892.950 790.950 895.050 791.400 ;
        RECT 916.950 790.950 919.050 791.400 ;
        RECT 418.950 789.600 421.050 790.050 ;
        RECT 356.400 788.400 421.050 789.600 ;
        RECT 250.950 787.950 253.050 788.400 ;
        RECT 352.950 787.950 355.050 788.400 ;
        RECT 418.950 787.950 421.050 788.400 ;
        RECT 436.950 789.600 439.050 790.050 ;
        RECT 442.950 789.600 445.050 790.050 ;
        RECT 520.950 789.600 523.050 790.050 ;
        RECT 436.950 788.400 523.050 789.600 ;
        RECT 436.950 787.950 439.050 788.400 ;
        RECT 442.950 787.950 445.050 788.400 ;
        RECT 520.950 787.950 523.050 788.400 ;
        RECT 529.950 789.600 532.050 790.050 ;
        RECT 541.950 789.600 544.050 790.050 ;
        RECT 529.950 788.400 544.050 789.600 ;
        RECT 529.950 787.950 532.050 788.400 ;
        RECT 541.950 787.950 544.050 788.400 ;
        RECT 595.950 789.600 598.050 790.050 ;
        RECT 661.800 789.600 663.900 790.050 ;
        RECT 595.950 788.400 663.900 789.600 ;
        RECT 595.950 787.950 598.050 788.400 ;
        RECT 661.800 787.950 663.900 788.400 ;
        RECT 664.950 789.600 667.050 790.050 ;
        RECT 766.950 789.600 769.050 790.050 ;
        RECT 664.950 788.400 769.050 789.600 ;
        RECT 664.950 787.950 667.050 788.400 ;
        RECT 766.950 787.950 769.050 788.400 ;
        RECT 919.950 789.600 922.050 790.050 ;
        RECT 925.950 789.600 928.050 790.050 ;
        RECT 919.950 788.400 928.050 789.600 ;
        RECT 919.950 787.950 922.050 788.400 ;
        RECT 925.950 787.950 928.050 788.400 ;
        RECT 253.950 786.600 256.050 787.050 ;
        RECT 376.950 786.600 379.050 787.050 ;
        RECT 421.950 786.600 424.050 787.050 ;
        RECT 253.950 785.400 300.600 786.600 ;
        RECT 253.950 784.950 256.050 785.400 ;
        RECT 299.400 783.600 300.600 785.400 ;
        RECT 376.950 785.400 424.050 786.600 ;
        RECT 376.950 784.950 379.050 785.400 ;
        RECT 421.950 784.950 424.050 785.400 ;
        RECT 439.950 786.600 442.050 787.050 ;
        RECT 541.950 786.600 544.050 786.900 ;
        RECT 439.950 785.400 544.050 786.600 ;
        RECT 439.950 784.950 442.050 785.400 ;
        RECT 541.950 784.800 544.050 785.400 ;
        RECT 580.950 786.600 583.050 787.050 ;
        RECT 580.950 785.400 633.600 786.600 ;
        RECT 580.950 784.950 583.050 785.400 ;
        RECT 451.950 783.600 454.050 784.050 ;
        RECT 547.950 783.600 550.050 784.050 ;
        RECT 299.400 782.400 441.600 783.600 ;
        RECT 136.950 780.600 139.050 781.050 ;
        RECT 253.950 780.600 256.050 781.050 ;
        RECT 136.950 779.400 256.050 780.600 ;
        RECT 136.950 778.950 139.050 779.400 ;
        RECT 253.950 778.950 256.050 779.400 ;
        RECT 274.950 780.600 277.050 781.050 ;
        RECT 280.950 780.600 283.050 781.050 ;
        RECT 292.950 780.600 295.050 781.050 ;
        RECT 412.950 780.600 415.050 781.050 ;
        RECT 274.950 779.400 295.050 780.600 ;
        RECT 274.950 778.950 277.050 779.400 ;
        RECT 280.950 778.950 283.050 779.400 ;
        RECT 292.950 778.950 295.050 779.400 ;
        RECT 335.400 779.400 415.050 780.600 ;
        RECT 440.400 780.600 441.600 782.400 ;
        RECT 451.950 782.400 550.050 783.600 ;
        RECT 632.400 783.600 633.600 785.400 ;
        RECT 691.950 783.600 694.050 784.050 ;
        RECT 742.950 783.600 745.050 784.050 ;
        RECT 632.400 782.400 694.050 783.600 ;
        RECT 451.950 781.950 454.050 782.400 ;
        RECT 547.950 781.950 550.050 782.400 ;
        RECT 691.950 781.950 694.050 782.400 ;
        RECT 695.400 782.400 745.050 783.600 ;
        RECT 460.950 780.600 463.050 781.050 ;
        RECT 484.950 780.600 487.050 781.050 ;
        RECT 440.400 779.400 487.050 780.600 ;
        RECT 133.950 777.600 136.050 778.050 ;
        RECT 262.950 777.600 265.050 778.050 ;
        RECT 133.950 776.400 265.050 777.600 ;
        RECT 133.950 775.950 136.050 776.400 ;
        RECT 262.950 775.950 265.050 776.400 ;
        RECT 301.950 777.600 304.050 778.050 ;
        RECT 335.400 777.600 336.600 779.400 ;
        RECT 412.950 778.950 415.050 779.400 ;
        RECT 460.950 778.950 463.050 779.400 ;
        RECT 484.950 778.950 487.050 779.400 ;
        RECT 514.950 780.600 517.050 781.050 ;
        RECT 532.950 780.600 535.050 781.050 ;
        RECT 514.950 779.400 535.050 780.600 ;
        RECT 514.950 778.950 517.050 779.400 ;
        RECT 532.950 778.950 535.050 779.400 ;
        RECT 583.950 780.600 586.050 781.050 ;
        RECT 695.400 780.600 696.600 782.400 ;
        RECT 742.950 781.950 745.050 782.400 ;
        RECT 802.950 783.600 805.050 784.050 ;
        RECT 808.950 783.600 811.050 784.050 ;
        RECT 802.950 782.400 811.050 783.600 ;
        RECT 802.950 781.950 805.050 782.400 ;
        RECT 808.950 781.950 811.050 782.400 ;
        RECT 583.950 779.400 696.600 780.600 ;
        RECT 718.950 780.600 721.050 781.050 ;
        RECT 739.950 780.600 742.050 781.050 ;
        RECT 814.950 780.600 817.050 781.050 ;
        RECT 916.950 780.600 919.050 781.050 ;
        RECT 718.950 779.400 817.050 780.600 ;
        RECT 583.950 778.950 586.050 779.400 ;
        RECT 718.950 778.950 721.050 779.400 ;
        RECT 739.950 778.950 742.050 779.400 ;
        RECT 814.950 778.950 817.050 779.400 ;
        RECT 821.400 779.400 919.050 780.600 ;
        RECT 301.950 776.400 336.600 777.600 ;
        RECT 427.950 777.600 430.050 778.050 ;
        RECT 580.950 777.600 583.050 778.050 ;
        RECT 427.950 776.400 583.050 777.600 ;
        RECT 301.950 775.950 304.050 776.400 ;
        RECT 427.950 775.950 430.050 776.400 ;
        RECT 580.950 775.950 583.050 776.400 ;
        RECT 601.950 777.600 604.050 778.050 ;
        RECT 643.950 777.600 646.050 778.050 ;
        RECT 661.950 777.600 664.050 778.050 ;
        RECT 727.950 777.600 730.050 778.050 ;
        RECT 601.950 776.400 730.050 777.600 ;
        RECT 601.950 775.950 604.050 776.400 ;
        RECT 643.950 775.950 646.050 776.400 ;
        RECT 661.950 775.950 664.050 776.400 ;
        RECT 727.950 775.950 730.050 776.400 ;
        RECT 742.950 777.600 745.050 778.050 ;
        RECT 821.400 777.600 822.600 779.400 ;
        RECT 916.950 778.950 919.050 779.400 ;
        RECT 742.950 776.400 822.600 777.600 ;
        RECT 826.950 777.600 829.050 778.050 ;
        RECT 847.950 777.600 850.050 778.050 ;
        RECT 826.950 776.400 850.050 777.600 ;
        RECT 742.950 775.950 745.050 776.400 ;
        RECT 826.950 775.950 829.050 776.400 ;
        RECT 847.950 775.950 850.050 776.400 ;
        RECT 94.950 774.600 97.050 775.050 ;
        RECT 124.950 774.600 127.050 775.050 ;
        RECT 94.950 773.400 127.050 774.600 ;
        RECT 94.950 772.950 97.050 773.400 ;
        RECT 124.950 772.950 127.050 773.400 ;
        RECT 232.950 774.600 235.050 775.050 ;
        RECT 277.950 774.600 280.050 775.050 ;
        RECT 430.950 774.600 433.050 775.050 ;
        RECT 232.950 773.400 280.050 774.600 ;
        RECT 232.950 772.950 235.050 773.400 ;
        RECT 277.950 772.950 280.050 773.400 ;
        RECT 404.400 773.400 433.050 774.600 ;
        RECT 404.400 772.050 405.600 773.400 ;
        RECT 430.950 772.950 433.050 773.400 ;
        RECT 484.950 774.600 487.050 775.050 ;
        RECT 520.950 774.600 523.050 775.050 ;
        RECT 529.950 774.600 532.050 775.050 ;
        RECT 484.950 773.400 532.050 774.600 ;
        RECT 484.950 772.950 487.050 773.400 ;
        RECT 520.950 772.950 523.050 773.400 ;
        RECT 529.950 772.950 532.050 773.400 ;
        RECT 535.950 774.600 538.050 775.050 ;
        RECT 583.950 774.600 586.050 775.050 ;
        RECT 535.950 773.400 586.050 774.600 ;
        RECT 535.950 772.950 538.050 773.400 ;
        RECT 583.950 772.950 586.050 773.400 ;
        RECT 760.950 774.600 763.050 775.050 ;
        RECT 799.950 774.600 802.050 775.050 ;
        RECT 760.950 773.400 802.050 774.600 ;
        RECT 760.950 772.950 763.050 773.400 ;
        RECT 799.950 772.950 802.050 773.400 ;
        RECT 814.950 774.600 817.050 775.050 ;
        RECT 823.950 774.600 826.050 775.050 ;
        RECT 859.950 774.600 862.050 775.050 ;
        RECT 814.950 773.400 862.050 774.600 ;
        RECT 814.950 772.950 817.050 773.400 ;
        RECT 823.950 772.950 826.050 773.400 ;
        RECT 859.950 772.950 862.050 773.400 ;
        RECT 49.950 771.600 52.050 772.050 ;
        RECT 133.950 771.600 136.050 772.050 ;
        RECT 49.950 770.400 136.050 771.600 ;
        RECT 49.950 769.950 52.050 770.400 ;
        RECT 133.950 769.950 136.050 770.400 ;
        RECT 193.950 771.600 196.050 772.050 ;
        RECT 202.950 771.600 205.050 772.050 ;
        RECT 193.950 770.400 205.050 771.600 ;
        RECT 193.950 769.950 196.050 770.400 ;
        RECT 202.950 769.950 205.050 770.400 ;
        RECT 343.950 771.600 346.050 772.050 ;
        RECT 355.950 771.600 358.050 772.050 ;
        RECT 403.950 771.600 406.050 772.050 ;
        RECT 343.950 770.400 406.050 771.600 ;
        RECT 343.950 769.950 346.050 770.400 ;
        RECT 355.950 769.950 358.050 770.400 ;
        RECT 403.950 769.950 406.050 770.400 ;
        RECT 421.950 771.600 424.050 772.050 ;
        RECT 481.950 771.600 484.050 772.050 ;
        RECT 421.950 770.400 484.050 771.600 ;
        RECT 421.950 769.950 424.050 770.400 ;
        RECT 481.950 769.950 484.050 770.400 ;
        RECT 649.950 771.600 652.050 772.050 ;
        RECT 703.950 771.600 706.050 772.050 ;
        RECT 796.950 771.600 799.050 772.050 ;
        RECT 649.950 770.400 706.050 771.600 ;
        RECT 649.950 769.950 652.050 770.400 ;
        RECT 703.950 769.950 706.050 770.400 ;
        RECT 779.400 770.400 799.050 771.600 ;
        RECT 79.950 768.600 82.050 769.050 ;
        RECT 88.950 768.600 91.050 769.050 ;
        RECT 79.950 767.400 91.050 768.600 ;
        RECT 79.950 766.950 82.050 767.400 ;
        RECT 88.950 766.950 91.050 767.400 ;
        RECT 103.950 768.600 106.050 769.050 ;
        RECT 115.950 768.600 118.050 769.050 ;
        RECT 103.950 767.400 118.050 768.600 ;
        RECT 103.950 766.950 106.050 767.400 ;
        RECT 115.950 766.950 118.050 767.400 ;
        RECT 142.950 768.600 145.050 769.050 ;
        RECT 154.950 768.600 157.050 769.050 ;
        RECT 142.950 767.400 157.050 768.600 ;
        RECT 142.950 766.950 145.050 767.400 ;
        RECT 154.950 766.950 157.050 767.400 ;
        RECT 244.950 768.600 247.050 769.050 ;
        RECT 256.950 768.600 259.050 769.050 ;
        RECT 289.950 768.600 292.050 769.050 ;
        RECT 244.950 767.400 292.050 768.600 ;
        RECT 244.950 766.950 247.050 767.400 ;
        RECT 256.950 766.950 259.050 767.400 ;
        RECT 289.950 766.950 292.050 767.400 ;
        RECT 370.950 768.600 373.050 769.050 ;
        RECT 511.950 768.600 514.050 769.050 ;
        RECT 532.950 768.600 535.050 769.050 ;
        RECT 538.950 768.600 541.050 769.050 ;
        RECT 370.950 767.400 402.600 768.600 ;
        RECT 370.950 766.950 373.050 767.400 ;
        RECT 118.950 765.600 121.050 766.050 ;
        RECT 68.400 764.400 121.050 765.600 ;
        RECT 68.400 763.200 69.600 764.400 ;
        RECT 118.950 763.950 121.050 764.400 ;
        RECT 190.950 765.600 193.050 766.050 ;
        RECT 214.950 765.600 217.050 766.050 ;
        RECT 190.950 764.400 217.050 765.600 ;
        RECT 401.400 765.600 402.600 767.400 ;
        RECT 511.950 767.400 541.050 768.600 ;
        RECT 511.950 766.950 514.050 767.400 ;
        RECT 532.950 766.950 535.050 767.400 ;
        RECT 538.950 766.950 541.050 767.400 ;
        RECT 595.950 768.600 598.050 769.050 ;
        RECT 604.950 768.600 607.050 769.050 ;
        RECT 595.950 767.400 607.050 768.600 ;
        RECT 595.950 766.950 598.050 767.400 ;
        RECT 604.950 766.950 607.050 767.400 ;
        RECT 616.950 768.600 621.000 769.050 ;
        RECT 715.950 768.600 718.050 769.050 ;
        RECT 779.400 768.600 780.600 770.400 ;
        RECT 796.950 769.950 799.050 770.400 ;
        RECT 616.950 766.950 621.600 768.600 ;
        RECT 715.950 767.400 780.600 768.600 ;
        RECT 784.950 768.600 787.050 769.050 ;
        RECT 793.950 768.600 796.050 769.050 ;
        RECT 784.950 767.400 796.050 768.600 ;
        RECT 715.950 766.950 718.050 767.400 ;
        RECT 784.950 766.950 787.050 767.400 ;
        RECT 793.950 766.950 796.050 767.400 ;
        RECT 805.950 768.600 808.050 769.050 ;
        RECT 868.950 768.600 871.050 769.050 ;
        RECT 805.950 767.400 871.050 768.600 ;
        RECT 805.950 766.950 808.050 767.400 ;
        RECT 868.950 766.950 871.050 767.400 ;
        RECT 889.950 768.600 892.050 769.050 ;
        RECT 925.950 768.600 928.050 769.050 ;
        RECT 889.950 767.400 928.050 768.600 ;
        RECT 889.950 766.950 892.050 767.400 ;
        RECT 925.950 766.950 928.050 767.400 ;
        RECT 415.950 765.600 418.050 766.050 ;
        RECT 401.400 764.400 418.050 765.600 ;
        RECT 190.950 763.950 193.050 764.400 ;
        RECT 214.950 763.950 217.050 764.400 ;
        RECT 415.950 763.950 418.050 764.400 ;
        RECT 457.950 765.600 460.050 766.200 ;
        RECT 466.950 765.600 469.050 766.050 ;
        RECT 457.950 764.400 469.050 765.600 ;
        RECT 457.950 764.100 460.050 764.400 ;
        RECT 466.950 763.950 469.050 764.400 ;
        RECT 481.950 765.600 484.050 766.050 ;
        RECT 607.950 765.600 610.050 766.050 ;
        RECT 481.950 764.400 610.050 765.600 ;
        RECT 481.950 763.950 484.050 764.400 ;
        RECT 4.950 762.750 7.050 763.200 ;
        RECT 13.950 762.750 16.050 763.200 ;
        RECT 4.950 761.550 16.050 762.750 ;
        RECT 4.950 761.100 7.050 761.550 ;
        RECT 13.950 761.100 16.050 761.550 ;
        RECT 19.950 761.100 22.050 763.200 ;
        RECT 49.950 762.750 52.050 763.200 ;
        RECT 55.950 762.750 58.050 763.200 ;
        RECT 49.950 761.550 58.050 762.750 ;
        RECT 49.950 761.100 52.050 761.550 ;
        RECT 55.950 761.100 58.050 761.550 ;
        RECT 61.950 762.750 64.050 763.200 ;
        RECT 67.950 762.750 70.050 763.200 ;
        RECT 61.950 761.550 70.050 762.750 ;
        RECT 61.950 761.100 64.050 761.550 ;
        RECT 67.950 761.100 70.050 761.550 ;
        RECT 76.950 761.100 79.050 763.200 ;
        RECT 82.950 762.600 85.050 763.200 ;
        RECT 97.950 762.600 100.050 763.200 ;
        RECT 82.950 761.400 100.050 762.600 ;
        RECT 82.950 761.100 85.050 761.400 ;
        RECT 97.950 761.100 100.050 761.400 ;
        RECT 20.400 757.050 21.600 761.100 ;
        RECT 7.950 756.450 10.050 756.900 ;
        RECT 16.950 756.450 19.050 756.900 ;
        RECT 7.950 755.250 19.050 756.450 ;
        RECT 20.400 755.400 25.050 757.050 ;
        RECT 7.950 754.800 10.050 755.250 ;
        RECT 16.950 754.800 19.050 755.250 ;
        RECT 21.000 754.950 25.050 755.400 ;
        RECT 56.400 753.600 57.600 761.100 ;
        RECT 58.950 756.600 61.050 756.900 ;
        RECT 77.400 756.600 78.600 761.100 ;
        RECT 58.950 755.400 78.600 756.600 ;
        RECT 83.400 757.050 84.600 761.100 ;
        RECT 109.950 760.950 112.050 763.050 ;
        RECT 118.950 762.600 121.050 763.200 ;
        RECT 148.950 762.600 151.050 763.200 ;
        RECT 118.950 761.400 151.050 762.600 ;
        RECT 118.950 761.100 121.050 761.400 ;
        RECT 148.950 761.100 151.050 761.400 ;
        RECT 166.950 761.100 169.050 763.200 ;
        RECT 172.950 761.100 175.050 763.200 ;
        RECT 178.950 762.750 181.050 763.200 ;
        RECT 190.950 762.750 193.050 763.200 ;
        RECT 178.950 761.550 193.050 762.750 ;
        RECT 178.950 761.100 181.050 761.550 ;
        RECT 190.950 761.100 193.050 761.550 ;
        RECT 196.950 762.750 199.050 763.200 ;
        RECT 205.950 762.750 208.050 763.200 ;
        RECT 196.950 761.550 208.050 762.750 ;
        RECT 196.950 761.100 199.050 761.550 ;
        RECT 205.950 761.100 208.050 761.550 ;
        RECT 220.950 762.750 223.050 763.200 ;
        RECT 226.950 762.750 229.050 763.200 ;
        RECT 220.950 762.600 229.050 762.750 ;
        RECT 235.950 762.600 238.050 763.200 ;
        RECT 220.950 761.550 238.050 762.600 ;
        RECT 220.950 761.100 223.050 761.550 ;
        RECT 226.950 761.400 238.050 761.550 ;
        RECT 226.950 761.100 229.050 761.400 ;
        RECT 235.950 761.100 238.050 761.400 ;
        RECT 241.950 762.600 244.050 763.200 ;
        RECT 253.950 762.750 256.050 763.200 ;
        RECT 259.950 762.750 262.050 763.200 ;
        RECT 253.950 762.600 262.050 762.750 ;
        RECT 241.950 761.550 262.050 762.600 ;
        RECT 241.950 761.400 256.050 761.550 ;
        RECT 241.950 761.100 244.050 761.400 ;
        RECT 253.950 761.100 256.050 761.400 ;
        RECT 259.950 761.100 262.050 761.550 ;
        RECT 295.950 762.750 298.050 763.200 ;
        RECT 304.800 762.750 306.900 763.200 ;
        RECT 295.950 761.550 306.900 762.750 ;
        RECT 295.950 761.100 298.050 761.550 ;
        RECT 304.800 761.100 306.900 761.550 ;
        RECT 83.400 755.400 88.050 757.050 ;
        RECT 58.950 754.800 61.050 755.400 ;
        RECT 84.000 754.950 88.050 755.400 ;
        RECT 106.950 756.600 109.050 756.900 ;
        RECT 110.400 756.600 111.600 760.950 ;
        RECT 121.950 756.600 124.050 756.900 ;
        RECT 106.950 755.400 111.600 756.600 ;
        RECT 116.400 756.000 124.050 756.600 ;
        RECT 115.950 755.400 124.050 756.000 ;
        RECT 106.950 754.800 109.050 755.400 ;
        RECT 76.950 753.600 79.050 754.050 ;
        RECT 56.400 752.400 79.050 753.600 ;
        RECT 76.950 751.950 79.050 752.400 ;
        RECT 82.950 753.600 85.050 754.050 ;
        RECT 88.950 753.600 91.050 754.050 ;
        RECT 82.950 752.400 91.050 753.600 ;
        RECT 82.950 751.950 85.050 752.400 ;
        RECT 88.950 751.950 91.050 752.400 ;
        RECT 115.950 751.950 118.050 755.400 ;
        RECT 121.950 754.800 124.050 755.400 ;
        RECT 127.950 756.600 130.050 756.900 ;
        RECT 139.950 756.600 142.050 756.900 ;
        RECT 127.950 755.400 142.050 756.600 ;
        RECT 127.950 754.800 130.050 755.400 ;
        RECT 139.950 754.800 142.050 755.400 ;
        RECT 145.950 756.600 148.050 756.900 ;
        RECT 167.400 756.600 168.600 761.100 ;
        RECT 145.950 755.400 168.600 756.600 ;
        RECT 173.400 757.050 174.600 761.100 ;
        RECT 307.950 759.600 310.050 763.050 ;
        RECT 319.950 762.750 322.050 763.200 ;
        RECT 325.950 762.750 328.050 763.200 ;
        RECT 319.950 761.550 328.050 762.750 ;
        RECT 319.950 761.100 322.050 761.550 ;
        RECT 325.950 761.100 328.050 761.550 ;
        RECT 337.950 761.100 340.050 763.200 ;
        RECT 370.950 762.600 373.050 763.200 ;
        RECT 382.950 762.600 385.050 763.050 ;
        RECT 370.950 761.400 385.050 762.600 ;
        RECT 370.950 761.100 373.050 761.400 ;
        RECT 302.400 759.000 310.050 759.600 ;
        RECT 338.400 759.600 339.600 761.100 ;
        RECT 382.950 760.950 385.050 761.400 ;
        RECT 388.950 762.600 391.050 763.200 ;
        RECT 397.950 762.600 400.050 762.900 ;
        RECT 424.950 762.600 427.050 763.200 ;
        RECT 388.950 761.400 400.050 762.600 ;
        RECT 388.950 761.100 391.050 761.400 ;
        RECT 397.950 760.800 400.050 761.400 ;
        RECT 416.400 761.400 427.050 762.600 ;
        RECT 302.400 758.400 309.600 759.000 ;
        RECT 338.400 758.400 366.600 759.600 ;
        RECT 173.400 755.400 178.050 757.050 ;
        RECT 145.950 754.800 148.050 755.400 ;
        RECT 174.000 754.950 178.050 755.400 ;
        RECT 181.950 756.450 184.050 756.900 ;
        RECT 187.950 756.450 190.050 756.900 ;
        RECT 181.950 755.250 190.050 756.450 ;
        RECT 181.950 754.800 184.050 755.250 ;
        RECT 187.950 754.800 190.050 755.250 ;
        RECT 205.950 756.600 208.050 757.050 ;
        RECT 211.950 756.600 214.050 756.900 ;
        RECT 205.950 755.400 214.050 756.600 ;
        RECT 205.950 754.950 208.050 755.400 ;
        RECT 211.950 754.800 214.050 755.400 ;
        RECT 238.950 756.600 241.050 756.900 ;
        RECT 256.950 756.600 259.050 757.050 ;
        RECT 238.950 755.400 259.050 756.600 ;
        RECT 238.950 754.800 241.050 755.400 ;
        RECT 256.950 754.950 259.050 755.400 ;
        RECT 274.800 754.800 276.900 756.900 ;
        RECT 277.950 756.600 280.050 757.050 ;
        RECT 286.950 756.600 289.050 756.900 ;
        RECT 277.950 755.400 289.050 756.600 ;
        RECT 277.950 754.950 280.050 755.400 ;
        RECT 286.950 754.800 289.050 755.400 ;
        RECT 154.950 753.600 157.050 754.050 ;
        RECT 163.950 753.600 166.050 754.050 ;
        RECT 169.950 753.600 172.050 754.050 ;
        RECT 275.400 753.600 276.600 754.800 ;
        RECT 302.400 754.050 303.600 758.400 ;
        RECT 304.950 756.600 307.050 757.050 ;
        RECT 310.950 756.600 313.050 756.900 ;
        RECT 304.950 755.400 313.050 756.600 ;
        RECT 304.950 754.950 307.050 755.400 ;
        RECT 310.950 754.800 313.050 755.400 ;
        RECT 325.950 756.600 328.050 757.050 ;
        RECT 334.950 756.600 337.050 756.900 ;
        RECT 325.950 755.400 337.050 756.600 ;
        RECT 325.950 754.950 328.050 755.400 ;
        RECT 334.950 754.800 337.050 755.400 ;
        RECT 349.950 756.450 352.050 756.900 ;
        RECT 358.950 756.450 361.050 756.900 ;
        RECT 349.950 755.250 361.050 756.450 ;
        RECT 365.400 756.600 366.600 758.400 ;
        RECT 373.950 756.600 376.050 756.900 ;
        RECT 365.400 755.400 376.050 756.600 ;
        RECT 349.950 754.800 352.050 755.250 ;
        RECT 358.950 754.800 361.050 755.250 ;
        RECT 373.950 754.800 376.050 755.400 ;
        RECT 406.950 756.600 409.050 756.900 ;
        RECT 416.400 756.600 417.600 761.400 ;
        RECT 424.950 761.100 427.050 761.400 ;
        RECT 439.950 762.750 442.050 763.200 ;
        RECT 445.950 762.750 448.050 763.200 ;
        RECT 439.950 761.550 448.050 762.750 ;
        RECT 439.950 761.100 442.050 761.550 ;
        RECT 445.950 761.100 448.050 761.550 ;
        RECT 502.950 762.600 505.050 763.050 ;
        RECT 502.950 761.400 522.600 762.600 ;
        RECT 502.950 760.950 505.050 761.400 ;
        RECT 481.950 759.600 484.050 760.200 ;
        RECT 467.400 758.400 484.050 759.600 ;
        RECT 521.400 759.600 522.600 761.400 ;
        RECT 530.400 760.050 531.600 764.400 ;
        RECT 607.950 763.950 610.050 764.400 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 521.400 758.400 528.600 759.600 ;
        RECT 406.950 755.400 417.600 756.600 ;
        RECT 418.950 756.600 421.050 757.050 ;
        RECT 442.950 756.600 445.050 757.050 ;
        RECT 418.950 755.400 445.050 756.600 ;
        RECT 406.950 754.800 409.050 755.400 ;
        RECT 418.950 754.950 421.050 755.400 ;
        RECT 442.950 754.950 445.050 755.400 ;
        RECT 154.950 752.400 172.050 753.600 ;
        RECT 154.950 751.950 157.050 752.400 ;
        RECT 163.950 751.950 166.050 752.400 ;
        RECT 169.950 751.950 172.050 752.400 ;
        RECT 245.400 752.400 276.600 753.600 ;
        RECT 298.950 752.400 303.600 754.050 ;
        RECT 379.950 753.600 382.050 754.050 ;
        RECT 394.950 753.600 397.050 753.900 ;
        RECT 379.950 752.400 397.050 753.600 ;
        RECT 245.400 751.050 246.600 752.400 ;
        RECT 298.950 751.950 303.000 752.400 ;
        RECT 379.950 751.950 382.050 752.400 ;
        RECT 394.950 751.800 397.050 752.400 ;
        RECT 427.950 753.600 430.050 754.050 ;
        RECT 467.400 753.600 468.600 758.400 ;
        RECT 481.950 758.100 484.050 758.400 ;
        RECT 527.400 756.600 528.600 758.400 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 562.950 758.100 565.050 760.200 ;
        RECT 538.950 756.600 541.050 757.050 ;
        RECT 527.400 755.400 541.050 756.600 ;
        RECT 538.950 754.950 541.050 755.400 ;
        RECT 427.950 752.400 468.600 753.600 ;
        RECT 511.950 753.600 514.050 754.050 ;
        RECT 517.950 753.600 520.050 754.050 ;
        RECT 511.950 752.400 520.050 753.600 ;
        RECT 427.950 751.950 430.050 752.400 ;
        RECT 511.950 751.950 514.050 752.400 ;
        RECT 517.950 751.950 520.050 752.400 ;
        RECT 535.950 753.600 538.050 754.050 ;
        RECT 563.400 753.600 564.600 758.100 ;
        RECT 607.950 756.600 610.050 757.050 ;
        RECT 617.400 756.600 618.600 761.100 ;
        RECT 620.400 756.900 621.600 766.950 ;
        RECT 622.950 765.600 625.050 766.050 ;
        RECT 640.950 765.600 643.050 766.050 ;
        RECT 622.950 764.400 643.050 765.600 ;
        RECT 622.950 763.950 625.050 764.400 ;
        RECT 640.950 763.950 643.050 764.400 ;
        RECT 652.950 765.600 655.050 766.050 ;
        RECT 667.950 765.600 670.050 766.050 ;
        RECT 652.950 764.400 670.050 765.600 ;
        RECT 652.950 763.950 655.050 764.400 ;
        RECT 667.950 763.950 670.050 764.400 ;
        RECT 682.950 765.600 685.050 766.050 ;
        RECT 688.950 765.600 691.050 766.050 ;
        RECT 682.950 764.400 691.050 765.600 ;
        RECT 682.950 763.950 685.050 764.400 ;
        RECT 688.950 763.950 691.050 764.400 ;
        RECT 643.950 762.600 646.050 763.200 ;
        RECT 641.400 761.400 646.050 762.600 ;
        RECT 641.400 759.600 642.600 761.400 ;
        RECT 643.950 761.100 646.050 761.400 ;
        RECT 679.950 762.600 682.050 763.050 ;
        RECT 724.950 762.600 727.050 763.200 ;
        RECT 679.950 761.400 727.050 762.600 ;
        RECT 679.950 760.950 682.050 761.400 ;
        RECT 724.950 761.100 727.050 761.400 ;
        RECT 730.950 762.600 733.050 763.050 ;
        RECT 748.950 762.600 751.050 763.050 ;
        RECT 781.950 762.600 784.050 763.050 ;
        RECT 730.950 761.400 784.050 762.600 ;
        RECT 629.400 759.000 642.600 759.600 ;
        RECT 628.950 758.400 642.600 759.000 ;
        RECT 725.400 759.600 726.600 761.100 ;
        RECT 730.950 760.950 733.050 761.400 ;
        RECT 748.950 760.950 751.050 761.400 ;
        RECT 781.950 760.950 784.050 761.400 ;
        RECT 814.950 762.750 817.050 763.200 ;
        RECT 820.950 762.750 823.050 763.200 ;
        RECT 814.950 761.550 823.050 762.750 ;
        RECT 814.950 761.100 817.050 761.550 ;
        RECT 820.950 761.100 823.050 761.550 ;
        RECT 826.950 760.950 829.050 763.050 ;
        RECT 832.950 761.100 835.050 763.200 ;
        RECT 838.950 762.750 841.050 763.200 ;
        RECT 844.950 762.750 847.050 763.200 ;
        RECT 838.950 761.550 847.050 762.750 ;
        RECT 838.950 761.100 841.050 761.550 ;
        RECT 844.950 761.100 847.050 761.550 ;
        RECT 853.950 761.100 856.050 763.200 ;
        RECT 874.950 761.100 877.050 763.200 ;
        RECT 907.950 762.750 910.050 763.200 ;
        RECT 934.950 762.750 937.050 763.200 ;
        RECT 907.950 761.550 937.050 762.750 ;
        RECT 907.950 761.100 910.050 761.550 ;
        RECT 934.950 761.100 937.050 761.550 ;
        RECT 725.400 758.400 768.600 759.600 ;
        RECT 607.950 755.400 618.600 756.600 ;
        RECT 607.950 754.950 610.050 755.400 ;
        RECT 619.950 754.800 622.050 756.900 ;
        RECT 628.950 754.950 631.050 758.400 ;
        RECT 640.950 756.600 643.050 756.900 ;
        RECT 652.950 756.600 655.050 757.050 ;
        RECT 737.400 756.900 738.600 758.400 ;
        RECT 640.950 755.400 655.050 756.600 ;
        RECT 640.950 754.800 643.050 755.400 ;
        RECT 652.950 754.950 655.050 755.400 ;
        RECT 736.950 754.800 739.050 756.900 ;
        RECT 742.950 756.450 745.050 756.900 ;
        RECT 748.950 756.450 751.050 756.900 ;
        RECT 742.950 755.250 751.050 756.450 ;
        RECT 742.950 754.800 745.050 755.250 ;
        RECT 748.950 754.800 751.050 755.250 ;
        RECT 754.950 756.450 757.050 756.900 ;
        RECT 763.950 756.450 766.050 756.900 ;
        RECT 754.950 755.250 766.050 756.450 ;
        RECT 767.400 756.600 768.600 758.400 ;
        RECT 827.400 757.050 828.600 760.950 ;
        RECT 778.950 756.600 781.050 756.900 ;
        RECT 767.400 755.400 781.050 756.600 ;
        RECT 754.950 754.800 757.050 755.250 ;
        RECT 763.950 754.800 766.050 755.250 ;
        RECT 778.950 754.800 781.050 755.400 ;
        RECT 796.950 756.450 799.050 756.900 ;
        RECT 811.950 756.450 814.050 756.900 ;
        RECT 796.950 755.250 814.050 756.450 ;
        RECT 796.950 754.800 799.050 755.250 ;
        RECT 811.950 754.800 814.050 755.250 ;
        RECT 826.950 754.950 829.050 757.050 ;
        RECT 535.950 752.400 564.600 753.600 ;
        RECT 601.950 753.600 604.050 754.050 ;
        RECT 613.950 753.600 616.050 754.050 ;
        RECT 601.950 752.400 616.050 753.600 ;
        RECT 535.950 751.950 538.050 752.400 ;
        RECT 601.950 751.950 604.050 752.400 ;
        RECT 613.950 751.950 616.050 752.400 ;
        RECT 661.950 753.600 664.050 754.050 ;
        RECT 715.950 753.600 718.050 754.050 ;
        RECT 661.950 752.400 718.050 753.600 ;
        RECT 749.400 753.600 750.600 754.800 ;
        RECT 787.950 753.600 790.050 754.050 ;
        RECT 749.400 752.400 790.050 753.600 ;
        RECT 661.950 751.950 664.050 752.400 ;
        RECT 715.950 751.950 718.050 752.400 ;
        RECT 787.950 751.950 790.050 752.400 ;
        RECT 814.950 753.600 817.050 754.050 ;
        RECT 820.950 753.600 823.050 754.050 ;
        RECT 814.950 752.400 823.050 753.600 ;
        RECT 833.400 753.600 834.600 761.100 ;
        RECT 854.400 757.050 855.600 761.100 ;
        RECT 850.950 755.400 855.600 757.050 ;
        RECT 850.950 754.950 855.000 755.400 ;
        RECT 875.400 754.050 876.600 761.100 ;
        RECT 919.950 756.600 922.050 757.050 ;
        RECT 928.950 756.600 931.050 756.900 ;
        RECT 919.950 755.400 931.050 756.600 ;
        RECT 919.950 754.950 922.050 755.400 ;
        RECT 928.950 754.800 931.050 755.400 ;
        RECT 838.950 753.600 841.050 754.050 ;
        RECT 833.400 752.400 841.050 753.600 ;
        RECT 814.950 751.950 817.050 752.400 ;
        RECT 820.950 751.950 823.050 752.400 ;
        RECT 838.950 751.950 841.050 752.400 ;
        RECT 859.950 753.600 862.050 754.050 ;
        RECT 859.950 752.400 873.600 753.600 ;
        RECT 859.950 751.950 862.050 752.400 ;
        RECT 4.950 750.600 7.050 751.050 ;
        RECT 16.950 750.600 19.050 751.050 ;
        RECT 4.950 749.400 19.050 750.600 ;
        RECT 4.950 748.950 7.050 749.400 ;
        RECT 16.950 748.950 19.050 749.400 ;
        RECT 52.950 750.600 55.050 751.050 ;
        RECT 217.950 750.600 220.050 751.050 ;
        RECT 244.950 750.600 247.050 751.050 ;
        RECT 52.950 749.400 90.600 750.600 ;
        RECT 52.950 748.950 55.050 749.400 ;
        RECT 55.950 747.600 58.050 748.050 ;
        RECT 85.950 747.600 88.050 748.050 ;
        RECT 55.950 746.400 88.050 747.600 ;
        RECT 89.400 747.600 90.600 749.400 ;
        RECT 217.950 749.400 247.050 750.600 ;
        RECT 217.950 748.950 220.050 749.400 ;
        RECT 244.950 748.950 247.050 749.400 ;
        RECT 268.950 750.600 271.050 751.050 ;
        RECT 280.950 750.600 283.050 751.050 ;
        RECT 268.950 749.400 283.050 750.600 ;
        RECT 268.950 748.950 271.050 749.400 ;
        RECT 280.950 748.950 283.050 749.400 ;
        RECT 295.950 750.600 298.050 751.050 ;
        RECT 322.950 750.600 325.050 751.050 ;
        RECT 295.950 749.400 325.050 750.600 ;
        RECT 295.950 748.950 298.050 749.400 ;
        RECT 322.950 748.950 325.050 749.400 ;
        RECT 442.950 750.600 445.050 751.050 ;
        RECT 512.400 750.600 513.600 751.950 ;
        RECT 442.950 749.400 513.600 750.600 ;
        RECT 619.950 750.600 622.050 751.050 ;
        RECT 634.950 750.600 637.050 751.050 ;
        RECT 619.950 749.400 637.050 750.600 ;
        RECT 442.950 748.950 445.050 749.400 ;
        RECT 619.950 748.950 622.050 749.400 ;
        RECT 634.950 748.950 637.050 749.400 ;
        RECT 664.950 750.600 667.050 751.050 ;
        RECT 670.950 750.600 673.050 751.050 ;
        RECT 664.950 749.400 673.050 750.600 ;
        RECT 664.950 748.950 667.050 749.400 ;
        RECT 670.950 748.950 673.050 749.400 ;
        RECT 697.950 750.600 700.050 751.050 ;
        RECT 721.950 750.600 724.050 751.050 ;
        RECT 697.950 749.400 724.050 750.600 ;
        RECT 697.950 748.950 700.050 749.400 ;
        RECT 721.950 748.950 724.050 749.400 ;
        RECT 805.950 750.600 808.050 751.050 ;
        RECT 826.950 750.600 829.050 751.050 ;
        RECT 805.950 749.400 829.050 750.600 ;
        RECT 805.950 748.950 808.050 749.400 ;
        RECT 826.950 748.950 829.050 749.400 ;
        RECT 844.950 750.600 847.050 751.050 ;
        RECT 856.950 750.600 859.050 751.050 ;
        RECT 844.950 749.400 859.050 750.600 ;
        RECT 872.400 750.600 873.600 752.400 ;
        RECT 874.950 751.950 877.050 754.050 ;
        RECT 886.950 753.600 889.050 754.050 ;
        RECT 895.950 753.600 898.050 754.050 ;
        RECT 886.950 752.400 898.050 753.600 ;
        RECT 886.950 751.950 889.050 752.400 ;
        RECT 895.950 751.950 898.050 752.400 ;
        RECT 883.950 750.600 886.050 751.050 ;
        RECT 872.400 749.400 886.050 750.600 ;
        RECT 844.950 748.950 847.050 749.400 ;
        RECT 856.950 748.950 859.050 749.400 ;
        RECT 883.950 748.950 886.050 749.400 ;
        RECT 904.950 750.600 907.050 751.050 ;
        RECT 916.950 750.600 919.050 751.050 ;
        RECT 904.950 749.400 919.050 750.600 ;
        RECT 904.950 748.950 907.050 749.400 ;
        RECT 916.950 748.950 919.050 749.400 ;
        RECT 925.950 750.600 928.050 751.050 ;
        RECT 934.950 750.600 937.050 751.050 ;
        RECT 925.950 749.400 937.050 750.600 ;
        RECT 925.950 748.950 928.050 749.400 ;
        RECT 934.950 748.950 937.050 749.400 ;
        RECT 184.950 747.600 187.050 748.050 ;
        RECT 89.400 746.400 187.050 747.600 ;
        RECT 55.950 745.950 58.050 746.400 ;
        RECT 85.950 745.950 88.050 746.400 ;
        RECT 184.950 745.950 187.050 746.400 ;
        RECT 193.950 747.600 196.050 748.050 ;
        RECT 226.950 747.600 229.050 748.050 ;
        RECT 193.950 746.400 229.050 747.600 ;
        RECT 193.950 745.950 196.050 746.400 ;
        RECT 226.950 745.950 229.050 746.400 ;
        RECT 346.950 747.600 349.050 748.050 ;
        RECT 406.950 747.600 409.050 748.050 ;
        RECT 346.950 746.400 409.050 747.600 ;
        RECT 346.950 745.950 349.050 746.400 ;
        RECT 406.950 745.950 409.050 746.400 ;
        RECT 415.950 747.600 418.050 748.050 ;
        RECT 430.950 747.600 433.050 748.050 ;
        RECT 415.950 746.400 433.050 747.600 ;
        RECT 415.950 745.950 418.050 746.400 ;
        RECT 430.950 745.950 433.050 746.400 ;
        RECT 460.950 747.600 463.050 748.050 ;
        RECT 514.950 747.600 517.050 748.050 ;
        RECT 460.950 746.400 517.050 747.600 ;
        RECT 460.950 745.950 463.050 746.400 ;
        RECT 514.950 745.950 517.050 746.400 ;
        RECT 538.950 747.600 541.050 748.050 ;
        RECT 577.950 747.600 580.050 748.050 ;
        RECT 538.950 746.400 580.050 747.600 ;
        RECT 538.950 745.950 541.050 746.400 ;
        RECT 577.950 745.950 580.050 746.400 ;
        RECT 595.950 747.600 598.050 748.050 ;
        RECT 862.950 747.600 865.050 748.050 ;
        RECT 595.950 746.400 865.050 747.600 ;
        RECT 595.950 745.950 598.050 746.400 ;
        RECT 862.950 745.950 865.050 746.400 ;
        RECT 37.950 744.600 40.050 745.050 ;
        RECT 32.400 743.400 40.050 744.600 ;
        RECT 4.950 741.600 7.050 742.050 ;
        RECT 32.400 741.600 33.600 743.400 ;
        RECT 37.950 742.950 40.050 743.400 ;
        RECT 73.950 744.600 76.050 745.050 ;
        RECT 91.950 744.600 94.050 745.050 ;
        RECT 73.950 743.400 94.050 744.600 ;
        RECT 73.950 742.950 76.050 743.400 ;
        RECT 91.950 742.950 94.050 743.400 ;
        RECT 118.950 744.600 121.050 745.050 ;
        RECT 160.950 744.600 163.050 745.050 ;
        RECT 118.950 743.400 163.050 744.600 ;
        RECT 118.950 742.950 121.050 743.400 ;
        RECT 160.950 742.950 163.050 743.400 ;
        RECT 178.950 744.600 181.050 745.050 ;
        RECT 190.950 744.600 193.050 745.050 ;
        RECT 178.950 743.400 193.050 744.600 ;
        RECT 178.950 742.950 181.050 743.400 ;
        RECT 190.950 742.950 193.050 743.400 ;
        RECT 244.950 744.600 247.050 745.050 ;
        RECT 274.950 744.600 277.050 745.050 ;
        RECT 244.950 743.400 277.050 744.600 ;
        RECT 244.950 742.950 247.050 743.400 ;
        RECT 274.950 742.950 277.050 743.400 ;
        RECT 283.950 744.600 286.050 745.050 ;
        RECT 316.950 744.600 319.050 745.050 ;
        RECT 283.950 743.400 319.050 744.600 ;
        RECT 283.950 742.950 286.050 743.400 ;
        RECT 316.950 742.950 319.050 743.400 ;
        RECT 322.950 744.600 325.050 745.050 ;
        RECT 445.950 744.600 448.050 745.050 ;
        RECT 322.950 743.400 448.050 744.600 ;
        RECT 322.950 742.950 325.050 743.400 ;
        RECT 445.950 742.950 448.050 743.400 ;
        RECT 481.950 744.600 484.050 745.050 ;
        RECT 502.950 744.600 505.050 745.050 ;
        RECT 481.950 743.400 505.050 744.600 ;
        RECT 481.950 742.950 484.050 743.400 ;
        RECT 502.950 742.950 505.050 743.400 ;
        RECT 520.950 744.600 523.050 745.050 ;
        RECT 574.950 744.600 577.050 745.050 ;
        RECT 520.950 743.400 577.050 744.600 ;
        RECT 520.950 742.950 523.050 743.400 ;
        RECT 574.950 742.950 577.050 743.400 ;
        RECT 598.950 744.600 601.050 745.050 ;
        RECT 610.950 744.600 613.050 745.050 ;
        RECT 598.950 743.400 613.050 744.600 ;
        RECT 598.950 742.950 601.050 743.400 ;
        RECT 610.950 742.950 613.050 743.400 ;
        RECT 622.950 744.600 625.050 745.050 ;
        RECT 661.950 744.600 664.050 745.050 ;
        RECT 622.950 743.400 664.050 744.600 ;
        RECT 622.950 742.950 625.050 743.400 ;
        RECT 661.950 742.950 664.050 743.400 ;
        RECT 691.950 744.600 694.050 745.050 ;
        RECT 835.950 744.600 838.050 745.050 ;
        RECT 691.950 743.400 838.050 744.600 ;
        RECT 691.950 742.950 694.050 743.400 ;
        RECT 835.950 742.950 838.050 743.400 ;
        RECT 847.950 744.600 850.050 745.050 ;
        RECT 859.950 744.600 862.050 745.050 ;
        RECT 847.950 743.400 862.050 744.600 ;
        RECT 847.950 742.950 850.050 743.400 ;
        RECT 859.950 742.950 862.050 743.400 ;
        RECT 865.950 744.600 868.050 745.050 ;
        RECT 937.950 744.600 940.050 745.050 ;
        RECT 865.950 743.400 940.050 744.600 ;
        RECT 865.950 742.950 868.050 743.400 ;
        RECT 937.950 742.950 940.050 743.400 ;
        RECT 4.950 740.400 33.600 741.600 ;
        RECT 109.950 741.600 112.050 742.050 ;
        RECT 130.950 741.600 133.050 742.050 ;
        RECT 109.950 740.400 133.050 741.600 ;
        RECT 4.950 739.950 7.050 740.400 ;
        RECT 109.950 739.950 112.050 740.400 ;
        RECT 130.950 739.950 133.050 740.400 ;
        RECT 208.950 741.600 211.050 742.050 ;
        RECT 229.950 741.600 232.050 742.050 ;
        RECT 208.950 740.400 232.050 741.600 ;
        RECT 208.950 739.950 211.050 740.400 ;
        RECT 229.950 739.950 232.050 740.400 ;
        RECT 319.950 741.600 322.050 742.050 ;
        RECT 367.950 741.600 370.050 742.050 ;
        RECT 466.950 741.600 469.050 742.050 ;
        RECT 319.950 740.400 370.050 741.600 ;
        RECT 319.950 739.950 322.050 740.400 ;
        RECT 367.950 739.950 370.050 740.400 ;
        RECT 449.400 740.400 469.050 741.600 ;
        RECT 265.950 738.600 268.050 739.050 ;
        RECT 292.950 738.600 295.050 739.050 ;
        RECT 265.950 737.400 295.050 738.600 ;
        RECT 265.950 736.950 268.050 737.400 ;
        RECT 292.950 736.950 295.050 737.400 ;
        RECT 307.950 738.600 310.050 739.050 ;
        RECT 316.950 738.600 319.050 739.050 ;
        RECT 307.950 737.400 319.050 738.600 ;
        RECT 307.950 736.950 310.050 737.400 ;
        RECT 316.950 736.950 319.050 737.400 ;
        RECT 337.950 738.600 340.050 739.050 ;
        RECT 343.950 738.600 346.050 739.050 ;
        RECT 337.950 737.400 346.050 738.600 ;
        RECT 337.950 736.950 340.050 737.400 ;
        RECT 343.950 736.950 346.050 737.400 ;
        RECT 352.950 738.600 355.050 739.050 ;
        RECT 361.950 738.600 364.050 739.050 ;
        RECT 373.950 738.600 376.050 739.050 ;
        RECT 352.950 737.400 376.050 738.600 ;
        RECT 352.950 736.950 355.050 737.400 ;
        RECT 361.950 736.950 364.050 737.400 ;
        RECT 373.950 736.950 376.050 737.400 ;
        RECT 388.950 738.600 391.050 739.050 ;
        RECT 403.950 738.600 406.050 739.050 ;
        RECT 388.950 737.400 406.050 738.600 ;
        RECT 388.950 736.950 391.050 737.400 ;
        RECT 403.950 736.950 406.050 737.400 ;
        RECT 433.950 738.600 436.050 739.050 ;
        RECT 449.400 738.600 450.600 740.400 ;
        RECT 466.950 739.950 469.050 740.400 ;
        RECT 502.950 741.600 505.050 741.900 ;
        RECT 538.950 741.600 541.050 742.050 ;
        RECT 502.950 740.400 541.050 741.600 ;
        RECT 502.950 739.800 505.050 740.400 ;
        RECT 538.950 739.950 541.050 740.400 ;
        RECT 556.950 741.600 559.050 742.050 ;
        RECT 616.950 741.600 619.050 742.050 ;
        RECT 556.950 740.400 619.050 741.600 ;
        RECT 556.950 739.950 559.050 740.400 ;
        RECT 616.950 739.950 619.050 740.400 ;
        RECT 628.950 741.600 631.050 742.050 ;
        RECT 634.950 741.600 637.050 742.050 ;
        RECT 649.950 741.600 652.050 742.050 ;
        RECT 628.950 740.400 652.050 741.600 ;
        RECT 628.950 739.950 631.050 740.400 ;
        RECT 634.950 739.950 637.050 740.400 ;
        RECT 649.950 739.950 652.050 740.400 ;
        RECT 433.950 737.400 450.600 738.600 ;
        RECT 466.950 738.600 469.050 738.900 ;
        RECT 553.950 738.600 556.050 739.050 ;
        RECT 658.950 738.600 661.050 742.050 ;
        RECT 706.950 741.600 709.050 742.050 ;
        RECT 772.950 741.600 775.050 742.050 ;
        RECT 706.950 740.400 775.050 741.600 ;
        RECT 706.950 739.950 709.050 740.400 ;
        RECT 772.950 739.950 775.050 740.400 ;
        RECT 820.950 741.600 823.050 742.050 ;
        RECT 829.950 741.600 832.050 742.050 ;
        RECT 820.950 740.400 832.050 741.600 ;
        RECT 820.950 739.950 823.050 740.400 ;
        RECT 829.950 739.950 832.050 740.400 ;
        RECT 466.950 737.400 556.050 738.600 ;
        RECT 433.950 736.950 436.050 737.400 ;
        RECT 466.950 736.800 469.050 737.400 ;
        RECT 553.950 736.950 556.050 737.400 ;
        RECT 632.400 738.000 661.050 738.600 ;
        RECT 736.950 738.600 739.050 739.050 ;
        RECT 760.950 738.600 763.050 739.050 ;
        RECT 632.400 737.400 660.600 738.000 ;
        RECT 736.950 737.400 763.050 738.600 ;
        RECT 632.400 736.050 633.600 737.400 ;
        RECT 736.950 736.950 739.050 737.400 ;
        RECT 760.950 736.950 763.050 737.400 ;
        RECT 784.950 738.600 787.050 739.050 ;
        RECT 805.950 738.600 808.050 739.050 ;
        RECT 835.950 738.600 838.050 739.050 ;
        RECT 850.950 738.600 853.050 739.050 ;
        RECT 784.950 737.400 853.050 738.600 ;
        RECT 784.950 736.950 787.050 737.400 ;
        RECT 805.950 736.950 808.050 737.400 ;
        RECT 835.950 736.950 838.050 737.400 ;
        RECT 850.950 736.950 853.050 737.400 ;
        RECT 892.950 738.600 895.050 739.050 ;
        RECT 919.950 738.600 922.050 739.050 ;
        RECT 892.950 737.400 922.050 738.600 ;
        RECT 892.950 736.950 895.050 737.400 ;
        RECT 919.950 736.950 922.050 737.400 ;
        RECT 34.950 735.600 37.050 736.050 ;
        RECT 64.950 735.600 67.050 736.050 ;
        RECT 118.950 735.600 121.050 736.050 ;
        RECT 34.950 734.400 121.050 735.600 ;
        RECT 34.950 733.950 37.050 734.400 ;
        RECT 64.950 733.950 67.050 734.400 ;
        RECT 118.950 733.950 121.050 734.400 ;
        RECT 124.950 735.600 127.050 736.050 ;
        RECT 133.950 735.600 136.050 736.050 ;
        RECT 124.950 734.400 136.050 735.600 ;
        RECT 124.950 733.950 127.050 734.400 ;
        RECT 133.950 733.950 136.050 734.400 ;
        RECT 172.950 735.600 175.050 736.050 ;
        RECT 205.950 735.600 208.050 736.050 ;
        RECT 172.950 734.400 208.050 735.600 ;
        RECT 172.950 733.950 175.050 734.400 ;
        RECT 205.950 733.950 208.050 734.400 ;
        RECT 223.950 735.600 226.050 736.050 ;
        RECT 238.950 735.600 241.050 736.050 ;
        RECT 223.950 734.400 241.050 735.600 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 238.950 733.950 241.050 734.400 ;
        RECT 280.950 735.600 283.050 736.050 ;
        RECT 301.950 735.600 304.050 736.050 ;
        RECT 280.950 734.400 304.050 735.600 ;
        RECT 280.950 733.950 283.050 734.400 ;
        RECT 301.950 733.950 304.050 734.400 ;
        RECT 328.950 735.600 331.050 736.050 ;
        RECT 340.950 735.600 343.050 736.050 ;
        RECT 328.950 734.400 343.050 735.600 ;
        RECT 328.950 733.950 331.050 734.400 ;
        RECT 340.950 733.950 343.050 734.400 ;
        RECT 529.950 735.600 532.050 736.050 ;
        RECT 550.950 735.600 553.050 736.050 ;
        RECT 631.950 735.600 634.050 736.050 ;
        RECT 529.950 734.400 553.050 735.600 ;
        RECT 529.950 733.950 532.050 734.400 ;
        RECT 550.950 733.950 553.050 734.400 ;
        RECT 593.400 734.400 634.050 735.600 ;
        RECT 593.400 733.050 594.600 734.400 ;
        RECT 631.950 733.950 634.050 734.400 ;
        RECT 712.950 735.600 715.050 736.050 ;
        RECT 733.950 735.600 736.050 736.050 ;
        RECT 712.950 734.400 736.050 735.600 ;
        RECT 712.950 733.950 715.050 734.400 ;
        RECT 733.950 733.950 736.050 734.400 ;
        RECT 811.950 735.600 814.050 736.050 ;
        RECT 826.950 735.600 829.050 736.050 ;
        RECT 811.950 734.400 829.050 735.600 ;
        RECT 811.950 733.950 814.050 734.400 ;
        RECT 826.950 733.950 829.050 734.400 ;
        RECT 862.950 735.600 865.050 736.050 ;
        RECT 880.950 735.600 883.050 736.050 ;
        RECT 862.950 734.400 883.050 735.600 ;
        RECT 862.950 733.950 865.050 734.400 ;
        RECT 880.950 733.950 883.050 734.400 ;
        RECT 43.950 732.600 46.050 733.050 ;
        RECT 211.950 732.600 214.050 733.050 ;
        RECT 220.950 732.600 223.050 733.050 ;
        RECT 43.950 731.400 63.600 732.600 ;
        RECT 43.950 730.950 46.050 731.400 ;
        RECT 22.950 729.750 25.050 730.200 ;
        RECT 31.950 729.750 34.050 730.200 ;
        RECT 22.950 729.600 34.050 729.750 ;
        RECT 58.950 729.600 61.050 730.200 ;
        RECT 22.950 728.550 61.050 729.600 ;
        RECT 22.950 728.100 25.050 728.550 ;
        RECT 31.950 728.400 61.050 728.550 ;
        RECT 62.400 729.600 63.600 731.400 ;
        RECT 211.950 731.400 223.050 732.600 ;
        RECT 211.950 730.950 214.050 731.400 ;
        RECT 220.950 730.950 223.050 731.400 ;
        RECT 277.950 732.600 280.050 733.050 ;
        RECT 283.950 732.600 286.050 732.900 ;
        RECT 319.950 732.600 322.050 733.050 ;
        RECT 352.950 732.600 355.050 733.050 ;
        RECT 277.950 731.400 322.050 732.600 ;
        RECT 277.950 730.950 280.050 731.400 ;
        RECT 283.950 730.800 286.050 731.400 ;
        RECT 319.950 730.950 322.050 731.400 ;
        RECT 332.400 731.400 355.050 732.600 ;
        RECT 70.950 729.750 73.050 730.200 ;
        RECT 76.950 729.750 79.050 730.200 ;
        RECT 62.400 728.400 69.600 729.600 ;
        RECT 31.950 728.100 34.050 728.400 ;
        RECT 58.950 728.100 61.050 728.400 ;
        RECT 68.400 726.600 69.600 728.400 ;
        RECT 70.950 728.550 79.050 729.750 ;
        RECT 70.950 728.100 73.050 728.550 ;
        RECT 76.950 728.100 79.050 728.550 ;
        RECT 88.950 729.600 91.050 730.200 ;
        RECT 106.950 729.600 109.050 730.200 ;
        RECT 88.950 728.400 109.050 729.600 ;
        RECT 88.950 728.100 91.050 728.400 ;
        RECT 106.950 728.100 109.050 728.400 ;
        RECT 112.950 729.600 115.050 730.200 ;
        RECT 118.950 729.600 121.050 730.050 ;
        RECT 112.950 728.400 121.050 729.600 ;
        RECT 112.950 728.100 115.050 728.400 ;
        RECT 118.950 727.950 121.050 728.400 ;
        RECT 124.950 729.750 127.050 730.200 ;
        RECT 130.950 729.750 133.050 730.200 ;
        RECT 124.950 728.550 133.050 729.750 ;
        RECT 124.950 728.100 127.050 728.550 ;
        RECT 130.950 728.100 133.050 728.550 ;
        RECT 139.950 729.750 142.050 730.200 ;
        RECT 178.950 729.750 181.050 730.200 ;
        RECT 139.950 728.550 181.050 729.750 ;
        RECT 139.950 728.100 142.050 728.550 ;
        RECT 178.950 728.100 181.050 728.550 ;
        RECT 196.950 728.100 199.050 730.200 ;
        RECT 68.400 725.400 75.600 726.600 ;
        RECT 31.950 723.600 34.050 724.050 ;
        RECT 37.950 723.600 40.050 723.900 ;
        RECT 31.950 722.400 40.050 723.600 ;
        RECT 74.400 723.600 75.600 725.400 ;
        RECT 79.950 723.600 82.050 723.900 ;
        RECT 74.400 722.400 82.050 723.600 ;
        RECT 31.950 721.950 34.050 722.400 ;
        RECT 37.950 721.800 40.050 722.400 ;
        RECT 79.950 721.800 82.050 722.400 ;
        RECT 100.950 723.600 103.050 724.050 ;
        RECT 109.950 723.600 112.050 723.900 ;
        RECT 127.950 723.600 130.050 723.900 ;
        RECT 100.950 722.400 130.050 723.600 ;
        RECT 100.950 721.950 103.050 722.400 ;
        RECT 109.950 721.800 112.050 722.400 ;
        RECT 127.950 721.800 130.050 722.400 ;
        RECT 136.950 723.450 139.050 723.900 ;
        RECT 142.950 723.450 145.050 723.900 ;
        RECT 136.950 722.250 145.050 723.450 ;
        RECT 136.950 721.800 139.050 722.250 ;
        RECT 142.950 721.800 145.050 722.250 ;
        RECT 175.950 723.600 178.050 723.900 ;
        RECT 197.400 723.600 198.600 728.100 ;
        RECT 202.950 727.950 205.050 730.050 ;
        RECT 229.950 729.750 232.050 730.200 ;
        RECT 244.950 729.750 247.050 730.200 ;
        RECT 229.950 728.550 247.050 729.750 ;
        RECT 229.950 728.100 232.050 728.550 ;
        RECT 244.950 728.100 247.050 728.550 ;
        RECT 203.400 724.050 204.600 727.950 ;
        RECT 274.950 726.600 277.050 727.050 ;
        RECT 280.950 726.600 283.050 730.050 ;
        RECT 292.950 729.600 295.050 730.050 ;
        RECT 313.950 729.600 316.050 730.050 ;
        RECT 292.950 728.400 316.050 729.600 ;
        RECT 292.950 727.950 295.050 728.400 ;
        RECT 313.950 727.950 316.050 728.400 ;
        RECT 332.400 726.600 333.600 731.400 ;
        RECT 352.950 730.950 355.050 731.400 ;
        RECT 373.950 732.600 376.050 733.050 ;
        RECT 421.950 732.600 424.050 733.050 ;
        RECT 439.950 732.600 442.050 733.050 ;
        RECT 466.950 732.600 469.050 733.050 ;
        RECT 525.000 732.600 529.050 733.050 ;
        RECT 373.950 731.400 469.050 732.600 ;
        RECT 373.950 730.950 376.050 731.400 ;
        RECT 421.950 730.950 424.050 731.400 ;
        RECT 439.950 730.950 442.050 731.400 ;
        RECT 466.950 730.950 469.050 731.400 ;
        RECT 524.400 730.950 529.050 732.600 ;
        RECT 553.950 732.600 556.050 733.050 ;
        RECT 592.950 732.600 595.050 733.050 ;
        RECT 553.950 731.400 595.050 732.600 ;
        RECT 553.950 730.950 556.050 731.400 ;
        RECT 592.950 730.950 595.050 731.400 ;
        RECT 616.950 732.600 619.050 733.050 ;
        RECT 745.950 732.600 748.050 732.900 ;
        RECT 754.950 732.600 757.050 733.050 ;
        RECT 616.950 731.400 684.600 732.600 ;
        RECT 616.950 730.950 619.050 731.400 ;
        RECT 340.950 729.600 345.000 730.050 ;
        RECT 370.950 729.600 373.050 730.200 ;
        RECT 382.800 729.600 384.900 730.050 ;
        RECT 340.950 727.950 345.600 729.600 ;
        RECT 370.950 728.400 384.900 729.600 ;
        RECT 370.950 728.100 373.050 728.400 ;
        RECT 382.800 727.950 384.900 728.400 ;
        RECT 274.950 726.000 283.050 726.600 ;
        RECT 302.400 726.000 333.600 726.600 ;
        RECT 274.950 725.400 282.600 726.000 ;
        RECT 301.950 725.400 333.600 726.000 ;
        RECT 274.950 724.950 277.050 725.400 ;
        RECT 175.950 722.400 198.600 723.600 ;
        RECT 175.950 721.800 178.050 722.400 ;
        RECT 202.950 721.950 205.050 724.050 ;
        RECT 226.950 723.450 229.050 723.900 ;
        RECT 235.950 723.450 238.050 723.900 ;
        RECT 226.950 722.250 238.050 723.450 ;
        RECT 226.950 721.800 229.050 722.250 ;
        RECT 235.950 721.800 238.050 722.250 ;
        RECT 301.950 721.950 304.050 725.400 ;
        RECT 319.950 723.600 322.050 724.050 ;
        RECT 332.400 723.900 333.600 725.400 ;
        RECT 344.400 723.900 345.600 727.950 ;
        RECT 385.950 726.600 388.050 730.050 ;
        RECT 415.950 729.600 418.050 730.200 ;
        RECT 374.400 726.000 388.050 726.600 ;
        RECT 398.400 728.400 418.050 729.600 ;
        RECT 374.400 725.400 387.600 726.000 ;
        RECT 374.400 723.900 375.600 725.400 ;
        RECT 398.400 723.900 399.600 728.400 ;
        RECT 415.950 728.100 418.050 728.400 ;
        RECT 436.950 729.600 439.050 730.200 ;
        RECT 481.950 729.600 484.050 730.200 ;
        RECT 524.400 729.600 525.600 730.950 ;
        RECT 532.800 729.600 534.900 730.050 ;
        RECT 436.950 728.400 484.050 729.600 ;
        RECT 436.950 728.100 439.050 728.400 ;
        RECT 481.950 728.100 484.050 728.400 ;
        RECT 509.400 728.400 525.600 729.600 ;
        RECT 527.400 728.400 534.900 729.600 ;
        RECT 325.950 723.600 328.050 723.900 ;
        RECT 319.950 722.400 328.050 723.600 ;
        RECT 319.950 721.950 322.050 722.400 ;
        RECT 325.950 721.800 328.050 722.400 ;
        RECT 331.950 721.800 334.050 723.900 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 373.950 721.800 376.050 723.900 ;
        RECT 397.950 721.800 400.050 723.900 ;
        RECT 448.950 723.450 451.050 723.900 ;
        RECT 457.950 723.450 460.050 723.900 ;
        RECT 448.950 722.250 460.050 723.450 ;
        RECT 448.950 721.800 451.050 722.250 ;
        RECT 457.950 721.800 460.050 722.250 ;
        RECT 487.950 723.600 490.050 723.900 ;
        RECT 499.950 723.600 502.050 723.900 ;
        RECT 487.950 722.400 502.050 723.600 ;
        RECT 487.950 721.800 490.050 722.400 ;
        RECT 499.950 721.800 502.050 722.400 ;
        RECT 505.950 723.600 508.050 723.900 ;
        RECT 509.400 723.600 510.600 728.400 ;
        RECT 527.400 723.900 528.600 728.400 ;
        RECT 532.800 727.950 534.900 728.400 ;
        RECT 535.950 729.600 538.050 729.900 ;
        RECT 541.950 729.600 544.050 730.050 ;
        RECT 535.950 728.400 544.050 729.600 ;
        RECT 535.950 727.800 538.050 728.400 ;
        RECT 541.950 727.950 544.050 728.400 ;
        RECT 547.950 729.600 550.050 730.200 ;
        RECT 559.950 729.600 562.050 730.050 ;
        RECT 547.950 728.400 562.050 729.600 ;
        RECT 547.950 728.100 550.050 728.400 ;
        RECT 559.950 727.950 562.050 728.400 ;
        RECT 565.950 729.750 568.050 730.200 ;
        RECT 577.950 729.750 580.050 730.200 ;
        RECT 565.950 728.550 580.050 729.750 ;
        RECT 565.950 728.100 568.050 728.550 ;
        RECT 577.950 728.100 580.050 728.550 ;
        RECT 595.950 729.750 598.050 730.200 ;
        RECT 607.950 729.750 610.050 730.200 ;
        RECT 595.950 728.550 610.050 729.750 ;
        RECT 595.950 728.100 598.050 728.550 ;
        RECT 607.950 728.100 610.050 728.550 ;
        RECT 683.400 729.600 684.600 731.400 ;
        RECT 745.950 731.400 757.050 732.600 ;
        RECT 745.950 730.800 748.050 731.400 ;
        RECT 754.950 730.950 757.050 731.400 ;
        RECT 820.800 730.950 822.900 733.050 ;
        RECT 823.950 732.600 828.000 733.050 ;
        RECT 850.950 732.600 853.050 733.050 ;
        RECT 865.950 732.600 868.050 733.050 ;
        RECT 823.950 730.950 828.600 732.600 ;
        RECT 850.950 731.400 868.050 732.600 ;
        RECT 850.950 730.950 853.050 731.400 ;
        RECT 865.950 730.950 868.050 731.400 ;
        RECT 721.950 729.600 724.050 730.200 ;
        RECT 727.950 729.600 730.050 730.200 ;
        RECT 683.400 728.400 724.050 729.600 ;
        RECT 721.950 728.100 724.050 728.400 ;
        RECT 725.400 728.400 730.050 729.600 ;
        RECT 619.950 725.100 622.050 727.200 ;
        RECT 658.950 726.600 661.050 727.050 ;
        RECT 670.950 726.600 673.050 727.050 ;
        RECT 725.400 726.600 726.600 728.400 ;
        RECT 727.950 728.100 730.050 728.400 ;
        RECT 757.950 729.600 760.050 730.050 ;
        RECT 766.950 729.600 769.050 730.200 ;
        RECT 757.950 728.400 769.050 729.600 ;
        RECT 757.950 727.950 760.050 728.400 ;
        RECT 766.950 728.100 769.050 728.400 ;
        RECT 775.950 729.750 778.050 730.200 ;
        RECT 787.950 729.750 790.050 730.200 ;
        RECT 775.950 728.550 790.050 729.750 ;
        RECT 775.950 728.100 778.050 728.550 ;
        RECT 787.950 728.100 790.050 728.550 ;
        RECT 799.950 729.600 802.050 730.050 ;
        RECT 811.950 729.600 814.050 730.050 ;
        RECT 799.950 728.400 814.050 729.600 ;
        RECT 799.950 727.950 802.050 728.400 ;
        RECT 811.950 727.950 814.050 728.400 ;
        RECT 658.950 725.400 673.050 726.600 ;
        RECT 505.950 722.400 510.600 723.600 ;
        RECT 514.950 723.450 517.050 723.900 ;
        RECT 520.950 723.450 523.050 723.900 ;
        RECT 505.950 721.800 508.050 722.400 ;
        RECT 514.950 722.250 523.050 723.450 ;
        RECT 514.950 721.800 517.050 722.250 ;
        RECT 520.950 721.800 523.050 722.250 ;
        RECT 526.950 721.800 529.050 723.900 ;
        RECT 538.950 723.450 541.050 723.900 ;
        RECT 544.950 723.450 547.050 723.900 ;
        RECT 538.950 722.250 547.050 723.450 ;
        RECT 538.950 721.800 541.050 722.250 ;
        RECT 544.950 721.800 547.050 722.250 ;
        RECT 550.950 723.600 553.050 723.900 ;
        RECT 562.950 723.600 565.050 724.050 ;
        RECT 571.950 723.600 574.050 723.900 ;
        RECT 550.950 722.400 574.050 723.600 ;
        RECT 620.400 723.600 621.600 725.100 ;
        RECT 658.950 724.950 661.050 725.400 ;
        RECT 670.950 724.950 673.050 725.400 ;
        RECT 704.400 725.400 726.600 726.600 ;
        RECT 655.950 723.600 658.050 724.050 ;
        RECT 704.400 723.900 705.600 725.400 ;
        RECT 821.400 724.050 822.600 730.950 ;
        RECT 620.400 722.400 658.050 723.600 ;
        RECT 550.950 721.800 553.050 722.400 ;
        RECT 562.950 721.950 565.050 722.400 ;
        RECT 571.950 721.800 574.050 722.400 ;
        RECT 655.950 721.950 658.050 722.400 ;
        RECT 703.950 721.800 706.050 723.900 ;
        RECT 712.950 723.450 715.050 723.900 ;
        RECT 718.950 723.450 721.050 723.900 ;
        RECT 712.950 722.250 721.050 723.450 ;
        RECT 712.950 721.800 715.050 722.250 ;
        RECT 718.950 721.800 721.050 722.250 ;
        RECT 730.950 723.600 733.050 723.900 ;
        RECT 748.950 723.600 751.050 723.900 ;
        RECT 730.950 722.400 751.050 723.600 ;
        RECT 730.950 721.800 733.050 722.400 ;
        RECT 748.950 721.800 751.050 722.400 ;
        RECT 784.950 723.600 787.050 723.900 ;
        RECT 784.950 722.400 789.600 723.600 ;
        RECT 784.950 721.800 787.050 722.400 ;
        RECT 7.950 720.600 10.050 721.050 ;
        RECT 19.950 720.600 22.050 721.050 ;
        RECT 7.950 719.400 22.050 720.600 ;
        RECT 7.950 718.950 10.050 719.400 ;
        RECT 19.950 718.950 22.050 719.400 ;
        RECT 139.950 720.600 142.050 721.050 ;
        RECT 148.950 720.600 151.050 721.050 ;
        RECT 139.950 719.400 151.050 720.600 ;
        RECT 139.950 718.950 142.050 719.400 ;
        RECT 148.950 718.950 151.050 719.400 ;
        RECT 382.950 720.600 385.050 721.050 ;
        RECT 391.800 720.600 393.900 721.050 ;
        RECT 382.950 719.400 393.900 720.600 ;
        RECT 382.950 718.950 385.050 719.400 ;
        RECT 391.800 718.950 393.900 719.400 ;
        RECT 394.950 720.600 397.050 721.050 ;
        RECT 418.800 720.600 420.900 721.050 ;
        RECT 394.950 719.400 420.900 720.600 ;
        RECT 394.950 718.950 397.050 719.400 ;
        RECT 418.800 718.950 420.900 719.400 ;
        RECT 421.950 720.600 424.050 721.050 ;
        RECT 430.950 720.600 433.050 721.050 ;
        RECT 421.950 719.400 433.050 720.600 ;
        RECT 421.950 718.950 424.050 719.400 ;
        RECT 430.950 718.950 433.050 719.400 ;
        RECT 463.950 720.600 466.050 721.050 ;
        RECT 484.950 720.600 487.050 721.050 ;
        RECT 697.950 720.600 700.050 721.050 ;
        RECT 463.950 719.400 487.050 720.600 ;
        RECT 463.950 718.950 466.050 719.400 ;
        RECT 484.950 718.950 487.050 719.400 ;
        RECT 689.400 719.400 700.050 720.600 ;
        RECT 13.950 717.600 16.050 718.050 ;
        RECT 34.950 717.600 37.050 718.050 ;
        RECT 13.950 716.400 37.050 717.600 ;
        RECT 13.950 715.950 16.050 716.400 ;
        RECT 34.950 715.950 37.050 716.400 ;
        RECT 64.950 717.600 67.050 718.050 ;
        RECT 70.950 717.600 73.050 718.050 ;
        RECT 103.950 717.600 106.050 718.050 ;
        RECT 115.950 717.600 118.050 718.050 ;
        RECT 133.950 717.600 136.050 718.050 ;
        RECT 64.950 716.400 136.050 717.600 ;
        RECT 149.400 717.600 150.600 718.950 ;
        RECT 199.950 717.600 202.050 718.050 ;
        RECT 149.400 716.400 202.050 717.600 ;
        RECT 64.950 715.950 67.050 716.400 ;
        RECT 70.950 715.950 73.050 716.400 ;
        RECT 103.950 715.950 106.050 716.400 ;
        RECT 115.950 715.950 118.050 716.400 ;
        RECT 133.950 715.950 136.050 716.400 ;
        RECT 199.950 715.950 202.050 716.400 ;
        RECT 235.950 717.600 238.050 718.050 ;
        RECT 295.950 717.600 298.050 718.050 ;
        RECT 235.950 716.400 298.050 717.600 ;
        RECT 235.950 715.950 238.050 716.400 ;
        RECT 295.950 715.950 298.050 716.400 ;
        RECT 328.950 717.600 331.050 718.050 ;
        RECT 337.950 717.600 340.050 718.050 ;
        RECT 402.000 717.600 405.900 718.050 ;
        RECT 328.950 716.400 340.050 717.600 ;
        RECT 328.950 715.950 331.050 716.400 ;
        RECT 337.950 715.950 340.050 716.400 ;
        RECT 401.400 715.950 405.900 717.600 ;
        RECT 406.950 717.600 409.050 718.050 ;
        RECT 689.400 717.600 690.600 719.400 ;
        RECT 697.950 718.950 700.050 719.400 ;
        RECT 769.950 720.600 772.050 721.050 ;
        RECT 781.950 720.600 784.050 721.050 ;
        RECT 769.950 719.400 784.050 720.600 ;
        RECT 788.400 720.600 789.600 722.400 ;
        RECT 820.950 721.950 823.050 724.050 ;
        RECT 827.400 723.900 828.600 730.950 ;
        RECT 834.000 729.600 838.050 730.050 ;
        RECT 833.400 727.950 838.050 729.600 ;
        RECT 841.950 729.600 844.050 730.050 ;
        RECT 856.950 729.600 859.050 730.200 ;
        RECT 892.950 729.600 895.050 730.200 ;
        RECT 898.950 729.600 901.050 730.200 ;
        RECT 841.950 728.400 859.050 729.600 ;
        RECT 841.950 727.950 844.050 728.400 ;
        RECT 856.950 728.100 859.050 728.400 ;
        RECT 869.400 728.400 895.050 729.600 ;
        RECT 833.400 723.900 834.600 727.950 ;
        RECT 869.400 726.600 870.600 728.400 ;
        RECT 892.950 728.100 895.050 728.400 ;
        RECT 896.400 728.400 901.050 729.600 ;
        RECT 896.400 726.600 897.600 728.400 ;
        RECT 898.950 728.100 901.050 728.400 ;
        RECT 910.950 727.950 913.050 730.050 ;
        RECT 928.950 729.750 931.050 730.200 ;
        RECT 943.950 729.750 946.050 730.200 ;
        RECT 928.950 728.550 946.050 729.750 ;
        RECT 928.950 728.100 931.050 728.550 ;
        RECT 943.950 728.100 946.050 728.550 ;
        RECT 860.400 726.000 870.600 726.600 ;
        RECT 859.950 725.400 870.600 726.000 ;
        RECT 872.400 725.400 897.600 726.600 ;
        RECT 826.950 721.800 829.050 723.900 ;
        RECT 832.950 721.800 835.050 723.900 ;
        RECT 859.950 721.950 862.050 725.400 ;
        RECT 872.400 723.600 873.600 725.400 ;
        RECT 863.400 722.400 873.600 723.600 ;
        RECT 901.950 723.600 904.050 723.900 ;
        RECT 907.950 723.600 910.050 724.050 ;
        RECT 901.950 722.400 910.050 723.600 ;
        RECT 802.950 720.600 805.050 721.050 ;
        RECT 788.400 719.400 805.050 720.600 ;
        RECT 769.950 718.950 772.050 719.400 ;
        RECT 781.950 718.950 784.050 719.400 ;
        RECT 802.950 718.950 805.050 719.400 ;
        RECT 853.950 720.600 856.050 721.050 ;
        RECT 863.400 720.600 864.600 722.400 ;
        RECT 901.950 721.800 904.050 722.400 ;
        RECT 907.950 721.950 910.050 722.400 ;
        RECT 853.950 719.400 864.600 720.600 ;
        RECT 889.950 720.600 892.050 721.050 ;
        RECT 901.950 720.600 904.050 721.050 ;
        RECT 889.950 719.400 904.050 720.600 ;
        RECT 853.950 718.950 856.050 719.400 ;
        RECT 889.950 718.950 892.050 719.400 ;
        RECT 901.950 718.950 904.050 719.400 ;
        RECT 406.950 716.400 690.600 717.600 ;
        RECT 808.950 717.600 811.050 718.050 ;
        RECT 847.950 717.600 850.050 718.050 ;
        RECT 808.950 716.400 850.050 717.600 ;
        RECT 406.950 715.950 409.050 716.400 ;
        RECT 808.950 715.950 811.050 716.400 ;
        RECT 847.950 715.950 850.050 716.400 ;
        RECT 862.950 717.600 865.050 718.050 ;
        RECT 904.950 717.600 907.050 718.050 ;
        RECT 862.950 716.400 907.050 717.600 ;
        RECT 911.400 717.600 912.600 727.950 ;
        RECT 916.950 723.600 919.050 723.900 ;
        RECT 934.950 723.600 937.050 723.900 ;
        RECT 916.950 722.400 937.050 723.600 ;
        RECT 916.950 721.800 919.050 722.400 ;
        RECT 934.950 721.800 937.050 722.400 ;
        RECT 940.950 723.450 943.050 723.900 ;
        RECT 946.950 723.450 949.050 723.900 ;
        RECT 940.950 722.250 949.050 723.450 ;
        RECT 940.950 721.800 943.050 722.250 ;
        RECT 946.950 721.800 949.050 722.250 ;
        RECT 919.950 717.600 922.050 718.050 ;
        RECT 911.400 716.400 922.050 717.600 ;
        RECT 862.950 715.950 865.050 716.400 ;
        RECT 904.950 715.950 907.050 716.400 ;
        RECT 919.950 715.950 922.050 716.400 ;
        RECT 1.950 714.600 4.050 715.050 ;
        RECT 61.950 714.600 64.050 715.050 ;
        RECT 1.950 713.400 64.050 714.600 ;
        RECT 1.950 712.950 4.050 713.400 ;
        RECT 61.950 712.950 64.050 713.400 ;
        RECT 76.950 714.600 79.050 715.050 ;
        RECT 85.950 714.600 88.050 715.050 ;
        RECT 76.950 713.400 88.050 714.600 ;
        RECT 76.950 712.950 79.050 713.400 ;
        RECT 85.950 712.950 88.050 713.400 ;
        RECT 163.950 714.600 166.050 715.050 ;
        RECT 172.950 714.600 175.050 715.050 ;
        RECT 163.950 713.400 175.050 714.600 ;
        RECT 163.950 712.950 166.050 713.400 ;
        RECT 172.950 712.950 175.050 713.400 ;
        RECT 187.950 714.600 190.050 715.050 ;
        RECT 226.800 714.600 228.900 715.050 ;
        RECT 187.950 713.400 228.900 714.600 ;
        RECT 187.950 712.950 190.050 713.400 ;
        RECT 226.800 712.950 228.900 713.400 ;
        RECT 229.950 714.600 232.050 715.050 ;
        RECT 313.950 714.600 316.050 715.050 ;
        RECT 229.950 713.400 316.050 714.600 ;
        RECT 229.950 712.950 232.050 713.400 ;
        RECT 313.950 712.950 316.050 713.400 ;
        RECT 328.950 714.600 331.050 714.900 ;
        RECT 349.950 714.600 352.050 715.050 ;
        RECT 328.950 713.400 352.050 714.600 ;
        RECT 328.950 712.800 331.050 713.400 ;
        RECT 349.950 712.950 352.050 713.400 ;
        RECT 391.950 714.600 394.050 715.050 ;
        RECT 401.400 714.600 402.600 715.950 ;
        RECT 391.950 713.400 402.600 714.600 ;
        RECT 409.950 714.600 412.050 715.050 ;
        RECT 529.950 714.600 532.050 715.050 ;
        RECT 409.950 713.400 532.050 714.600 ;
        RECT 391.950 712.950 394.050 713.400 ;
        RECT 409.950 712.950 412.050 713.400 ;
        RECT 529.950 712.950 532.050 713.400 ;
        RECT 541.950 714.600 544.050 715.050 ;
        RECT 559.950 714.600 562.050 715.050 ;
        RECT 541.950 713.400 562.050 714.600 ;
        RECT 541.950 712.950 544.050 713.400 ;
        RECT 559.950 712.950 562.050 713.400 ;
        RECT 820.950 714.600 823.050 715.050 ;
        RECT 871.950 714.600 874.050 715.050 ;
        RECT 820.950 713.400 874.050 714.600 ;
        RECT 820.950 712.950 823.050 713.400 ;
        RECT 871.950 712.950 874.050 713.400 ;
        RECT 250.950 711.600 253.050 712.050 ;
        RECT 259.950 711.600 262.050 712.050 ;
        RECT 250.950 710.400 262.050 711.600 ;
        RECT 250.950 709.950 253.050 710.400 ;
        RECT 259.950 709.950 262.050 710.400 ;
        RECT 286.950 711.600 289.050 712.050 ;
        RECT 316.950 711.600 319.050 712.050 ;
        RECT 286.950 710.400 319.050 711.600 ;
        RECT 286.950 709.950 289.050 710.400 ;
        RECT 316.950 709.950 319.050 710.400 ;
        RECT 430.950 711.600 433.050 712.050 ;
        RECT 496.800 711.600 498.900 712.050 ;
        RECT 430.950 710.400 498.900 711.600 ;
        RECT 430.950 709.950 433.050 710.400 ;
        RECT 496.800 709.950 498.900 710.400 ;
        RECT 535.950 711.600 538.050 712.050 ;
        RECT 568.950 711.600 571.050 712.050 ;
        RECT 535.950 710.400 571.050 711.600 ;
        RECT 535.950 709.950 538.050 710.400 ;
        RECT 568.950 709.950 571.050 710.400 ;
        RECT 634.950 711.600 637.050 712.050 ;
        RECT 670.950 711.600 673.050 712.050 ;
        RECT 634.950 710.400 673.050 711.600 ;
        RECT 634.950 709.950 637.050 710.400 ;
        RECT 670.950 709.950 673.050 710.400 ;
        RECT 688.950 711.600 691.050 712.050 ;
        RECT 817.950 711.600 820.050 712.050 ;
        RECT 688.950 710.400 820.050 711.600 ;
        RECT 688.950 709.950 691.050 710.400 ;
        RECT 817.950 709.950 820.050 710.400 ;
        RECT 823.950 711.600 826.050 712.050 ;
        RECT 838.950 711.600 841.050 712.050 ;
        RECT 823.950 710.400 841.050 711.600 ;
        RECT 823.950 709.950 826.050 710.400 ;
        RECT 838.950 709.950 841.050 710.400 ;
        RECT 7.950 708.600 10.050 709.050 ;
        RECT 52.950 708.600 55.050 709.050 ;
        RECT 7.950 707.400 55.050 708.600 ;
        RECT 7.950 706.950 10.050 707.400 ;
        RECT 52.950 706.950 55.050 707.400 ;
        RECT 85.950 708.600 88.050 709.050 ;
        RECT 97.950 708.600 100.050 709.050 ;
        RECT 85.950 707.400 100.050 708.600 ;
        RECT 85.950 706.950 88.050 707.400 ;
        RECT 97.950 706.950 100.050 707.400 ;
        RECT 133.950 708.600 136.050 709.050 ;
        RECT 178.950 708.600 181.050 709.050 ;
        RECT 133.950 707.400 181.050 708.600 ;
        RECT 133.950 706.950 136.050 707.400 ;
        RECT 178.950 706.950 181.050 707.400 ;
        RECT 199.950 708.600 202.050 709.050 ;
        RECT 400.950 708.600 403.050 709.050 ;
        RECT 199.950 707.400 403.050 708.600 ;
        RECT 199.950 706.950 202.050 707.400 ;
        RECT 400.950 706.950 403.050 707.400 ;
        RECT 418.950 708.600 421.050 709.050 ;
        RECT 424.950 708.600 427.050 709.050 ;
        RECT 418.950 707.400 427.050 708.600 ;
        RECT 418.950 706.950 421.050 707.400 ;
        RECT 424.950 706.950 427.050 707.400 ;
        RECT 442.950 708.600 445.050 709.050 ;
        RECT 457.950 708.600 460.050 709.050 ;
        RECT 442.950 707.400 460.050 708.600 ;
        RECT 442.950 706.950 445.050 707.400 ;
        RECT 457.950 706.950 460.050 707.400 ;
        RECT 478.950 708.600 481.050 709.050 ;
        RECT 595.950 708.600 598.050 709.050 ;
        RECT 478.950 707.400 598.050 708.600 ;
        RECT 478.950 706.950 481.050 707.400 ;
        RECT 595.950 706.950 598.050 707.400 ;
        RECT 775.950 708.600 778.050 709.050 ;
        RECT 784.950 708.600 787.050 709.050 ;
        RECT 775.950 707.400 787.050 708.600 ;
        RECT 775.950 706.950 778.050 707.400 ;
        RECT 784.950 706.950 787.050 707.400 ;
        RECT 109.950 705.600 112.050 706.050 ;
        RECT 124.950 705.600 127.050 706.050 ;
        RECT 109.950 704.400 127.050 705.600 ;
        RECT 109.950 703.950 112.050 704.400 ;
        RECT 124.950 703.950 127.050 704.400 ;
        RECT 184.950 705.600 187.050 706.050 ;
        RECT 235.950 705.600 238.050 706.050 ;
        RECT 184.950 704.400 238.050 705.600 ;
        RECT 184.950 703.950 187.050 704.400 ;
        RECT 235.950 703.950 238.050 704.400 ;
        RECT 403.950 705.600 406.050 706.050 ;
        RECT 424.950 705.600 427.050 705.900 ;
        RECT 442.950 705.600 445.050 705.900 ;
        RECT 487.950 705.600 490.050 706.050 ;
        RECT 403.950 704.400 490.050 705.600 ;
        RECT 403.950 703.950 406.050 704.400 ;
        RECT 424.950 703.800 427.050 704.400 ;
        RECT 442.950 703.800 445.050 704.400 ;
        RECT 487.950 703.950 490.050 704.400 ;
        RECT 613.950 705.600 616.050 706.050 ;
        RECT 634.950 705.600 637.050 706.050 ;
        RECT 679.950 705.600 682.050 706.050 ;
        RECT 613.950 704.400 682.050 705.600 ;
        RECT 613.950 703.950 616.050 704.400 ;
        RECT 634.950 703.950 637.050 704.400 ;
        RECT 679.950 703.950 682.050 704.400 ;
        RECT 799.950 705.600 802.050 706.050 ;
        RECT 820.950 705.600 823.050 706.050 ;
        RECT 799.950 704.400 823.050 705.600 ;
        RECT 799.950 703.950 802.050 704.400 ;
        RECT 820.950 703.950 823.050 704.400 ;
        RECT 847.950 705.600 850.050 706.050 ;
        RECT 877.950 705.600 880.050 706.050 ;
        RECT 847.950 704.400 880.050 705.600 ;
        RECT 847.950 703.950 850.050 704.400 ;
        RECT 877.950 703.950 880.050 704.400 ;
        RECT 907.950 705.600 910.050 706.050 ;
        RECT 928.950 705.600 931.050 706.050 ;
        RECT 907.950 704.400 931.050 705.600 ;
        RECT 907.950 703.950 910.050 704.400 ;
        RECT 928.950 703.950 931.050 704.400 ;
        RECT 73.950 702.600 76.050 703.050 ;
        RECT 103.950 702.600 106.050 703.050 ;
        RECT 73.950 701.400 106.050 702.600 ;
        RECT 73.950 700.950 76.050 701.400 ;
        RECT 103.950 700.950 106.050 701.400 ;
        RECT 118.950 702.600 121.050 703.050 ;
        RECT 145.950 702.600 148.050 703.050 ;
        RECT 118.950 701.400 148.050 702.600 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 145.950 700.950 148.050 701.400 ;
        RECT 175.950 702.600 178.050 703.050 ;
        RECT 277.950 702.600 280.050 703.050 ;
        RECT 289.950 702.600 292.050 703.050 ;
        RECT 304.950 702.600 307.050 703.050 ;
        RECT 175.950 701.400 307.050 702.600 ;
        RECT 175.950 700.950 178.050 701.400 ;
        RECT 277.950 700.950 280.050 701.400 ;
        RECT 289.950 700.950 292.050 701.400 ;
        RECT 304.950 700.950 307.050 701.400 ;
        RECT 313.950 702.600 316.050 703.050 ;
        RECT 400.950 702.600 403.050 703.050 ;
        RECT 313.950 701.400 403.050 702.600 ;
        RECT 313.950 700.950 316.050 701.400 ;
        RECT 400.950 700.950 403.050 701.400 ;
        RECT 445.950 702.600 448.050 703.050 ;
        RECT 523.950 702.600 526.050 703.050 ;
        RECT 445.950 701.400 526.050 702.600 ;
        RECT 445.950 700.950 448.050 701.400 ;
        RECT 523.950 700.950 526.050 701.400 ;
        RECT 529.950 702.600 532.050 703.050 ;
        RECT 580.950 702.600 583.050 702.900 ;
        RECT 529.950 701.400 583.050 702.600 ;
        RECT 529.950 700.950 532.050 701.400 ;
        RECT 580.950 700.800 583.050 701.400 ;
        RECT 712.950 702.600 715.050 703.050 ;
        RECT 724.950 702.600 727.050 703.050 ;
        RECT 712.950 701.400 727.050 702.600 ;
        RECT 712.950 700.950 715.050 701.400 ;
        RECT 724.950 700.950 727.050 701.400 ;
        RECT 892.950 702.600 895.050 703.050 ;
        RECT 925.950 702.600 928.050 703.050 ;
        RECT 892.950 701.400 928.050 702.600 ;
        RECT 892.950 700.950 895.050 701.400 ;
        RECT 925.950 700.950 928.050 701.400 ;
        RECT 178.950 699.600 181.050 700.050 ;
        RECT 187.950 699.600 190.050 700.050 ;
        RECT 178.950 698.400 190.050 699.600 ;
        RECT 178.950 697.950 181.050 698.400 ;
        RECT 187.950 697.950 190.050 698.400 ;
        RECT 196.950 699.600 199.050 700.050 ;
        RECT 262.950 699.600 265.050 700.050 ;
        RECT 598.950 699.600 601.050 700.050 ;
        RECT 196.950 698.400 265.050 699.600 ;
        RECT 196.950 697.950 199.050 698.400 ;
        RECT 262.950 697.950 265.050 698.400 ;
        RECT 443.400 698.400 601.050 699.600 ;
        RECT 136.950 696.600 139.050 697.050 ;
        RECT 142.950 696.600 145.050 697.050 ;
        RECT 148.950 696.600 151.050 697.050 ;
        RECT 187.950 696.600 190.050 696.900 ;
        RECT 136.950 695.400 190.050 696.600 ;
        RECT 136.950 694.950 139.050 695.400 ;
        RECT 142.950 694.950 145.050 695.400 ;
        RECT 148.950 694.950 151.050 695.400 ;
        RECT 187.950 694.800 190.050 695.400 ;
        RECT 358.950 696.600 361.050 697.050 ;
        RECT 373.950 696.600 376.050 697.050 ;
        RECT 443.400 696.600 444.600 698.400 ;
        RECT 598.950 697.950 601.050 698.400 ;
        RECT 769.950 699.600 772.050 700.050 ;
        RECT 781.950 699.600 784.050 700.050 ;
        RECT 799.950 699.600 802.050 700.050 ;
        RECT 769.950 698.400 802.050 699.600 ;
        RECT 769.950 697.950 772.050 698.400 ;
        RECT 781.950 697.950 784.050 698.400 ;
        RECT 799.950 697.950 802.050 698.400 ;
        RECT 358.950 695.400 444.600 696.600 ;
        RECT 607.950 696.600 610.050 697.050 ;
        RECT 625.950 696.600 628.050 697.050 ;
        RECT 607.950 695.400 628.050 696.600 ;
        RECT 358.950 694.950 361.050 695.400 ;
        RECT 373.950 694.950 376.050 695.400 ;
        RECT 607.950 694.950 610.050 695.400 ;
        RECT 625.950 694.950 628.050 695.400 ;
        RECT 655.950 696.600 658.050 697.050 ;
        RECT 697.950 696.600 700.050 697.050 ;
        RECT 655.950 695.400 700.050 696.600 ;
        RECT 655.950 694.950 658.050 695.400 ;
        RECT 697.950 694.950 700.050 695.400 ;
        RECT 196.950 693.600 199.050 693.900 ;
        RECT 229.950 693.600 232.050 694.050 ;
        RECT 241.950 693.600 244.050 694.050 ;
        RECT 196.950 692.400 244.050 693.600 ;
        RECT 196.950 691.800 199.050 692.400 ;
        RECT 229.950 691.950 232.050 692.400 ;
        RECT 241.950 691.950 244.050 692.400 ;
        RECT 382.950 693.600 385.050 694.050 ;
        RECT 409.950 693.600 412.050 694.050 ;
        RECT 382.950 692.400 412.050 693.600 ;
        RECT 382.950 691.950 385.050 692.400 ;
        RECT 409.950 691.950 412.050 692.400 ;
        RECT 418.950 693.600 421.050 693.900 ;
        RECT 424.950 693.600 427.050 694.050 ;
        RECT 418.950 692.400 427.050 693.600 ;
        RECT 418.950 691.800 421.050 692.400 ;
        RECT 424.950 691.950 427.050 692.400 ;
        RECT 775.950 693.600 778.050 694.050 ;
        RECT 793.950 693.600 796.050 694.050 ;
        RECT 775.950 692.400 796.050 693.600 ;
        RECT 775.950 691.950 778.050 692.400 ;
        RECT 793.950 691.950 796.050 692.400 ;
        RECT 877.950 693.600 880.050 694.050 ;
        RECT 907.950 693.600 910.050 694.050 ;
        RECT 877.950 692.400 910.050 693.600 ;
        RECT 877.950 691.950 880.050 692.400 ;
        RECT 907.950 691.950 910.050 692.400 ;
        RECT 13.950 690.600 16.050 691.050 ;
        RECT 22.950 690.600 25.050 691.050 ;
        RECT 13.950 689.400 25.050 690.600 ;
        RECT 13.950 688.950 16.050 689.400 ;
        RECT 22.950 688.950 25.050 689.400 ;
        RECT 127.950 690.600 130.050 691.050 ;
        RECT 178.950 690.600 181.050 691.050 ;
        RECT 190.950 690.600 193.050 691.050 ;
        RECT 217.950 690.600 220.050 691.050 ;
        RECT 127.950 689.400 193.050 690.600 ;
        RECT 127.950 688.950 130.050 689.400 ;
        RECT 178.950 688.950 181.050 689.400 ;
        RECT 190.950 688.950 193.050 689.400 ;
        RECT 209.400 689.400 220.050 690.600 ;
        RECT 94.950 687.600 97.050 688.050 ;
        RECT 118.950 687.600 121.050 688.050 ;
        RECT 94.950 686.400 121.050 687.600 ;
        RECT 94.950 685.950 97.050 686.400 ;
        RECT 118.950 685.950 121.050 686.400 ;
        RECT 145.950 687.600 148.050 688.050 ;
        RECT 154.950 687.600 157.050 688.050 ;
        RECT 209.400 687.600 210.600 689.400 ;
        RECT 217.950 688.950 220.050 689.400 ;
        RECT 244.950 690.600 247.050 691.050 ;
        RECT 265.950 690.600 268.050 691.050 ;
        RECT 244.950 689.400 268.050 690.600 ;
        RECT 244.950 688.950 247.050 689.400 ;
        RECT 265.950 688.950 268.050 689.400 ;
        RECT 292.950 690.600 295.050 691.050 ;
        RECT 307.950 690.600 310.050 691.050 ;
        RECT 292.950 689.400 310.050 690.600 ;
        RECT 292.950 688.950 295.050 689.400 ;
        RECT 307.950 688.950 310.050 689.400 ;
        RECT 400.950 690.600 403.050 691.050 ;
        RECT 427.950 690.600 430.050 691.050 ;
        RECT 400.950 689.400 430.050 690.600 ;
        RECT 400.950 688.950 403.050 689.400 ;
        RECT 427.950 688.950 430.050 689.400 ;
        RECT 742.950 690.600 745.050 691.050 ;
        RECT 769.950 690.600 772.050 691.050 ;
        RECT 742.950 689.400 772.050 690.600 ;
        RECT 742.950 688.950 745.050 689.400 ;
        RECT 769.950 688.950 772.050 689.400 ;
        RECT 832.950 690.600 835.050 691.050 ;
        RECT 844.950 690.600 847.050 691.050 ;
        RECT 832.950 689.400 847.050 690.600 ;
        RECT 832.950 688.950 835.050 689.400 ;
        RECT 844.950 688.950 847.050 689.400 ;
        RECT 145.950 686.400 157.050 687.600 ;
        RECT 145.950 685.950 148.050 686.400 ;
        RECT 154.950 685.950 157.050 686.400 ;
        RECT 206.400 686.400 210.600 687.600 ;
        RECT 304.950 687.600 307.050 688.050 ;
        RECT 454.950 687.600 457.050 688.050 ;
        RECT 304.950 686.400 333.600 687.600 ;
        RECT 206.400 685.200 207.600 686.400 ;
        RECT 304.950 685.950 307.050 686.400 ;
        RECT 82.950 683.100 85.050 685.200 ;
        RECT 83.400 679.050 84.600 683.100 ;
        RECT 103.950 682.950 106.050 685.050 ;
        RECT 126.000 684.600 130.050 685.050 ;
        RECT 125.400 682.950 130.050 684.600 ;
        RECT 133.950 684.600 136.050 685.050 ;
        RECT 139.950 684.600 142.050 685.200 ;
        RECT 133.950 683.400 142.050 684.600 ;
        RECT 133.950 682.950 136.050 683.400 ;
        RECT 139.950 683.100 142.050 683.400 ;
        RECT 163.950 684.750 166.050 685.200 ;
        RECT 169.950 684.750 172.050 685.200 ;
        RECT 163.950 683.550 172.050 684.750 ;
        RECT 163.950 683.100 166.050 683.550 ;
        RECT 169.950 683.100 172.050 683.550 ;
        RECT 199.950 683.100 202.050 685.200 ;
        RECT 205.950 683.100 208.050 685.200 ;
        RECT 211.950 684.750 214.050 685.200 ;
        RECT 217.950 684.750 220.050 685.200 ;
        RECT 211.950 683.550 220.050 684.750 ;
        RECT 211.950 683.100 214.050 683.550 ;
        RECT 217.950 683.100 220.050 683.550 ;
        RECT 226.950 683.100 229.050 685.200 ;
        RECT 241.950 684.750 244.050 685.200 ;
        RECT 250.950 684.750 253.050 685.200 ;
        RECT 241.950 683.550 253.050 684.750 ;
        RECT 241.950 683.100 244.050 683.550 ;
        RECT 250.950 683.100 253.050 683.550 ;
        RECT 262.950 684.600 265.050 685.050 ;
        RECT 274.950 684.600 277.050 685.050 ;
        RECT 262.950 683.400 277.050 684.600 ;
        RECT 332.400 684.600 333.600 686.400 ;
        RECT 434.400 686.400 457.050 687.600 ;
        RECT 358.950 684.600 361.050 685.050 ;
        RECT 332.400 683.400 361.050 684.600 ;
        RECT 16.950 678.600 19.050 678.900 ;
        RECT 22.950 678.600 25.050 679.050 ;
        RECT 28.950 678.600 31.050 679.050 ;
        RECT 16.950 677.400 31.050 678.600 ;
        RECT 16.950 676.800 19.050 677.400 ;
        RECT 22.950 676.950 25.050 677.400 ;
        RECT 28.950 676.950 31.050 677.400 ;
        RECT 34.950 678.600 37.050 678.900 ;
        RECT 49.950 678.600 52.050 678.900 ;
        RECT 64.950 678.600 67.050 679.050 ;
        RECT 34.950 677.400 67.050 678.600 ;
        RECT 83.400 677.400 88.050 679.050 ;
        RECT 34.950 676.800 37.050 677.400 ;
        RECT 49.950 676.800 52.050 677.400 ;
        RECT 64.950 676.950 67.050 677.400 ;
        RECT 84.000 676.950 88.050 677.400 ;
        RECT 97.950 678.600 100.050 678.900 ;
        RECT 104.400 678.600 105.600 682.950 ;
        RECT 125.400 678.900 126.600 682.950 ;
        RECT 97.950 677.400 105.600 678.600 ;
        RECT 97.950 676.800 100.050 677.400 ;
        RECT 124.950 676.800 127.050 678.900 ;
        RECT 166.950 678.600 169.050 679.050 ;
        RECT 200.400 678.600 201.600 683.100 ;
        RECT 227.400 681.600 228.600 683.100 ;
        RECT 262.950 682.950 265.050 683.400 ;
        RECT 274.950 682.950 277.050 683.400 ;
        RECT 358.950 682.950 361.050 683.400 ;
        RECT 409.950 683.100 412.050 685.200 ;
        RECT 415.950 684.600 418.050 685.050 ;
        RECT 434.400 684.600 435.600 686.400 ;
        RECT 454.950 685.950 457.050 686.400 ;
        RECT 613.950 687.600 616.050 688.050 ;
        RECT 625.950 687.600 628.050 688.050 ;
        RECT 613.950 686.400 628.050 687.600 ;
        RECT 613.950 685.950 616.050 686.400 ;
        RECT 625.950 685.950 628.050 686.400 ;
        RECT 679.950 687.600 682.050 688.200 ;
        RECT 688.950 687.600 691.050 688.200 ;
        RECT 679.950 686.400 691.050 687.600 ;
        RECT 679.950 686.100 682.050 686.400 ;
        RECT 688.950 686.100 691.050 686.400 ;
        RECT 760.950 687.600 763.050 688.050 ;
        RECT 775.950 687.600 778.050 688.050 ;
        RECT 760.950 686.400 778.050 687.600 ;
        RECT 760.950 685.950 763.050 686.400 ;
        RECT 775.950 685.950 778.050 686.400 ;
        RECT 886.950 687.600 889.050 688.050 ;
        RECT 901.950 687.600 904.050 688.050 ;
        RECT 886.950 686.400 904.050 687.600 ;
        RECT 886.950 685.950 889.050 686.400 ;
        RECT 901.950 685.950 904.050 686.400 ;
        RECT 457.950 684.600 460.050 685.050 ;
        RECT 415.950 683.400 435.600 684.600 ;
        RECT 437.400 684.000 460.050 684.600 ;
        RECT 436.950 683.400 460.050 684.000 ;
        RECT 280.950 681.600 283.050 681.900 ;
        RECT 328.950 681.600 331.050 682.050 ;
        RECT 227.400 680.400 234.600 681.600 ;
        RECT 166.950 677.400 201.600 678.600 ;
        RECT 220.950 678.600 223.050 679.050 ;
        RECT 229.950 678.600 232.050 678.900 ;
        RECT 220.950 677.400 232.050 678.600 ;
        RECT 166.950 676.950 169.050 677.400 ;
        RECT 220.950 676.950 223.050 677.400 ;
        RECT 229.950 676.800 232.050 677.400 ;
        RECT 4.950 675.600 7.050 676.050 ;
        RECT 10.950 675.600 13.050 676.050 ;
        RECT 4.950 674.400 13.050 675.600 ;
        RECT 4.950 673.950 7.050 674.400 ;
        RECT 10.950 673.950 13.050 674.400 ;
        RECT 169.950 675.600 172.050 676.050 ;
        RECT 178.950 675.600 181.050 676.050 ;
        RECT 169.950 674.400 181.050 675.600 ;
        RECT 233.400 675.600 234.600 680.400 ;
        RECT 280.950 680.400 331.050 681.600 ;
        RECT 280.950 679.800 283.050 680.400 ;
        RECT 328.950 679.950 331.050 680.400 ;
        RECT 268.950 678.450 271.050 678.900 ;
        RECT 277.950 678.450 280.050 679.050 ;
        RECT 268.950 677.250 280.050 678.450 ;
        RECT 268.950 676.800 271.050 677.250 ;
        RECT 277.950 676.950 280.050 677.250 ;
        RECT 304.950 678.450 307.050 678.900 ;
        RECT 310.950 678.450 313.050 678.900 ;
        RECT 304.950 677.250 313.050 678.450 ;
        RECT 304.950 676.800 307.050 677.250 ;
        RECT 310.950 676.800 313.050 677.250 ;
        RECT 316.950 678.600 319.050 678.900 ;
        RECT 400.950 678.600 403.050 678.900 ;
        RECT 316.950 677.400 403.050 678.600 ;
        RECT 410.400 678.600 411.600 683.100 ;
        RECT 415.950 682.950 418.050 683.400 ;
        RECT 436.950 679.950 439.050 683.400 ;
        RECT 457.950 682.950 460.050 683.400 ;
        RECT 499.950 684.600 502.050 685.050 ;
        RECT 514.950 684.600 517.050 685.200 ;
        RECT 499.950 683.400 517.050 684.600 ;
        RECT 499.950 682.950 502.050 683.400 ;
        RECT 514.950 683.100 517.050 683.400 ;
        RECT 538.950 684.600 541.050 685.050 ;
        RECT 553.950 684.600 556.050 685.200 ;
        RECT 538.950 683.400 556.050 684.600 ;
        RECT 538.950 682.950 541.050 683.400 ;
        RECT 553.950 683.100 556.050 683.400 ;
        RECT 589.950 684.750 592.050 685.200 ;
        RECT 595.800 684.750 597.900 685.200 ;
        RECT 589.950 683.550 597.900 684.750 ;
        RECT 589.950 683.100 592.050 683.550 ;
        RECT 595.800 683.100 597.900 683.550 ;
        RECT 598.950 684.600 601.050 685.050 ;
        RECT 655.950 684.600 658.050 685.050 ;
        RECT 598.950 683.400 658.050 684.600 ;
        RECT 598.950 682.950 601.050 683.400 ;
        RECT 655.950 682.950 658.050 683.400 ;
        RECT 763.950 682.950 766.050 685.050 ;
        RECT 811.950 684.600 814.050 685.200 ;
        RECT 797.400 683.400 814.050 684.600 ;
        RECT 682.950 681.600 685.050 682.050 ;
        RECT 590.400 680.400 685.050 681.600 ;
        RECT 424.950 678.600 427.050 678.900 ;
        RECT 410.400 677.400 427.050 678.600 ;
        RECT 316.950 676.800 319.050 677.400 ;
        RECT 400.950 676.800 403.050 677.400 ;
        RECT 424.950 676.800 427.050 677.400 ;
        RECT 508.950 678.600 511.050 679.050 ;
        RECT 565.950 678.600 568.050 679.050 ;
        RECT 508.950 677.400 568.050 678.600 ;
        RECT 508.950 676.950 511.050 677.400 ;
        RECT 565.950 676.950 568.050 677.400 ;
        RECT 580.950 678.450 583.050 678.900 ;
        RECT 586.950 678.450 589.050 678.900 ;
        RECT 580.950 677.250 589.050 678.450 ;
        RECT 580.950 676.800 583.050 677.250 ;
        RECT 586.950 676.800 589.050 677.250 ;
        RECT 244.950 675.600 247.050 676.050 ;
        RECT 233.400 674.400 247.050 675.600 ;
        RECT 169.950 673.950 172.050 674.400 ;
        RECT 178.950 673.950 181.050 674.400 ;
        RECT 244.950 673.950 247.050 674.400 ;
        RECT 250.950 675.600 253.050 676.050 ;
        RECT 259.950 675.600 262.050 676.050 ;
        RECT 250.950 674.400 262.050 675.600 ;
        RECT 250.950 673.950 253.050 674.400 ;
        RECT 259.950 673.950 262.050 674.400 ;
        RECT 271.950 675.600 274.050 676.050 ;
        RECT 280.950 675.600 283.050 676.050 ;
        RECT 271.950 674.400 283.050 675.600 ;
        RECT 271.950 673.950 274.050 674.400 ;
        RECT 280.950 673.950 283.050 674.400 ;
        RECT 484.950 675.600 487.050 676.050 ;
        RECT 511.950 675.600 514.050 676.050 ;
        RECT 538.950 675.600 541.050 676.050 ;
        RECT 484.950 674.400 541.050 675.600 ;
        RECT 484.950 673.950 487.050 674.400 ;
        RECT 511.950 673.950 514.050 674.400 ;
        RECT 538.950 673.950 541.050 674.400 ;
        RECT 568.950 675.600 571.050 676.050 ;
        RECT 590.400 675.600 591.600 680.400 ;
        RECT 682.950 679.950 685.050 680.400 ;
        RECT 748.950 681.450 751.050 681.900 ;
        RECT 754.950 681.450 757.050 681.900 ;
        RECT 748.950 680.250 757.050 681.450 ;
        RECT 748.950 679.800 751.050 680.250 ;
        RECT 754.950 679.800 757.050 680.250 ;
        RECT 595.950 678.600 598.050 679.050 ;
        RECT 604.950 678.600 607.050 678.900 ;
        RECT 595.950 677.400 607.050 678.600 ;
        RECT 764.400 678.600 765.600 682.950 ;
        RECT 797.400 678.900 798.600 683.400 ;
        RECT 811.950 683.100 814.050 683.400 ;
        RECT 838.950 683.100 841.050 685.200 ;
        RECT 853.950 684.600 856.050 685.200 ;
        RECT 865.950 684.750 868.050 685.200 ;
        RECT 871.950 684.750 874.050 685.200 ;
        RECT 853.950 683.400 858.600 684.600 ;
        RECT 853.950 683.100 856.050 683.400 ;
        RECT 766.950 678.600 769.050 678.900 ;
        RECT 764.400 677.400 769.050 678.600 ;
        RECT 595.950 676.950 598.050 677.400 ;
        RECT 604.950 676.800 607.050 677.400 ;
        RECT 766.950 676.800 769.050 677.400 ;
        RECT 772.950 678.450 775.050 678.900 ;
        RECT 778.950 678.450 781.050 678.900 ;
        RECT 772.950 677.250 781.050 678.450 ;
        RECT 772.950 676.800 775.050 677.250 ;
        RECT 778.950 676.800 781.050 677.250 ;
        RECT 796.950 676.800 799.050 678.900 ;
        RECT 814.950 678.600 817.050 678.900 ;
        RECT 817.950 678.600 820.050 679.050 ;
        RECT 835.950 678.600 838.050 678.900 ;
        RECT 814.950 677.400 838.050 678.600 ;
        RECT 839.400 678.600 840.600 683.100 ;
        RECT 857.400 681.600 858.600 683.400 ;
        RECT 865.950 683.550 874.050 684.750 ;
        RECT 865.950 683.100 868.050 683.550 ;
        RECT 871.950 683.100 874.050 683.550 ;
        RECT 895.950 684.600 898.050 685.200 ;
        RECT 913.950 684.600 916.050 685.200 ;
        RECT 895.950 683.400 916.050 684.600 ;
        RECT 895.950 683.100 898.050 683.400 ;
        RECT 913.950 683.100 916.050 683.400 ;
        RECT 925.950 684.600 928.050 685.200 ;
        RECT 931.950 684.750 934.050 685.200 ;
        RECT 937.950 684.750 940.050 685.200 ;
        RECT 931.950 684.600 940.050 684.750 ;
        RECT 925.950 683.550 940.050 684.600 ;
        RECT 925.950 683.400 934.050 683.550 ;
        RECT 925.950 683.100 928.050 683.400 ;
        RECT 931.950 683.100 934.050 683.400 ;
        RECT 937.950 683.100 940.050 683.550 ;
        RECT 943.800 683.100 945.900 685.200 ;
        RECT 889.950 681.600 892.050 682.050 ;
        RECT 857.400 680.400 892.050 681.600 ;
        RECT 889.950 679.950 892.050 680.400 ;
        RECT 856.950 678.600 859.050 678.900 ;
        RECT 839.400 677.400 859.050 678.600 ;
        RECT 814.950 676.800 817.050 677.400 ;
        RECT 817.950 676.950 820.050 677.400 ;
        RECT 835.950 676.800 838.050 677.400 ;
        RECT 856.950 676.800 859.050 677.400 ;
        RECT 568.950 674.400 591.600 675.600 ;
        RECT 628.950 675.600 631.050 676.050 ;
        RECT 670.950 675.600 673.050 676.050 ;
        RECT 739.950 675.600 742.050 676.050 ;
        RECT 628.950 674.400 742.050 675.600 ;
        RECT 568.950 673.950 571.050 674.400 ;
        RECT 628.950 673.950 631.050 674.400 ;
        RECT 670.950 673.950 673.050 674.400 ;
        RECT 739.950 673.950 742.050 674.400 ;
        RECT 784.950 675.600 787.050 676.050 ;
        RECT 790.950 675.600 793.050 676.050 ;
        RECT 784.950 674.400 793.050 675.600 ;
        RECT 784.950 673.950 787.050 674.400 ;
        RECT 790.950 673.950 793.050 674.400 ;
        RECT 847.950 675.600 850.050 676.050 ;
        RECT 853.950 675.600 856.050 676.050 ;
        RECT 847.950 674.400 856.050 675.600 ;
        RECT 847.950 673.950 850.050 674.400 ;
        RECT 853.950 673.950 856.050 674.400 ;
        RECT 880.950 675.600 883.050 676.050 ;
        RECT 896.400 675.600 897.600 683.100 ;
        RECT 944.400 681.600 945.600 683.100 ;
        RECT 946.950 682.950 949.050 685.050 ;
        RECT 938.400 680.400 945.600 681.600 ;
        RECT 898.950 678.600 901.050 678.900 ;
        RECT 907.950 678.600 910.050 679.050 ;
        RECT 898.950 677.400 910.050 678.600 ;
        RECT 898.950 676.800 901.050 677.400 ;
        RECT 907.950 676.950 910.050 677.400 ;
        RECT 922.950 678.600 925.050 678.900 ;
        RECT 938.400 678.600 939.600 680.400 ;
        RECT 922.950 677.400 939.600 678.600 ;
        RECT 940.950 678.600 943.050 678.900 ;
        RECT 947.400 678.600 948.600 682.950 ;
        RECT 940.950 677.400 948.600 678.600 ;
        RECT 922.950 676.800 925.050 677.400 ;
        RECT 940.950 676.800 943.050 677.400 ;
        RECT 880.950 674.400 897.600 675.600 ;
        RECT 880.950 673.950 883.050 674.400 ;
        RECT 55.950 672.600 58.050 673.050 ;
        RECT 91.950 672.600 94.050 673.050 ;
        RECT 55.950 671.400 94.050 672.600 ;
        RECT 55.950 670.950 58.050 671.400 ;
        RECT 91.950 670.950 94.050 671.400 ;
        RECT 217.950 672.600 220.050 673.050 ;
        RECT 247.950 672.600 250.050 673.050 ;
        RECT 217.950 671.400 250.050 672.600 ;
        RECT 217.950 670.950 220.050 671.400 ;
        RECT 247.950 670.950 250.050 671.400 ;
        RECT 256.950 672.600 259.050 673.050 ;
        RECT 313.950 672.600 316.050 673.050 ;
        RECT 256.950 671.400 316.050 672.600 ;
        RECT 256.950 670.950 259.050 671.400 ;
        RECT 313.950 670.950 316.050 671.400 ;
        RECT 406.950 672.600 409.050 673.050 ;
        RECT 415.950 672.600 418.050 673.050 ;
        RECT 508.950 672.600 511.050 673.050 ;
        RECT 406.950 671.400 418.050 672.600 ;
        RECT 406.950 670.950 409.050 671.400 ;
        RECT 415.950 670.950 418.050 671.400 ;
        RECT 473.400 671.400 511.050 672.600 ;
        RECT 58.950 669.600 61.050 670.050 ;
        RECT 94.950 669.600 97.050 670.050 ;
        RECT 175.950 669.600 178.050 670.050 ;
        RECT 208.950 669.600 211.050 670.050 ;
        RECT 58.950 668.400 97.050 669.600 ;
        RECT 58.950 667.950 61.050 668.400 ;
        RECT 94.950 667.950 97.050 668.400 ;
        RECT 98.400 668.400 144.600 669.600 ;
        RECT 82.950 666.600 85.050 667.050 ;
        RECT 88.950 666.600 91.050 667.050 ;
        RECT 98.400 666.600 99.600 668.400 ;
        RECT 143.400 667.050 144.600 668.400 ;
        RECT 175.950 668.400 211.050 669.600 ;
        RECT 175.950 667.950 178.050 668.400 ;
        RECT 208.950 667.950 211.050 668.400 ;
        RECT 229.950 669.600 232.050 670.050 ;
        RECT 238.950 669.600 241.050 670.050 ;
        RECT 229.950 668.400 241.050 669.600 ;
        RECT 229.950 667.950 232.050 668.400 ;
        RECT 238.950 667.950 241.050 668.400 ;
        RECT 280.950 669.600 283.050 670.050 ;
        RECT 298.950 669.600 301.050 670.050 ;
        RECT 280.950 668.400 301.050 669.600 ;
        RECT 280.950 667.950 283.050 668.400 ;
        RECT 298.950 667.950 301.050 668.400 ;
        RECT 319.950 669.600 322.050 670.050 ;
        RECT 394.950 669.600 397.050 670.050 ;
        RECT 424.950 669.600 427.050 670.050 ;
        RECT 319.950 669.000 372.600 669.600 ;
        RECT 319.950 668.400 373.050 669.000 ;
        RECT 319.950 667.950 322.050 668.400 ;
        RECT 82.950 665.400 99.600 666.600 ;
        RECT 142.950 666.600 145.050 667.050 ;
        RECT 163.950 666.600 166.050 667.050 ;
        RECT 142.950 665.400 166.050 666.600 ;
        RECT 82.950 664.950 85.050 665.400 ;
        RECT 88.950 664.950 91.050 665.400 ;
        RECT 142.950 664.950 145.050 665.400 ;
        RECT 163.950 664.950 166.050 665.400 ;
        RECT 202.950 666.600 205.050 667.050 ;
        RECT 268.950 666.600 271.050 667.050 ;
        RECT 202.950 665.400 271.050 666.600 ;
        RECT 202.950 664.950 205.050 665.400 ;
        RECT 268.950 664.950 271.050 665.400 ;
        RECT 295.950 666.600 298.050 667.050 ;
        RECT 322.950 666.600 325.050 667.050 ;
        RECT 295.950 665.400 325.050 666.600 ;
        RECT 295.950 664.950 298.050 665.400 ;
        RECT 322.950 664.950 325.050 665.400 ;
        RECT 337.950 666.600 340.050 667.050 ;
        RECT 343.950 666.600 346.050 667.050 ;
        RECT 337.950 665.400 346.050 666.600 ;
        RECT 337.950 664.950 340.050 665.400 ;
        RECT 343.950 664.950 346.050 665.400 ;
        RECT 370.950 664.950 373.050 668.400 ;
        RECT 394.950 668.400 427.050 669.600 ;
        RECT 394.950 667.950 397.050 668.400 ;
        RECT 424.950 667.950 427.050 668.400 ;
        RECT 430.950 669.600 433.050 670.050 ;
        RECT 473.400 669.600 474.600 671.400 ;
        RECT 508.950 670.950 511.050 671.400 ;
        RECT 598.950 672.600 601.050 673.050 ;
        RECT 610.800 672.600 612.900 673.050 ;
        RECT 598.950 671.400 612.900 672.600 ;
        RECT 598.950 670.950 601.050 671.400 ;
        RECT 610.800 670.950 612.900 671.400 ;
        RECT 613.950 672.600 616.050 673.050 ;
        RECT 670.950 672.600 673.050 672.900 ;
        RECT 613.950 671.400 673.050 672.600 ;
        RECT 613.950 670.950 616.050 671.400 ;
        RECT 670.950 670.800 673.050 671.400 ;
        RECT 688.950 672.600 691.050 673.050 ;
        RECT 697.950 672.600 700.050 673.050 ;
        RECT 688.950 671.400 700.050 672.600 ;
        RECT 688.950 670.950 691.050 671.400 ;
        RECT 697.950 670.950 700.050 671.400 ;
        RECT 805.950 672.600 808.050 673.050 ;
        RECT 811.950 672.600 814.050 673.050 ;
        RECT 805.950 671.400 814.050 672.600 ;
        RECT 805.950 670.950 808.050 671.400 ;
        RECT 811.950 670.950 814.050 671.400 ;
        RECT 865.950 672.600 868.050 673.050 ;
        RECT 877.950 672.600 880.050 673.050 ;
        RECT 865.950 671.400 880.050 672.600 ;
        RECT 865.950 670.950 868.050 671.400 ;
        RECT 877.950 670.950 880.050 671.400 ;
        RECT 886.950 672.600 889.050 673.050 ;
        RECT 904.950 672.600 907.050 673.050 ;
        RECT 916.950 672.600 919.050 673.050 ;
        RECT 886.950 671.400 919.050 672.600 ;
        RECT 886.950 670.950 889.050 671.400 ;
        RECT 904.950 670.950 907.050 671.400 ;
        RECT 916.950 670.950 919.050 671.400 ;
        RECT 931.950 672.600 934.050 673.050 ;
        RECT 940.950 672.600 943.050 673.050 ;
        RECT 931.950 671.400 943.050 672.600 ;
        RECT 931.950 670.950 934.050 671.400 ;
        RECT 940.950 670.950 943.050 671.400 ;
        RECT 430.950 668.400 474.600 669.600 ;
        RECT 484.950 669.600 487.050 670.050 ;
        RECT 502.950 669.600 505.050 670.050 ;
        RECT 484.950 668.400 505.050 669.600 ;
        RECT 430.950 667.950 433.050 668.400 ;
        RECT 484.950 667.950 487.050 668.400 ;
        RECT 502.950 667.950 505.050 668.400 ;
        RECT 463.950 666.600 466.050 667.050 ;
        RECT 380.400 665.400 466.050 666.600 ;
        RECT 19.950 663.600 22.050 664.050 ;
        RECT 49.950 663.600 52.050 664.050 ;
        RECT 73.950 663.600 76.050 664.050 ;
        RECT 19.950 662.400 42.600 663.600 ;
        RECT 19.950 661.950 22.050 662.400 ;
        RECT 41.400 661.050 42.600 662.400 ;
        RECT 49.950 662.400 76.050 663.600 ;
        RECT 49.950 661.950 52.050 662.400 ;
        RECT 73.950 661.950 76.050 662.400 ;
        RECT 79.950 663.600 82.050 664.050 ;
        RECT 109.950 663.600 112.050 664.050 ;
        RECT 79.950 662.400 112.050 663.600 ;
        RECT 79.950 661.950 82.050 662.400 ;
        RECT 109.950 661.950 112.050 662.400 ;
        RECT 178.950 663.600 181.050 664.050 ;
        RECT 256.950 663.600 259.050 664.050 ;
        RECT 178.950 662.400 259.050 663.600 ;
        RECT 178.950 661.950 181.050 662.400 ;
        RECT 256.950 661.950 259.050 662.400 ;
        RECT 331.950 663.600 334.050 664.050 ;
        RECT 364.950 663.600 367.050 664.050 ;
        RECT 331.950 662.400 367.050 663.600 ;
        RECT 331.950 661.950 334.050 662.400 ;
        RECT 364.950 661.950 367.050 662.400 ;
        RECT 40.950 660.600 43.050 661.050 ;
        RECT 88.950 660.600 91.050 661.050 ;
        RECT 40.950 659.400 91.050 660.600 ;
        RECT 40.950 658.950 43.050 659.400 ;
        RECT 88.950 658.950 91.050 659.400 ;
        RECT 148.950 660.600 151.050 661.050 ;
        RECT 169.950 660.600 172.050 661.050 ;
        RECT 259.950 660.600 262.050 661.050 ;
        RECT 380.400 660.600 381.600 665.400 ;
        RECT 463.950 664.950 466.050 665.400 ;
        RECT 565.950 666.600 568.050 667.050 ;
        RECT 613.950 666.600 616.050 667.050 ;
        RECT 565.950 665.400 616.050 666.600 ;
        RECT 565.950 664.950 568.050 665.400 ;
        RECT 613.950 664.950 616.050 665.400 ;
        RECT 619.950 666.600 622.050 667.050 ;
        RECT 640.950 666.600 643.050 667.050 ;
        RECT 619.950 665.400 643.050 666.600 ;
        RECT 619.950 664.950 622.050 665.400 ;
        RECT 640.950 664.950 643.050 665.400 ;
        RECT 682.950 666.600 685.050 667.050 ;
        RECT 706.950 666.600 709.050 667.050 ;
        RECT 682.950 665.400 709.050 666.600 ;
        RECT 682.950 664.950 685.050 665.400 ;
        RECT 706.950 664.950 709.050 665.400 ;
        RECT 718.950 666.600 721.050 667.050 ;
        RECT 733.950 666.600 736.050 667.050 ;
        RECT 718.950 665.400 736.050 666.600 ;
        RECT 718.950 664.950 721.050 665.400 ;
        RECT 733.950 664.950 736.050 665.400 ;
        RECT 778.950 666.600 781.050 667.050 ;
        RECT 796.950 666.600 799.050 667.050 ;
        RECT 778.950 665.400 799.050 666.600 ;
        RECT 778.950 664.950 781.050 665.400 ;
        RECT 796.950 664.950 799.050 665.400 ;
        RECT 802.950 666.600 805.050 667.050 ;
        RECT 820.950 666.600 823.050 667.050 ;
        RECT 802.950 665.400 823.050 666.600 ;
        RECT 802.950 664.950 805.050 665.400 ;
        RECT 820.950 664.950 823.050 665.400 ;
        RECT 841.950 666.600 844.050 667.050 ;
        RECT 889.950 666.600 892.050 667.050 ;
        RECT 841.950 665.400 892.050 666.600 ;
        RECT 841.950 664.950 844.050 665.400 ;
        RECT 889.950 664.950 892.050 665.400 ;
        RECT 148.950 659.400 165.600 660.600 ;
        RECT 148.950 658.950 151.050 659.400 ;
        RECT 164.400 658.050 165.600 659.400 ;
        RECT 169.950 659.400 381.600 660.600 ;
        RECT 391.950 660.600 394.050 664.050 ;
        RECT 418.950 663.600 421.050 664.050 ;
        RECT 427.950 663.600 430.050 664.050 ;
        RECT 418.950 662.400 430.050 663.600 ;
        RECT 418.950 661.950 421.050 662.400 ;
        RECT 427.950 661.950 430.050 662.400 ;
        RECT 508.950 663.600 511.050 664.050 ;
        RECT 544.950 663.600 547.050 664.050 ;
        RECT 508.950 662.400 547.050 663.600 ;
        RECT 508.950 661.950 511.050 662.400 ;
        RECT 544.950 661.950 547.050 662.400 ;
        RECT 562.950 663.600 565.050 664.050 ;
        RECT 601.950 663.600 604.050 664.050 ;
        RECT 562.950 662.400 604.050 663.600 ;
        RECT 562.950 661.950 565.050 662.400 ;
        RECT 601.950 661.950 604.050 662.400 ;
        RECT 625.950 663.600 628.050 664.050 ;
        RECT 652.950 663.600 655.050 664.050 ;
        RECT 625.950 662.400 655.050 663.600 ;
        RECT 625.950 661.950 628.050 662.400 ;
        RECT 652.950 661.950 655.050 662.400 ;
        RECT 676.950 663.600 679.050 664.050 ;
        RECT 751.950 663.600 754.050 664.050 ;
        RECT 676.950 662.400 754.050 663.600 ;
        RECT 676.950 661.950 679.050 662.400 ;
        RECT 751.950 661.950 754.050 662.400 ;
        RECT 760.950 663.600 763.050 664.050 ;
        RECT 925.950 663.600 928.050 664.050 ;
        RECT 760.950 662.400 928.050 663.600 ;
        RECT 760.950 661.950 763.050 662.400 ;
        RECT 925.950 661.950 928.050 662.400 ;
        RECT 409.950 660.600 412.050 661.050 ;
        RECT 391.950 660.000 412.050 660.600 ;
        RECT 392.400 659.400 412.050 660.000 ;
        RECT 169.950 658.950 172.050 659.400 ;
        RECT 259.950 658.950 262.050 659.400 ;
        RECT 409.950 658.950 412.050 659.400 ;
        RECT 472.950 660.600 475.050 661.050 ;
        RECT 499.950 660.600 502.050 661.050 ;
        RECT 472.950 659.400 502.050 660.600 ;
        RECT 472.950 658.950 475.050 659.400 ;
        RECT 499.950 658.950 502.050 659.400 ;
        RECT 517.950 660.600 520.050 661.050 ;
        RECT 535.950 660.600 538.050 661.050 ;
        RECT 517.950 659.400 538.050 660.600 ;
        RECT 517.950 658.950 520.050 659.400 ;
        RECT 535.950 658.950 538.050 659.400 ;
        RECT 61.950 657.600 64.050 658.050 ;
        RECT 67.950 657.600 70.050 658.050 ;
        RECT 61.950 656.400 70.050 657.600 ;
        RECT 61.950 655.950 64.050 656.400 ;
        RECT 67.950 655.950 70.050 656.400 ;
        RECT 85.950 657.600 88.050 658.050 ;
        RECT 121.950 657.600 124.050 658.050 ;
        RECT 85.950 656.400 124.050 657.600 ;
        RECT 164.400 656.400 169.050 658.050 ;
        RECT 85.950 655.950 88.050 656.400 ;
        RECT 121.950 655.950 124.050 656.400 ;
        RECT 165.000 655.950 169.050 656.400 ;
        RECT 181.950 657.600 184.050 658.050 ;
        RECT 187.950 657.600 190.050 658.050 ;
        RECT 181.950 656.400 190.050 657.600 ;
        RECT 181.950 655.950 184.050 656.400 ;
        RECT 187.950 655.950 190.050 656.400 ;
        RECT 262.950 657.600 265.050 658.050 ;
        RECT 268.950 657.600 271.050 658.050 ;
        RECT 262.950 656.400 271.050 657.600 ;
        RECT 262.950 655.950 265.050 656.400 ;
        RECT 268.950 655.950 271.050 656.400 ;
        RECT 286.950 657.600 289.050 658.050 ;
        RECT 298.950 657.600 301.050 658.050 ;
        RECT 286.950 656.400 301.050 657.600 ;
        RECT 286.950 655.950 289.050 656.400 ;
        RECT 298.950 655.950 301.050 656.400 ;
        RECT 439.950 657.600 442.050 658.050 ;
        RECT 448.950 657.600 451.050 658.050 ;
        RECT 439.950 656.400 451.050 657.600 ;
        RECT 439.950 655.950 442.050 656.400 ;
        RECT 448.950 655.950 451.050 656.400 ;
        RECT 505.950 657.600 508.050 658.050 ;
        RECT 529.950 657.600 532.050 658.050 ;
        RECT 505.950 656.400 532.050 657.600 ;
        RECT 505.950 655.950 508.050 656.400 ;
        RECT 529.950 655.950 532.050 656.400 ;
        RECT 622.950 657.600 625.050 658.050 ;
        RECT 634.950 657.600 637.050 658.050 ;
        RECT 622.950 656.400 637.050 657.600 ;
        RECT 622.950 655.950 625.050 656.400 ;
        RECT 634.950 655.950 637.050 656.400 ;
        RECT 772.950 657.600 775.050 658.050 ;
        RECT 850.950 657.600 853.050 658.050 ;
        RECT 772.950 656.400 853.050 657.600 ;
        RECT 772.950 655.950 775.050 656.400 ;
        RECT 850.950 655.950 853.050 656.400 ;
        RECT 856.950 657.600 859.050 658.050 ;
        RECT 868.950 657.600 871.050 658.050 ;
        RECT 874.950 657.600 877.050 658.050 ;
        RECT 856.950 656.400 877.050 657.600 ;
        RECT 856.950 655.950 859.050 656.400 ;
        RECT 868.950 655.950 871.050 656.400 ;
        RECT 874.950 655.950 877.050 656.400 ;
        RECT 127.950 654.600 130.050 655.050 ;
        RECT 74.400 653.400 130.050 654.600 ;
        RECT 74.400 645.900 75.600 653.400 ;
        RECT 127.950 652.950 130.050 653.400 ;
        RECT 139.950 654.600 142.050 655.050 ;
        RECT 148.950 654.600 151.050 655.050 ;
        RECT 220.950 654.600 223.050 655.050 ;
        RECT 139.950 653.400 151.050 654.600 ;
        RECT 139.950 652.950 142.050 653.400 ;
        RECT 148.950 652.950 151.050 653.400 ;
        RECT 188.400 653.400 223.050 654.600 ;
        RECT 88.950 649.950 91.050 652.050 ;
        RECT 160.950 651.600 163.050 652.050 ;
        RECT 184.950 651.600 187.050 652.050 ;
        RECT 160.950 650.400 187.050 651.600 ;
        RECT 160.950 649.950 163.050 650.400 ;
        RECT 184.950 649.950 187.050 650.400 ;
        RECT 89.400 646.050 90.600 649.950 ;
        RECT 188.400 649.050 189.600 653.400 ;
        RECT 220.950 652.950 223.050 653.400 ;
        RECT 301.950 654.600 304.050 655.050 ;
        RECT 313.950 654.600 316.050 655.050 ;
        RECT 319.950 654.600 322.050 655.050 ;
        RECT 301.950 653.400 322.050 654.600 ;
        RECT 301.950 652.950 304.050 653.400 ;
        RECT 313.950 652.950 316.050 653.400 ;
        RECT 319.950 652.950 322.050 653.400 ;
        RECT 436.950 654.600 439.050 655.050 ;
        RECT 451.950 654.600 454.050 655.050 ;
        RECT 436.950 653.400 454.050 654.600 ;
        RECT 436.950 652.950 439.050 653.400 ;
        RECT 451.950 652.950 454.050 653.400 ;
        RECT 460.950 654.600 463.050 655.050 ;
        RECT 478.950 654.600 481.050 655.050 ;
        RECT 460.950 653.400 481.050 654.600 ;
        RECT 460.950 652.950 463.050 653.400 ;
        RECT 478.950 652.950 481.050 653.400 ;
        RECT 490.950 654.600 493.050 655.050 ;
        RECT 499.950 654.600 502.050 655.050 ;
        RECT 490.950 653.400 502.050 654.600 ;
        RECT 490.950 652.950 493.050 653.400 ;
        RECT 499.950 652.950 502.050 653.400 ;
        RECT 541.950 654.600 544.050 655.050 ;
        RECT 613.950 654.600 616.050 655.050 ;
        RECT 541.950 653.400 616.050 654.600 ;
        RECT 541.950 652.950 544.050 653.400 ;
        RECT 613.950 652.950 616.050 653.400 ;
        RECT 643.950 654.600 646.050 655.050 ;
        RECT 676.950 654.600 679.050 655.050 ;
        RECT 643.950 653.400 679.050 654.600 ;
        RECT 643.950 652.950 646.050 653.400 ;
        RECT 676.950 652.950 679.050 653.400 ;
        RECT 781.950 654.600 784.050 655.050 ;
        RECT 790.950 654.600 793.050 655.050 ;
        RECT 781.950 653.400 793.050 654.600 ;
        RECT 781.950 652.950 784.050 653.400 ;
        RECT 790.950 652.950 793.050 653.400 ;
        RECT 136.950 648.600 139.050 649.050 ;
        RECT 186.000 648.900 189.600 649.050 ;
        RECT 104.400 647.400 139.050 648.600 ;
        RECT 73.950 643.800 76.050 645.900 ;
        RECT 88.950 643.950 91.050 646.050 ;
        RECT 94.950 645.450 97.050 645.900 ;
        RECT 100.950 645.450 103.050 645.900 ;
        RECT 94.950 644.250 103.050 645.450 ;
        RECT 94.950 643.800 97.050 644.250 ;
        RECT 100.950 643.800 103.050 644.250 ;
        RECT 43.950 642.600 46.050 643.050 ;
        RECT 104.400 642.600 105.600 647.400 ;
        RECT 136.950 646.950 139.050 647.400 ;
        RECT 184.950 647.400 189.600 648.900 ;
        RECT 190.950 648.600 193.050 652.050 ;
        RECT 202.950 651.600 205.050 652.200 ;
        RECT 238.950 651.600 241.050 652.200 ;
        RECT 202.950 650.400 241.050 651.600 ;
        RECT 202.950 650.100 205.050 650.400 ;
        RECT 238.950 650.100 241.050 650.400 ;
        RECT 244.950 650.100 247.050 652.200 ;
        RECT 286.950 650.100 289.050 652.200 ;
        RECT 304.950 650.100 307.050 652.200 ;
        RECT 322.950 650.100 325.050 652.200 ;
        RECT 444.000 651.600 448.050 652.050 ;
        RECT 190.950 648.000 204.600 648.600 ;
        RECT 191.400 647.400 204.600 648.000 ;
        RECT 184.950 646.950 189.000 647.400 ;
        RECT 184.950 646.800 187.050 646.950 ;
        RECT 115.950 645.450 118.050 645.900 ;
        RECT 124.950 645.450 127.050 645.900 ;
        RECT 115.950 644.250 127.050 645.450 ;
        RECT 115.950 643.800 118.050 644.250 ;
        RECT 124.950 643.800 127.050 644.250 ;
        RECT 130.950 645.450 133.050 645.900 ;
        RECT 142.950 645.450 145.050 645.900 ;
        RECT 130.950 644.250 145.050 645.450 ;
        RECT 130.950 643.800 133.050 644.250 ;
        RECT 142.950 643.800 145.050 644.250 ;
        RECT 172.950 645.600 175.050 645.900 ;
        RECT 199.950 645.600 202.050 645.900 ;
        RECT 172.950 644.400 202.050 645.600 ;
        RECT 203.400 645.600 204.600 647.400 ;
        RECT 214.950 645.600 217.050 646.050 ;
        RECT 203.400 644.400 217.050 645.600 ;
        RECT 172.950 643.800 175.050 644.400 ;
        RECT 199.950 643.800 202.050 644.400 ;
        RECT 214.950 643.950 217.050 644.400 ;
        RECT 229.950 645.450 232.050 645.900 ;
        RECT 235.950 645.450 238.050 645.900 ;
        RECT 229.950 644.250 238.050 645.450 ;
        RECT 229.950 643.800 232.050 644.250 ;
        RECT 235.950 643.800 238.050 644.250 ;
        RECT 43.950 641.400 105.600 642.600 ;
        RECT 187.950 642.600 190.050 643.050 ;
        RECT 193.950 642.600 196.050 643.050 ;
        RECT 187.950 641.400 196.050 642.600 ;
        RECT 43.950 640.950 46.050 641.400 ;
        RECT 187.950 640.950 190.050 641.400 ;
        RECT 193.950 640.950 196.050 641.400 ;
        RECT 217.950 642.600 220.050 643.050 ;
        RECT 245.400 642.600 246.600 650.100 ;
        RECT 287.400 648.600 288.600 650.100 ;
        RECT 305.400 648.600 306.600 650.100 ;
        RECT 323.400 648.600 324.600 650.100 ;
        RECT 443.400 649.950 448.050 651.600 ;
        RECT 481.950 651.600 484.050 652.200 ;
        RECT 505.950 651.600 508.050 652.050 ;
        RECT 481.950 650.400 508.050 651.600 ;
        RECT 481.950 650.100 484.050 650.400 ;
        RECT 505.950 649.950 508.050 650.400 ;
        RECT 511.950 649.950 514.050 652.050 ;
        RECT 523.950 650.100 526.050 652.200 ;
        RECT 631.950 651.600 634.050 652.200 ;
        RECT 617.400 650.400 634.050 651.600 ;
        RECT 358.950 648.600 361.050 649.200 ;
        RECT 287.400 647.400 306.600 648.600 ;
        RECT 311.400 648.000 324.600 648.600 ;
        RECT 329.400 648.000 361.050 648.600 ;
        RECT 310.950 647.400 324.600 648.000 ;
        RECT 328.950 647.400 361.050 648.000 ;
        RECT 247.950 645.600 250.050 646.050 ;
        RECT 253.950 645.600 256.050 646.050 ;
        RECT 247.950 644.400 256.050 645.600 ;
        RECT 287.400 645.600 288.600 647.400 ;
        RECT 292.950 645.600 295.050 646.050 ;
        RECT 287.400 644.400 295.050 645.600 ;
        RECT 247.950 643.950 250.050 644.400 ;
        RECT 253.950 643.950 256.050 644.400 ;
        RECT 292.950 643.950 295.050 644.400 ;
        RECT 301.950 645.450 304.050 645.900 ;
        RECT 307.800 645.450 309.900 645.900 ;
        RECT 301.950 644.250 309.900 645.450 ;
        RECT 301.950 643.800 304.050 644.250 ;
        RECT 307.800 643.800 309.900 644.250 ;
        RECT 310.950 643.950 313.050 647.400 ;
        RECT 328.950 643.950 331.050 647.400 ;
        RECT 358.950 647.100 361.050 647.400 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 371.400 643.050 372.600 646.950 ;
        RECT 443.400 645.900 444.600 649.950 ;
        RECT 463.950 648.600 466.050 649.050 ;
        RECT 463.950 647.400 498.600 648.600 ;
        RECT 463.950 646.950 466.050 647.400 ;
        RECT 476.400 645.900 477.600 647.400 ;
        RECT 497.400 645.900 498.600 647.400 ;
        RECT 512.400 646.050 513.600 649.950 ;
        RECT 524.400 646.050 525.600 650.100 ;
        RECT 529.950 647.100 532.050 649.200 ;
        RECT 442.950 643.800 445.050 645.900 ;
        RECT 475.950 643.800 478.050 645.900 ;
        RECT 496.950 643.800 499.050 645.900 ;
        RECT 511.950 643.950 514.050 646.050 ;
        RECT 524.400 644.400 529.050 646.050 ;
        RECT 525.000 643.950 529.050 644.400 ;
        RECT 262.950 642.600 265.050 643.050 ;
        RECT 217.950 641.400 265.050 642.600 ;
        RECT 217.950 640.950 220.050 641.400 ;
        RECT 262.950 640.950 265.050 641.400 ;
        RECT 277.950 642.600 280.050 643.050 ;
        RECT 283.950 642.600 286.050 643.050 ;
        RECT 277.950 641.400 286.050 642.600 ;
        RECT 277.950 640.950 280.050 641.400 ;
        RECT 283.950 640.950 286.050 641.400 ;
        RECT 370.950 640.950 373.050 643.050 ;
        RECT 418.950 642.450 421.050 642.900 ;
        RECT 439.950 642.450 442.050 643.050 ;
        RECT 454.950 642.450 457.050 642.900 ;
        RECT 418.950 641.250 457.050 642.450 ;
        RECT 418.950 640.800 421.050 641.250 ;
        RECT 439.950 640.950 442.050 641.250 ;
        RECT 454.950 640.800 457.050 641.250 ;
        RECT 478.950 642.600 481.050 643.050 ;
        RECT 487.950 642.600 490.050 643.050 ;
        RECT 478.950 641.400 490.050 642.600 ;
        RECT 478.950 640.950 481.050 641.400 ;
        RECT 487.950 640.950 490.050 641.400 ;
        RECT 517.950 642.600 520.050 643.050 ;
        RECT 530.400 642.600 531.600 647.100 ;
        RECT 541.800 646.950 543.900 649.050 ;
        RECT 568.950 648.600 571.050 649.050 ;
        RECT 586.950 648.600 589.050 649.050 ;
        RECT 568.950 647.400 589.050 648.600 ;
        RECT 568.950 646.950 571.050 647.400 ;
        RECT 586.950 646.950 589.050 647.400 ;
        RECT 542.250 643.050 543.450 646.950 ;
        RECT 601.950 645.450 604.050 646.050 ;
        RECT 617.400 645.900 618.600 650.400 ;
        RECT 631.950 650.100 634.050 650.400 ;
        RECT 679.950 651.600 682.050 652.200 ;
        RECT 685.950 651.600 688.050 652.050 ;
        RECT 694.950 651.600 697.050 652.200 ;
        RECT 679.950 650.400 697.050 651.600 ;
        RECT 679.950 650.100 682.050 650.400 ;
        RECT 685.950 649.950 688.050 650.400 ;
        RECT 694.950 650.100 697.050 650.400 ;
        RECT 700.950 651.600 703.050 652.200 ;
        RECT 862.950 651.600 865.050 652.200 ;
        RECT 895.950 651.600 898.050 652.200 ;
        RECT 910.950 651.600 913.050 652.200 ;
        RECT 700.950 650.400 717.600 651.600 ;
        RECT 700.950 650.100 703.050 650.400 ;
        RECT 716.400 645.900 717.600 650.400 ;
        RECT 815.400 650.400 865.050 651.600 ;
        RECT 610.950 645.450 613.050 645.900 ;
        RECT 601.950 644.250 613.050 645.450 ;
        RECT 601.950 643.950 604.050 644.250 ;
        RECT 610.950 643.800 613.050 644.250 ;
        RECT 616.950 643.800 619.050 645.900 ;
        RECT 676.950 645.600 679.050 645.900 ;
        RECT 691.950 645.600 694.050 645.900 ;
        RECT 676.950 644.400 694.050 645.600 ;
        RECT 676.950 643.800 679.050 644.400 ;
        RECT 691.950 643.800 694.050 644.400 ;
        RECT 715.950 643.800 718.050 645.900 ;
        RECT 787.950 645.600 790.050 646.050 ;
        RECT 802.950 645.600 805.050 646.050 ;
        RECT 815.400 645.900 816.600 650.400 ;
        RECT 862.950 650.100 865.050 650.400 ;
        RECT 866.400 650.400 913.050 651.600 ;
        RECT 866.400 645.900 867.600 650.400 ;
        RECT 895.950 650.100 898.050 650.400 ;
        RECT 910.950 650.100 913.050 650.400 ;
        RECT 931.950 650.100 934.050 652.200 ;
        RECT 787.950 644.400 805.050 645.600 ;
        RECT 787.950 643.950 790.050 644.400 ;
        RECT 802.950 643.950 805.050 644.400 ;
        RECT 814.950 643.800 817.050 645.900 ;
        RECT 865.950 643.800 868.050 645.900 ;
        RECT 913.950 645.600 916.050 645.900 ;
        RECT 932.400 645.600 933.600 650.100 ;
        RECT 913.950 644.400 933.600 645.600 ;
        RECT 913.950 643.800 916.050 644.400 ;
        RECT 517.950 641.400 531.600 642.600 ;
        RECT 517.950 640.950 520.050 641.400 ;
        RECT 541.800 640.950 543.900 643.050 ;
        RECT 544.950 642.600 547.050 643.050 ;
        RECT 589.950 642.600 592.050 642.900 ;
        RECT 544.950 642.450 592.050 642.600 ;
        RECT 622.950 642.450 625.050 642.900 ;
        RECT 544.950 641.400 625.050 642.450 ;
        RECT 544.950 640.950 547.050 641.400 ;
        RECT 589.950 641.250 625.050 641.400 ;
        RECT 589.950 640.800 592.050 641.250 ;
        RECT 622.950 640.800 625.050 641.250 ;
        RECT 631.950 642.600 634.050 643.050 ;
        RECT 658.950 642.600 661.050 643.050 ;
        RECT 631.950 641.400 661.050 642.600 ;
        RECT 631.950 640.950 634.050 641.400 ;
        RECT 658.950 640.950 661.050 641.400 ;
        RECT 856.950 642.600 859.050 643.050 ;
        RECT 868.950 642.600 871.050 643.050 ;
        RECT 856.950 641.400 871.050 642.600 ;
        RECT 856.950 640.950 859.050 641.400 ;
        RECT 868.950 640.950 871.050 641.400 ;
        RECT 28.950 639.600 31.050 640.050 ;
        RECT 64.800 639.600 66.900 640.050 ;
        RECT 28.950 638.400 66.900 639.600 ;
        RECT 28.950 637.950 31.050 638.400 ;
        RECT 64.800 637.950 66.900 638.400 ;
        RECT 67.950 639.600 70.050 640.050 ;
        RECT 127.950 639.600 130.050 640.050 ;
        RECT 67.950 638.400 130.050 639.600 ;
        RECT 67.950 637.950 70.050 638.400 ;
        RECT 127.950 637.950 130.050 638.400 ;
        RECT 148.950 639.600 151.050 640.050 ;
        RECT 220.800 639.600 222.900 640.050 ;
        RECT 148.950 638.400 222.900 639.600 ;
        RECT 148.950 637.950 151.050 638.400 ;
        RECT 220.800 637.950 222.900 638.400 ;
        RECT 223.950 639.600 226.050 640.050 ;
        RECT 241.950 639.600 244.050 640.050 ;
        RECT 256.950 639.600 259.050 640.050 ;
        RECT 223.950 638.400 259.050 639.600 ;
        RECT 223.950 637.950 226.050 638.400 ;
        RECT 241.950 637.950 244.050 638.400 ;
        RECT 256.950 637.950 259.050 638.400 ;
        RECT 286.950 639.600 289.050 640.050 ;
        RECT 319.950 639.600 322.050 640.050 ;
        RECT 334.950 639.600 337.050 640.050 ;
        RECT 286.950 638.400 337.050 639.600 ;
        RECT 286.950 637.950 289.050 638.400 ;
        RECT 319.950 637.950 322.050 638.400 ;
        RECT 334.950 637.950 337.050 638.400 ;
        RECT 490.950 639.600 493.050 640.050 ;
        RECT 514.950 639.600 517.050 640.050 ;
        RECT 490.950 638.400 517.050 639.600 ;
        RECT 490.950 637.950 493.050 638.400 ;
        RECT 514.950 637.950 517.050 638.400 ;
        RECT 70.950 636.600 73.050 637.050 ;
        RECT 154.950 636.600 157.050 637.050 ;
        RECT 70.950 635.400 157.050 636.600 ;
        RECT 70.950 634.950 73.050 635.400 ;
        RECT 154.950 634.950 157.050 635.400 ;
        RECT 163.950 636.600 166.050 637.050 ;
        RECT 214.950 636.600 217.050 637.050 ;
        RECT 265.950 636.600 268.050 637.050 ;
        RECT 163.950 635.400 195.600 636.600 ;
        RECT 163.950 634.950 166.050 635.400 ;
        RECT 19.950 633.600 22.050 634.050 ;
        RECT 58.950 633.600 61.050 634.050 ;
        RECT 19.950 632.400 61.050 633.600 ;
        RECT 19.950 631.950 22.050 632.400 ;
        RECT 58.950 631.950 61.050 632.400 ;
        RECT 79.950 633.600 82.050 634.050 ;
        RECT 106.950 633.600 109.050 634.050 ;
        RECT 79.950 632.400 109.050 633.600 ;
        RECT 79.950 631.950 82.050 632.400 ;
        RECT 106.950 631.950 109.050 632.400 ;
        RECT 115.950 633.600 118.050 634.050 ;
        RECT 139.950 633.600 142.050 634.050 ;
        RECT 166.950 633.600 169.050 634.050 ;
        RECT 115.950 632.400 169.050 633.600 ;
        RECT 194.400 633.600 195.600 635.400 ;
        RECT 214.950 635.400 268.050 636.600 ;
        RECT 214.950 634.950 217.050 635.400 ;
        RECT 265.950 634.950 268.050 635.400 ;
        RECT 289.950 636.600 292.050 637.050 ;
        RECT 310.950 636.600 313.050 637.050 ;
        RECT 289.950 635.400 313.050 636.600 ;
        RECT 289.950 634.950 292.050 635.400 ;
        RECT 310.950 634.950 313.050 635.400 ;
        RECT 328.950 636.600 331.050 637.050 ;
        RECT 358.950 636.600 361.050 637.050 ;
        RECT 328.950 635.400 361.050 636.600 ;
        RECT 328.950 634.950 331.050 635.400 ;
        RECT 358.950 634.950 361.050 635.400 ;
        RECT 436.950 636.600 439.050 637.050 ;
        RECT 457.950 636.600 460.050 637.050 ;
        RECT 436.950 635.400 460.050 636.600 ;
        RECT 436.950 634.950 439.050 635.400 ;
        RECT 457.950 634.950 460.050 635.400 ;
        RECT 535.950 636.600 538.050 637.050 ;
        RECT 565.950 636.600 568.050 637.050 ;
        RECT 535.950 635.400 568.050 636.600 ;
        RECT 568.950 636.600 571.050 640.050 ;
        RECT 610.950 639.600 613.050 640.050 ;
        RECT 628.950 639.600 631.050 640.050 ;
        RECT 610.950 638.400 631.050 639.600 ;
        RECT 610.950 637.950 613.050 638.400 ;
        RECT 628.950 637.950 631.050 638.400 ;
        RECT 667.950 639.600 670.050 640.050 ;
        RECT 685.950 639.600 688.050 640.050 ;
        RECT 721.950 639.600 724.050 640.050 ;
        RECT 667.950 638.400 724.050 639.600 ;
        RECT 667.950 637.950 670.050 638.400 ;
        RECT 685.950 637.950 688.050 638.400 ;
        RECT 721.950 637.950 724.050 638.400 ;
        RECT 811.950 639.600 814.050 640.050 ;
        RECT 829.950 639.600 832.050 640.050 ;
        RECT 811.950 638.400 832.050 639.600 ;
        RECT 811.950 637.950 814.050 638.400 ;
        RECT 829.950 637.950 832.050 638.400 ;
        RECT 919.950 639.600 922.050 640.050 ;
        RECT 934.950 639.600 937.050 640.050 ;
        RECT 919.950 638.400 937.050 639.600 ;
        RECT 919.950 637.950 922.050 638.400 ;
        RECT 934.950 637.950 937.050 638.400 ;
        RECT 595.950 636.600 598.050 637.050 ;
        RECT 568.950 636.000 598.050 636.600 ;
        RECT 569.400 635.400 598.050 636.000 ;
        RECT 535.950 634.950 538.050 635.400 ;
        RECT 565.950 634.950 568.050 635.400 ;
        RECT 595.950 634.950 598.050 635.400 ;
        RECT 607.950 636.600 610.050 637.050 ;
        RECT 640.950 636.600 643.050 637.050 ;
        RECT 649.950 636.600 652.050 637.050 ;
        RECT 607.950 635.400 652.050 636.600 ;
        RECT 607.950 634.950 610.050 635.400 ;
        RECT 640.950 634.950 643.050 635.400 ;
        RECT 649.950 634.950 652.050 635.400 ;
        RECT 748.950 636.600 751.050 637.050 ;
        RECT 760.950 636.600 763.050 637.050 ;
        RECT 748.950 635.400 763.050 636.600 ;
        RECT 748.950 634.950 751.050 635.400 ;
        RECT 760.950 634.950 763.050 635.400 ;
        RECT 823.950 636.600 826.050 637.050 ;
        RECT 832.950 636.600 835.050 637.050 ;
        RECT 823.950 635.400 835.050 636.600 ;
        RECT 823.950 634.950 826.050 635.400 ;
        RECT 832.950 634.950 835.050 635.400 ;
        RECT 856.950 636.600 859.050 637.050 ;
        RECT 871.950 636.600 874.050 637.050 ;
        RECT 877.950 636.600 880.050 637.050 ;
        RECT 856.950 635.400 880.050 636.600 ;
        RECT 856.950 634.950 859.050 635.400 ;
        RECT 871.950 634.950 874.050 635.400 ;
        RECT 877.950 634.950 880.050 635.400 ;
        RECT 280.950 633.600 283.050 634.050 ;
        RECT 194.400 632.400 283.050 633.600 ;
        RECT 115.950 631.950 118.050 632.400 ;
        RECT 139.950 631.950 142.050 632.400 ;
        RECT 166.950 631.950 169.050 632.400 ;
        RECT 280.950 631.950 283.050 632.400 ;
        RECT 421.950 633.600 424.050 634.050 ;
        RECT 493.950 633.600 496.050 634.050 ;
        RECT 586.950 633.600 589.050 634.050 ;
        RECT 421.950 632.400 486.600 633.600 ;
        RECT 421.950 631.950 424.050 632.400 ;
        RECT 49.950 630.600 52.050 631.050 ;
        RECT 73.950 630.600 76.050 631.050 ;
        RECT 49.950 629.400 76.050 630.600 ;
        RECT 49.950 628.950 52.050 629.400 ;
        RECT 73.950 628.950 76.050 629.400 ;
        RECT 217.950 630.600 220.050 631.050 ;
        RECT 355.950 630.600 358.050 631.050 ;
        RECT 364.950 630.600 367.050 631.050 ;
        RECT 454.950 630.600 457.050 631.050 ;
        RECT 217.950 629.400 339.600 630.600 ;
        RECT 217.950 628.950 220.050 629.400 ;
        RECT 79.950 627.600 82.050 628.050 ;
        RECT 91.950 627.600 94.050 628.050 ;
        RECT 79.950 626.400 94.050 627.600 ;
        RECT 79.950 625.950 82.050 626.400 ;
        RECT 91.950 625.950 94.050 626.400 ;
        RECT 124.950 627.600 127.050 628.050 ;
        RECT 199.950 627.600 202.050 628.050 ;
        RECT 205.950 627.600 208.050 628.050 ;
        RECT 124.950 626.400 208.050 627.600 ;
        RECT 124.950 625.950 127.050 626.400 ;
        RECT 199.950 625.950 202.050 626.400 ;
        RECT 205.950 625.950 208.050 626.400 ;
        RECT 220.950 627.600 223.050 628.050 ;
        RECT 271.950 627.600 274.050 628.050 ;
        RECT 220.950 626.400 274.050 627.600 ;
        RECT 220.950 625.950 223.050 626.400 ;
        RECT 271.950 625.950 274.050 626.400 ;
        RECT 280.950 627.600 283.050 628.050 ;
        RECT 328.950 627.600 331.050 628.050 ;
        RECT 280.950 626.400 331.050 627.600 ;
        RECT 338.400 627.600 339.600 629.400 ;
        RECT 355.950 629.400 457.050 630.600 ;
        RECT 485.400 630.600 486.600 632.400 ;
        RECT 493.950 632.400 589.050 633.600 ;
        RECT 493.950 631.950 496.050 632.400 ;
        RECT 586.950 631.950 589.050 632.400 ;
        RECT 604.950 633.600 607.050 634.050 ;
        RECT 610.950 633.600 613.050 634.050 ;
        RECT 604.950 632.400 613.050 633.600 ;
        RECT 604.950 631.950 607.050 632.400 ;
        RECT 610.950 631.950 613.050 632.400 ;
        RECT 622.950 633.600 625.050 634.050 ;
        RECT 643.950 633.600 646.050 634.050 ;
        RECT 622.950 632.400 646.050 633.600 ;
        RECT 622.950 631.950 625.050 632.400 ;
        RECT 643.950 631.950 646.050 632.400 ;
        RECT 592.950 630.600 595.050 631.050 ;
        RECT 640.950 630.600 643.050 631.050 ;
        RECT 485.400 629.400 643.050 630.600 ;
        RECT 355.950 628.950 358.050 629.400 ;
        RECT 364.950 628.950 367.050 629.400 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 592.950 628.950 595.050 629.400 ;
        RECT 640.950 628.950 643.050 629.400 ;
        RECT 694.950 630.600 697.050 631.050 ;
        RECT 730.950 630.600 733.050 631.050 ;
        RECT 694.950 629.400 733.050 630.600 ;
        RECT 694.950 628.950 697.050 629.400 ;
        RECT 730.950 628.950 733.050 629.400 ;
        RECT 871.950 630.600 874.050 631.050 ;
        RECT 886.950 630.600 889.050 631.050 ;
        RECT 907.950 630.600 910.050 631.050 ;
        RECT 871.950 629.400 910.050 630.600 ;
        RECT 871.950 628.950 874.050 629.400 ;
        RECT 886.950 628.950 889.050 629.400 ;
        RECT 907.950 628.950 910.050 629.400 ;
        RECT 436.950 627.600 439.050 628.050 ;
        RECT 338.400 626.400 439.050 627.600 ;
        RECT 280.950 625.950 283.050 626.400 ;
        RECT 328.950 625.950 331.050 626.400 ;
        RECT 436.950 625.950 439.050 626.400 ;
        RECT 634.950 627.600 637.050 628.050 ;
        RECT 652.950 627.600 655.050 628.050 ;
        RECT 634.950 626.400 655.050 627.600 ;
        RECT 634.950 625.950 637.050 626.400 ;
        RECT 652.950 625.950 655.050 626.400 ;
        RECT 715.950 627.600 718.050 628.050 ;
        RECT 781.950 627.600 784.050 628.050 ;
        RECT 715.950 626.400 784.050 627.600 ;
        RECT 715.950 625.950 718.050 626.400 ;
        RECT 781.950 625.950 784.050 626.400 ;
        RECT 121.950 624.600 124.050 625.050 ;
        RECT 136.950 624.600 139.050 625.050 ;
        RECT 207.000 624.600 211.050 625.050 ;
        RECT 121.950 623.400 139.050 624.600 ;
        RECT 121.950 622.950 124.050 623.400 ;
        RECT 136.950 622.950 139.050 623.400 ;
        RECT 206.400 622.950 211.050 624.600 ;
        RECT 307.950 624.600 310.050 625.050 ;
        RECT 313.950 624.600 316.050 625.050 ;
        RECT 307.950 623.400 316.050 624.600 ;
        RECT 307.950 622.950 310.050 623.400 ;
        RECT 313.950 622.950 316.050 623.400 ;
        RECT 400.950 624.600 403.050 625.050 ;
        RECT 409.950 624.600 412.050 625.050 ;
        RECT 400.950 623.400 412.050 624.600 ;
        RECT 400.950 622.950 403.050 623.400 ;
        RECT 409.950 622.950 412.050 623.400 ;
        RECT 418.950 624.600 421.050 625.050 ;
        RECT 502.950 624.600 505.050 625.050 ;
        RECT 520.950 624.600 523.050 625.050 ;
        RECT 655.950 624.600 658.050 625.050 ;
        RECT 418.950 623.400 658.050 624.600 ;
        RECT 418.950 622.950 421.050 623.400 ;
        RECT 502.950 622.950 505.050 623.400 ;
        RECT 520.950 622.950 523.050 623.400 ;
        RECT 655.950 622.950 658.050 623.400 ;
        RECT 706.950 624.600 709.050 625.050 ;
        RECT 730.950 624.600 733.050 625.050 ;
        RECT 706.950 623.400 733.050 624.600 ;
        RECT 706.950 622.950 709.050 623.400 ;
        RECT 730.950 622.950 733.050 623.400 ;
        RECT 73.950 621.600 76.050 622.050 ;
        RECT 184.950 621.600 187.050 622.050 ;
        RECT 206.400 621.600 207.600 622.950 ;
        RECT 73.950 620.400 207.600 621.600 ;
        RECT 211.950 621.600 214.050 622.050 ;
        RECT 232.950 621.600 235.050 622.050 ;
        RECT 211.950 620.400 235.050 621.600 ;
        RECT 73.950 619.950 76.050 620.400 ;
        RECT 184.950 619.950 187.050 620.400 ;
        RECT 211.950 619.950 214.050 620.400 ;
        RECT 232.950 619.950 235.050 620.400 ;
        RECT 274.950 621.600 277.050 622.050 ;
        RECT 280.950 621.600 283.050 622.050 ;
        RECT 274.950 620.400 283.050 621.600 ;
        RECT 274.950 619.950 277.050 620.400 ;
        RECT 280.950 619.950 283.050 620.400 ;
        RECT 415.950 621.600 418.050 621.900 ;
        RECT 427.950 621.600 430.050 622.050 ;
        RECT 415.950 620.400 430.050 621.600 ;
        RECT 415.950 619.800 418.050 620.400 ;
        RECT 427.950 619.950 430.050 620.400 ;
        RECT 436.950 621.600 439.050 622.050 ;
        RECT 448.950 621.600 451.050 622.050 ;
        RECT 436.950 620.400 451.050 621.600 ;
        RECT 436.950 619.950 439.050 620.400 ;
        RECT 448.950 619.950 451.050 620.400 ;
        RECT 454.950 621.600 457.050 622.050 ;
        RECT 472.950 621.600 475.050 622.050 ;
        RECT 454.950 620.400 475.050 621.600 ;
        RECT 454.950 619.950 457.050 620.400 ;
        RECT 472.950 619.950 475.050 620.400 ;
        RECT 541.950 621.600 544.050 622.050 ;
        RECT 547.950 621.600 550.050 622.050 ;
        RECT 541.950 620.400 550.050 621.600 ;
        RECT 541.950 619.950 544.050 620.400 ;
        RECT 547.950 619.950 550.050 620.400 ;
        RECT 31.950 618.600 34.050 619.050 ;
        RECT 61.800 618.600 63.900 619.050 ;
        RECT 31.950 617.400 63.900 618.600 ;
        RECT 31.950 616.950 34.050 617.400 ;
        RECT 61.800 616.950 63.900 617.400 ;
        RECT 64.950 618.600 67.050 619.050 ;
        RECT 106.950 618.600 109.050 619.050 ;
        RECT 121.950 618.600 124.050 619.050 ;
        RECT 208.950 618.600 211.050 619.050 ;
        RECT 64.950 617.400 124.050 618.600 ;
        RECT 64.950 616.950 67.050 617.400 ;
        RECT 106.950 616.950 109.050 617.400 ;
        RECT 121.950 616.950 124.050 617.400 ;
        RECT 149.400 617.400 211.050 618.600 ;
        RECT 149.400 615.600 150.600 617.400 ;
        RECT 208.950 616.950 211.050 617.400 ;
        RECT 295.950 618.600 298.050 619.050 ;
        RECT 313.950 618.600 316.050 619.050 ;
        RECT 295.950 617.400 316.050 618.600 ;
        RECT 295.950 616.950 298.050 617.400 ;
        RECT 313.950 616.950 316.050 617.400 ;
        RECT 337.950 618.600 340.050 619.050 ;
        RECT 373.950 618.600 376.050 619.050 ;
        RECT 337.950 617.400 376.050 618.600 ;
        RECT 337.950 616.950 340.050 617.400 ;
        RECT 373.950 616.950 376.050 617.400 ;
        RECT 433.950 618.600 436.050 619.050 ;
        RECT 451.950 618.600 454.050 619.050 ;
        RECT 433.950 617.400 454.050 618.600 ;
        RECT 433.950 616.950 436.050 617.400 ;
        RECT 451.950 616.950 454.050 617.400 ;
        RECT 562.950 618.600 565.050 619.050 ;
        RECT 598.950 618.600 601.050 619.050 ;
        RECT 562.950 617.400 601.050 618.600 ;
        RECT 562.950 616.950 565.050 617.400 ;
        RECT 598.950 616.950 601.050 617.400 ;
        RECT 137.400 614.400 150.600 615.600 ;
        RECT 322.950 615.600 325.050 616.050 ;
        RECT 334.950 615.600 337.050 616.050 ;
        RECT 346.950 615.600 349.050 616.050 ;
        RECT 322.950 614.400 349.050 615.600 ;
        RECT 25.950 610.950 28.050 613.050 ;
        RECT 58.950 612.600 61.050 613.050 ;
        RECT 70.950 612.600 73.050 613.050 ;
        RECT 94.950 612.600 97.050 613.050 ;
        RECT 58.950 611.400 97.050 612.600 ;
        RECT 58.950 610.950 61.050 611.400 ;
        RECT 70.950 610.950 73.050 611.400 ;
        RECT 94.950 610.950 97.050 611.400 ;
        RECT 22.950 604.950 25.050 607.050 ;
        RECT 16.950 600.600 19.050 600.900 ;
        RECT 23.400 600.600 24.600 604.950 ;
        RECT 16.950 599.400 24.600 600.600 ;
        RECT 26.400 600.600 27.600 610.950 ;
        RECT 82.950 609.600 85.050 610.050 ;
        RECT 115.950 609.600 118.050 610.050 ;
        RECT 82.950 608.400 118.050 609.600 ;
        RECT 37.950 604.950 40.050 607.050 ;
        RECT 79.950 606.600 82.050 607.200 ;
        RECT 68.400 605.400 82.050 606.600 ;
        RECT 82.950 606.600 85.050 608.400 ;
        RECT 115.950 607.950 118.050 608.400 ;
        RECT 88.950 606.600 91.050 606.900 ;
        RECT 82.950 606.000 91.050 606.600 ;
        RECT 83.400 605.400 91.050 606.000 ;
        RECT 38.400 603.600 39.600 604.950 ;
        RECT 46.950 603.600 49.050 604.050 ;
        RECT 38.400 602.400 49.050 603.600 ;
        RECT 46.950 601.950 49.050 602.400 ;
        RECT 68.400 601.050 69.600 605.400 ;
        RECT 79.950 605.100 82.050 605.400 ;
        RECT 88.950 604.800 91.050 605.400 ;
        RECT 100.950 605.100 103.050 607.200 ;
        RECT 118.950 606.600 121.050 607.200 ;
        RECT 133.950 606.600 136.050 607.200 ;
        RECT 118.950 605.400 136.050 606.600 ;
        RECT 118.950 605.100 121.050 605.400 ;
        RECT 133.950 605.100 136.050 605.400 ;
        RECT 34.950 600.600 37.050 600.900 ;
        RECT 26.400 599.400 37.050 600.600 ;
        RECT 16.950 598.800 19.050 599.400 ;
        RECT 34.950 598.800 37.050 599.400 ;
        RECT 67.950 598.950 70.050 601.050 ;
        RECT 101.400 598.050 102.600 605.100 ;
        RECT 137.400 600.900 138.600 614.400 ;
        RECT 322.950 613.950 325.050 614.400 ;
        RECT 334.950 613.950 337.050 614.400 ;
        RECT 346.950 613.950 349.050 614.400 ;
        RECT 424.950 615.600 427.050 616.050 ;
        RECT 604.950 615.600 607.050 616.050 ;
        RECT 424.950 614.400 607.050 615.600 ;
        RECT 424.950 613.950 427.050 614.400 ;
        RECT 604.950 613.950 607.050 614.400 ;
        RECT 763.950 615.600 766.050 616.050 ;
        RECT 817.950 615.600 820.050 616.050 ;
        RECT 844.950 615.600 847.050 616.050 ;
        RECT 763.950 614.400 847.050 615.600 ;
        RECT 763.950 613.950 766.050 614.400 ;
        RECT 817.950 613.950 820.050 614.400 ;
        RECT 844.950 613.950 847.050 614.400 ;
        RECT 145.950 612.600 148.050 613.050 ;
        RECT 151.950 612.600 154.050 613.050 ;
        RECT 145.950 611.400 154.050 612.600 ;
        RECT 145.950 610.950 148.050 611.400 ;
        RECT 151.950 610.950 154.050 611.400 ;
        RECT 220.950 612.600 223.050 613.050 ;
        RECT 226.950 612.600 229.050 613.050 ;
        RECT 220.950 611.400 229.050 612.600 ;
        RECT 220.950 610.950 223.050 611.400 ;
        RECT 226.950 610.950 229.050 611.400 ;
        RECT 259.950 612.600 262.050 613.050 ;
        RECT 325.950 612.600 328.050 613.050 ;
        RECT 352.950 612.600 355.050 613.050 ;
        RECT 259.950 611.400 355.050 612.600 ;
        RECT 259.950 610.950 262.050 611.400 ;
        RECT 325.950 610.950 328.050 611.400 ;
        RECT 352.950 610.950 355.050 611.400 ;
        RECT 358.950 612.600 361.050 613.050 ;
        RECT 448.950 612.600 451.050 613.050 ;
        RECT 358.950 611.400 451.050 612.600 ;
        RECT 358.950 610.950 361.050 611.400 ;
        RECT 448.950 610.950 451.050 611.400 ;
        RECT 511.950 612.600 514.050 613.050 ;
        RECT 526.950 612.600 529.050 613.050 ;
        RECT 511.950 611.400 529.050 612.600 ;
        RECT 511.950 610.950 514.050 611.400 ;
        RECT 526.950 610.950 529.050 611.400 ;
        RECT 580.950 612.600 583.050 613.050 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 631.950 612.600 634.050 613.050 ;
        RECT 676.950 612.600 679.050 613.050 ;
        RECT 580.950 611.400 634.050 612.600 ;
        RECT 580.950 610.950 583.050 611.400 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 631.950 610.950 634.050 611.400 ;
        RECT 647.400 611.400 679.050 612.600 ;
        RECT 169.950 609.600 172.050 610.050 ;
        RECT 178.950 609.600 181.050 610.050 ;
        RECT 169.950 608.400 181.050 609.600 ;
        RECT 169.950 607.950 172.050 608.400 ;
        RECT 178.950 607.950 181.050 608.400 ;
        RECT 205.950 609.600 208.050 609.900 ;
        RECT 235.950 609.600 238.050 610.050 ;
        RECT 241.950 609.600 244.050 610.050 ;
        RECT 205.950 608.400 244.050 609.600 ;
        RECT 205.950 607.800 208.050 608.400 ;
        RECT 235.950 607.950 238.050 608.400 ;
        RECT 241.950 607.950 244.050 608.400 ;
        RECT 250.950 607.950 253.050 610.050 ;
        RECT 316.950 609.600 319.050 610.050 ;
        RECT 367.800 609.600 369.900 610.050 ;
        RECT 316.950 608.400 369.900 609.600 ;
        RECT 316.950 607.950 319.050 608.400 ;
        RECT 367.800 607.950 369.900 608.400 ;
        RECT 370.950 609.600 373.050 610.050 ;
        RECT 388.950 609.600 391.050 610.050 ;
        RECT 370.950 608.400 391.050 609.600 ;
        RECT 370.950 607.950 373.050 608.400 ;
        RECT 388.950 607.950 391.050 608.400 ;
        RECT 151.950 606.600 154.050 607.050 ;
        RECT 143.400 605.400 154.050 606.600 ;
        RECT 143.400 600.900 144.600 605.400 ;
        RECT 151.950 604.950 154.050 605.400 ;
        RECT 160.950 605.100 163.050 607.200 ;
        RECT 166.950 606.750 169.050 607.200 ;
        RECT 172.950 606.750 175.050 607.200 ;
        RECT 166.950 605.550 175.050 606.750 ;
        RECT 166.950 605.100 169.050 605.550 ;
        RECT 172.950 605.100 175.050 605.550 ;
        RECT 190.950 606.750 193.050 607.200 ;
        RECT 205.950 606.750 208.050 607.200 ;
        RECT 190.950 605.550 208.050 606.750 ;
        RECT 190.950 605.100 193.050 605.550 ;
        RECT 205.950 605.100 208.050 605.550 ;
        RECT 214.950 606.750 217.050 607.200 ;
        RECT 220.950 606.750 223.050 607.200 ;
        RECT 214.950 605.550 223.050 606.750 ;
        RECT 214.950 605.100 217.050 605.550 ;
        RECT 220.950 605.100 223.050 605.550 ;
        RECT 161.400 603.600 162.600 605.100 ;
        RECT 161.400 603.000 171.600 603.600 ;
        RECT 161.400 602.400 172.050 603.000 ;
        RECT 136.950 598.800 139.050 600.900 ;
        RECT 142.950 598.800 145.050 600.900 ;
        RECT 157.950 600.600 160.050 600.900 ;
        RECT 166.800 600.600 168.900 601.050 ;
        RECT 157.950 599.400 168.900 600.600 ;
        RECT 157.950 598.800 160.050 599.400 ;
        RECT 166.800 598.950 168.900 599.400 ;
        RECT 169.950 598.950 172.050 602.400 ;
        RECT 175.950 600.600 178.050 600.900 ;
        RECT 190.950 600.600 193.050 601.050 ;
        RECT 175.950 599.400 193.050 600.600 ;
        RECT 175.950 598.800 178.050 599.400 ;
        RECT 190.950 598.950 193.050 599.400 ;
        RECT 202.950 600.600 205.050 600.900 ;
        RECT 214.950 600.600 217.050 601.050 ;
        RECT 202.950 599.400 217.050 600.600 ;
        RECT 202.950 598.800 205.050 599.400 ;
        RECT 214.950 598.950 217.050 599.400 ;
        RECT 229.950 600.450 232.050 600.900 ;
        RECT 235.950 600.450 238.050 600.900 ;
        RECT 229.950 599.250 238.050 600.450 ;
        RECT 229.950 598.800 232.050 599.250 ;
        RECT 235.950 598.800 238.050 599.250 ;
        RECT 251.400 598.050 252.600 607.950 ;
        RECT 253.950 606.750 256.050 607.200 ;
        RECT 259.950 606.750 262.050 607.200 ;
        RECT 253.950 605.550 262.050 606.750 ;
        RECT 268.950 606.600 271.050 607.200 ;
        RECT 253.950 605.100 256.050 605.550 ;
        RECT 259.950 605.100 262.050 605.550 ;
        RECT 266.400 605.400 271.050 606.600 ;
        RECT 266.400 601.050 267.600 605.400 ;
        RECT 268.950 605.100 271.050 605.400 ;
        RECT 289.950 606.600 292.050 607.200 ;
        RECT 289.950 605.400 297.600 606.600 ;
        RECT 289.950 605.100 292.050 605.400 ;
        RECT 296.400 603.600 297.600 605.400 ;
        RECT 340.950 605.100 343.050 607.200 ;
        RECT 346.950 606.600 349.050 607.200 ;
        RECT 361.950 606.600 364.050 607.200 ;
        RECT 346.950 605.400 364.050 606.600 ;
        RECT 346.950 605.100 349.050 605.400 ;
        RECT 361.950 605.100 364.050 605.400 ;
        RECT 367.950 606.600 370.050 607.200 ;
        RECT 382.950 606.600 385.050 607.200 ;
        RECT 367.950 605.400 385.050 606.600 ;
        RECT 367.950 605.100 370.050 605.400 ;
        RECT 382.950 605.100 385.050 605.400 ;
        RECT 403.950 606.600 406.050 607.050 ;
        RECT 430.950 606.600 433.050 607.050 ;
        RECT 433.950 606.600 436.050 610.050 ;
        RECT 453.000 609.600 457.050 610.050 ;
        RECT 452.400 607.950 457.050 609.600 ;
        RECT 502.950 609.750 505.050 610.200 ;
        RECT 508.950 609.750 511.050 610.200 ;
        RECT 502.950 608.550 511.050 609.750 ;
        RECT 502.950 608.100 505.050 608.550 ;
        RECT 508.950 608.100 511.050 608.550 ;
        RECT 523.950 607.950 526.050 610.050 ;
        RECT 571.950 609.750 574.050 610.200 ;
        RECT 589.950 609.750 592.050 610.200 ;
        RECT 571.950 608.550 592.050 609.750 ;
        RECT 571.950 608.100 574.050 608.550 ;
        RECT 589.950 608.100 592.050 608.550 ;
        RECT 598.950 609.600 601.050 610.050 ;
        RECT 616.950 609.600 619.050 610.050 ;
        RECT 647.400 609.600 648.600 611.400 ;
        RECT 676.950 610.950 679.050 611.400 ;
        RECT 757.950 612.600 760.050 613.050 ;
        RECT 775.950 612.600 778.050 613.050 ;
        RECT 757.950 611.400 778.050 612.600 ;
        RECT 757.950 610.950 760.050 611.400 ;
        RECT 775.950 610.950 778.050 611.400 ;
        RECT 598.950 608.400 648.600 609.600 ;
        RECT 700.950 609.600 703.050 610.050 ;
        RECT 715.950 609.600 718.050 610.050 ;
        RECT 700.950 608.400 718.050 609.600 ;
        RECT 598.950 607.950 601.050 608.400 ;
        RECT 616.950 607.950 619.050 608.400 ;
        RECT 700.950 607.950 703.050 608.400 ;
        RECT 715.950 607.950 718.050 608.400 ;
        RECT 403.950 606.000 436.050 606.600 ;
        RECT 403.950 605.400 435.600 606.000 ;
        RECT 341.400 603.600 342.600 605.100 ;
        RECT 403.950 604.950 406.050 605.400 ;
        RECT 430.950 604.950 433.050 605.400 ;
        RECT 296.400 602.400 312.600 603.600 ;
        RECT 265.950 598.950 268.050 601.050 ;
        RECT 280.950 600.600 283.050 601.050 ;
        RECT 292.950 600.600 295.050 601.050 ;
        RECT 280.950 599.400 295.050 600.600 ;
        RECT 311.400 600.600 312.600 602.400 ;
        RECT 326.400 602.400 342.600 603.600 ;
        RECT 439.950 603.600 442.050 607.050 ;
        RECT 445.950 603.600 448.050 604.050 ;
        RECT 452.400 603.900 453.600 607.950 ;
        RECT 439.950 603.000 448.050 603.600 ;
        RECT 440.400 602.400 448.050 603.000 ;
        RECT 326.400 600.900 327.600 602.400 ;
        RECT 445.950 601.950 448.050 602.400 ;
        RECT 451.950 601.800 454.050 603.900 ;
        RECT 478.800 602.100 480.900 604.200 ;
        RECT 524.400 604.050 525.600 607.950 ;
        RECT 481.950 603.600 484.050 604.050 ;
        RECT 514.950 603.600 517.050 604.050 ;
        RECT 481.950 602.400 517.050 603.600 ;
        RECT 311.400 599.400 315.600 600.600 ;
        RECT 280.950 598.950 283.050 599.400 ;
        RECT 292.950 598.950 295.050 599.400 ;
        RECT 82.950 597.600 85.050 598.050 ;
        RECT 91.950 597.600 94.050 598.050 ;
        RECT 82.950 596.400 94.050 597.600 ;
        RECT 82.950 595.950 85.050 596.400 ;
        RECT 91.950 595.950 94.050 596.400 ;
        RECT 100.950 595.950 103.050 598.050 ;
        RECT 112.950 597.600 115.050 598.050 ;
        RECT 127.950 597.600 130.050 598.050 ;
        RECT 196.950 597.600 199.050 598.050 ;
        RECT 112.950 596.400 199.050 597.600 ;
        RECT 251.400 596.400 256.050 598.050 ;
        RECT 112.950 595.950 115.050 596.400 ;
        RECT 127.950 595.950 130.050 596.400 ;
        RECT 196.950 595.950 199.050 596.400 ;
        RECT 252.000 595.950 256.050 596.400 ;
        RECT 262.950 597.600 265.050 598.050 ;
        RECT 274.950 597.600 277.050 597.900 ;
        RECT 262.950 596.400 277.050 597.600 ;
        RECT 262.950 595.950 265.050 596.400 ;
        RECT 274.950 595.800 277.050 596.400 ;
        RECT 286.950 597.600 289.050 598.050 ;
        RECT 298.950 597.600 301.050 598.050 ;
        RECT 286.950 596.400 301.050 597.600 ;
        RECT 314.400 597.600 315.600 599.400 ;
        RECT 325.950 598.800 328.050 600.900 ;
        RECT 391.950 600.600 394.050 600.900 ;
        RECT 400.950 600.600 403.050 601.050 ;
        RECT 391.950 599.400 403.050 600.600 ;
        RECT 391.950 598.800 394.050 599.400 ;
        RECT 400.950 598.950 403.050 599.400 ;
        RECT 406.950 600.600 409.050 600.900 ;
        RECT 421.950 600.600 424.050 601.050 ;
        RECT 406.950 599.400 424.050 600.600 ;
        RECT 406.950 598.800 409.050 599.400 ;
        RECT 421.950 598.950 424.050 599.400 ;
        RECT 454.950 600.600 457.050 601.050 ;
        RECT 479.400 600.600 480.600 602.100 ;
        RECT 481.950 601.950 484.050 602.400 ;
        RECT 514.950 601.950 517.050 602.400 ;
        RECT 523.950 601.950 526.050 604.050 ;
        RECT 601.950 603.600 604.050 607.050 ;
        RECT 622.950 604.950 625.050 607.050 ;
        RECT 640.950 606.600 643.050 607.200 ;
        RECT 629.400 605.400 643.050 606.600 ;
        RECT 593.400 603.000 604.050 603.600 ;
        RECT 593.400 602.400 603.600 603.000 ;
        RECT 454.950 599.400 480.600 600.600 ;
        RECT 520.950 600.600 523.050 601.050 ;
        RECT 526.950 600.600 529.050 601.050 ;
        RECT 520.950 599.400 529.050 600.600 ;
        RECT 454.950 598.950 457.050 599.400 ;
        RECT 520.950 598.950 523.050 599.400 ;
        RECT 526.950 598.950 529.050 599.400 ;
        RECT 568.950 600.600 571.050 601.050 ;
        RECT 580.950 600.600 583.050 601.050 ;
        RECT 568.950 599.400 583.050 600.600 ;
        RECT 568.950 598.950 571.050 599.400 ;
        RECT 580.950 598.950 583.050 599.400 ;
        RECT 586.950 600.600 589.050 601.050 ;
        RECT 593.400 600.600 594.600 602.400 ;
        RECT 586.950 599.400 594.600 600.600 ;
        RECT 595.950 600.600 598.050 600.900 ;
        RECT 623.400 600.600 624.600 604.950 ;
        RECT 629.400 601.050 630.600 605.400 ;
        RECT 640.950 605.100 643.050 605.400 ;
        RECT 649.950 606.750 652.050 607.200 ;
        RECT 658.950 606.750 661.050 607.200 ;
        RECT 649.950 605.550 661.050 606.750 ;
        RECT 649.950 605.100 652.050 605.550 ;
        RECT 658.950 605.100 661.050 605.550 ;
        RECT 673.950 606.600 676.050 607.050 ;
        RECT 682.950 606.600 685.050 607.050 ;
        RECT 673.950 605.400 685.050 606.600 ;
        RECT 673.950 604.950 676.050 605.400 ;
        RECT 682.950 604.950 685.050 605.400 ;
        RECT 688.950 605.100 691.050 607.200 ;
        RECT 706.950 606.600 709.050 607.200 ;
        RECT 724.950 606.600 727.050 607.200 ;
        RECT 706.950 605.400 727.050 606.600 ;
        RECT 706.950 605.100 709.050 605.400 ;
        RECT 724.950 605.100 727.050 605.400 ;
        RECT 739.950 606.600 742.050 607.200 ;
        RECT 769.950 606.600 772.050 607.200 ;
        RECT 739.950 605.400 772.050 606.600 ;
        RECT 739.950 605.100 742.050 605.400 ;
        RECT 769.950 605.100 772.050 605.400 ;
        RECT 793.950 605.100 796.050 607.200 ;
        RECT 823.950 606.750 826.050 607.200 ;
        RECT 829.950 606.750 832.050 607.200 ;
        RECT 823.950 605.550 832.050 606.750 ;
        RECT 823.950 605.100 826.050 605.550 ;
        RECT 829.950 605.100 832.050 605.550 ;
        RECT 838.950 605.100 841.050 607.200 ;
        RECT 880.950 606.750 883.050 607.200 ;
        RECT 895.950 606.750 898.050 607.200 ;
        RECT 880.950 605.550 898.050 606.750 ;
        RECT 880.950 605.100 883.050 605.550 ;
        RECT 895.950 605.100 898.050 605.550 ;
        RECT 901.950 606.750 904.050 607.200 ;
        RECT 913.950 606.750 916.050 607.200 ;
        RECT 901.950 605.550 916.050 606.750 ;
        RECT 901.950 605.100 904.050 605.550 ;
        RECT 913.950 605.100 916.050 605.550 ;
        RECT 689.400 603.600 690.600 605.100 ;
        RECT 689.400 602.400 699.600 603.600 ;
        RECT 595.950 599.400 624.600 600.600 ;
        RECT 586.950 598.950 589.050 599.400 ;
        RECT 595.950 598.800 598.050 599.400 ;
        RECT 628.950 598.950 631.050 601.050 ;
        RECT 637.950 600.600 640.050 600.900 ;
        RECT 649.950 600.600 652.050 601.050 ;
        RECT 637.950 599.400 652.050 600.600 ;
        RECT 637.950 598.800 640.050 599.400 ;
        RECT 649.950 598.950 652.050 599.400 ;
        RECT 685.950 600.600 688.050 600.900 ;
        RECT 694.950 600.600 697.050 601.050 ;
        RECT 685.950 599.400 697.050 600.600 ;
        RECT 698.400 600.600 699.600 602.400 ;
        RECT 703.950 600.600 706.050 600.900 ;
        RECT 698.400 599.400 706.050 600.600 ;
        RECT 685.950 598.800 688.050 599.400 ;
        RECT 694.950 598.950 697.050 599.400 ;
        RECT 703.950 598.800 706.050 599.400 ;
        RECT 721.950 600.600 724.050 600.900 ;
        RECT 748.950 600.600 751.050 601.050 ;
        RECT 721.950 599.400 751.050 600.600 ;
        RECT 721.950 598.800 724.050 599.400 ;
        RECT 748.950 598.950 751.050 599.400 ;
        RECT 763.950 600.600 766.050 601.050 ;
        RECT 772.950 600.600 775.050 600.900 ;
        RECT 763.950 599.400 775.050 600.600 ;
        RECT 763.950 598.950 766.050 599.400 ;
        RECT 772.950 598.800 775.050 599.400 ;
        RECT 322.950 597.600 325.050 598.050 ;
        RECT 314.400 596.400 325.050 597.600 ;
        RECT 286.950 595.950 289.050 596.400 ;
        RECT 298.950 595.950 301.050 596.400 ;
        RECT 322.950 595.950 325.050 596.400 ;
        RECT 331.950 597.600 334.050 598.050 ;
        RECT 346.950 597.600 349.050 598.050 ;
        RECT 355.950 597.600 358.050 598.050 ;
        RECT 331.950 596.400 358.050 597.600 ;
        RECT 331.950 595.950 334.050 596.400 ;
        RECT 346.950 595.950 349.050 596.400 ;
        RECT 355.950 595.950 358.050 596.400 ;
        RECT 607.950 597.600 610.050 598.050 ;
        RECT 616.950 597.600 619.050 598.050 ;
        RECT 607.950 596.400 619.050 597.600 ;
        RECT 607.950 595.950 610.050 596.400 ;
        RECT 616.950 595.950 619.050 596.400 ;
        RECT 634.950 597.600 637.050 598.050 ;
        RECT 670.950 597.600 673.050 598.050 ;
        RECT 634.950 596.400 673.050 597.600 ;
        RECT 634.950 595.950 637.050 596.400 ;
        RECT 670.950 595.950 673.050 596.400 ;
        RECT 784.950 597.600 787.050 598.050 ;
        RECT 794.400 597.600 795.600 605.100 ;
        RECT 839.400 601.050 840.600 605.100 ;
        RECT 870.000 603.600 874.050 604.050 ;
        RECT 802.950 600.600 805.050 600.900 ;
        RECT 811.950 600.600 814.050 601.050 ;
        RECT 802.950 599.400 814.050 600.600 ;
        RECT 802.950 598.800 805.050 599.400 ;
        RECT 811.950 598.950 814.050 599.400 ;
        RECT 835.950 599.400 840.600 601.050 ;
        RECT 869.400 601.950 874.050 603.600 ;
        RECT 847.950 600.600 850.050 600.900 ;
        RECT 869.400 600.600 870.600 601.950 ;
        RECT 847.950 599.400 870.600 600.600 ;
        RECT 889.950 600.450 892.050 600.900 ;
        RECT 910.950 600.450 913.050 600.900 ;
        RECT 835.950 598.950 840.000 599.400 ;
        RECT 847.950 598.800 850.050 599.400 ;
        RECT 889.950 599.250 913.050 600.450 ;
        RECT 889.950 598.800 892.050 599.250 ;
        RECT 910.950 598.800 913.050 599.250 ;
        RECT 784.950 596.400 795.600 597.600 ;
        RECT 823.950 597.600 826.050 598.050 ;
        RECT 829.950 597.600 832.050 598.050 ;
        RECT 841.950 597.600 844.050 598.050 ;
        RECT 823.950 596.400 844.050 597.600 ;
        RECT 784.950 595.950 787.050 596.400 ;
        RECT 823.950 595.950 826.050 596.400 ;
        RECT 829.950 595.950 832.050 596.400 ;
        RECT 841.950 595.950 844.050 596.400 ;
        RECT 865.950 597.600 868.050 598.050 ;
        RECT 901.950 597.600 904.050 598.050 ;
        RECT 865.950 596.400 904.050 597.600 ;
        RECT 40.950 594.600 43.050 595.050 ;
        RECT 46.950 594.600 49.050 595.050 ;
        RECT 40.950 593.400 49.050 594.600 ;
        RECT 40.950 592.950 43.050 593.400 ;
        RECT 46.950 592.950 49.050 593.400 ;
        RECT 103.950 594.600 106.050 595.050 ;
        RECT 115.950 594.600 118.050 595.050 ;
        RECT 124.950 594.600 127.050 595.050 ;
        RECT 103.950 593.400 127.050 594.600 ;
        RECT 103.950 592.950 106.050 593.400 ;
        RECT 115.950 592.950 118.050 593.400 ;
        RECT 124.950 592.950 127.050 593.400 ;
        RECT 157.950 594.600 160.050 595.050 ;
        RECT 163.950 594.600 166.050 595.050 ;
        RECT 157.950 593.400 166.050 594.600 ;
        RECT 157.950 592.950 160.050 593.400 ;
        RECT 163.950 592.950 166.050 593.400 ;
        RECT 181.950 594.600 184.050 595.050 ;
        RECT 193.950 594.600 196.050 595.050 ;
        RECT 181.950 593.400 196.050 594.600 ;
        RECT 181.950 592.950 184.050 593.400 ;
        RECT 193.950 592.950 196.050 593.400 ;
        RECT 199.950 594.600 202.050 595.050 ;
        RECT 208.950 594.600 211.050 595.050 ;
        RECT 199.950 593.400 211.050 594.600 ;
        RECT 199.950 592.950 202.050 593.400 ;
        RECT 208.950 592.950 211.050 593.400 ;
        RECT 217.950 594.600 220.050 595.050 ;
        RECT 244.950 594.600 247.050 595.050 ;
        RECT 217.950 593.400 247.050 594.600 ;
        RECT 217.950 592.950 220.050 593.400 ;
        RECT 244.950 592.950 247.050 593.400 ;
        RECT 343.950 594.600 346.050 595.050 ;
        RECT 397.950 594.600 400.050 595.050 ;
        RECT 427.950 594.600 430.050 595.050 ;
        RECT 343.950 593.400 400.050 594.600 ;
        RECT 343.950 592.950 346.050 593.400 ;
        RECT 397.950 592.950 400.050 593.400 ;
        RECT 416.400 593.400 430.050 594.600 ;
        RECT 10.950 591.600 13.050 592.050 ;
        RECT 22.950 591.600 25.050 592.050 ;
        RECT 43.950 591.600 46.050 592.050 ;
        RECT 61.950 591.600 64.050 592.050 ;
        RECT 10.950 590.400 39.600 591.600 ;
        RECT 10.950 589.950 13.050 590.400 ;
        RECT 22.950 589.950 25.050 590.400 ;
        RECT 38.400 588.600 39.600 590.400 ;
        RECT 43.950 590.400 64.050 591.600 ;
        RECT 43.950 589.950 46.050 590.400 ;
        RECT 61.950 589.950 64.050 590.400 ;
        RECT 250.950 591.600 253.050 592.050 ;
        RECT 259.950 591.600 262.050 592.050 ;
        RECT 250.950 590.400 262.050 591.600 ;
        RECT 250.950 589.950 253.050 590.400 ;
        RECT 259.950 589.950 262.050 590.400 ;
        RECT 322.950 591.600 325.050 592.050 ;
        RECT 349.950 591.600 352.050 592.050 ;
        RECT 416.400 591.600 417.600 593.400 ;
        RECT 427.950 592.950 430.050 593.400 ;
        RECT 589.950 594.600 592.050 595.050 ;
        RECT 601.950 594.600 604.050 595.050 ;
        RECT 589.950 593.400 604.050 594.600 ;
        RECT 589.950 592.950 592.050 593.400 ;
        RECT 601.950 592.950 604.050 593.400 ;
        RECT 625.950 594.600 628.050 595.050 ;
        RECT 652.950 594.600 655.050 595.050 ;
        RECT 625.950 593.400 655.050 594.600 ;
        RECT 625.950 592.950 628.050 593.400 ;
        RECT 652.950 592.950 655.050 593.400 ;
        RECT 661.950 594.600 664.050 595.050 ;
        RECT 673.950 594.600 676.050 595.050 ;
        RECT 697.950 594.600 700.050 595.050 ;
        RECT 661.950 593.400 700.050 594.600 ;
        RECT 661.950 592.950 664.050 593.400 ;
        RECT 673.950 592.950 676.050 593.400 ;
        RECT 697.950 592.950 700.050 593.400 ;
        RECT 724.950 594.600 727.050 595.050 ;
        RECT 736.950 594.600 739.050 595.050 ;
        RECT 724.950 593.400 739.050 594.600 ;
        RECT 724.950 592.950 727.050 593.400 ;
        RECT 736.950 592.950 739.050 593.400 ;
        RECT 754.950 594.600 757.050 595.050 ;
        RECT 796.950 594.600 799.050 595.050 ;
        RECT 814.950 594.600 817.050 595.050 ;
        RECT 754.950 593.400 817.050 594.600 ;
        RECT 754.950 592.950 757.050 593.400 ;
        RECT 796.950 592.950 799.050 593.400 ;
        RECT 814.950 592.950 817.050 593.400 ;
        RECT 847.950 594.600 850.050 595.050 ;
        RECT 865.950 594.600 868.050 596.400 ;
        RECT 901.950 595.950 904.050 596.400 ;
        RECT 847.950 594.000 868.050 594.600 ;
        RECT 847.950 593.400 867.600 594.000 ;
        RECT 847.950 592.950 850.050 593.400 ;
        RECT 322.950 590.400 417.600 591.600 ;
        RECT 433.950 591.600 436.050 592.050 ;
        RECT 454.950 591.600 457.050 592.050 ;
        RECT 586.950 591.600 589.050 592.050 ;
        RECT 433.950 590.400 457.050 591.600 ;
        RECT 322.950 589.950 325.050 590.400 ;
        RECT 349.950 589.950 352.050 590.400 ;
        RECT 433.950 589.950 436.050 590.400 ;
        RECT 454.950 589.950 457.050 590.400 ;
        RECT 578.400 590.400 589.050 591.600 ;
        RECT 602.400 591.600 603.600 592.950 ;
        RECT 631.950 591.600 634.050 592.050 ;
        RECT 602.400 590.400 634.050 591.600 ;
        RECT 55.950 588.600 58.050 589.050 ;
        RECT 38.400 587.400 58.050 588.600 ;
        RECT 55.950 586.950 58.050 587.400 ;
        RECT 76.950 588.600 79.050 589.050 ;
        RECT 106.950 588.600 109.050 589.050 ;
        RECT 151.950 588.600 154.050 589.050 ;
        RECT 76.950 587.400 109.050 588.600 ;
        RECT 76.950 586.950 79.050 587.400 ;
        RECT 106.950 586.950 109.050 587.400 ;
        RECT 110.400 587.400 154.050 588.600 ;
        RECT 64.950 585.600 67.050 586.050 ;
        RECT 88.800 585.600 90.900 586.050 ;
        RECT 64.950 584.400 90.900 585.600 ;
        RECT 64.950 583.950 67.050 584.400 ;
        RECT 88.800 583.950 90.900 584.400 ;
        RECT 91.950 585.600 94.050 586.050 ;
        RECT 110.400 585.600 111.600 587.400 ;
        RECT 151.950 586.950 154.050 587.400 ;
        RECT 181.950 588.600 184.050 589.050 ;
        RECT 211.950 588.600 214.050 589.050 ;
        RECT 181.950 587.400 214.050 588.600 ;
        RECT 181.950 586.950 184.050 587.400 ;
        RECT 211.950 586.950 214.050 587.400 ;
        RECT 313.950 588.600 316.050 589.050 ;
        RECT 349.950 588.600 352.050 588.900 ;
        RECT 313.950 587.400 352.050 588.600 ;
        RECT 313.950 586.950 316.050 587.400 ;
        RECT 349.950 586.800 352.050 587.400 ;
        RECT 418.950 588.600 421.050 589.050 ;
        RECT 427.950 588.600 430.050 589.050 ;
        RECT 418.950 587.400 430.050 588.600 ;
        RECT 418.950 586.950 421.050 587.400 ;
        RECT 427.950 586.950 430.050 587.400 ;
        RECT 457.950 588.600 460.050 589.050 ;
        RECT 466.950 588.600 469.050 589.050 ;
        RECT 457.950 587.400 469.050 588.600 ;
        RECT 457.950 586.950 460.050 587.400 ;
        RECT 466.950 586.950 469.050 587.400 ;
        RECT 523.950 588.600 526.050 589.050 ;
        RECT 544.950 588.600 547.050 589.050 ;
        RECT 523.950 587.400 547.050 588.600 ;
        RECT 523.950 586.950 526.050 587.400 ;
        RECT 544.950 586.950 547.050 587.400 ;
        RECT 559.950 588.600 562.050 589.050 ;
        RECT 578.400 588.600 579.600 590.400 ;
        RECT 586.950 589.950 589.050 590.400 ;
        RECT 631.950 589.950 634.050 590.400 ;
        RECT 706.950 591.600 709.050 592.050 ;
        RECT 721.950 591.600 724.050 592.050 ;
        RECT 706.950 590.400 724.050 591.600 ;
        RECT 706.950 589.950 709.050 590.400 ;
        RECT 721.950 589.950 724.050 590.400 ;
        RECT 856.950 591.600 859.050 592.050 ;
        RECT 865.950 591.600 868.050 591.900 ;
        RECT 856.950 590.400 868.050 591.600 ;
        RECT 856.950 589.950 859.050 590.400 ;
        RECT 865.950 589.800 868.050 590.400 ;
        RECT 559.950 587.400 579.600 588.600 ;
        RECT 598.950 588.600 601.050 589.050 ;
        RECT 613.950 588.600 616.050 589.050 ;
        RECT 598.950 587.400 616.050 588.600 ;
        RECT 559.950 586.950 562.050 587.400 ;
        RECT 598.950 586.950 601.050 587.400 ;
        RECT 613.950 586.950 616.050 587.400 ;
        RECT 730.950 588.600 733.050 589.050 ;
        RECT 850.950 588.600 853.050 589.050 ;
        RECT 730.950 587.400 853.050 588.600 ;
        RECT 730.950 586.950 733.050 587.400 ;
        RECT 850.950 586.950 853.050 587.400 ;
        RECT 862.950 588.600 865.050 589.050 ;
        RECT 892.950 588.600 895.050 589.050 ;
        RECT 862.950 587.400 895.050 588.600 ;
        RECT 862.950 586.950 865.050 587.400 ;
        RECT 892.950 586.950 895.050 587.400 ;
        RECT 91.950 584.400 111.600 585.600 ;
        RECT 154.950 585.600 157.050 586.050 ;
        RECT 235.950 585.600 238.050 586.050 ;
        RECT 154.950 584.400 238.050 585.600 ;
        RECT 91.950 583.950 94.050 584.400 ;
        RECT 154.950 583.950 157.050 584.400 ;
        RECT 235.950 583.950 238.050 584.400 ;
        RECT 259.950 585.600 262.050 586.050 ;
        RECT 277.950 585.600 280.050 586.050 ;
        RECT 259.950 584.400 280.050 585.600 ;
        RECT 259.950 583.950 262.050 584.400 ;
        RECT 277.950 583.950 280.050 584.400 ;
        RECT 364.950 585.600 367.050 586.050 ;
        RECT 400.950 585.600 403.050 586.050 ;
        RECT 364.950 584.400 403.050 585.600 ;
        RECT 364.950 583.950 367.050 584.400 ;
        RECT 400.950 583.950 403.050 584.400 ;
        RECT 442.950 585.600 447.000 586.050 ;
        RECT 442.950 583.950 447.600 585.600 ;
        RECT 85.950 582.600 88.050 583.050 ;
        RECT 97.950 582.600 100.050 583.050 ;
        RECT 115.950 582.600 118.050 583.050 ;
        RECT 151.950 582.600 154.050 583.050 ;
        RECT 85.950 581.400 154.050 582.600 ;
        RECT 85.950 580.950 88.050 581.400 ;
        RECT 97.950 580.950 100.050 581.400 ;
        RECT 115.950 580.950 118.050 581.400 ;
        RECT 151.950 580.950 154.050 581.400 ;
        RECT 211.950 582.600 214.050 583.050 ;
        RECT 226.950 582.600 229.050 583.050 ;
        RECT 211.950 581.400 229.050 582.600 ;
        RECT 211.950 580.950 214.050 581.400 ;
        RECT 226.950 580.950 229.050 581.400 ;
        RECT 238.950 582.600 241.050 583.050 ;
        RECT 295.950 582.600 298.050 583.050 ;
        RECT 238.950 581.400 298.050 582.600 ;
        RECT 446.400 582.600 447.600 583.950 ;
        RECT 454.950 582.600 457.050 583.050 ;
        RECT 463.950 582.600 466.050 583.050 ;
        RECT 446.400 581.400 466.050 582.600 ;
        RECT 511.950 582.600 514.050 586.050 ;
        RECT 614.400 585.600 615.600 586.950 ;
        RECT 643.950 585.600 646.050 586.050 ;
        RECT 661.950 585.600 664.050 586.050 ;
        RECT 614.400 584.400 664.050 585.600 ;
        RECT 643.950 583.950 646.050 584.400 ;
        RECT 661.950 583.950 664.050 584.400 ;
        RECT 853.950 585.600 856.050 586.050 ;
        RECT 883.950 585.600 886.050 586.050 ;
        RECT 853.950 584.400 886.050 585.600 ;
        RECT 853.950 583.950 856.050 584.400 ;
        RECT 883.950 583.950 886.050 584.400 ;
        RECT 565.950 582.600 568.050 583.050 ;
        RECT 511.950 582.000 568.050 582.600 ;
        RECT 512.400 581.400 568.050 582.000 ;
        RECT 238.950 580.950 241.050 581.400 ;
        RECT 295.950 580.950 298.050 581.400 ;
        RECT 454.950 580.950 457.050 581.400 ;
        RECT 463.950 580.950 466.050 581.400 ;
        RECT 565.950 580.950 568.050 581.400 ;
        RECT 619.950 582.600 622.050 583.050 ;
        RECT 628.950 582.600 631.050 583.050 ;
        RECT 619.950 581.400 631.050 582.600 ;
        RECT 619.950 580.950 622.050 581.400 ;
        RECT 628.950 580.950 631.050 581.400 ;
        RECT 667.950 582.600 670.050 583.050 ;
        RECT 694.950 582.600 697.050 583.050 ;
        RECT 667.950 581.400 697.050 582.600 ;
        RECT 667.950 580.950 670.050 581.400 ;
        RECT 694.950 580.950 697.050 581.400 ;
        RECT 820.950 582.600 823.050 583.050 ;
        RECT 844.950 582.600 847.050 583.050 ;
        RECT 820.950 581.400 847.050 582.600 ;
        RECT 820.950 580.950 823.050 581.400 ;
        RECT 844.950 580.950 847.050 581.400 ;
        RECT 859.950 582.600 862.050 583.050 ;
        RECT 877.950 582.600 880.050 583.050 ;
        RECT 859.950 581.400 880.050 582.600 ;
        RECT 859.950 580.950 862.050 581.400 ;
        RECT 877.950 580.950 880.050 581.400 ;
        RECT 895.950 582.600 898.050 583.050 ;
        RECT 916.950 582.600 919.050 583.050 ;
        RECT 895.950 581.400 919.050 582.600 ;
        RECT 895.950 580.950 898.050 581.400 ;
        RECT 916.950 580.950 919.050 581.400 ;
        RECT 58.950 579.600 61.050 580.050 ;
        RECT 82.950 579.600 85.050 580.050 ;
        RECT 88.950 579.600 91.050 580.050 ;
        RECT 58.950 578.400 91.050 579.600 ;
        RECT 58.950 577.950 61.050 578.400 ;
        RECT 82.950 577.950 85.050 578.400 ;
        RECT 88.950 577.950 91.050 578.400 ;
        RECT 106.950 579.600 109.050 580.050 ;
        RECT 148.950 579.600 151.050 580.050 ;
        RECT 106.950 578.400 151.050 579.600 ;
        RECT 106.950 577.950 109.050 578.400 ;
        RECT 148.950 577.950 151.050 578.400 ;
        RECT 172.950 579.600 175.050 580.050 ;
        RECT 232.800 579.600 234.900 580.050 ;
        RECT 172.950 578.400 234.900 579.600 ;
        RECT 172.950 577.950 175.050 578.400 ;
        RECT 232.800 577.950 234.900 578.400 ;
        RECT 235.950 579.600 238.050 580.050 ;
        RECT 274.950 579.600 277.050 580.050 ;
        RECT 235.950 578.400 277.050 579.600 ;
        RECT 235.950 577.950 238.050 578.400 ;
        RECT 274.950 577.950 277.050 578.400 ;
        RECT 304.950 579.600 307.050 580.050 ;
        RECT 310.950 579.600 313.050 580.050 ;
        RECT 304.950 578.400 313.050 579.600 ;
        RECT 304.950 577.950 307.050 578.400 ;
        RECT 310.950 577.950 313.050 578.400 ;
        RECT 334.950 579.600 337.050 580.050 ;
        RECT 340.950 579.600 343.050 580.050 ;
        RECT 334.950 578.400 343.050 579.600 ;
        RECT 334.950 577.950 337.050 578.400 ;
        RECT 340.950 577.950 343.050 578.400 ;
        RECT 406.950 579.600 409.050 580.050 ;
        RECT 421.950 579.600 424.050 580.050 ;
        RECT 433.950 579.600 436.050 580.050 ;
        RECT 406.950 578.400 436.050 579.600 ;
        RECT 406.950 577.950 409.050 578.400 ;
        RECT 421.950 577.950 424.050 578.400 ;
        RECT 433.950 577.950 436.050 578.400 ;
        RECT 538.950 579.600 541.050 580.050 ;
        RECT 559.950 579.600 562.050 580.050 ;
        RECT 538.950 578.400 562.050 579.600 ;
        RECT 538.950 577.950 541.050 578.400 ;
        RECT 559.950 577.950 562.050 578.400 ;
        RECT 913.950 579.600 916.050 580.050 ;
        RECT 919.950 579.600 922.050 580.050 ;
        RECT 913.950 578.400 922.050 579.600 ;
        RECT 913.950 577.950 916.050 578.400 ;
        RECT 919.950 577.950 922.050 578.400 ;
        RECT 931.950 579.600 934.050 580.050 ;
        RECT 943.950 579.600 946.050 580.050 ;
        RECT 931.950 578.400 946.050 579.600 ;
        RECT 931.950 577.950 934.050 578.400 ;
        RECT 943.950 577.950 946.050 578.400 ;
        RECT 52.950 576.600 55.050 577.050 ;
        RECT 76.950 576.600 79.050 577.050 ;
        RECT 82.950 576.600 85.050 576.900 ;
        RECT 52.950 575.400 85.050 576.600 ;
        RECT 52.950 574.950 55.050 575.400 ;
        RECT 76.950 574.950 79.050 575.400 ;
        RECT 82.950 574.800 85.050 575.400 ;
        RECT 151.950 576.600 154.050 577.050 ;
        RECT 181.950 576.600 184.050 577.050 ;
        RECT 151.950 575.400 184.050 576.600 ;
        RECT 151.950 574.950 154.050 575.400 ;
        RECT 181.950 574.950 184.050 575.400 ;
        RECT 391.950 576.600 394.050 577.050 ;
        RECT 415.950 576.600 418.050 577.050 ;
        RECT 391.950 575.400 418.050 576.600 ;
        RECT 391.950 574.950 394.050 575.400 ;
        RECT 415.950 574.950 418.050 575.400 ;
        RECT 439.950 576.600 442.050 577.050 ;
        RECT 472.950 576.600 475.050 577.050 ;
        RECT 439.950 575.400 475.050 576.600 ;
        RECT 439.950 574.950 442.050 575.400 ;
        RECT 472.950 574.950 475.050 575.400 ;
        RECT 565.950 576.600 568.050 577.050 ;
        RECT 625.950 576.600 628.050 577.050 ;
        RECT 565.950 575.400 628.050 576.600 ;
        RECT 565.950 574.950 568.050 575.400 ;
        RECT 625.950 574.950 628.050 575.400 ;
        RECT 676.950 576.600 679.050 577.050 ;
        RECT 685.950 576.600 688.050 577.050 ;
        RECT 676.950 575.400 688.050 576.600 ;
        RECT 676.950 574.950 679.050 575.400 ;
        RECT 685.950 574.950 688.050 575.400 ;
        RECT 883.950 576.600 886.050 577.050 ;
        RECT 889.950 576.600 892.050 577.050 ;
        RECT 883.950 575.400 892.050 576.600 ;
        RECT 883.950 574.950 886.050 575.400 ;
        RECT 889.950 574.950 892.050 575.400 ;
        RECT 904.950 576.600 907.050 577.050 ;
        RECT 922.950 576.600 925.050 577.050 ;
        RECT 904.950 575.400 925.050 576.600 ;
        RECT 904.950 574.950 907.050 575.400 ;
        RECT 922.950 574.950 925.050 575.400 ;
        RECT 31.950 573.600 34.050 574.200 ;
        RECT 31.950 572.400 39.450 573.600 ;
        RECT 31.950 572.100 34.050 572.400 ;
        RECT 38.250 568.050 39.450 572.400 ;
        RECT 64.800 571.950 66.900 574.050 ;
        RECT 70.950 573.750 73.050 574.200 ;
        RECT 94.950 573.750 97.050 574.200 ;
        RECT 70.950 572.550 97.050 573.750 ;
        RECT 70.950 572.100 73.050 572.550 ;
        RECT 94.950 572.100 97.050 572.550 ;
        RECT 112.950 571.950 115.050 574.050 ;
        RECT 142.950 573.600 145.050 574.050 ;
        RECT 163.950 573.600 166.050 574.200 ;
        RECT 196.950 573.600 199.050 573.900 ;
        RECT 205.950 573.600 208.050 574.200 ;
        RECT 142.950 572.400 162.600 573.600 ;
        RECT 142.950 571.950 145.050 572.400 ;
        RECT 4.950 567.450 7.050 567.900 ;
        RECT 13.950 567.450 16.050 567.900 ;
        RECT 4.950 566.250 16.050 567.450 ;
        RECT 4.950 565.800 7.050 566.250 ;
        RECT 13.950 565.800 16.050 566.250 ;
        RECT 22.950 567.600 25.050 568.050 ;
        RECT 28.950 567.600 31.050 567.900 ;
        RECT 22.950 566.400 31.050 567.600 ;
        RECT 22.950 565.950 25.050 566.400 ;
        RECT 28.950 565.800 31.050 566.400 ;
        RECT 37.800 565.950 39.900 568.050 ;
        RECT 40.950 567.600 43.050 568.050 ;
        RECT 55.950 567.600 58.050 567.900 ;
        RECT 40.950 566.400 58.050 567.600 ;
        RECT 40.950 565.950 43.050 566.400 ;
        RECT 55.950 565.800 58.050 566.400 ;
        RECT 61.950 567.600 64.050 567.900 ;
        RECT 65.250 567.600 66.450 571.950 ;
        RECT 113.400 568.050 114.600 571.950 ;
        RECT 61.950 566.400 66.450 567.600 ;
        RECT 85.950 567.450 88.050 567.900 ;
        RECT 97.950 567.450 100.050 567.900 ;
        RECT 61.950 565.800 64.050 566.400 ;
        RECT 85.950 566.250 100.050 567.450 ;
        RECT 85.950 565.800 88.050 566.250 ;
        RECT 97.950 565.800 100.050 566.250 ;
        RECT 112.950 565.950 115.050 568.050 ;
        RECT 127.950 567.600 130.050 567.900 ;
        RECT 148.950 567.600 151.050 567.900 ;
        RECT 127.950 567.450 151.050 567.600 ;
        RECT 154.950 567.450 157.050 567.900 ;
        RECT 127.950 566.400 157.050 567.450 ;
        RECT 161.400 567.600 162.600 572.400 ;
        RECT 163.950 572.400 171.600 573.600 ;
        RECT 163.950 572.100 166.050 572.400 ;
        RECT 166.950 567.600 169.050 568.050 ;
        RECT 161.400 566.400 169.050 567.600 ;
        RECT 170.400 567.600 171.600 572.400 ;
        RECT 196.950 572.400 208.050 573.600 ;
        RECT 196.950 571.800 199.050 572.400 ;
        RECT 205.950 572.100 208.050 572.400 ;
        RECT 223.950 573.600 226.050 574.050 ;
        RECT 271.950 573.600 274.050 574.050 ;
        RECT 223.950 572.400 274.050 573.600 ;
        RECT 223.950 571.950 226.050 572.400 ;
        RECT 271.950 571.950 274.050 572.400 ;
        RECT 310.950 571.950 313.050 574.050 ;
        RECT 424.950 571.950 427.050 574.050 ;
        RECT 478.950 573.600 481.050 574.050 ;
        RECT 517.950 573.600 520.050 574.050 ;
        RECT 478.950 572.400 520.050 573.600 ;
        RECT 478.950 571.950 481.050 572.400 ;
        RECT 517.950 571.950 520.050 572.400 ;
        RECT 535.950 573.600 538.050 574.050 ;
        RECT 550.950 573.600 553.050 574.200 ;
        RECT 571.950 573.600 574.050 574.200 ;
        RECT 535.950 572.400 553.050 573.600 ;
        RECT 535.950 571.950 538.050 572.400 ;
        RECT 550.950 572.100 553.050 572.400 ;
        RECT 554.400 572.400 574.050 573.600 ;
        RECT 311.400 568.050 312.600 571.950 ;
        RECT 313.950 570.750 316.050 571.200 ;
        RECT 334.950 570.750 337.050 571.200 ;
        RECT 313.950 569.550 337.050 570.750 ;
        RECT 313.950 569.100 316.050 569.550 ;
        RECT 334.950 569.100 337.050 569.550 ;
        RECT 370.950 570.600 373.050 570.900 ;
        RECT 391.950 570.600 394.050 571.050 ;
        RECT 370.950 569.400 394.050 570.600 ;
        RECT 370.950 568.800 373.050 569.400 ;
        RECT 391.950 568.950 394.050 569.400 ;
        RECT 170.400 566.400 183.600 567.600 ;
        RECT 127.950 565.800 130.050 566.400 ;
        RECT 148.950 566.250 157.050 566.400 ;
        RECT 148.950 565.800 151.050 566.250 ;
        RECT 154.950 565.800 157.050 566.250 ;
        RECT 166.950 565.950 169.050 566.400 ;
        RECT 34.950 564.600 37.050 565.050 ;
        RECT 43.950 564.600 46.050 565.050 ;
        RECT 34.950 563.400 46.050 564.600 ;
        RECT 182.400 564.600 183.600 566.400 ;
        RECT 190.950 567.450 193.050 567.900 ;
        RECT 196.800 567.450 198.900 567.900 ;
        RECT 190.950 566.250 198.900 567.450 ;
        RECT 190.950 565.800 193.050 566.250 ;
        RECT 196.800 565.800 198.900 566.250 ;
        RECT 199.950 567.600 202.050 568.050 ;
        RECT 208.950 567.600 211.050 567.900 ;
        RECT 199.950 566.400 211.050 567.600 ;
        RECT 199.950 565.950 202.050 566.400 ;
        RECT 208.950 565.800 211.050 566.400 ;
        RECT 220.950 567.450 223.050 567.900 ;
        RECT 229.950 567.450 232.050 567.900 ;
        RECT 220.950 566.250 232.050 567.450 ;
        RECT 220.950 565.800 223.050 566.250 ;
        RECT 229.950 565.800 232.050 566.250 ;
        RECT 250.950 567.600 253.050 568.050 ;
        RECT 256.950 567.600 259.050 568.050 ;
        RECT 250.950 566.400 259.050 567.600 ;
        RECT 250.950 565.950 253.050 566.400 ;
        RECT 256.950 565.950 259.050 566.400 ;
        RECT 274.950 567.450 277.050 567.900 ;
        RECT 283.950 567.450 286.050 567.900 ;
        RECT 274.950 566.250 286.050 567.450 ;
        RECT 274.950 565.800 277.050 566.250 ;
        RECT 283.950 565.800 286.050 566.250 ;
        RECT 310.950 565.950 313.050 568.050 ;
        RECT 322.950 567.600 325.050 567.900 ;
        RECT 340.950 567.600 343.050 568.050 ;
        RECT 322.950 566.400 343.050 567.600 ;
        RECT 322.950 565.800 325.050 566.400 ;
        RECT 340.950 565.950 343.050 566.400 ;
        RECT 400.950 567.450 403.050 568.050 ;
        RECT 412.950 567.450 415.050 567.900 ;
        RECT 400.950 566.250 415.050 567.450 ;
        RECT 425.400 567.600 426.600 571.950 ;
        RECT 430.950 567.600 433.050 568.050 ;
        RECT 425.400 566.400 433.050 567.600 ;
        RECT 400.950 565.950 403.050 566.250 ;
        RECT 412.950 565.800 415.050 566.250 ;
        RECT 430.950 565.950 433.050 566.400 ;
        RECT 457.950 567.600 460.050 567.900 ;
        RECT 466.950 567.600 469.050 571.050 ;
        RECT 472.950 570.450 475.050 570.900 ;
        RECT 493.950 570.450 496.050 570.900 ;
        RECT 472.950 569.250 496.050 570.450 ;
        RECT 472.950 568.800 475.050 569.250 ;
        RECT 493.950 568.800 496.050 569.250 ;
        RECT 535.950 567.600 538.050 568.050 ;
        RECT 554.400 567.900 555.600 572.400 ;
        RECT 571.950 572.100 574.050 572.400 ;
        RECT 589.950 572.100 592.050 574.200 ;
        RECT 631.950 572.100 634.050 574.200 ;
        RECT 637.950 573.750 640.050 574.200 ;
        RECT 643.950 573.750 646.050 574.200 ;
        RECT 637.950 572.550 646.050 573.750 ;
        RECT 637.950 572.100 640.050 572.550 ;
        RECT 643.950 572.100 646.050 572.550 ;
        RECT 580.950 570.600 583.050 571.050 ;
        RECT 590.400 570.600 591.600 572.100 ;
        RECT 632.400 570.600 633.600 572.100 ;
        RECT 679.950 571.950 682.050 574.050 ;
        RECT 733.950 573.600 736.050 574.200 ;
        RECT 745.950 573.600 748.050 574.050 ;
        RECT 760.950 573.600 763.050 574.050 ;
        RECT 733.950 572.400 763.050 573.600 ;
        RECT 733.950 572.100 736.050 572.400 ;
        RECT 745.950 571.950 748.050 572.400 ;
        RECT 760.950 571.950 763.050 572.400 ;
        RECT 775.950 573.600 778.050 574.200 ;
        RECT 793.950 573.600 796.050 574.200 ;
        RECT 775.950 572.400 796.050 573.600 ;
        RECT 775.950 572.100 778.050 572.400 ;
        RECT 793.950 572.100 796.050 572.400 ;
        RECT 826.950 573.750 829.050 574.200 ;
        RECT 856.950 573.750 859.050 574.200 ;
        RECT 826.950 572.550 859.050 573.750 ;
        RECT 826.950 572.100 829.050 572.550 ;
        RECT 856.950 572.100 859.050 572.550 ;
        RECT 580.950 569.400 591.600 570.600 ;
        RECT 620.400 569.400 633.600 570.600 ;
        RECT 580.950 568.950 583.050 569.400 ;
        RECT 457.950 567.000 469.050 567.600 ;
        RECT 518.400 567.000 538.050 567.600 ;
        RECT 457.950 566.400 468.600 567.000 ;
        RECT 517.950 566.400 538.050 567.000 ;
        RECT 457.950 565.800 460.050 566.400 ;
        RECT 193.950 564.600 196.050 565.050 ;
        RECT 182.400 563.400 196.050 564.600 ;
        RECT 34.950 562.950 37.050 563.400 ;
        RECT 43.950 562.950 46.050 563.400 ;
        RECT 193.950 562.950 196.050 563.400 ;
        RECT 316.950 564.600 319.050 565.050 ;
        RECT 322.950 564.600 325.050 564.750 ;
        RECT 316.950 563.400 325.050 564.600 ;
        RECT 316.950 562.950 319.050 563.400 ;
        RECT 322.950 562.650 325.050 563.400 ;
        RECT 397.950 564.600 400.050 565.050 ;
        RECT 406.950 564.600 409.050 564.900 ;
        RECT 397.950 563.400 409.050 564.600 ;
        RECT 397.950 562.950 400.050 563.400 ;
        RECT 406.950 562.800 409.050 563.400 ;
        RECT 418.950 564.600 421.050 565.050 ;
        RECT 427.950 564.600 430.050 565.050 ;
        RECT 418.950 563.400 430.050 564.600 ;
        RECT 418.950 562.950 421.050 563.400 ;
        RECT 427.950 562.950 430.050 563.400 ;
        RECT 517.950 562.950 520.050 566.400 ;
        RECT 535.950 565.950 538.050 566.400 ;
        RECT 553.950 565.800 556.050 567.900 ;
        RECT 562.950 567.450 565.050 567.900 ;
        RECT 574.950 567.450 577.050 567.900 ;
        RECT 562.950 566.250 577.050 567.450 ;
        RECT 562.950 565.800 565.050 566.250 ;
        RECT 574.950 565.800 577.050 566.250 ;
        RECT 595.950 567.600 598.050 568.050 ;
        RECT 620.400 567.600 621.600 569.400 ;
        RECT 595.950 566.400 621.600 567.600 ;
        RECT 622.950 567.600 625.050 568.050 ;
        RECT 628.950 567.600 631.050 567.900 ;
        RECT 622.950 566.400 631.050 567.600 ;
        RECT 595.950 565.950 598.050 566.400 ;
        RECT 622.950 565.950 625.050 566.400 ;
        RECT 628.950 565.800 631.050 566.400 ;
        RECT 646.950 567.600 649.050 567.900 ;
        RECT 664.950 567.600 667.050 567.900 ;
        RECT 646.950 566.400 667.050 567.600 ;
        RECT 646.950 565.800 649.050 566.400 ;
        RECT 664.950 565.800 667.050 566.400 ;
        RECT 670.950 567.450 673.050 567.900 ;
        RECT 676.950 567.450 679.050 567.900 ;
        RECT 670.950 566.250 679.050 567.450 ;
        RECT 680.400 567.600 681.600 571.950 ;
        RECT 763.950 570.600 766.050 571.050 ;
        RECT 776.400 570.600 777.600 572.100 ;
        RECT 865.950 571.950 868.050 574.050 ;
        RECT 892.950 573.750 895.050 574.200 ;
        RECT 898.950 573.750 901.050 574.200 ;
        RECT 892.950 572.550 901.050 573.750 ;
        RECT 892.950 572.100 895.050 572.550 ;
        RECT 898.950 572.100 901.050 572.550 ;
        RECT 913.950 573.600 918.000 574.050 ;
        RECT 922.950 573.750 925.050 574.200 ;
        RECT 934.800 573.750 936.900 574.200 ;
        RECT 913.950 571.950 918.600 573.600 ;
        RECT 922.950 572.550 936.900 573.750 ;
        RECT 922.950 572.100 925.050 572.550 ;
        RECT 934.800 572.100 936.900 572.550 ;
        RECT 763.950 569.400 777.600 570.600 ;
        RECT 763.950 568.950 766.050 569.400 ;
        RECT 715.950 567.600 718.050 567.900 ;
        RECT 730.950 567.600 733.050 567.900 ;
        RECT 680.400 566.400 733.050 567.600 ;
        RECT 670.950 565.800 673.050 566.250 ;
        RECT 676.950 565.800 679.050 566.250 ;
        RECT 715.950 565.800 718.050 566.400 ;
        RECT 730.950 565.800 733.050 566.400 ;
        RECT 745.950 567.450 748.050 567.900 ;
        RECT 751.950 567.450 754.050 567.900 ;
        RECT 745.950 566.250 754.050 567.450 ;
        RECT 745.950 565.800 748.050 566.250 ;
        RECT 751.950 565.800 754.050 566.250 ;
        RECT 772.950 567.600 775.050 567.900 ;
        RECT 781.950 567.600 784.050 568.050 ;
        RECT 772.950 566.400 784.050 567.600 ;
        RECT 772.950 565.800 775.050 566.400 ;
        RECT 781.950 565.950 784.050 566.400 ;
        RECT 838.950 567.600 841.050 567.900 ;
        RECT 853.950 567.600 856.050 567.900 ;
        RECT 838.950 566.400 856.050 567.600 ;
        RECT 866.400 567.600 867.600 571.950 ;
        RECT 871.950 567.600 874.050 568.050 ;
        RECT 866.400 566.400 874.050 567.600 ;
        RECT 838.950 565.800 841.050 566.400 ;
        RECT 853.950 565.800 856.050 566.400 ;
        RECT 871.950 565.950 874.050 566.400 ;
        RECT 880.950 567.600 883.050 567.900 ;
        RECT 901.950 567.600 904.050 567.900 ;
        RECT 880.950 566.400 904.050 567.600 ;
        RECT 917.400 567.600 918.600 571.950 ;
        RECT 937.950 570.600 940.050 574.050 ;
        RECT 937.950 570.000 945.600 570.600 ;
        RECT 938.400 569.400 945.600 570.000 ;
        RECT 944.400 568.050 945.600 569.400 ;
        RECT 919.950 567.600 922.050 567.900 ;
        RECT 917.400 566.400 922.050 567.600 ;
        RECT 880.950 565.800 883.050 566.400 ;
        RECT 901.950 565.800 904.050 566.400 ;
        RECT 919.950 565.800 922.050 566.400 ;
        RECT 934.950 567.600 937.050 568.050 ;
        RECT 940.950 567.600 943.050 567.900 ;
        RECT 934.950 566.400 943.050 567.600 ;
        RECT 944.400 566.400 949.050 568.050 ;
        RECT 934.950 565.950 937.050 566.400 ;
        RECT 940.950 565.800 943.050 566.400 ;
        RECT 945.000 565.950 949.050 566.400 ;
        RECT 547.950 564.600 550.050 565.050 ;
        RECT 563.400 564.600 564.600 565.800 ;
        RECT 547.950 563.400 564.600 564.600 ;
        RECT 757.950 564.600 760.050 565.050 ;
        RECT 763.950 564.600 766.050 565.050 ;
        RECT 769.950 564.600 772.050 565.050 ;
        RECT 757.950 563.400 772.050 564.600 ;
        RECT 547.950 562.950 550.050 563.400 ;
        RECT 757.950 562.950 760.050 563.400 ;
        RECT 763.950 562.950 766.050 563.400 ;
        RECT 769.950 562.950 772.050 563.400 ;
        RECT 337.950 561.600 340.050 562.050 ;
        RECT 469.950 561.600 472.050 562.050 ;
        RECT 337.950 560.400 472.050 561.600 ;
        RECT 337.950 559.950 340.050 560.400 ;
        RECT 469.950 559.950 472.050 560.400 ;
        RECT 475.950 561.600 478.050 562.050 ;
        RECT 532.950 561.600 535.050 562.050 ;
        RECT 592.950 561.600 595.050 562.050 ;
        RECT 598.950 561.600 601.050 562.050 ;
        RECT 475.950 560.400 549.600 561.600 ;
        RECT 475.950 559.950 478.050 560.400 ;
        RECT 532.950 559.950 535.050 560.400 ;
        RECT 61.950 558.600 64.050 559.050 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 115.950 558.600 118.050 559.050 ;
        RECT 61.950 557.400 81.600 558.600 ;
        RECT 61.950 556.950 64.050 557.400 ;
        RECT 80.400 556.050 81.600 557.400 ;
        RECT 88.950 557.400 118.050 558.600 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 115.950 556.950 118.050 557.400 ;
        RECT 139.950 558.600 142.050 559.050 ;
        RECT 160.950 558.600 163.050 559.050 ;
        RECT 139.950 557.400 163.050 558.600 ;
        RECT 139.950 556.950 142.050 557.400 ;
        RECT 160.950 556.950 163.050 557.400 ;
        RECT 178.950 558.600 181.050 559.050 ;
        RECT 187.800 558.600 189.900 559.050 ;
        RECT 178.950 557.400 189.900 558.600 ;
        RECT 178.950 556.950 181.050 557.400 ;
        RECT 187.800 556.950 189.900 557.400 ;
        RECT 190.950 558.600 193.050 559.050 ;
        RECT 220.950 558.600 223.050 559.050 ;
        RECT 190.950 557.400 223.050 558.600 ;
        RECT 190.950 556.950 193.050 557.400 ;
        RECT 220.950 556.950 223.050 557.400 ;
        RECT 229.950 558.600 232.050 559.050 ;
        RECT 286.950 558.600 289.050 559.050 ;
        RECT 229.950 557.400 289.050 558.600 ;
        RECT 229.950 556.950 232.050 557.400 ;
        RECT 286.950 556.950 289.050 557.400 ;
        RECT 295.950 558.600 298.050 559.050 ;
        RECT 316.950 558.600 319.050 559.050 ;
        RECT 295.950 557.400 319.050 558.600 ;
        RECT 295.950 556.950 298.050 557.400 ;
        RECT 316.950 556.950 319.050 557.400 ;
        RECT 406.950 558.600 409.050 559.050 ;
        RECT 424.950 558.600 427.050 559.050 ;
        RECT 406.950 557.400 427.050 558.600 ;
        RECT 406.950 556.950 409.050 557.400 ;
        RECT 424.950 556.950 427.050 557.400 ;
        RECT 451.950 558.600 454.050 559.050 ;
        RECT 466.950 558.600 469.050 559.050 ;
        RECT 451.950 557.400 469.050 558.600 ;
        RECT 451.950 556.950 454.050 557.400 ;
        RECT 466.950 556.950 469.050 557.400 ;
        RECT 472.950 558.600 475.050 559.050 ;
        RECT 538.950 558.600 541.050 559.050 ;
        RECT 472.950 557.400 541.050 558.600 ;
        RECT 548.400 558.600 549.600 560.400 ;
        RECT 592.950 560.400 601.050 561.600 ;
        RECT 592.950 559.950 595.050 560.400 ;
        RECT 598.950 559.950 601.050 560.400 ;
        RECT 613.950 561.600 616.050 562.050 ;
        RECT 655.950 561.600 658.050 562.050 ;
        RECT 613.950 560.400 658.050 561.600 ;
        RECT 613.950 559.950 616.050 560.400 ;
        RECT 655.950 559.950 658.050 560.400 ;
        RECT 859.950 561.600 862.050 561.900 ;
        RECT 868.950 561.600 871.050 562.050 ;
        RECT 859.950 560.400 871.050 561.600 ;
        RECT 859.950 559.800 862.050 560.400 ;
        RECT 868.950 559.950 871.050 560.400 ;
        RECT 889.950 561.600 892.050 562.050 ;
        RECT 907.950 561.600 910.050 562.050 ;
        RECT 889.950 560.400 910.050 561.600 ;
        RECT 889.950 559.950 892.050 560.400 ;
        RECT 907.950 559.950 910.050 560.400 ;
        RECT 583.950 558.600 586.050 559.050 ;
        RECT 548.400 557.400 586.050 558.600 ;
        RECT 472.950 556.950 475.050 557.400 ;
        RECT 538.950 556.950 541.050 557.400 ;
        RECT 583.950 556.950 586.050 557.400 ;
        RECT 706.950 558.600 709.050 559.050 ;
        RECT 718.950 558.600 721.050 559.050 ;
        RECT 706.950 557.400 721.050 558.600 ;
        RECT 706.950 556.950 709.050 557.400 ;
        RECT 718.950 556.950 721.050 557.400 ;
        RECT 751.950 558.600 754.050 559.050 ;
        RECT 790.950 558.600 793.050 559.050 ;
        RECT 751.950 557.400 793.050 558.600 ;
        RECT 751.950 556.950 754.050 557.400 ;
        RECT 790.950 556.950 793.050 557.400 ;
        RECT 79.950 555.600 82.050 556.050 ;
        RECT 136.950 555.600 139.050 556.050 ;
        RECT 79.950 554.400 139.050 555.600 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 136.950 553.950 139.050 554.400 ;
        RECT 193.950 555.600 196.050 556.050 ;
        RECT 223.950 555.600 226.050 555.900 ;
        RECT 262.950 555.600 265.050 556.050 ;
        RECT 289.950 555.600 292.050 556.050 ;
        RECT 193.950 554.400 213.600 555.600 ;
        RECT 193.950 553.950 196.050 554.400 ;
        RECT 212.400 553.050 213.600 554.400 ;
        RECT 223.950 554.400 292.050 555.600 ;
        RECT 223.950 553.800 226.050 554.400 ;
        RECT 262.950 553.950 265.050 554.400 ;
        RECT 289.950 553.950 292.050 554.400 ;
        RECT 415.950 555.600 418.050 556.050 ;
        RECT 430.950 555.600 433.050 556.050 ;
        RECT 415.950 554.400 433.050 555.600 ;
        RECT 415.950 553.950 418.050 554.400 ;
        RECT 430.950 553.950 433.050 554.400 ;
        RECT 448.950 555.600 451.050 556.050 ;
        RECT 604.950 555.600 607.050 556.050 ;
        RECT 748.950 555.600 751.050 556.050 ;
        RECT 448.950 554.400 600.600 555.600 ;
        RECT 448.950 553.950 451.050 554.400 ;
        RECT 599.400 553.050 600.600 554.400 ;
        RECT 604.950 554.400 751.050 555.600 ;
        RECT 604.950 553.950 607.050 554.400 ;
        RECT 748.950 553.950 751.050 554.400 ;
        RECT 793.950 555.600 796.050 556.050 ;
        RECT 838.950 555.600 841.050 556.050 ;
        RECT 793.950 554.400 841.050 555.600 ;
        RECT 793.950 553.950 796.050 554.400 ;
        RECT 838.950 553.950 841.050 554.400 ;
        RECT 847.950 555.600 850.050 556.050 ;
        RECT 862.950 555.600 865.050 556.050 ;
        RECT 847.950 554.400 865.050 555.600 ;
        RECT 847.950 553.950 850.050 554.400 ;
        RECT 862.950 553.950 865.050 554.400 ;
        RECT 892.950 555.600 895.050 556.050 ;
        RECT 928.950 555.600 931.050 556.050 ;
        RECT 892.950 554.400 931.050 555.600 ;
        RECT 892.950 553.950 895.050 554.400 ;
        RECT 928.950 553.950 931.050 554.400 ;
        RECT 106.950 552.600 109.050 553.050 ;
        RECT 124.950 552.600 127.050 553.050 ;
        RECT 106.950 551.400 127.050 552.600 ;
        RECT 106.950 550.950 109.050 551.400 ;
        RECT 124.950 550.950 127.050 551.400 ;
        RECT 130.950 552.600 133.050 553.050 ;
        RECT 169.950 552.600 172.050 553.050 ;
        RECT 130.950 551.400 172.050 552.600 ;
        RECT 130.950 550.950 133.050 551.400 ;
        RECT 169.950 550.950 172.050 551.400 ;
        RECT 211.950 552.600 214.050 553.050 ;
        RECT 232.950 552.600 235.050 553.050 ;
        RECT 211.950 551.400 235.050 552.600 ;
        RECT 211.950 550.950 214.050 551.400 ;
        RECT 232.950 550.950 235.050 551.400 ;
        RECT 286.950 552.600 289.050 553.050 ;
        RECT 292.950 552.600 295.050 553.050 ;
        RECT 286.950 551.400 295.050 552.600 ;
        RECT 286.950 550.950 289.050 551.400 ;
        RECT 292.950 550.950 295.050 551.400 ;
        RECT 307.950 552.600 310.050 553.050 ;
        RECT 397.950 552.600 400.050 553.050 ;
        RECT 307.950 551.400 400.050 552.600 ;
        RECT 307.950 550.950 310.050 551.400 ;
        RECT 397.950 550.950 400.050 551.400 ;
        RECT 406.950 552.600 409.050 553.050 ;
        RECT 436.950 552.600 439.050 553.050 ;
        RECT 406.950 551.400 439.050 552.600 ;
        RECT 406.950 550.950 409.050 551.400 ;
        RECT 436.950 550.950 439.050 551.400 ;
        RECT 466.950 552.600 469.050 553.050 ;
        RECT 493.950 552.600 496.050 553.050 ;
        RECT 466.950 551.400 496.050 552.600 ;
        RECT 466.950 550.950 469.050 551.400 ;
        RECT 493.950 550.950 496.050 551.400 ;
        RECT 523.950 552.600 526.050 553.050 ;
        RECT 547.950 552.600 550.050 553.050 ;
        RECT 523.950 551.400 550.050 552.600 ;
        RECT 523.950 550.950 526.050 551.400 ;
        RECT 547.950 550.950 550.050 551.400 ;
        RECT 562.950 552.600 565.050 553.050 ;
        RECT 589.950 552.600 592.050 553.050 ;
        RECT 562.950 551.400 592.050 552.600 ;
        RECT 562.950 550.950 565.050 551.400 ;
        RECT 589.950 550.950 592.050 551.400 ;
        RECT 598.950 552.600 601.050 553.050 ;
        RECT 637.800 552.600 639.900 553.050 ;
        RECT 598.950 551.400 639.900 552.600 ;
        RECT 598.950 550.950 601.050 551.400 ;
        RECT 637.800 550.950 639.900 551.400 ;
        RECT 640.950 552.600 643.050 553.050 ;
        RECT 682.950 552.600 685.050 553.050 ;
        RECT 640.950 551.400 685.050 552.600 ;
        RECT 640.950 550.950 643.050 551.400 ;
        RECT 682.950 550.950 685.050 551.400 ;
        RECT 694.950 552.600 697.050 553.050 ;
        RECT 736.950 552.600 739.050 553.050 ;
        RECT 694.950 551.400 739.050 552.600 ;
        RECT 694.950 550.950 697.050 551.400 ;
        RECT 736.950 550.950 739.050 551.400 ;
        RECT 277.950 549.600 280.050 550.050 ;
        RECT 295.950 549.600 298.050 550.050 ;
        RECT 277.950 548.400 298.050 549.600 ;
        RECT 277.950 547.950 280.050 548.400 ;
        RECT 295.950 547.950 298.050 548.400 ;
        RECT 403.950 549.600 406.050 550.050 ;
        RECT 442.950 549.600 445.050 550.050 ;
        RECT 403.950 548.400 445.050 549.600 ;
        RECT 403.950 547.950 406.050 548.400 ;
        RECT 442.950 547.950 445.050 548.400 ;
        RECT 487.950 549.600 490.050 550.050 ;
        RECT 514.950 549.600 517.050 550.050 ;
        RECT 487.950 548.400 517.050 549.600 ;
        RECT 487.950 547.950 490.050 548.400 ;
        RECT 514.950 547.950 517.050 548.400 ;
        RECT 556.950 549.600 559.050 550.050 ;
        RECT 616.950 549.600 619.050 550.050 ;
        RECT 556.950 548.400 619.050 549.600 ;
        RECT 556.950 547.950 559.050 548.400 ;
        RECT 616.950 547.950 619.050 548.400 ;
        RECT 688.950 549.600 691.050 550.050 ;
        RECT 694.950 549.600 697.050 549.900 ;
        RECT 688.950 548.400 697.050 549.600 ;
        RECT 688.950 547.950 691.050 548.400 ;
        RECT 694.950 547.800 697.050 548.400 ;
        RECT 703.950 549.600 706.050 550.050 ;
        RECT 730.950 549.600 733.050 550.050 ;
        RECT 703.950 548.400 733.050 549.600 ;
        RECT 703.950 547.950 706.050 548.400 ;
        RECT 730.950 547.950 733.050 548.400 ;
        RECT 766.950 549.600 769.050 550.050 ;
        RECT 844.950 549.600 847.050 550.050 ;
        RECT 766.950 548.400 847.050 549.600 ;
        RECT 766.950 547.950 769.050 548.400 ;
        RECT 844.950 547.950 847.050 548.400 ;
        RECT 925.950 549.600 928.050 550.050 ;
        RECT 931.950 549.600 934.050 550.050 ;
        RECT 925.950 548.400 934.050 549.600 ;
        RECT 925.950 547.950 928.050 548.400 ;
        RECT 931.950 547.950 934.050 548.400 ;
        RECT 4.950 546.600 7.050 547.050 ;
        RECT 64.950 546.600 67.050 547.050 ;
        RECT 4.950 545.400 67.050 546.600 ;
        RECT 4.950 544.950 7.050 545.400 ;
        RECT 64.950 544.950 67.050 545.400 ;
        RECT 73.950 546.600 76.050 547.050 ;
        RECT 103.950 546.600 106.050 547.050 ;
        RECT 73.950 545.400 106.050 546.600 ;
        RECT 73.950 544.950 76.050 545.400 ;
        RECT 103.950 544.950 106.050 545.400 ;
        RECT 118.950 546.600 121.050 547.050 ;
        RECT 208.950 546.600 211.050 547.050 ;
        RECT 247.950 546.600 250.050 547.050 ;
        RECT 118.950 545.400 250.050 546.600 ;
        RECT 118.950 544.950 121.050 545.400 ;
        RECT 208.950 544.950 211.050 545.400 ;
        RECT 247.950 544.950 250.050 545.400 ;
        RECT 280.950 546.600 283.050 547.050 ;
        RECT 385.950 546.600 388.050 547.050 ;
        RECT 400.950 546.600 403.050 547.050 ;
        RECT 280.950 545.400 403.050 546.600 ;
        RECT 280.950 544.950 283.050 545.400 ;
        RECT 385.950 544.950 388.050 545.400 ;
        RECT 400.950 544.950 403.050 545.400 ;
        RECT 430.950 546.600 433.050 547.050 ;
        RECT 472.950 546.600 475.050 547.050 ;
        RECT 430.950 545.400 475.050 546.600 ;
        RECT 430.950 544.950 433.050 545.400 ;
        RECT 472.950 544.950 475.050 545.400 ;
        RECT 46.950 543.600 49.050 544.050 ;
        RECT 100.950 543.600 103.050 544.050 ;
        RECT 178.950 543.600 181.050 544.050 ;
        RECT 46.950 542.400 103.050 543.600 ;
        RECT 46.950 541.950 49.050 542.400 ;
        RECT 100.950 541.950 103.050 542.400 ;
        RECT 143.400 542.400 181.050 543.600 ;
        RECT 49.950 540.600 52.050 541.050 ;
        RECT 112.950 540.600 115.050 541.050 ;
        RECT 124.950 540.600 127.050 541.050 ;
        RECT 49.950 539.400 96.600 540.600 ;
        RECT 49.950 538.950 52.050 539.400 ;
        RECT 67.950 537.600 70.050 538.050 ;
        RECT 79.950 537.600 82.050 538.050 ;
        RECT 67.950 536.400 82.050 537.600 ;
        RECT 95.400 537.600 96.600 539.400 ;
        RECT 112.950 539.400 127.050 540.600 ;
        RECT 112.950 538.950 115.050 539.400 ;
        RECT 124.950 538.950 127.050 539.400 ;
        RECT 136.950 540.600 139.050 541.050 ;
        RECT 143.400 540.600 144.600 542.400 ;
        RECT 178.950 541.950 181.050 542.400 ;
        RECT 202.950 543.600 205.050 544.050 ;
        RECT 235.950 543.600 238.050 544.050 ;
        RECT 202.950 542.400 238.050 543.600 ;
        RECT 202.950 541.950 205.050 542.400 ;
        RECT 235.950 541.950 238.050 542.400 ;
        RECT 292.950 543.600 295.050 544.050 ;
        RECT 385.950 543.600 388.050 543.900 ;
        RECT 292.950 542.400 388.050 543.600 ;
        RECT 292.950 541.950 295.050 542.400 ;
        RECT 385.950 541.800 388.050 542.400 ;
        RECT 412.950 543.600 415.050 544.050 ;
        RECT 418.950 543.600 421.050 544.050 ;
        RECT 412.950 542.400 421.050 543.600 ;
        RECT 412.950 541.950 415.050 542.400 ;
        RECT 418.950 541.950 421.050 542.400 ;
        RECT 433.950 543.600 436.050 544.050 ;
        RECT 454.950 543.600 457.050 544.050 ;
        RECT 433.950 542.400 457.050 543.600 ;
        RECT 433.950 541.950 436.050 542.400 ;
        RECT 454.950 541.950 457.050 542.400 ;
        RECT 502.950 543.600 505.050 544.050 ;
        RECT 523.950 543.600 526.050 544.050 ;
        RECT 502.950 542.400 526.050 543.600 ;
        RECT 502.950 541.950 505.050 542.400 ;
        RECT 523.950 541.950 526.050 542.400 ;
        RECT 601.950 543.600 604.050 544.050 ;
        RECT 643.950 543.600 646.050 544.050 ;
        RECT 601.950 542.400 646.050 543.600 ;
        RECT 601.950 541.950 604.050 542.400 ;
        RECT 643.950 541.950 646.050 542.400 ;
        RECT 724.950 543.600 727.050 544.050 ;
        RECT 784.950 543.600 787.050 544.050 ;
        RECT 811.950 543.600 814.050 544.050 ;
        RECT 724.950 542.400 814.050 543.600 ;
        RECT 724.950 541.950 727.050 542.400 ;
        RECT 784.950 541.950 787.050 542.400 ;
        RECT 811.950 541.950 814.050 542.400 ;
        RECT 136.950 539.400 144.600 540.600 ;
        RECT 148.950 540.600 151.050 541.050 ;
        RECT 184.950 540.600 187.050 541.050 ;
        RECT 196.950 540.600 199.050 541.050 ;
        RECT 148.950 539.400 199.050 540.600 ;
        RECT 136.950 538.950 139.050 539.400 ;
        RECT 148.950 538.950 151.050 539.400 ;
        RECT 184.950 538.950 187.050 539.400 ;
        RECT 196.950 538.950 199.050 539.400 ;
        RECT 268.950 540.600 271.050 541.050 ;
        RECT 289.950 540.600 292.050 541.050 ;
        RECT 268.950 539.400 292.050 540.600 ;
        RECT 268.950 538.950 271.050 539.400 ;
        RECT 289.950 538.950 292.050 539.400 ;
        RECT 424.950 540.600 427.050 541.050 ;
        RECT 451.950 540.600 454.050 541.050 ;
        RECT 424.950 539.400 454.050 540.600 ;
        RECT 424.950 538.950 427.050 539.400 ;
        RECT 451.950 538.950 454.050 539.400 ;
        RECT 469.950 540.600 472.050 541.050 ;
        RECT 490.950 540.600 493.050 541.050 ;
        RECT 469.950 539.400 493.050 540.600 ;
        RECT 469.950 538.950 472.050 539.400 ;
        RECT 490.950 538.950 493.050 539.400 ;
        RECT 106.950 537.600 109.050 538.050 ;
        RECT 95.400 536.400 109.050 537.600 ;
        RECT 67.950 535.950 70.050 536.400 ;
        RECT 79.950 535.950 82.050 536.400 ;
        RECT 106.950 535.950 109.050 536.400 ;
        RECT 160.950 537.600 163.050 538.050 ;
        RECT 202.950 537.600 205.050 538.050 ;
        RECT 160.950 536.400 205.050 537.600 ;
        RECT 160.950 535.950 163.050 536.400 ;
        RECT 202.950 535.950 205.050 536.400 ;
        RECT 331.950 537.600 334.050 538.050 ;
        RECT 349.950 537.600 352.050 538.050 ;
        RECT 331.950 536.400 352.050 537.600 ;
        RECT 331.950 535.950 334.050 536.400 ;
        RECT 349.950 535.950 352.050 536.400 ;
        RECT 409.950 537.600 412.050 538.050 ;
        RECT 448.950 537.600 451.050 538.050 ;
        RECT 409.950 536.400 451.050 537.600 ;
        RECT 409.950 535.950 412.050 536.400 ;
        RECT 448.950 535.950 451.050 536.400 ;
        RECT 550.950 537.600 553.050 538.050 ;
        RECT 568.950 537.600 571.050 538.050 ;
        RECT 550.950 536.400 571.050 537.600 ;
        RECT 550.950 535.950 553.050 536.400 ;
        RECT 568.950 535.950 571.050 536.400 ;
        RECT 619.950 537.600 622.050 538.050 ;
        RECT 664.950 537.600 667.050 538.050 ;
        RECT 619.950 536.400 667.050 537.600 ;
        RECT 619.950 535.950 622.050 536.400 ;
        RECT 664.950 535.950 667.050 536.400 ;
        RECT 91.950 534.600 94.050 535.050 ;
        RECT 106.950 534.600 109.050 534.900 ;
        RECT 91.950 533.400 109.050 534.600 ;
        RECT 91.950 532.950 94.050 533.400 ;
        RECT 106.950 532.800 109.050 533.400 ;
        RECT 115.950 534.600 118.050 535.050 ;
        RECT 145.950 534.600 148.050 535.050 ;
        RECT 115.950 533.400 148.050 534.600 ;
        RECT 115.950 532.950 118.050 533.400 ;
        RECT 145.950 532.950 148.050 533.400 ;
        RECT 154.950 534.600 157.050 535.050 ;
        RECT 205.950 534.600 208.050 535.050 ;
        RECT 154.950 533.400 208.050 534.600 ;
        RECT 154.950 532.950 157.050 533.400 ;
        RECT 205.950 532.950 208.050 533.400 ;
        RECT 412.950 534.600 415.050 535.050 ;
        RECT 430.950 534.600 433.050 535.050 ;
        RECT 475.950 534.600 478.050 535.050 ;
        RECT 412.950 533.400 433.050 534.600 ;
        RECT 412.950 532.950 415.050 533.400 ;
        RECT 430.950 532.950 433.050 533.400 ;
        RECT 434.400 533.400 478.050 534.600 ;
        RECT 19.950 531.600 22.050 532.050 ;
        RECT 64.950 531.600 67.050 532.050 ;
        RECT 73.950 531.600 76.050 532.050 ;
        RECT 19.950 530.400 76.050 531.600 ;
        RECT 19.950 529.950 22.050 530.400 ;
        RECT 64.950 529.950 67.050 530.400 ;
        RECT 73.950 529.950 76.050 530.400 ;
        RECT 169.950 531.600 172.050 532.050 ;
        RECT 178.950 531.600 181.050 532.050 ;
        RECT 222.000 531.600 226.050 532.050 ;
        RECT 169.950 530.400 181.050 531.600 ;
        RECT 169.950 529.950 172.050 530.400 ;
        RECT 178.950 529.950 181.050 530.400 ;
        RECT 221.400 529.950 226.050 531.600 ;
        RECT 229.950 531.600 232.050 532.050 ;
        RECT 271.950 531.600 274.050 532.050 ;
        RECT 229.950 530.400 240.600 531.600 ;
        RECT 229.950 529.950 232.050 530.400 ;
        RECT 31.950 528.600 34.050 529.050 ;
        RECT 37.950 528.600 40.050 529.200 ;
        RECT 55.950 528.600 58.050 529.200 ;
        RECT 31.950 527.400 40.050 528.600 ;
        RECT 31.950 526.950 34.050 527.400 ;
        RECT 37.950 527.100 40.050 527.400 ;
        RECT 53.400 527.400 58.050 528.600 ;
        RECT 53.400 523.050 54.600 527.400 ;
        RECT 55.950 527.100 58.050 527.400 ;
        RECT 94.950 527.100 97.050 529.200 ;
        RECT 127.950 528.750 130.050 529.200 ;
        RECT 136.950 528.750 139.050 529.200 ;
        RECT 127.950 527.550 139.050 528.750 ;
        RECT 127.950 527.100 130.050 527.550 ;
        RECT 136.950 527.100 139.050 527.550 ;
        RECT 142.950 528.600 145.050 529.200 ;
        RECT 142.950 527.400 147.600 528.600 ;
        RECT 142.950 527.100 145.050 527.400 ;
        RECT 52.950 520.950 55.050 523.050 ;
        RECT 82.950 522.600 85.050 522.900 ;
        RECT 95.400 522.600 96.600 527.100 ;
        RECT 146.400 522.900 147.600 527.400 ;
        RECT 166.950 526.950 169.050 529.050 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 207.000 528.600 211.050 529.050 ;
        RECT 206.400 526.950 211.050 528.600 ;
        RECT 167.400 523.050 168.600 526.950 ;
        RECT 82.950 521.400 96.600 522.600 ;
        RECT 124.950 522.450 127.050 522.900 ;
        RECT 133.950 522.450 136.050 522.900 ;
        RECT 82.950 520.800 85.050 521.400 ;
        RECT 124.950 521.250 136.050 522.450 ;
        RECT 124.950 520.800 127.050 521.250 ;
        RECT 133.950 520.800 136.050 521.250 ;
        RECT 145.950 522.450 148.050 522.900 ;
        RECT 157.950 522.450 160.050 522.900 ;
        RECT 145.950 521.250 160.050 522.450 ;
        RECT 145.950 520.800 148.050 521.250 ;
        RECT 157.950 520.800 160.050 521.250 ;
        RECT 166.950 520.950 169.050 523.050 ;
        RECT 40.950 519.600 43.050 520.050 ;
        RECT 58.950 519.600 61.050 520.050 ;
        RECT 40.950 518.400 61.050 519.600 ;
        RECT 40.950 517.950 43.050 518.400 ;
        RECT 58.950 517.950 61.050 518.400 ;
        RECT 103.950 519.600 106.050 520.050 ;
        RECT 127.950 519.600 130.050 520.050 ;
        RECT 103.950 518.400 130.050 519.600 ;
        RECT 173.400 519.600 174.600 526.950 ;
        RECT 181.950 522.600 184.050 522.900 ;
        RECT 190.950 522.600 193.050 523.050 ;
        RECT 206.400 522.900 207.600 526.950 ;
        RECT 221.400 522.900 222.600 529.950 ;
        RECT 226.950 526.950 229.050 529.050 ;
        RECT 235.950 526.950 238.050 529.050 ;
        RECT 239.400 528.600 240.600 530.400 ;
        RECT 271.950 530.400 321.600 531.600 ;
        RECT 271.950 529.950 274.050 530.400 ;
        RECT 241.950 528.600 244.050 529.200 ;
        RECT 239.400 527.400 244.050 528.600 ;
        RECT 241.950 527.100 244.050 527.400 ;
        RECT 256.950 526.950 259.050 529.050 ;
        RECT 262.950 528.600 265.050 529.200 ;
        RECT 283.950 528.600 286.050 529.200 ;
        RECT 301.950 528.600 304.050 529.200 ;
        RECT 262.950 527.400 282.600 528.600 ;
        RECT 262.950 527.100 265.050 527.400 ;
        RECT 227.400 523.050 228.600 526.950 ;
        RECT 181.950 521.400 193.050 522.600 ;
        RECT 181.950 520.800 184.050 521.400 ;
        RECT 190.950 520.950 193.050 521.400 ;
        RECT 205.950 520.800 208.050 522.900 ;
        RECT 220.950 520.800 223.050 522.900 ;
        RECT 226.950 520.950 229.050 523.050 ;
        RECT 236.400 522.600 237.600 526.950 ;
        RECT 238.950 522.600 241.050 522.900 ;
        RECT 236.400 521.400 241.050 522.600 ;
        RECT 238.950 520.800 241.050 521.400 ;
        RECT 250.950 522.600 253.050 523.050 ;
        RECT 257.400 522.600 258.600 526.950 ;
        RECT 281.400 522.900 282.600 527.400 ;
        RECT 283.950 527.400 304.050 528.600 ;
        RECT 283.950 527.100 286.050 527.400 ;
        RECT 301.950 527.100 304.050 527.400 ;
        RECT 307.950 527.100 310.050 529.200 ;
        RECT 250.950 521.400 258.600 522.600 ;
        RECT 250.950 520.950 253.050 521.400 ;
        RECT 280.950 520.800 283.050 522.900 ;
        RECT 308.400 522.600 309.600 527.100 ;
        RECT 320.400 525.600 321.600 530.400 ;
        RECT 337.950 529.950 340.050 532.050 ;
        RECT 322.950 528.600 325.050 529.200 ;
        RECT 331.950 528.600 334.050 529.050 ;
        RECT 322.950 527.400 334.050 528.600 ;
        RECT 322.950 527.100 325.050 527.400 ;
        RECT 331.950 526.950 334.050 527.400 ;
        RECT 338.400 526.050 339.600 529.950 ;
        RECT 346.950 528.600 349.050 532.050 ;
        RECT 397.950 531.600 400.050 532.050 ;
        RECT 406.950 531.600 409.050 532.050 ;
        RECT 415.800 531.600 417.900 532.050 ;
        RECT 397.950 530.400 405.600 531.600 ;
        RECT 397.950 529.950 400.050 530.400 ;
        RECT 344.400 528.000 349.050 528.600 ;
        RECT 404.400 528.600 405.600 530.400 ;
        RECT 406.950 530.400 417.900 531.600 ;
        RECT 406.950 529.950 409.050 530.400 ;
        RECT 415.800 529.950 417.900 530.400 ;
        RECT 418.950 531.600 421.050 532.050 ;
        RECT 434.400 531.600 435.600 533.400 ;
        RECT 475.950 532.950 478.050 533.400 ;
        RECT 538.950 534.600 541.050 534.900 ;
        RECT 574.950 534.600 577.050 535.050 ;
        RECT 595.950 534.600 598.050 535.050 ;
        RECT 538.950 533.400 598.050 534.600 ;
        RECT 538.950 532.800 541.050 533.400 ;
        RECT 574.950 532.950 577.050 533.400 ;
        RECT 595.950 532.950 598.050 533.400 ;
        RECT 889.950 534.600 892.050 535.050 ;
        RECT 934.950 534.600 937.050 535.050 ;
        RECT 889.950 533.400 937.050 534.600 ;
        RECT 889.950 532.950 892.050 533.400 ;
        RECT 934.950 532.950 937.050 533.400 ;
        RECT 418.950 530.400 435.600 531.600 ;
        RECT 490.950 531.600 493.050 532.050 ;
        RECT 539.400 531.600 540.600 532.800 ;
        RECT 490.950 530.400 540.600 531.600 ;
        RECT 418.950 529.950 421.050 530.400 ;
        RECT 490.950 529.950 493.050 530.400 ;
        RECT 550.950 529.950 553.050 532.050 ;
        RECT 715.950 531.600 718.050 532.050 ;
        RECT 727.950 531.600 730.050 532.050 ;
        RECT 715.950 530.400 730.050 531.600 ;
        RECT 715.950 529.950 718.050 530.400 ;
        RECT 727.950 529.950 730.050 530.400 ;
        RECT 742.950 531.600 745.050 532.050 ;
        RECT 757.950 531.600 760.050 532.050 ;
        RECT 742.950 530.400 760.050 531.600 ;
        RECT 742.950 529.950 745.050 530.400 ;
        RECT 757.950 529.950 760.050 530.400 ;
        RECT 829.950 531.600 832.050 532.050 ;
        RECT 835.950 531.600 838.050 532.050 ;
        RECT 829.950 530.400 838.050 531.600 ;
        RECT 829.950 529.950 832.050 530.400 ;
        RECT 835.950 529.950 838.050 530.400 ;
        RECT 412.950 528.600 415.050 529.050 ;
        RECT 433.950 528.600 436.050 529.050 ;
        RECT 344.400 527.400 348.600 528.000 ;
        RECT 404.400 527.400 423.600 528.600 ;
        RECT 428.400 528.000 436.050 528.600 ;
        RECT 334.800 525.600 336.900 525.900 ;
        RECT 320.400 524.400 336.900 525.600 ;
        RECT 334.800 523.800 336.900 524.400 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 344.400 525.600 345.600 527.400 ;
        RECT 412.950 526.950 415.050 527.400 ;
        RECT 370.950 525.600 373.050 526.200 ;
        RECT 341.400 524.400 345.600 525.600 ;
        RECT 347.400 525.000 373.050 525.600 ;
        RECT 346.950 524.400 373.050 525.000 ;
        RECT 284.400 522.000 309.600 522.600 ;
        RECT 283.950 521.400 309.600 522.000 ;
        RECT 313.950 522.600 316.050 523.050 ;
        RECT 328.950 522.600 331.050 522.900 ;
        RECT 313.950 521.400 331.050 522.600 ;
        RECT 178.950 519.600 181.050 520.050 ;
        RECT 173.400 518.400 181.050 519.600 ;
        RECT 103.950 517.950 106.050 518.400 ;
        RECT 127.950 517.950 130.050 518.400 ;
        RECT 178.950 517.950 181.050 518.400 ;
        RECT 262.950 519.600 265.050 520.050 ;
        RECT 268.950 519.600 271.050 520.050 ;
        RECT 262.950 518.400 271.050 519.600 ;
        RECT 262.950 517.950 265.050 518.400 ;
        RECT 268.950 517.950 271.050 518.400 ;
        RECT 283.950 517.950 286.050 521.400 ;
        RECT 313.950 520.950 316.050 521.400 ;
        RECT 328.950 520.800 331.050 521.400 ;
        RECT 341.400 520.050 342.600 524.400 ;
        RECT 346.950 520.950 349.050 524.400 ;
        RECT 370.950 524.100 373.050 524.400 ;
        RECT 391.950 525.600 394.050 526.050 ;
        RECT 400.950 525.600 403.050 526.050 ;
        RECT 391.950 524.400 403.050 525.600 ;
        RECT 391.950 523.950 394.050 524.400 ;
        RECT 400.950 523.950 403.050 524.400 ;
        RECT 422.400 523.050 423.600 527.400 ;
        RECT 427.950 527.400 436.050 528.000 ;
        RECT 427.950 523.950 430.050 527.400 ;
        RECT 433.950 526.950 436.050 527.400 ;
        RECT 475.950 525.450 478.050 525.900 ;
        RECT 502.950 525.450 505.050 525.900 ;
        RECT 475.950 524.250 505.050 525.450 ;
        RECT 475.950 523.800 478.050 524.250 ;
        RECT 502.950 523.800 505.050 524.250 ;
        RECT 541.950 525.450 544.050 525.900 ;
        RECT 551.400 525.450 552.600 529.950 ;
        RECT 580.950 528.750 583.050 529.200 ;
        RECT 595.950 528.750 598.050 529.200 ;
        RECT 580.950 527.550 598.050 528.750 ;
        RECT 580.950 527.100 583.050 527.550 ;
        RECT 595.950 527.100 598.050 527.550 ;
        RECT 607.950 527.100 610.050 529.200 ;
        RECT 619.950 528.750 622.050 529.200 ;
        RECT 634.950 528.750 637.050 529.200 ;
        RECT 619.950 527.550 637.050 528.750 ;
        RECT 619.950 527.100 622.050 527.550 ;
        RECT 634.950 527.100 637.050 527.550 ;
        RECT 646.950 528.750 649.050 529.200 ;
        RECT 652.950 528.750 655.050 529.200 ;
        RECT 646.950 527.550 655.050 528.750 ;
        RECT 646.950 527.100 649.050 527.550 ;
        RECT 652.950 527.100 655.050 527.550 ;
        RECT 658.950 527.100 661.050 529.200 ;
        RECT 679.950 528.750 682.050 529.200 ;
        RECT 694.950 528.750 697.050 529.200 ;
        RECT 679.950 527.550 697.050 528.750 ;
        RECT 679.950 527.100 682.050 527.550 ;
        RECT 694.950 527.100 697.050 527.550 ;
        RECT 721.950 527.100 724.050 529.200 ;
        RECT 730.950 528.750 733.050 529.200 ;
        RECT 736.950 528.750 739.050 529.200 ;
        RECT 730.950 527.550 739.050 528.750 ;
        RECT 730.950 527.100 733.050 527.550 ;
        RECT 736.950 527.100 739.050 527.550 ;
        RECT 766.950 528.750 769.050 529.200 ;
        RECT 772.950 528.750 775.050 529.200 ;
        RECT 766.950 527.550 775.050 528.750 ;
        RECT 766.950 527.100 769.050 527.550 ;
        RECT 772.950 527.100 775.050 527.550 ;
        RECT 805.950 528.750 808.050 529.200 ;
        RECT 820.950 528.750 823.050 529.200 ;
        RECT 805.950 527.550 823.050 528.750 ;
        RECT 805.950 527.100 808.050 527.550 ;
        RECT 820.950 527.100 823.050 527.550 ;
        RECT 850.950 527.100 853.050 529.200 ;
        RECT 868.950 528.750 871.050 529.200 ;
        RECT 889.950 528.750 892.050 529.200 ;
        RECT 868.950 527.550 892.050 528.750 ;
        RECT 868.950 527.100 871.050 527.550 ;
        RECT 889.950 527.100 892.050 527.550 ;
        RECT 940.950 527.100 943.050 529.200 ;
        RECT 553.950 525.450 556.050 525.900 ;
        RECT 541.950 524.250 556.050 525.450 ;
        RECT 541.950 523.800 544.050 524.250 ;
        RECT 553.950 523.800 556.050 524.250 ;
        RECT 559.950 525.600 562.050 526.050 ;
        RECT 608.400 525.600 609.600 527.100 ;
        RECT 559.950 524.400 609.600 525.600 ;
        RECT 559.950 523.950 562.050 524.400 ;
        RECT 385.950 522.600 388.050 523.050 ;
        RECT 409.950 522.600 412.050 523.050 ;
        RECT 385.950 521.400 412.050 522.600 ;
        RECT 385.950 520.950 388.050 521.400 ;
        RECT 409.950 520.950 412.050 521.400 ;
        RECT 421.950 520.950 424.050 523.050 ;
        RECT 433.950 522.600 436.050 523.050 ;
        RECT 484.950 522.600 487.050 523.050 ;
        RECT 433.950 521.400 487.050 522.600 ;
        RECT 433.950 520.950 436.050 521.400 ;
        RECT 484.950 520.950 487.050 521.400 ;
        RECT 571.950 522.600 574.050 522.900 ;
        RECT 631.950 522.600 634.050 522.900 ;
        RECT 640.950 522.600 643.050 523.050 ;
        RECT 571.950 521.400 627.600 522.600 ;
        RECT 571.950 520.800 574.050 521.400 ;
        RECT 626.400 520.050 627.600 521.400 ;
        RECT 631.950 521.400 643.050 522.600 ;
        RECT 631.950 520.800 634.050 521.400 ;
        RECT 640.950 520.950 643.050 521.400 ;
        RECT 341.400 518.400 346.050 520.050 ;
        RECT 342.000 517.950 346.050 518.400 ;
        RECT 493.950 519.600 496.050 520.050 ;
        RECT 541.950 519.600 544.050 520.050 ;
        RECT 493.950 518.400 544.050 519.600 ;
        RECT 493.950 517.950 496.050 518.400 ;
        RECT 541.950 517.950 544.050 518.400 ;
        RECT 580.950 519.600 583.050 520.050 ;
        RECT 589.950 519.600 592.050 520.050 ;
        RECT 580.950 518.400 592.050 519.600 ;
        RECT 626.400 518.400 631.050 520.050 ;
        RECT 580.950 517.950 583.050 518.400 ;
        RECT 589.950 517.950 592.050 518.400 ;
        RECT 627.000 517.950 631.050 518.400 ;
        RECT 652.950 519.600 655.050 520.050 ;
        RECT 659.400 519.600 660.600 527.100 ;
        RECT 722.400 525.600 723.600 527.100 ;
        RECT 751.950 525.600 754.050 526.050 ;
        RECT 722.400 524.400 729.600 525.600 ;
        RECT 682.950 522.450 685.050 522.900 ;
        RECT 691.950 522.450 694.050 522.900 ;
        RECT 682.950 521.250 694.050 522.450 ;
        RECT 682.950 520.800 685.050 521.250 ;
        RECT 691.950 520.800 694.050 521.250 ;
        RECT 718.950 522.600 721.050 522.900 ;
        RECT 724.950 522.600 727.050 523.050 ;
        RECT 718.950 521.400 727.050 522.600 ;
        RECT 728.400 522.600 729.600 524.400 ;
        RECT 751.950 525.000 765.600 525.600 ;
        RECT 751.950 524.400 766.050 525.000 ;
        RECT 751.950 523.950 754.050 524.400 ;
        RECT 733.950 522.600 736.050 523.050 ;
        RECT 728.400 521.400 736.050 522.600 ;
        RECT 718.950 520.800 721.050 521.400 ;
        RECT 724.950 520.950 727.050 521.400 ;
        RECT 733.950 520.950 736.050 521.400 ;
        RECT 763.950 520.950 766.050 524.400 ;
        RECT 790.950 522.600 793.050 526.050 ;
        RECT 802.950 522.600 805.050 522.900 ;
        RECT 790.950 522.000 805.050 522.600 ;
        RECT 791.400 521.400 805.050 522.000 ;
        RECT 652.950 518.400 660.600 519.600 ;
        RECT 703.950 519.600 706.050 520.050 ;
        RECT 712.950 519.600 715.050 520.050 ;
        RECT 730.800 519.600 732.900 520.050 ;
        RECT 703.950 518.400 732.900 519.600 ;
        RECT 734.400 519.600 735.600 520.950 ;
        RECT 802.950 520.800 805.050 521.400 ;
        RECT 841.950 522.600 844.050 523.050 ;
        RECT 851.400 522.600 852.600 527.100 ;
        RECT 941.400 523.050 942.600 527.100 ;
        RECT 841.950 521.400 852.600 522.600 ;
        RECT 853.950 522.600 856.050 522.900 ;
        RECT 859.950 522.600 862.050 523.050 ;
        RECT 853.950 521.400 862.050 522.600 ;
        RECT 841.950 520.950 844.050 521.400 ;
        RECT 853.950 520.800 856.050 521.400 ;
        RECT 859.950 520.950 862.050 521.400 ;
        RECT 865.950 522.450 868.050 522.900 ;
        RECT 877.950 522.450 880.050 522.900 ;
        RECT 865.950 521.250 880.050 522.450 ;
        RECT 865.950 520.800 868.050 521.250 ;
        RECT 877.950 520.800 880.050 521.250 ;
        RECT 913.950 522.600 916.050 523.050 ;
        RECT 925.950 522.600 928.050 523.050 ;
        RECT 913.950 521.400 928.050 522.600 ;
        RECT 941.400 521.400 946.050 523.050 ;
        RECT 913.950 520.950 916.050 521.400 ;
        RECT 925.950 520.950 928.050 521.400 ;
        RECT 942.000 520.950 946.050 521.400 ;
        RECT 751.950 519.600 754.050 520.050 ;
        RECT 734.400 518.400 754.050 519.600 ;
        RECT 652.950 517.950 655.050 518.400 ;
        RECT 703.950 517.950 706.050 518.400 ;
        RECT 712.950 517.950 715.050 518.400 ;
        RECT 730.800 517.950 732.900 518.400 ;
        RECT 751.950 517.950 754.050 518.400 ;
        RECT 760.950 519.600 763.050 520.050 ;
        RECT 766.950 519.600 769.050 520.050 ;
        RECT 760.950 518.400 769.050 519.600 ;
        RECT 760.950 517.950 763.050 518.400 ;
        RECT 766.950 517.950 769.050 518.400 ;
        RECT 808.950 519.600 811.050 520.050 ;
        RECT 829.950 519.600 832.050 520.050 ;
        RECT 808.950 518.400 832.050 519.600 ;
        RECT 808.950 517.950 811.050 518.400 ;
        RECT 829.950 517.950 832.050 518.400 ;
        RECT 22.950 516.600 25.050 517.050 ;
        RECT 31.950 516.600 34.050 517.050 ;
        RECT 22.950 515.400 34.050 516.600 ;
        RECT 22.950 514.950 25.050 515.400 ;
        RECT 31.950 514.950 34.050 515.400 ;
        RECT 61.950 516.600 64.050 517.050 ;
        RECT 76.950 516.600 79.050 517.050 ;
        RECT 61.950 515.400 79.050 516.600 ;
        RECT 61.950 514.950 64.050 515.400 ;
        RECT 76.950 514.950 79.050 515.400 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 136.950 516.600 139.050 517.050 ;
        RECT 130.950 515.400 139.050 516.600 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 136.950 514.950 139.050 515.400 ;
        RECT 160.950 516.600 163.050 517.050 ;
        RECT 184.950 516.600 187.050 517.050 ;
        RECT 160.950 515.400 187.050 516.600 ;
        RECT 160.950 514.950 163.050 515.400 ;
        RECT 184.950 514.950 187.050 515.400 ;
        RECT 199.950 516.600 202.050 517.050 ;
        RECT 211.950 516.600 214.050 517.050 ;
        RECT 199.950 515.400 214.050 516.600 ;
        RECT 199.950 514.950 202.050 515.400 ;
        RECT 211.950 514.950 214.050 515.400 ;
        RECT 256.950 516.600 259.050 517.050 ;
        RECT 277.950 516.600 280.050 517.050 ;
        RECT 256.950 515.400 280.050 516.600 ;
        RECT 256.950 514.950 259.050 515.400 ;
        RECT 277.950 514.950 280.050 515.400 ;
        RECT 403.950 516.600 406.050 517.050 ;
        RECT 415.950 516.600 418.050 517.050 ;
        RECT 403.950 515.400 418.050 516.600 ;
        RECT 403.950 514.950 406.050 515.400 ;
        RECT 415.950 514.950 418.050 515.400 ;
        RECT 481.950 516.600 484.050 517.050 ;
        RECT 544.950 516.600 547.050 517.050 ;
        RECT 559.950 516.600 562.050 517.050 ;
        RECT 481.950 515.400 562.050 516.600 ;
        RECT 481.950 514.950 484.050 515.400 ;
        RECT 544.950 514.950 547.050 515.400 ;
        RECT 559.950 514.950 562.050 515.400 ;
        RECT 574.950 516.600 577.050 517.050 ;
        RECT 592.950 516.600 595.050 517.050 ;
        RECT 622.950 516.600 625.050 517.050 ;
        RECT 574.950 515.400 625.050 516.600 ;
        RECT 574.950 514.950 577.050 515.400 ;
        RECT 592.950 514.950 595.050 515.400 ;
        RECT 622.950 514.950 625.050 515.400 ;
        RECT 739.950 516.600 742.050 517.050 ;
        RECT 745.950 516.600 748.050 517.050 ;
        RECT 739.950 515.400 748.050 516.600 ;
        RECT 739.950 514.950 742.050 515.400 ;
        RECT 745.950 514.950 748.050 515.400 ;
        RECT 832.950 516.600 835.050 517.050 ;
        RECT 856.950 516.600 859.050 517.050 ;
        RECT 832.950 515.400 859.050 516.600 ;
        RECT 832.950 514.950 835.050 515.400 ;
        RECT 856.950 514.950 859.050 515.400 ;
        RECT 862.950 516.600 867.000 517.050 ;
        RECT 871.950 516.600 874.050 517.050 ;
        RECT 940.950 516.600 943.050 517.050 ;
        RECT 862.950 514.950 867.600 516.600 ;
        RECT 871.950 515.400 943.050 516.600 ;
        RECT 871.950 514.950 874.050 515.400 ;
        RECT 940.950 514.950 943.050 515.400 ;
        RECT 46.950 513.600 49.050 514.050 ;
        RECT 62.400 513.600 63.600 514.950 ;
        RECT 46.950 512.400 63.600 513.600 ;
        RECT 100.950 513.600 103.050 514.050 ;
        RECT 115.950 513.600 118.050 514.050 ;
        RECT 100.950 512.400 118.050 513.600 ;
        RECT 46.950 511.950 49.050 512.400 ;
        RECT 100.950 511.950 103.050 512.400 ;
        RECT 115.950 511.950 118.050 512.400 ;
        RECT 139.950 513.600 142.050 514.050 ;
        RECT 148.950 513.600 151.050 514.050 ;
        RECT 139.950 512.400 151.050 513.600 ;
        RECT 139.950 511.950 142.050 512.400 ;
        RECT 148.950 511.950 151.050 512.400 ;
        RECT 157.950 513.600 160.050 514.050 ;
        RECT 187.950 513.600 190.050 514.050 ;
        RECT 157.950 512.400 190.050 513.600 ;
        RECT 157.950 511.950 160.050 512.400 ;
        RECT 187.950 511.950 190.050 512.400 ;
        RECT 250.950 513.600 253.050 514.050 ;
        RECT 286.950 513.600 289.050 514.050 ;
        RECT 250.950 512.400 289.050 513.600 ;
        RECT 250.950 511.950 253.050 512.400 ;
        RECT 286.950 511.950 289.050 512.400 ;
        RECT 295.950 513.600 298.050 514.050 ;
        RECT 385.950 513.600 388.050 514.050 ;
        RECT 295.950 512.400 388.050 513.600 ;
        RECT 295.950 511.950 298.050 512.400 ;
        RECT 385.950 511.950 388.050 512.400 ;
        RECT 412.950 513.600 415.050 514.050 ;
        RECT 478.950 513.600 481.050 514.050 ;
        RECT 412.950 512.400 481.050 513.600 ;
        RECT 412.950 511.950 415.050 512.400 ;
        RECT 478.950 511.950 481.050 512.400 ;
        RECT 502.950 513.600 505.050 514.050 ;
        RECT 556.950 513.600 559.050 514.050 ;
        RECT 625.950 513.600 628.050 514.050 ;
        RECT 634.950 513.600 637.050 514.050 ;
        RECT 502.950 512.400 559.050 513.600 ;
        RECT 502.950 511.950 505.050 512.400 ;
        RECT 556.950 511.950 559.050 512.400 ;
        RECT 584.400 512.400 637.050 513.600 ;
        RECT 139.950 510.600 142.050 510.900 ;
        RECT 151.950 510.600 154.050 511.050 ;
        RECT 139.950 509.400 154.050 510.600 ;
        RECT 139.950 508.800 142.050 509.400 ;
        RECT 151.950 508.950 154.050 509.400 ;
        RECT 190.950 510.600 193.050 511.050 ;
        RECT 211.950 510.600 214.050 511.050 ;
        RECT 262.950 510.600 265.050 511.050 ;
        RECT 190.950 509.400 214.050 510.600 ;
        RECT 190.950 508.950 193.050 509.400 ;
        RECT 211.950 508.950 214.050 509.400 ;
        RECT 257.400 509.400 265.050 510.600 ;
        RECT 7.950 507.600 10.050 508.050 ;
        RECT 28.950 507.600 31.050 508.050 ;
        RECT 7.950 506.400 31.050 507.600 ;
        RECT 7.950 505.950 10.050 506.400 ;
        RECT 28.950 505.950 31.050 506.400 ;
        RECT 67.950 507.600 70.050 508.050 ;
        RECT 100.950 507.600 103.050 508.050 ;
        RECT 67.950 506.400 103.050 507.600 ;
        RECT 67.950 505.950 70.050 506.400 ;
        RECT 100.950 505.950 103.050 506.400 ;
        RECT 145.950 507.600 148.050 508.050 ;
        RECT 175.950 507.600 178.050 508.050 ;
        RECT 257.400 507.600 258.600 509.400 ;
        RECT 262.950 508.950 265.050 509.400 ;
        RECT 298.950 510.600 301.050 511.050 ;
        RECT 337.950 510.600 340.050 511.050 ;
        RECT 298.950 509.400 340.050 510.600 ;
        RECT 298.950 508.950 301.050 509.400 ;
        RECT 337.950 508.950 340.050 509.400 ;
        RECT 373.950 510.600 376.050 511.050 ;
        RECT 400.950 510.600 403.050 511.050 ;
        RECT 373.950 509.400 403.050 510.600 ;
        RECT 373.950 508.950 376.050 509.400 ;
        RECT 400.950 508.950 403.050 509.400 ;
        RECT 496.950 510.600 499.050 511.050 ;
        RECT 562.950 510.600 565.050 511.050 ;
        RECT 584.400 510.600 585.600 512.400 ;
        RECT 625.950 511.950 628.050 512.400 ;
        RECT 634.950 511.950 637.050 512.400 ;
        RECT 655.950 513.600 658.050 514.050 ;
        RECT 679.950 513.600 682.050 514.050 ;
        RECT 655.950 512.400 682.050 513.600 ;
        RECT 655.950 511.950 658.050 512.400 ;
        RECT 679.950 511.950 682.050 512.400 ;
        RECT 685.950 513.600 688.050 514.050 ;
        RECT 706.950 513.600 709.050 514.050 ;
        RECT 685.950 512.400 709.050 513.600 ;
        RECT 685.950 511.950 688.050 512.400 ;
        RECT 706.950 511.950 709.050 512.400 ;
        RECT 790.950 513.600 793.050 514.050 ;
        RECT 802.950 513.600 805.050 514.050 ;
        RECT 790.950 512.400 805.050 513.600 ;
        RECT 790.950 511.950 793.050 512.400 ;
        RECT 802.950 511.950 805.050 512.400 ;
        RECT 841.950 513.600 844.050 514.050 ;
        RECT 859.950 513.600 862.050 514.050 ;
        RECT 841.950 512.400 862.050 513.600 ;
        RECT 866.400 513.600 867.600 514.950 ;
        RECT 895.950 513.600 898.050 514.050 ;
        RECT 919.950 513.600 922.050 514.050 ;
        RECT 866.400 512.400 922.050 513.600 ;
        RECT 841.950 511.950 844.050 512.400 ;
        RECT 859.950 511.950 862.050 512.400 ;
        RECT 895.950 511.950 898.050 512.400 ;
        RECT 919.950 511.950 922.050 512.400 ;
        RECT 496.950 509.400 585.600 510.600 ;
        RECT 589.950 510.600 592.050 511.050 ;
        RECT 607.950 510.600 610.050 511.050 ;
        RECT 589.950 509.400 610.050 510.600 ;
        RECT 496.950 508.950 499.050 509.400 ;
        RECT 562.950 508.950 565.050 509.400 ;
        RECT 589.950 508.950 592.050 509.400 ;
        RECT 607.950 508.950 610.050 509.400 ;
        RECT 664.950 510.600 667.050 511.050 ;
        RECT 676.950 510.600 679.050 511.050 ;
        RECT 664.950 509.400 679.050 510.600 ;
        RECT 664.950 508.950 667.050 509.400 ;
        RECT 676.950 508.950 679.050 509.400 ;
        RECT 712.950 510.600 715.050 511.050 ;
        RECT 727.950 510.600 730.050 511.050 ;
        RECT 742.950 510.600 745.050 511.050 ;
        RECT 712.950 509.400 745.050 510.600 ;
        RECT 712.950 508.950 715.050 509.400 ;
        RECT 727.950 508.950 730.050 509.400 ;
        RECT 742.950 508.950 745.050 509.400 ;
        RECT 754.950 510.600 757.050 511.050 ;
        RECT 781.950 510.600 784.050 511.050 ;
        RECT 754.950 509.400 784.050 510.600 ;
        RECT 754.950 508.950 757.050 509.400 ;
        RECT 781.950 508.950 784.050 509.400 ;
        RECT 901.950 510.600 904.050 511.050 ;
        RECT 913.950 510.600 916.050 511.050 ;
        RECT 901.950 509.400 916.050 510.600 ;
        RECT 901.950 508.950 904.050 509.400 ;
        RECT 913.950 508.950 916.050 509.400 ;
        RECT 145.950 506.400 178.050 507.600 ;
        RECT 145.950 505.950 148.050 506.400 ;
        RECT 175.950 505.950 178.050 506.400 ;
        RECT 251.400 506.400 258.600 507.600 ;
        RECT 274.950 507.600 277.050 508.050 ;
        RECT 304.950 507.600 307.050 508.050 ;
        RECT 274.950 506.400 307.050 507.600 ;
        RECT 251.400 505.050 252.600 506.400 ;
        RECT 274.950 505.950 277.050 506.400 ;
        RECT 304.950 505.950 307.050 506.400 ;
        RECT 382.950 507.600 385.050 508.050 ;
        RECT 391.950 507.600 394.050 508.050 ;
        RECT 382.950 506.400 394.050 507.600 ;
        RECT 382.950 505.950 385.050 506.400 ;
        RECT 391.950 505.950 394.050 506.400 ;
        RECT 433.950 507.600 436.050 508.050 ;
        RECT 442.950 507.600 445.050 508.050 ;
        RECT 433.950 506.400 445.050 507.600 ;
        RECT 433.950 505.950 436.050 506.400 ;
        RECT 442.950 505.950 445.050 506.400 ;
        RECT 448.950 507.600 451.050 508.050 ;
        RECT 481.950 507.600 484.050 508.050 ;
        RECT 448.950 506.400 484.050 507.600 ;
        RECT 448.950 505.950 451.050 506.400 ;
        RECT 481.950 505.950 484.050 506.400 ;
        RECT 514.950 507.600 517.050 508.050 ;
        RECT 586.950 507.600 589.050 508.050 ;
        RECT 514.950 506.400 589.050 507.600 ;
        RECT 514.950 505.950 517.050 506.400 ;
        RECT 586.950 505.950 589.050 506.400 ;
        RECT 628.950 507.600 631.050 508.050 ;
        RECT 703.950 507.600 706.050 508.050 ;
        RECT 628.950 506.400 706.050 507.600 ;
        RECT 628.950 505.950 631.050 506.400 ;
        RECT 703.950 505.950 706.050 506.400 ;
        RECT 847.950 507.600 850.050 508.050 ;
        RECT 886.950 507.600 889.050 508.050 ;
        RECT 847.950 506.400 889.050 507.600 ;
        RECT 847.950 505.950 850.050 506.400 ;
        RECT 886.950 505.950 889.050 506.400 ;
        RECT 895.950 507.600 898.050 508.050 ;
        RECT 946.950 507.600 949.050 508.050 ;
        RECT 895.950 506.400 949.050 507.600 ;
        RECT 895.950 505.950 898.050 506.400 ;
        RECT 946.950 505.950 949.050 506.400 ;
        RECT 37.950 504.600 40.050 505.050 ;
        RECT 79.950 504.600 82.050 505.050 ;
        RECT 94.950 504.600 97.050 505.050 ;
        RECT 37.950 503.400 97.050 504.600 ;
        RECT 37.950 502.950 40.050 503.400 ;
        RECT 79.950 502.950 82.050 503.400 ;
        RECT 94.950 502.950 97.050 503.400 ;
        RECT 127.950 504.600 130.050 505.050 ;
        RECT 163.950 504.600 166.050 505.050 ;
        RECT 169.950 504.600 172.050 505.050 ;
        RECT 127.950 503.400 172.050 504.600 ;
        RECT 127.950 502.950 130.050 503.400 ;
        RECT 163.950 502.950 166.050 503.400 ;
        RECT 169.950 502.950 172.050 503.400 ;
        RECT 181.950 504.600 184.050 505.050 ;
        RECT 211.950 504.600 214.050 505.050 ;
        RECT 181.950 503.400 214.050 504.600 ;
        RECT 181.950 502.950 184.050 503.400 ;
        RECT 211.950 502.950 214.050 503.400 ;
        RECT 244.950 504.600 247.050 505.050 ;
        RECT 250.950 504.600 253.050 505.050 ;
        RECT 244.950 503.400 253.050 504.600 ;
        RECT 244.950 502.950 247.050 503.400 ;
        RECT 250.950 502.950 253.050 503.400 ;
        RECT 259.950 504.600 262.050 505.050 ;
        RECT 277.950 504.600 280.050 505.050 ;
        RECT 259.950 503.400 280.050 504.600 ;
        RECT 259.950 502.950 262.050 503.400 ;
        RECT 277.950 502.950 280.050 503.400 ;
        RECT 304.950 504.600 307.050 504.900 ;
        RECT 316.950 504.600 319.050 505.050 ;
        RECT 304.950 503.400 319.050 504.600 ;
        RECT 304.950 502.800 307.050 503.400 ;
        RECT 316.950 502.950 319.050 503.400 ;
        RECT 385.950 504.600 388.050 505.050 ;
        RECT 403.950 504.600 406.050 505.050 ;
        RECT 385.950 503.400 406.050 504.600 ;
        RECT 385.950 502.950 388.050 503.400 ;
        RECT 403.950 502.950 406.050 503.400 ;
        RECT 409.950 504.600 412.050 505.050 ;
        RECT 484.950 504.600 487.050 505.050 ;
        RECT 409.950 503.400 487.050 504.600 ;
        RECT 409.950 502.950 412.050 503.400 ;
        RECT 484.950 502.950 487.050 503.400 ;
        RECT 526.950 504.600 529.050 505.050 ;
        RECT 538.950 504.600 541.050 505.050 ;
        RECT 526.950 503.400 541.050 504.600 ;
        RECT 526.950 502.950 529.050 503.400 ;
        RECT 538.950 502.950 541.050 503.400 ;
        RECT 592.950 504.600 595.050 505.050 ;
        RECT 601.950 504.600 604.050 505.050 ;
        RECT 610.950 504.600 613.050 505.050 ;
        RECT 592.950 503.400 613.050 504.600 ;
        RECT 592.950 502.950 595.050 503.400 ;
        RECT 601.950 502.950 604.050 503.400 ;
        RECT 610.950 502.950 613.050 503.400 ;
        RECT 820.950 504.600 823.050 505.050 ;
        RECT 844.950 504.600 847.050 505.050 ;
        RECT 820.950 503.400 847.050 504.600 ;
        RECT 820.950 502.950 823.050 503.400 ;
        RECT 844.950 502.950 847.050 503.400 ;
        RECT 190.950 501.600 193.050 502.050 ;
        RECT 202.950 501.600 205.050 502.050 ;
        RECT 190.950 500.400 205.050 501.600 ;
        RECT 190.950 499.950 193.050 500.400 ;
        RECT 202.950 499.950 205.050 500.400 ;
        RECT 214.950 501.600 217.050 502.050 ;
        RECT 289.950 501.600 292.050 502.050 ;
        RECT 214.950 500.400 292.050 501.600 ;
        RECT 214.950 499.950 217.050 500.400 ;
        RECT 289.950 499.950 292.050 500.400 ;
        RECT 295.950 501.600 298.050 502.050 ;
        RECT 310.950 501.600 313.050 502.050 ;
        RECT 295.950 500.400 313.050 501.600 ;
        RECT 295.950 499.950 298.050 500.400 ;
        RECT 310.950 499.950 313.050 500.400 ;
        RECT 451.950 501.600 454.050 502.050 ;
        RECT 487.950 501.600 490.050 502.050 ;
        RECT 451.950 500.400 490.050 501.600 ;
        RECT 451.950 499.950 454.050 500.400 ;
        RECT 487.950 499.950 490.050 500.400 ;
        RECT 553.950 501.600 556.050 502.050 ;
        RECT 568.950 501.600 571.050 502.050 ;
        RECT 553.950 500.400 571.050 501.600 ;
        RECT 553.950 499.950 556.050 500.400 ;
        RECT 568.950 499.950 571.050 500.400 ;
        RECT 628.950 501.600 631.050 502.050 ;
        RECT 670.950 501.600 673.050 502.050 ;
        RECT 628.950 500.400 673.050 501.600 ;
        RECT 628.950 499.950 631.050 500.400 ;
        RECT 670.950 499.950 673.050 500.400 ;
        RECT 739.950 501.600 742.050 502.050 ;
        RECT 757.950 501.600 760.050 502.050 ;
        RECT 739.950 500.400 760.050 501.600 ;
        RECT 739.950 499.950 742.050 500.400 ;
        RECT 757.950 499.950 760.050 500.400 ;
        RECT 769.950 501.600 772.050 502.050 ;
        RECT 781.950 501.600 784.050 502.050 ;
        RECT 769.950 500.400 784.050 501.600 ;
        RECT 769.950 499.950 772.050 500.400 ;
        RECT 781.950 499.950 784.050 500.400 ;
        RECT 886.950 501.600 889.050 502.050 ;
        RECT 907.950 501.600 910.050 502.050 ;
        RECT 886.950 500.400 910.050 501.600 ;
        RECT 886.950 499.950 889.050 500.400 ;
        RECT 907.950 499.950 910.050 500.400 ;
        RECT 31.950 498.600 34.050 499.200 ;
        RECT 46.950 498.600 49.050 499.050 ;
        RECT 31.950 497.400 49.050 498.600 ;
        RECT 31.950 497.100 34.050 497.400 ;
        RECT 46.950 496.950 49.050 497.400 ;
        RECT 82.950 496.950 85.050 499.050 ;
        RECT 133.950 498.600 136.050 499.050 ;
        RECT 163.950 498.600 166.050 499.050 ;
        RECT 181.950 498.600 184.050 499.050 ;
        RECT 229.950 498.600 232.050 499.050 ;
        RECT 262.950 498.600 265.050 499.050 ;
        RECT 271.950 498.600 274.050 499.050 ;
        RECT 133.950 497.400 184.050 498.600 ;
        RECT 133.950 496.950 136.050 497.400 ;
        RECT 163.950 496.950 166.050 497.400 ;
        RECT 181.950 496.950 184.050 497.400 ;
        RECT 215.400 497.400 274.050 498.600 ;
        RECT 25.950 495.600 28.050 496.050 ;
        RECT 31.950 495.600 34.050 496.050 ;
        RECT 25.950 494.400 34.050 495.600 ;
        RECT 25.950 493.950 28.050 494.400 ;
        RECT 31.950 493.950 34.050 494.400 ;
        RECT 58.950 495.600 61.050 496.200 ;
        RECT 58.950 494.400 75.600 495.600 ;
        RECT 58.950 494.100 61.050 494.400 ;
        RECT 74.400 490.050 75.600 494.400 ;
        RECT 73.950 487.950 76.050 490.050 ;
        RECT 83.400 487.050 84.600 496.950 ;
        RECT 85.950 495.600 88.050 496.200 ;
        RECT 94.950 495.600 97.050 496.050 ;
        RECT 106.950 495.600 109.050 496.200 ;
        RECT 127.950 495.600 130.050 496.200 ;
        RECT 145.800 495.600 147.900 496.050 ;
        RECT 85.950 494.400 93.600 495.600 ;
        RECT 85.950 494.100 88.050 494.400 ;
        RECT 92.400 489.600 93.600 494.400 ;
        RECT 94.950 494.400 102.600 495.600 ;
        RECT 94.950 493.950 97.050 494.400 ;
        RECT 97.950 489.600 100.050 489.900 ;
        RECT 92.400 488.400 100.050 489.600 ;
        RECT 101.400 489.600 102.600 494.400 ;
        RECT 106.950 494.400 130.050 495.600 ;
        RECT 106.950 494.100 109.050 494.400 ;
        RECT 127.950 494.100 130.050 494.400 ;
        RECT 137.400 494.400 147.900 495.600 ;
        RECT 137.400 490.050 138.600 494.400 ;
        RECT 145.800 493.950 147.900 494.400 ;
        RECT 148.950 495.600 151.050 496.200 ;
        RECT 154.950 495.600 157.050 496.050 ;
        RECT 148.950 494.400 157.050 495.600 ;
        RECT 148.950 494.100 151.050 494.400 ;
        RECT 154.950 493.950 157.050 494.400 ;
        RECT 169.950 495.600 172.050 496.200 ;
        RECT 175.950 495.600 178.050 496.050 ;
        RECT 169.950 494.400 178.050 495.600 ;
        RECT 169.950 494.100 172.050 494.400 ;
        RECT 175.950 493.950 178.050 494.400 ;
        RECT 196.950 495.600 199.050 496.200 ;
        RECT 215.400 495.600 216.600 497.400 ;
        RECT 229.950 496.950 232.050 497.400 ;
        RECT 262.950 496.950 265.050 497.400 ;
        RECT 271.950 496.950 274.050 497.400 ;
        RECT 196.950 494.400 216.600 495.600 ;
        RECT 217.950 495.600 220.050 496.200 ;
        RECT 235.950 495.600 238.050 496.200 ;
        RECT 217.950 494.400 238.050 495.600 ;
        RECT 196.950 494.100 199.050 494.400 ;
        RECT 217.950 494.100 220.050 494.400 ;
        RECT 235.950 494.100 238.050 494.400 ;
        RECT 244.950 494.100 247.050 496.200 ;
        RECT 277.950 495.600 280.050 496.200 ;
        RECT 310.950 495.750 313.050 496.200 ;
        RECT 316.950 495.750 319.050 496.200 ;
        RECT 277.950 494.400 282.600 495.600 ;
        RECT 277.950 494.100 280.050 494.400 ;
        RECT 155.400 490.050 156.600 493.950 ;
        RECT 245.400 492.600 246.600 494.100 ;
        RECT 221.400 491.400 246.600 492.600 ;
        RECT 124.950 489.600 127.050 489.900 ;
        RECT 101.400 488.400 127.050 489.600 ;
        RECT 97.950 487.800 100.050 488.400 ;
        RECT 124.950 487.800 127.050 488.400 ;
        RECT 136.950 487.950 139.050 490.050 ;
        RECT 154.950 487.950 157.050 490.050 ;
        RECT 160.950 489.600 163.050 490.050 ;
        RECT 178.800 489.600 180.900 490.050 ;
        RECT 221.400 489.900 222.600 491.400 ;
        RECT 160.950 488.400 180.900 489.600 ;
        RECT 160.950 487.950 163.050 488.400 ;
        RECT 178.800 487.950 180.900 488.400 ;
        RECT 181.950 489.450 184.050 489.900 ;
        RECT 187.950 489.450 190.050 489.900 ;
        RECT 181.950 488.250 190.050 489.450 ;
        RECT 181.950 487.800 184.050 488.250 ;
        RECT 187.950 487.800 190.050 488.250 ;
        RECT 220.950 487.800 223.050 489.900 ;
        RECT 226.950 489.600 229.050 490.050 ;
        RECT 238.950 489.600 241.050 489.900 ;
        RECT 226.950 488.400 241.050 489.600 ;
        RECT 245.400 489.600 246.600 491.400 ;
        RECT 250.950 492.600 253.050 493.050 ;
        RECT 281.400 492.600 282.600 494.400 ;
        RECT 310.950 494.550 319.050 495.750 ;
        RECT 310.950 494.100 313.050 494.550 ;
        RECT 316.950 494.100 319.050 494.550 ;
        RECT 292.950 492.600 295.050 493.050 ;
        RECT 331.950 492.600 334.050 496.050 ;
        RECT 340.950 492.600 343.050 496.050 ;
        RECT 343.950 495.600 346.050 499.050 ;
        RECT 484.950 498.600 487.050 499.050 ;
        RECT 502.950 498.600 505.050 499.050 ;
        RECT 484.950 497.400 505.050 498.600 ;
        RECT 484.950 496.950 487.050 497.400 ;
        RECT 502.950 496.950 505.050 497.400 ;
        RECT 535.950 498.600 538.050 499.050 ;
        RECT 565.950 498.600 568.050 499.050 ;
        RECT 535.950 497.400 568.050 498.600 ;
        RECT 535.950 496.950 538.050 497.400 ;
        RECT 565.950 496.950 568.050 497.400 ;
        RECT 355.950 495.600 358.050 496.050 ;
        RECT 367.950 495.600 370.050 496.200 ;
        RECT 343.950 495.000 354.600 495.600 ;
        RECT 344.400 494.400 354.600 495.000 ;
        RECT 250.950 491.400 270.600 492.600 ;
        RECT 281.400 492.000 291.600 492.600 ;
        RECT 292.950 492.000 334.050 492.600 ;
        RECT 281.400 491.400 292.050 492.000 ;
        RECT 250.950 490.950 253.050 491.400 ;
        RECT 259.950 489.600 262.050 489.900 ;
        RECT 245.400 488.400 262.050 489.600 ;
        RECT 226.950 487.950 229.050 488.400 ;
        RECT 238.950 487.800 241.050 488.400 ;
        RECT 259.950 487.800 262.050 488.400 ;
        RECT 34.950 486.600 37.050 487.050 ;
        RECT 46.950 486.600 49.050 487.050 ;
        RECT 34.950 485.400 49.050 486.600 ;
        RECT 83.400 485.400 88.050 487.050 ;
        RECT 256.950 486.600 259.050 487.050 ;
        RECT 34.950 484.950 37.050 485.400 ;
        RECT 46.950 484.950 49.050 485.400 ;
        RECT 84.000 484.950 88.050 485.400 ;
        RECT 245.400 485.400 259.050 486.600 ;
        RECT 269.400 486.600 270.600 491.400 ;
        RECT 271.950 489.450 274.050 489.900 ;
        RECT 280.950 489.450 283.050 489.900 ;
        RECT 271.950 488.250 283.050 489.450 ;
        RECT 271.950 487.800 274.050 488.250 ;
        RECT 280.950 487.800 283.050 488.250 ;
        RECT 289.950 487.950 292.050 491.400 ;
        RECT 292.950 491.400 333.600 492.000 ;
        RECT 335.400 491.400 351.600 492.600 ;
        RECT 292.950 490.950 295.050 491.400 ;
        RECT 295.950 489.450 298.050 489.900 ;
        RECT 301.950 489.450 304.050 489.900 ;
        RECT 295.950 488.250 304.050 489.450 ;
        RECT 295.950 487.800 298.050 488.250 ;
        RECT 301.950 487.800 304.050 488.250 ;
        RECT 322.950 489.600 325.050 489.900 ;
        RECT 335.400 489.600 336.600 491.400 ;
        RECT 350.400 489.900 351.600 491.400 ;
        RECT 353.400 490.050 354.600 494.400 ;
        RECT 355.950 494.400 370.050 495.600 ;
        RECT 355.950 493.950 358.050 494.400 ;
        RECT 367.950 494.100 370.050 494.400 ;
        RECT 385.950 495.600 388.050 496.050 ;
        RECT 394.950 495.600 397.050 496.200 ;
        RECT 385.950 494.400 397.050 495.600 ;
        RECT 385.950 493.950 388.050 494.400 ;
        RECT 394.950 494.100 397.050 494.400 ;
        RECT 427.950 495.750 430.050 496.200 ;
        RECT 439.950 495.750 442.050 496.200 ;
        RECT 427.950 495.600 442.050 495.750 ;
        RECT 454.950 495.600 457.050 496.200 ;
        RECT 472.950 495.600 475.050 496.200 ;
        RECT 427.950 494.550 475.050 495.600 ;
        RECT 427.950 494.100 430.050 494.550 ;
        RECT 439.950 494.400 475.050 494.550 ;
        RECT 439.950 494.100 442.050 494.400 ;
        RECT 454.950 494.100 457.050 494.400 ;
        RECT 472.950 494.100 475.050 494.400 ;
        RECT 505.950 495.600 508.050 496.050 ;
        RECT 523.950 495.600 526.050 496.050 ;
        RECT 505.950 494.400 526.050 495.600 ;
        RECT 505.950 493.950 508.050 494.400 ;
        RECT 523.950 493.950 526.050 494.400 ;
        RECT 559.950 493.950 562.050 496.050 ;
        RECT 598.950 495.600 601.050 496.200 ;
        RECT 604.950 495.600 607.050 499.050 ;
        RECT 610.950 498.600 613.050 499.050 ;
        RECT 616.950 498.600 619.050 499.050 ;
        RECT 610.950 497.400 619.050 498.600 ;
        RECT 610.950 496.950 613.050 497.400 ;
        RECT 616.950 496.950 619.050 497.400 ;
        RECT 658.950 498.600 661.050 499.050 ;
        RECT 664.950 498.600 667.050 499.050 ;
        RECT 658.950 497.400 667.050 498.600 ;
        RECT 658.950 496.950 661.050 497.400 ;
        RECT 664.950 496.950 667.050 497.400 ;
        RECT 730.950 498.600 733.050 499.050 ;
        RECT 745.950 498.600 748.050 499.050 ;
        RECT 730.950 497.400 748.050 498.600 ;
        RECT 730.950 496.950 733.050 497.400 ;
        RECT 745.950 496.950 748.050 497.400 ;
        RECT 796.950 498.600 799.050 499.050 ;
        RECT 823.950 498.600 826.050 499.050 ;
        RECT 832.950 498.600 835.050 499.050 ;
        RECT 796.950 497.400 835.050 498.600 ;
        RECT 796.950 496.950 799.050 497.400 ;
        RECT 823.950 496.950 826.050 497.400 ;
        RECT 832.950 496.950 835.050 497.400 ;
        RECT 931.950 498.600 934.050 499.050 ;
        RECT 937.950 498.600 940.050 499.050 ;
        RECT 931.950 497.400 940.050 498.600 ;
        RECT 931.950 496.950 934.050 497.400 ;
        RECT 937.950 496.950 940.050 497.400 ;
        RECT 598.950 495.000 607.050 495.600 ;
        RECT 625.950 495.600 628.050 496.200 ;
        RECT 673.950 495.600 676.050 496.050 ;
        RECT 751.950 495.600 754.050 496.200 ;
        RECT 763.950 495.600 766.050 496.050 ;
        RECT 598.950 494.400 606.600 495.000 ;
        RECT 625.950 494.400 678.600 495.600 ;
        RECT 751.950 494.400 766.050 495.600 ;
        RECT 598.950 494.100 601.050 494.400 ;
        RECT 625.950 494.100 628.050 494.400 ;
        RECT 560.400 490.050 561.600 493.950 ;
        RECT 626.400 492.600 627.600 494.100 ;
        RECT 673.950 493.950 676.050 494.400 ;
        RECT 751.950 494.100 754.050 494.400 ;
        RECT 596.400 491.400 627.600 492.600 ;
        RECT 322.950 488.400 336.600 489.600 ;
        RECT 337.950 489.450 340.050 489.900 ;
        RECT 343.950 489.450 346.050 489.900 ;
        RECT 322.950 487.800 325.050 488.400 ;
        RECT 337.950 488.250 346.050 489.450 ;
        RECT 337.950 487.800 340.050 488.250 ;
        RECT 343.950 487.800 346.050 488.250 ;
        RECT 349.950 487.800 352.050 489.900 ;
        RECT 353.400 488.400 358.050 490.050 ;
        RECT 354.000 487.950 358.050 488.400 ;
        RECT 376.950 489.450 379.050 489.900 ;
        RECT 385.950 489.450 388.050 489.900 ;
        RECT 376.950 488.250 388.050 489.450 ;
        RECT 376.950 487.800 379.050 488.250 ;
        RECT 385.950 487.800 388.050 488.250 ;
        RECT 397.950 489.450 400.050 489.900 ;
        RECT 421.950 489.450 424.050 489.900 ;
        RECT 397.950 488.250 424.050 489.450 ;
        RECT 397.950 487.800 400.050 488.250 ;
        RECT 421.950 487.800 424.050 488.250 ;
        RECT 487.950 489.600 490.050 490.050 ;
        RECT 517.950 489.600 520.050 489.900 ;
        RECT 487.950 488.400 520.050 489.600 ;
        RECT 487.950 487.950 490.050 488.400 ;
        RECT 517.950 487.800 520.050 488.400 ;
        RECT 559.950 487.950 562.050 490.050 ;
        RECT 583.950 489.600 586.050 490.050 ;
        RECT 589.950 489.600 592.050 490.050 ;
        RECT 596.400 489.900 597.600 491.400 ;
        RECT 583.950 488.400 592.050 489.600 ;
        RECT 583.950 487.950 586.050 488.400 ;
        RECT 589.950 487.950 592.050 488.400 ;
        RECT 595.950 487.800 598.050 489.900 ;
        RECT 622.950 489.600 625.050 489.900 ;
        RECT 658.950 489.600 661.050 489.900 ;
        RECT 682.950 489.600 685.050 489.900 ;
        RECT 622.950 488.400 685.050 489.600 ;
        RECT 622.950 487.800 625.050 488.400 ;
        RECT 658.950 487.800 661.050 488.400 ;
        RECT 682.950 487.800 685.050 488.400 ;
        RECT 730.950 489.600 733.050 489.900 ;
        RECT 748.950 489.600 751.050 489.900 ;
        RECT 730.950 488.400 751.050 489.600 ;
        RECT 755.400 489.600 756.600 494.400 ;
        RECT 763.950 493.950 766.050 494.400 ;
        RECT 775.950 495.600 778.050 496.200 ;
        RECT 790.950 495.600 793.050 496.200 ;
        RECT 775.950 494.400 793.050 495.600 ;
        RECT 775.950 494.100 778.050 494.400 ;
        RECT 790.950 494.100 793.050 494.400 ;
        RECT 805.950 495.600 808.050 496.050 ;
        RECT 814.950 495.600 817.050 496.200 ;
        RECT 805.950 494.400 817.050 495.600 ;
        RECT 805.950 493.950 808.050 494.400 ;
        RECT 814.950 494.100 817.050 494.400 ;
        RECT 838.950 495.600 841.050 496.200 ;
        RECT 838.950 494.400 843.600 495.600 ;
        RECT 838.950 494.100 841.050 494.400 ;
        RECT 842.400 490.050 843.600 494.400 ;
        RECT 850.950 494.100 853.050 496.200 ;
        RECT 851.400 490.050 852.600 494.100 ;
        RECT 859.950 493.950 862.050 496.050 ;
        RECT 865.950 493.950 868.050 496.050 ;
        RECT 877.950 495.600 880.050 496.200 ;
        RECT 883.950 495.600 886.050 496.050 ;
        RECT 877.950 494.400 886.050 495.600 ;
        RECT 877.950 494.100 880.050 494.400 ;
        RECT 883.950 493.950 886.050 494.400 ;
        RECT 889.950 495.600 892.050 496.050 ;
        RECT 907.950 495.600 910.050 496.050 ;
        RECT 889.950 494.400 910.050 495.600 ;
        RECT 889.950 493.950 892.050 494.400 ;
        RECT 907.950 493.950 910.050 494.400 ;
        RECT 913.950 493.950 916.050 496.050 ;
        RECT 925.950 493.950 928.050 496.050 ;
        RECT 766.950 489.600 769.050 489.900 ;
        RECT 755.400 488.400 769.050 489.600 ;
        RECT 730.950 487.800 733.050 488.400 ;
        RECT 748.950 487.800 751.050 488.400 ;
        RECT 766.950 487.800 769.050 488.400 ;
        RECT 817.950 489.450 820.050 489.900 ;
        RECT 823.950 489.450 826.050 489.900 ;
        RECT 817.950 488.250 826.050 489.450 ;
        RECT 817.950 487.800 820.050 488.250 ;
        RECT 823.950 487.800 826.050 488.250 ;
        RECT 841.950 487.950 844.050 490.050 ;
        RECT 847.950 488.400 852.600 490.050 ;
        RECT 853.950 489.600 856.050 489.900 ;
        RECT 860.400 489.600 861.600 493.950 ;
        RECT 866.400 490.050 867.600 493.950 ;
        RECT 853.950 488.400 861.600 489.600 ;
        RECT 847.950 487.950 852.000 488.400 ;
        RECT 853.950 487.800 856.050 488.400 ;
        RECT 865.950 487.950 868.050 490.050 ;
        RECT 286.950 486.600 289.050 487.050 ;
        RECT 269.400 485.400 289.050 486.600 ;
        RECT 46.950 483.600 49.050 483.900 ;
        RECT 61.950 483.600 64.050 484.050 ;
        RECT 46.950 482.400 64.050 483.600 ;
        RECT 46.950 481.800 49.050 482.400 ;
        RECT 61.950 481.950 64.050 482.400 ;
        RECT 124.950 483.600 127.050 484.050 ;
        RECT 136.950 483.600 139.050 484.050 ;
        RECT 124.950 482.400 139.050 483.600 ;
        RECT 124.950 481.950 127.050 482.400 ;
        RECT 136.950 481.950 139.050 482.400 ;
        RECT 175.950 483.600 178.050 484.050 ;
        RECT 245.400 483.600 246.600 485.400 ;
        RECT 256.950 484.950 259.050 485.400 ;
        RECT 286.950 484.950 289.050 485.400 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 394.950 486.600 397.050 487.050 ;
        RECT 370.950 485.400 397.050 486.600 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 394.950 484.950 397.050 485.400 ;
        RECT 418.950 486.600 421.050 487.050 ;
        RECT 472.950 486.600 475.050 487.050 ;
        RECT 511.950 486.600 514.050 487.050 ;
        RECT 418.950 485.400 514.050 486.600 ;
        RECT 418.950 484.950 421.050 485.400 ;
        RECT 472.950 484.950 475.050 485.400 ;
        RECT 511.950 484.950 514.050 485.400 ;
        RECT 520.950 486.600 523.050 487.050 ;
        RECT 526.950 486.600 529.050 487.050 ;
        RECT 532.950 486.600 535.050 487.050 ;
        RECT 520.950 485.400 535.050 486.600 ;
        RECT 520.950 484.950 523.050 485.400 ;
        RECT 526.950 484.950 529.050 485.400 ;
        RECT 532.950 484.950 535.050 485.400 ;
        RECT 778.950 486.600 781.050 487.050 ;
        RECT 793.950 486.600 796.050 487.050 ;
        RECT 778.950 485.400 796.050 486.600 ;
        RECT 778.950 484.950 781.050 485.400 ;
        RECT 793.950 484.950 796.050 485.400 ;
        RECT 868.950 486.600 871.050 487.050 ;
        RECT 889.950 486.600 892.050 486.900 ;
        RECT 907.950 486.600 910.050 487.050 ;
        RECT 868.950 485.400 910.050 486.600 ;
        RECT 914.400 486.600 915.600 493.950 ;
        RECT 926.400 489.600 927.600 493.950 ;
        RECT 937.950 489.600 940.050 489.900 ;
        RECT 926.400 488.400 940.050 489.600 ;
        RECT 937.950 487.800 940.050 488.400 ;
        RECT 919.950 486.600 922.050 487.050 ;
        RECT 914.400 485.400 922.050 486.600 ;
        RECT 868.950 484.950 871.050 485.400 ;
        RECT 889.950 484.800 892.050 485.400 ;
        RECT 907.950 484.950 910.050 485.400 ;
        RECT 919.950 484.950 922.050 485.400 ;
        RECT 175.950 482.400 246.600 483.600 ;
        RECT 247.950 483.600 250.050 484.050 ;
        RECT 253.950 483.600 256.050 484.050 ;
        RECT 247.950 482.400 256.050 483.600 ;
        RECT 175.950 481.950 178.050 482.400 ;
        RECT 247.950 481.950 250.050 482.400 ;
        RECT 253.950 481.950 256.050 482.400 ;
        RECT 286.950 483.600 289.050 483.900 ;
        RECT 292.950 483.600 295.050 484.050 ;
        RECT 406.950 483.600 409.050 484.050 ;
        RECT 286.950 482.400 295.050 483.600 ;
        RECT 286.950 481.800 289.050 482.400 ;
        RECT 292.950 481.950 295.050 482.400 ;
        RECT 389.400 482.400 409.050 483.600 ;
        RECT 16.950 480.600 19.050 481.050 ;
        RECT 67.950 480.600 70.050 481.050 ;
        RECT 214.950 480.600 217.050 481.050 ;
        RECT 16.950 479.400 70.050 480.600 ;
        RECT 16.950 478.950 19.050 479.400 ;
        RECT 67.950 478.950 70.050 479.400 ;
        RECT 173.400 479.400 217.050 480.600 ;
        RECT 173.400 478.050 174.600 479.400 ;
        RECT 214.950 478.950 217.050 479.400 ;
        RECT 340.950 480.600 343.050 481.050 ;
        RECT 389.400 480.600 390.600 482.400 ;
        RECT 406.950 481.950 409.050 482.400 ;
        RECT 460.950 483.600 463.050 484.050 ;
        RECT 466.950 483.600 469.050 484.050 ;
        RECT 493.950 483.600 496.050 484.050 ;
        RECT 505.950 483.600 508.050 484.050 ;
        RECT 460.950 482.400 508.050 483.600 ;
        RECT 460.950 481.950 463.050 482.400 ;
        RECT 466.950 481.950 469.050 482.400 ;
        RECT 493.950 481.950 496.050 482.400 ;
        RECT 505.950 481.950 508.050 482.400 ;
        RECT 544.950 483.600 547.050 484.050 ;
        RECT 556.950 483.600 559.050 484.050 ;
        RECT 571.950 483.600 574.050 484.050 ;
        RECT 544.950 482.400 574.050 483.600 ;
        RECT 544.950 481.950 547.050 482.400 ;
        RECT 556.950 481.950 559.050 482.400 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 580.950 483.600 583.050 484.050 ;
        RECT 601.950 483.600 604.050 484.050 ;
        RECT 622.950 483.600 625.050 484.050 ;
        RECT 580.950 482.400 625.050 483.600 ;
        RECT 580.950 481.950 583.050 482.400 ;
        RECT 601.950 481.950 604.050 482.400 ;
        RECT 622.950 481.950 625.050 482.400 ;
        RECT 631.950 483.600 634.050 484.050 ;
        RECT 637.950 483.600 640.050 484.050 ;
        RECT 631.950 482.400 640.050 483.600 ;
        RECT 631.950 481.950 634.050 482.400 ;
        RECT 637.950 481.950 640.050 482.400 ;
        RECT 667.950 483.600 670.050 484.050 ;
        RECT 724.950 483.600 727.050 484.050 ;
        RECT 667.950 482.400 727.050 483.600 ;
        RECT 667.950 481.950 670.050 482.400 ;
        RECT 724.950 481.950 727.050 482.400 ;
        RECT 811.950 483.600 814.050 484.050 ;
        RECT 820.950 483.600 823.050 484.050 ;
        RECT 811.950 482.400 823.050 483.600 ;
        RECT 890.400 483.600 891.600 484.800 ;
        RECT 916.950 483.600 919.050 484.050 ;
        RECT 890.400 482.400 919.050 483.600 ;
        RECT 811.950 481.950 814.050 482.400 ;
        RECT 820.950 481.950 823.050 482.400 ;
        RECT 916.950 481.950 919.050 482.400 ;
        RECT 340.950 479.400 390.600 480.600 ;
        RECT 391.950 480.600 394.050 481.050 ;
        RECT 442.950 480.600 445.050 481.050 ;
        RECT 391.950 479.400 445.050 480.600 ;
        RECT 340.950 478.950 343.050 479.400 ;
        RECT 391.950 478.950 394.050 479.400 ;
        RECT 442.950 478.950 445.050 479.400 ;
        RECT 523.950 480.600 526.050 481.050 ;
        RECT 538.950 480.600 541.050 481.050 ;
        RECT 523.950 479.400 541.050 480.600 ;
        RECT 523.950 478.950 526.050 479.400 ;
        RECT 538.950 478.950 541.050 479.400 ;
        RECT 565.950 480.600 568.050 481.050 ;
        RECT 628.950 480.600 631.050 481.050 ;
        RECT 565.950 479.400 631.050 480.600 ;
        RECT 565.950 478.950 568.050 479.400 ;
        RECT 628.950 478.950 631.050 479.400 ;
        RECT 670.950 480.600 673.050 481.050 ;
        RECT 691.950 480.600 694.050 481.050 ;
        RECT 670.950 479.400 694.050 480.600 ;
        RECT 670.950 478.950 673.050 479.400 ;
        RECT 691.950 478.950 694.050 479.400 ;
        RECT 841.950 480.600 844.050 481.050 ;
        RECT 922.950 480.600 925.050 481.050 ;
        RECT 943.950 480.600 946.050 481.050 ;
        RECT 841.950 479.400 946.050 480.600 ;
        RECT 841.950 478.950 844.050 479.400 ;
        RECT 922.950 478.950 925.050 479.400 ;
        RECT 943.950 478.950 946.050 479.400 ;
        RECT 70.950 477.600 73.050 478.050 ;
        RECT 130.950 477.600 133.050 478.050 ;
        RECT 70.950 476.400 133.050 477.600 ;
        RECT 70.950 475.950 73.050 476.400 ;
        RECT 130.950 475.950 133.050 476.400 ;
        RECT 145.950 477.600 148.050 478.050 ;
        RECT 172.950 477.600 175.050 478.050 ;
        RECT 145.950 476.400 175.050 477.600 ;
        RECT 145.950 475.950 148.050 476.400 ;
        RECT 172.950 475.950 175.050 476.400 ;
        RECT 232.950 477.600 235.050 478.050 ;
        RECT 280.950 477.600 283.050 478.050 ;
        RECT 232.950 476.400 283.050 477.600 ;
        RECT 232.950 475.950 235.050 476.400 ;
        RECT 280.950 475.950 283.050 476.400 ;
        RECT 460.950 477.600 463.050 478.050 ;
        RECT 514.950 477.600 517.050 478.050 ;
        RECT 460.950 476.400 517.050 477.600 ;
        RECT 460.950 475.950 463.050 476.400 ;
        RECT 514.950 475.950 517.050 476.400 ;
        RECT 610.950 477.600 613.050 478.050 ;
        RECT 637.950 477.600 640.050 478.050 ;
        RECT 610.950 476.400 640.050 477.600 ;
        RECT 610.950 475.950 613.050 476.400 ;
        RECT 637.950 475.950 640.050 476.400 ;
        RECT 646.950 477.600 649.050 478.050 ;
        RECT 655.950 477.600 658.050 478.050 ;
        RECT 688.950 477.600 691.050 478.050 ;
        RECT 862.950 477.600 865.050 478.050 ;
        RECT 646.950 476.400 691.050 477.600 ;
        RECT 646.950 475.950 649.050 476.400 ;
        RECT 655.950 475.950 658.050 476.400 ;
        RECT 688.950 475.950 691.050 476.400 ;
        RECT 845.400 476.400 865.050 477.600 ;
        RECT 67.950 474.600 70.050 475.050 ;
        RECT 91.950 474.600 94.050 475.050 ;
        RECT 67.950 473.400 94.050 474.600 ;
        RECT 67.950 472.950 70.050 473.400 ;
        RECT 91.950 472.950 94.050 473.400 ;
        RECT 136.950 474.600 139.050 475.050 ;
        RECT 175.950 474.600 178.050 475.050 ;
        RECT 136.950 473.400 178.050 474.600 ;
        RECT 136.950 472.950 139.050 473.400 ;
        RECT 175.950 472.950 178.050 473.400 ;
        RECT 187.950 474.600 190.050 475.050 ;
        RECT 358.950 474.600 361.050 475.050 ;
        RECT 187.950 473.400 361.050 474.600 ;
        RECT 187.950 472.950 190.050 473.400 ;
        RECT 358.950 472.950 361.050 473.400 ;
        RECT 463.950 474.600 466.050 475.050 ;
        RECT 517.950 474.600 520.050 475.050 ;
        RECT 559.950 474.600 562.050 475.050 ;
        RECT 583.950 474.600 586.050 475.050 ;
        RECT 463.950 473.400 513.600 474.600 ;
        RECT 463.950 472.950 466.050 473.400 ;
        RECT 64.950 471.600 67.050 472.050 ;
        RECT 109.950 471.600 112.050 472.050 ;
        RECT 64.950 470.400 112.050 471.600 ;
        RECT 64.950 469.950 67.050 470.400 ;
        RECT 109.950 469.950 112.050 470.400 ;
        RECT 205.950 471.600 208.050 472.050 ;
        RECT 226.950 471.600 229.050 472.050 ;
        RECT 205.950 470.400 229.050 471.600 ;
        RECT 205.950 469.950 208.050 470.400 ;
        RECT 226.950 469.950 229.050 470.400 ;
        RECT 241.950 471.600 244.050 472.050 ;
        RECT 295.950 471.600 298.050 472.050 ;
        RECT 241.950 470.400 298.050 471.600 ;
        RECT 241.950 469.950 244.050 470.400 ;
        RECT 295.950 469.950 298.050 470.400 ;
        RECT 364.950 471.600 367.050 472.050 ;
        RECT 469.950 471.600 472.050 472.050 ;
        RECT 364.950 470.400 472.050 471.600 ;
        RECT 512.400 471.600 513.600 473.400 ;
        RECT 517.950 473.400 586.050 474.600 ;
        RECT 517.950 472.950 520.050 473.400 ;
        RECT 559.950 472.950 562.050 473.400 ;
        RECT 583.950 472.950 586.050 473.400 ;
        RECT 772.950 474.600 775.050 475.050 ;
        RECT 790.950 474.600 793.050 475.050 ;
        RECT 772.950 473.400 793.050 474.600 ;
        RECT 772.950 472.950 775.050 473.400 ;
        RECT 790.950 472.950 793.050 473.400 ;
        RECT 817.950 474.600 820.050 475.050 ;
        RECT 845.400 474.600 846.600 476.400 ;
        RECT 862.950 475.950 865.050 476.400 ;
        RECT 904.950 477.600 907.050 478.050 ;
        RECT 916.950 477.600 919.050 478.050 ;
        RECT 904.950 476.400 919.050 477.600 ;
        RECT 904.950 475.950 907.050 476.400 ;
        RECT 916.950 475.950 919.050 476.400 ;
        RECT 817.950 473.400 846.600 474.600 ;
        RECT 892.950 474.600 895.050 475.050 ;
        RECT 928.950 474.600 931.050 475.050 ;
        RECT 892.950 473.400 931.050 474.600 ;
        RECT 817.950 472.950 820.050 473.400 ;
        RECT 892.950 472.950 895.050 473.400 ;
        RECT 928.950 472.950 931.050 473.400 ;
        RECT 568.950 471.600 571.050 472.050 ;
        RECT 760.950 471.600 763.050 472.050 ;
        RECT 910.950 471.600 913.050 472.050 ;
        RECT 512.400 470.400 516.600 471.600 ;
        RECT 364.950 469.950 367.050 470.400 ;
        RECT 469.950 469.950 472.050 470.400 ;
        RECT 7.950 468.600 10.050 469.050 ;
        RECT 106.950 468.600 109.050 469.050 ;
        RECT 178.950 468.600 181.050 469.050 ;
        RECT 7.950 467.400 109.050 468.600 ;
        RECT 7.950 466.950 10.050 467.400 ;
        RECT 106.950 466.950 109.050 467.400 ;
        RECT 131.400 467.400 181.050 468.600 ;
        RECT 131.400 466.050 132.600 467.400 ;
        RECT 178.950 466.950 181.050 467.400 ;
        RECT 196.950 468.600 199.050 469.050 ;
        RECT 202.950 468.600 205.050 469.050 ;
        RECT 238.950 468.600 241.050 469.050 ;
        RECT 328.950 468.600 331.050 469.050 ;
        RECT 196.950 467.400 331.050 468.600 ;
        RECT 196.950 466.950 199.050 467.400 ;
        RECT 202.950 466.950 205.050 467.400 ;
        RECT 238.950 466.950 241.050 467.400 ;
        RECT 328.950 466.950 331.050 467.400 ;
        RECT 484.950 468.600 487.050 469.050 ;
        RECT 490.950 468.600 493.050 469.050 ;
        RECT 484.950 467.400 493.050 468.600 ;
        RECT 515.400 468.600 516.600 470.400 ;
        RECT 568.950 470.400 913.050 471.600 ;
        RECT 568.950 469.950 571.050 470.400 ;
        RECT 760.950 469.950 763.050 470.400 ;
        RECT 910.950 469.950 913.050 470.400 ;
        RECT 916.950 471.600 919.050 472.050 ;
        RECT 937.950 471.600 940.050 472.050 ;
        RECT 916.950 470.400 940.050 471.600 ;
        RECT 916.950 469.950 919.050 470.400 ;
        RECT 937.950 469.950 940.050 470.400 ;
        RECT 553.950 468.600 556.050 469.050 ;
        RECT 515.400 467.400 556.050 468.600 ;
        RECT 484.950 466.950 487.050 467.400 ;
        RECT 490.950 466.950 493.050 467.400 ;
        RECT 553.950 466.950 556.050 467.400 ;
        RECT 802.950 468.600 805.050 469.050 ;
        RECT 871.950 468.600 874.050 469.050 ;
        RECT 802.950 467.400 874.050 468.600 ;
        RECT 802.950 466.950 805.050 467.400 ;
        RECT 871.950 466.950 874.050 467.400 ;
        RECT 913.950 468.600 916.050 469.050 ;
        RECT 946.950 468.600 949.050 469.050 ;
        RECT 913.950 467.400 949.050 468.600 ;
        RECT 913.950 466.950 916.050 467.400 ;
        RECT 946.950 466.950 949.050 467.400 ;
        RECT 4.950 465.600 7.050 466.050 ;
        RECT 19.950 465.600 22.050 466.050 ;
        RECT 4.950 464.400 22.050 465.600 ;
        RECT 4.950 463.950 7.050 464.400 ;
        RECT 19.950 463.950 22.050 464.400 ;
        RECT 115.950 465.600 118.050 466.050 ;
        RECT 130.950 465.600 133.050 466.050 ;
        RECT 115.950 464.400 133.050 465.600 ;
        RECT 115.950 463.950 118.050 464.400 ;
        RECT 130.950 463.950 133.050 464.400 ;
        RECT 154.950 465.600 157.050 466.050 ;
        RECT 223.800 465.600 225.900 466.050 ;
        RECT 154.950 464.400 225.900 465.600 ;
        RECT 154.950 463.950 157.050 464.400 ;
        RECT 223.800 463.950 225.900 464.400 ;
        RECT 226.950 465.600 229.050 466.050 ;
        RECT 241.950 465.600 244.050 466.050 ;
        RECT 226.950 464.400 244.050 465.600 ;
        RECT 226.950 463.950 229.050 464.400 ;
        RECT 241.950 463.950 244.050 464.400 ;
        RECT 250.950 465.600 253.050 466.050 ;
        RECT 271.950 465.600 274.050 466.050 ;
        RECT 289.950 465.600 292.050 466.050 ;
        RECT 250.950 464.400 292.050 465.600 ;
        RECT 250.950 463.950 253.050 464.400 ;
        RECT 271.950 463.950 274.050 464.400 ;
        RECT 289.950 463.950 292.050 464.400 ;
        RECT 295.950 465.600 298.050 466.050 ;
        RECT 364.950 465.600 367.050 466.050 ;
        RECT 295.950 464.400 367.050 465.600 ;
        RECT 295.950 463.950 298.050 464.400 ;
        RECT 364.950 463.950 367.050 464.400 ;
        RECT 373.950 465.600 376.050 466.050 ;
        RECT 409.950 465.600 412.050 466.050 ;
        RECT 373.950 464.400 412.050 465.600 ;
        RECT 373.950 463.950 376.050 464.400 ;
        RECT 409.950 463.950 412.050 464.400 ;
        RECT 415.950 465.600 418.050 466.050 ;
        RECT 448.950 465.600 451.050 466.050 ;
        RECT 415.950 464.400 451.050 465.600 ;
        RECT 415.950 463.950 418.050 464.400 ;
        RECT 448.950 463.950 451.050 464.400 ;
        RECT 475.950 465.600 478.050 466.050 ;
        RECT 508.950 465.600 511.050 466.050 ;
        RECT 475.950 464.400 511.050 465.600 ;
        RECT 475.950 463.950 478.050 464.400 ;
        RECT 508.950 463.950 511.050 464.400 ;
        RECT 514.950 465.600 517.050 466.050 ;
        RECT 526.800 465.600 528.900 466.050 ;
        RECT 514.950 464.400 528.900 465.600 ;
        RECT 514.950 463.950 517.050 464.400 ;
        RECT 526.800 463.950 528.900 464.400 ;
        RECT 529.950 465.600 532.050 466.050 ;
        RECT 538.950 465.600 541.050 466.050 ;
        RECT 529.950 464.400 541.050 465.600 ;
        RECT 529.950 463.950 532.050 464.400 ;
        RECT 538.950 463.950 541.050 464.400 ;
        RECT 607.950 465.600 610.050 466.050 ;
        RECT 649.950 465.600 652.050 466.050 ;
        RECT 607.950 464.400 652.050 465.600 ;
        RECT 607.950 463.950 610.050 464.400 ;
        RECT 649.950 463.950 652.050 464.400 ;
        RECT 775.950 465.600 778.050 466.050 ;
        RECT 781.950 465.600 784.050 466.050 ;
        RECT 793.950 465.600 796.050 466.050 ;
        RECT 775.950 464.400 796.050 465.600 ;
        RECT 775.950 463.950 778.050 464.400 ;
        RECT 781.950 463.950 784.050 464.400 ;
        RECT 793.950 463.950 796.050 464.400 ;
        RECT 76.950 462.600 79.050 463.050 ;
        RECT 94.950 462.600 97.050 463.050 ;
        RECT 76.950 461.400 97.050 462.600 ;
        RECT 76.950 460.950 79.050 461.400 ;
        RECT 94.950 460.950 97.050 461.400 ;
        RECT 106.950 462.600 109.050 463.050 ;
        RECT 367.950 462.600 370.050 463.050 ;
        RECT 385.950 462.600 388.050 463.050 ;
        RECT 106.950 461.400 141.600 462.600 ;
        RECT 106.950 460.950 109.050 461.400 ;
        RECT 4.950 459.600 7.050 460.050 ;
        RECT 40.950 459.600 43.050 460.050 ;
        RECT 4.950 458.400 43.050 459.600 ;
        RECT 4.950 457.950 7.050 458.400 ;
        RECT 40.950 457.950 43.050 458.400 ;
        RECT 103.950 459.600 106.050 460.050 ;
        RECT 136.950 459.600 139.050 460.050 ;
        RECT 103.950 458.400 139.050 459.600 ;
        RECT 140.400 459.600 141.600 461.400 ;
        RECT 367.950 461.400 388.050 462.600 ;
        RECT 367.950 460.950 370.050 461.400 ;
        RECT 385.950 460.950 388.050 461.400 ;
        RECT 511.950 462.600 514.050 463.050 ;
        RECT 550.950 462.600 553.050 463.050 ;
        RECT 565.950 462.600 568.050 463.050 ;
        RECT 646.950 462.600 649.050 463.050 ;
        RECT 652.950 462.600 655.050 463.050 ;
        RECT 511.950 461.400 568.050 462.600 ;
        RECT 511.950 460.950 514.050 461.400 ;
        RECT 550.950 460.950 553.050 461.400 ;
        RECT 565.950 460.950 568.050 461.400 ;
        RECT 620.400 461.400 655.050 462.600 ;
        RECT 620.400 460.050 621.600 461.400 ;
        RECT 646.950 460.950 649.050 461.400 ;
        RECT 652.950 460.950 655.050 461.400 ;
        RECT 700.950 462.600 703.050 463.050 ;
        RECT 712.950 462.600 715.050 463.050 ;
        RECT 700.950 461.400 715.050 462.600 ;
        RECT 700.950 460.950 703.050 461.400 ;
        RECT 712.950 460.950 715.050 461.400 ;
        RECT 760.950 462.600 763.050 463.050 ;
        RECT 766.950 462.600 769.050 463.050 ;
        RECT 760.950 461.400 769.050 462.600 ;
        RECT 760.950 460.950 763.050 461.400 ;
        RECT 766.950 460.950 769.050 461.400 ;
        RECT 886.950 462.600 889.050 463.050 ;
        RECT 907.950 462.600 910.050 463.050 ;
        RECT 886.950 461.400 910.050 462.600 ;
        RECT 886.950 460.950 889.050 461.400 ;
        RECT 907.950 460.950 910.050 461.400 ;
        RECT 205.800 459.600 207.900 460.050 ;
        RECT 140.400 458.400 207.900 459.600 ;
        RECT 103.950 457.950 106.050 458.400 ;
        RECT 136.950 457.950 139.050 458.400 ;
        RECT 205.800 457.950 207.900 458.400 ;
        RECT 208.950 459.600 211.050 460.050 ;
        RECT 250.950 459.600 253.050 460.050 ;
        RECT 208.950 458.400 253.050 459.600 ;
        RECT 208.950 457.950 211.050 458.400 ;
        RECT 250.950 457.950 253.050 458.400 ;
        RECT 379.950 459.600 382.050 460.050 ;
        RECT 463.950 459.600 466.050 460.050 ;
        RECT 379.950 458.400 466.050 459.600 ;
        RECT 379.950 457.950 382.050 458.400 ;
        RECT 463.950 457.950 466.050 458.400 ;
        RECT 469.950 459.600 472.050 460.050 ;
        RECT 487.950 459.600 490.050 460.050 ;
        RECT 469.950 458.400 490.050 459.600 ;
        RECT 469.950 457.950 472.050 458.400 ;
        RECT 487.950 457.950 490.050 458.400 ;
        RECT 514.950 459.600 517.050 460.050 ;
        RECT 535.950 459.600 538.050 460.050 ;
        RECT 514.950 458.400 538.050 459.600 ;
        RECT 514.950 457.950 517.050 458.400 ;
        RECT 535.950 457.950 538.050 458.400 ;
        RECT 586.950 459.600 589.050 460.050 ;
        RECT 619.950 459.600 622.050 460.050 ;
        RECT 586.950 458.400 622.050 459.600 ;
        RECT 586.950 457.950 589.050 458.400 ;
        RECT 619.950 457.950 622.050 458.400 ;
        RECT 628.950 459.600 631.050 460.050 ;
        RECT 658.950 459.600 661.050 460.050 ;
        RECT 628.950 458.400 661.050 459.600 ;
        RECT 628.950 457.950 631.050 458.400 ;
        RECT 658.950 457.950 661.050 458.400 ;
        RECT 673.950 459.600 676.050 460.050 ;
        RECT 787.950 459.600 790.050 460.050 ;
        RECT 796.950 459.600 799.050 460.050 ;
        RECT 673.950 458.400 799.050 459.600 ;
        RECT 673.950 457.950 676.050 458.400 ;
        RECT 787.950 457.950 790.050 458.400 ;
        RECT 796.950 457.950 799.050 458.400 ;
        RECT 805.950 459.600 808.050 460.050 ;
        RECT 880.950 459.600 883.050 460.050 ;
        RECT 900.000 459.600 904.050 460.050 ;
        RECT 805.950 458.400 883.050 459.600 ;
        RECT 805.950 457.950 808.050 458.400 ;
        RECT 880.950 457.950 883.050 458.400 ;
        RECT 899.400 457.950 904.050 459.600 ;
        RECT 166.950 456.600 169.050 457.050 ;
        RECT 196.950 456.600 199.050 457.050 ;
        RECT 166.950 455.400 199.050 456.600 ;
        RECT 166.950 454.950 169.050 455.400 ;
        RECT 196.950 454.950 199.050 455.400 ;
        RECT 358.950 456.600 361.050 457.050 ;
        RECT 382.800 456.600 384.900 457.050 ;
        RECT 358.950 455.400 384.900 456.600 ;
        RECT 358.950 454.950 361.050 455.400 ;
        RECT 382.800 454.950 384.900 455.400 ;
        RECT 385.950 456.600 388.050 457.050 ;
        RECT 412.950 456.600 415.050 457.050 ;
        RECT 385.950 455.400 415.050 456.600 ;
        RECT 385.950 454.950 388.050 455.400 ;
        RECT 412.950 454.950 415.050 455.400 ;
        RECT 508.950 456.600 511.050 457.050 ;
        RECT 568.950 456.600 571.050 457.050 ;
        RECT 508.950 455.400 571.050 456.600 ;
        RECT 508.950 454.950 511.050 455.400 ;
        RECT 568.950 454.950 571.050 455.400 ;
        RECT 577.950 456.600 580.050 457.050 ;
        RECT 592.950 456.600 595.050 457.050 ;
        RECT 577.950 455.400 595.050 456.600 ;
        RECT 577.950 454.950 580.050 455.400 ;
        RECT 592.950 454.950 595.050 455.400 ;
        RECT 598.950 456.600 601.050 457.050 ;
        RECT 625.950 456.600 628.050 457.050 ;
        RECT 598.950 455.400 628.050 456.600 ;
        RECT 598.950 454.950 601.050 455.400 ;
        RECT 625.950 454.950 628.050 455.400 ;
        RECT 706.950 456.600 709.050 457.050 ;
        RECT 739.950 456.600 742.050 457.050 ;
        RECT 706.950 455.400 742.050 456.600 ;
        RECT 706.950 454.950 709.050 455.400 ;
        RECT 739.950 454.950 742.050 455.400 ;
        RECT 745.950 456.600 748.050 457.050 ;
        RECT 766.950 456.600 769.050 457.050 ;
        RECT 745.950 455.400 769.050 456.600 ;
        RECT 745.950 454.950 748.050 455.400 ;
        RECT 766.950 454.950 769.050 455.400 ;
        RECT 853.950 456.600 856.050 457.050 ;
        RECT 899.400 456.600 900.600 457.950 ;
        RECT 853.950 455.400 900.600 456.600 ;
        RECT 853.950 454.950 856.050 455.400 ;
        RECT 13.950 453.600 16.050 454.050 ;
        RECT 25.950 453.600 28.050 454.050 ;
        RECT 13.950 452.400 28.050 453.600 ;
        RECT 13.950 451.950 16.050 452.400 ;
        RECT 25.950 451.950 28.050 452.400 ;
        RECT 40.950 453.600 43.050 454.050 ;
        RECT 49.950 453.600 52.050 454.050 ;
        RECT 100.950 453.600 103.050 454.050 ;
        RECT 40.950 452.400 52.050 453.600 ;
        RECT 40.950 451.950 43.050 452.400 ;
        RECT 49.950 451.950 52.050 452.400 ;
        RECT 83.400 452.400 103.050 453.600 ;
        RECT 19.950 450.600 22.050 451.200 ;
        RECT 28.950 450.750 31.050 451.200 ;
        RECT 34.950 450.750 37.050 451.200 ;
        RECT 19.950 449.400 27.600 450.600 ;
        RECT 19.950 449.100 22.050 449.400 ;
        RECT 26.400 447.600 27.600 449.400 ;
        RECT 28.950 449.550 37.050 450.750 ;
        RECT 28.950 449.100 31.050 449.550 ;
        RECT 34.950 449.100 37.050 449.550 ;
        RECT 58.950 450.750 61.050 451.200 ;
        RECT 67.950 450.750 70.050 451.200 ;
        RECT 58.950 449.550 70.050 450.750 ;
        RECT 58.950 449.100 61.050 449.550 ;
        RECT 67.950 449.100 70.050 449.550 ;
        RECT 83.400 447.600 84.600 452.400 ;
        RECT 100.950 451.950 103.050 452.400 ;
        RECT 118.950 453.600 121.050 454.050 ;
        RECT 118.950 452.400 138.600 453.600 ;
        RECT 118.950 451.950 121.050 452.400 ;
        RECT 137.400 451.200 138.600 452.400 ;
        RECT 250.950 451.950 253.050 454.050 ;
        RECT 421.950 453.600 424.050 454.050 ;
        RECT 436.950 453.600 439.050 454.050 ;
        RECT 421.950 452.400 439.050 453.600 ;
        RECT 421.950 451.950 424.050 452.400 ;
        RECT 436.950 451.950 439.050 452.400 ;
        RECT 526.950 453.600 529.050 454.050 ;
        RECT 547.950 453.600 550.050 454.050 ;
        RECT 526.950 452.400 550.050 453.600 ;
        RECT 526.950 451.950 529.050 452.400 ;
        RECT 547.950 451.950 550.050 452.400 ;
        RECT 622.950 451.950 625.050 454.050 ;
        RECT 916.950 453.600 919.050 454.050 ;
        RECT 916.950 452.400 924.600 453.600 ;
        RECT 916.950 451.950 919.050 452.400 ;
        RECT 85.950 450.600 88.050 451.050 ;
        RECT 118.950 450.600 121.050 451.200 ;
        RECT 124.950 450.600 127.050 451.200 ;
        RECT 85.950 449.400 121.050 450.600 ;
        RECT 85.950 448.950 88.050 449.400 ;
        RECT 118.950 449.100 121.050 449.400 ;
        RECT 122.400 449.400 127.050 450.600 ;
        RECT 26.400 446.400 81.600 447.600 ;
        RECT 83.400 447.000 87.600 447.600 ;
        RECT 83.400 446.400 88.050 447.000 ;
        RECT 16.950 444.600 19.050 444.900 ;
        RECT 28.950 444.600 31.050 445.050 ;
        RECT 16.950 443.400 31.050 444.600 ;
        RECT 16.950 442.800 19.050 443.400 ;
        RECT 28.950 442.950 31.050 443.400 ;
        RECT 46.950 444.600 49.050 445.050 ;
        RECT 55.950 444.600 58.050 444.900 ;
        RECT 46.950 443.400 58.050 444.600 ;
        RECT 46.950 442.950 49.050 443.400 ;
        RECT 55.950 442.800 58.050 443.400 ;
        RECT 67.950 444.600 70.050 445.050 ;
        RECT 80.400 444.900 81.600 446.400 ;
        RECT 73.950 444.600 76.050 444.900 ;
        RECT 67.950 443.400 76.050 444.600 ;
        RECT 67.950 442.950 70.050 443.400 ;
        RECT 73.950 442.800 76.050 443.400 ;
        RECT 79.950 442.800 82.050 444.900 ;
        RECT 85.950 442.950 88.050 446.400 ;
        RECT 97.950 444.600 100.050 444.900 ;
        RECT 112.950 444.600 115.050 448.050 ;
        RECT 122.400 447.600 123.600 449.400 ;
        RECT 124.950 449.100 127.050 449.400 ;
        RECT 136.950 450.750 139.050 451.200 ;
        RECT 145.950 450.750 148.050 451.200 ;
        RECT 136.950 449.550 148.050 450.750 ;
        RECT 202.950 450.600 205.050 451.200 ;
        RECT 136.950 449.100 139.050 449.550 ;
        RECT 145.950 449.100 148.050 449.550 ;
        RECT 182.400 449.400 205.050 450.600 ;
        RECT 97.950 444.000 115.050 444.600 ;
        RECT 116.400 446.400 123.600 447.600 ;
        RECT 157.950 447.600 160.050 448.050 ;
        RECT 182.400 447.600 183.600 449.400 ;
        RECT 202.950 449.100 205.050 449.400 ;
        RECT 214.950 450.750 217.050 451.200 ;
        RECT 220.800 450.750 222.900 451.200 ;
        RECT 214.950 449.550 222.900 450.750 ;
        RECT 214.950 449.100 217.050 449.550 ;
        RECT 220.800 449.100 222.900 449.550 ;
        RECT 223.950 450.750 226.050 451.200 ;
        RECT 229.950 450.750 232.050 451.200 ;
        RECT 223.950 449.550 232.050 450.750 ;
        RECT 223.950 449.100 226.050 449.550 ;
        RECT 229.950 449.100 232.050 449.550 ;
        RECT 235.950 450.750 238.050 451.200 ;
        RECT 241.950 450.750 244.050 451.200 ;
        RECT 235.950 449.550 244.050 450.750 ;
        RECT 235.950 449.100 238.050 449.550 ;
        RECT 241.950 449.100 244.050 449.550 ;
        RECT 247.950 447.600 250.050 451.050 ;
        RECT 157.950 446.400 183.600 447.600 ;
        RECT 218.400 447.000 250.050 447.600 ;
        RECT 218.400 446.400 249.600 447.000 ;
        RECT 97.950 443.400 114.600 444.000 ;
        RECT 97.950 442.800 100.050 443.400 ;
        RECT 103.950 441.600 106.050 442.050 ;
        RECT 116.400 441.600 117.600 446.400 ;
        RECT 157.950 445.950 160.050 446.400 ;
        RECT 127.950 444.600 130.050 444.900 ;
        RECT 148.950 444.600 151.050 444.900 ;
        RECT 127.950 443.400 151.050 444.600 ;
        RECT 127.950 442.800 130.050 443.400 ;
        RECT 148.950 442.800 151.050 443.400 ;
        RECT 169.950 444.600 172.050 444.900 ;
        RECT 173.400 444.600 174.600 446.400 ;
        RECT 169.950 443.400 174.600 444.600 ;
        RECT 196.950 444.450 199.050 444.900 ;
        RECT 205.950 444.450 208.050 444.900 ;
        RECT 169.950 442.800 172.050 443.400 ;
        RECT 196.950 443.250 208.050 444.450 ;
        RECT 196.950 442.800 199.050 443.250 ;
        RECT 205.950 442.800 208.050 443.250 ;
        RECT 218.400 442.050 219.600 446.400 ;
        RECT 220.950 444.600 223.050 445.050 ;
        RECT 251.400 444.900 252.600 451.950 ;
        RECT 259.950 450.750 262.050 451.200 ;
        RECT 265.950 450.750 268.050 451.200 ;
        RECT 259.950 449.550 268.050 450.750 ;
        RECT 259.950 449.100 262.050 449.550 ;
        RECT 265.950 449.100 268.050 449.550 ;
        RECT 271.950 448.950 274.050 451.050 ;
        RECT 322.950 449.100 325.050 451.200 ;
        RECT 226.950 444.600 229.050 444.900 ;
        RECT 220.950 443.400 229.050 444.600 ;
        RECT 220.950 442.950 223.050 443.400 ;
        RECT 226.950 442.800 229.050 443.400 ;
        RECT 232.950 444.450 235.050 444.900 ;
        RECT 238.950 444.450 241.050 444.900 ;
        RECT 232.950 443.250 241.050 444.450 ;
        RECT 232.950 442.800 235.050 443.250 ;
        RECT 238.950 442.800 241.050 443.250 ;
        RECT 250.950 442.800 253.050 444.900 ;
        RECT 256.950 444.600 259.050 444.900 ;
        RECT 272.400 444.600 273.600 448.950 ;
        RECT 323.400 447.600 324.600 449.100 ;
        RECT 379.950 448.950 382.050 451.050 ;
        RECT 391.950 450.750 394.050 451.200 ;
        RECT 397.950 450.750 400.050 451.200 ;
        RECT 391.950 449.550 400.050 450.750 ;
        RECT 391.950 449.100 394.050 449.550 ;
        RECT 397.950 449.100 400.050 449.550 ;
        RECT 403.950 449.100 406.050 451.200 ;
        RECT 290.400 446.400 324.600 447.600 ;
        RECT 256.950 443.400 273.600 444.600 ;
        RECT 283.950 444.600 286.050 445.050 ;
        RECT 290.400 444.600 291.600 446.400 ;
        RECT 302.400 444.900 303.600 446.400 ;
        RECT 283.950 443.400 291.600 444.600 ;
        RECT 256.950 442.800 259.050 443.400 ;
        RECT 283.950 442.950 286.050 443.400 ;
        RECT 301.950 442.800 304.050 444.900 ;
        RECT 313.950 444.600 316.050 445.050 ;
        RECT 325.950 444.600 328.050 444.900 ;
        RECT 313.950 443.400 328.050 444.600 ;
        RECT 313.950 442.950 316.050 443.400 ;
        RECT 325.950 442.800 328.050 443.400 ;
        RECT 355.950 444.600 358.050 445.050 ;
        RECT 361.950 444.600 364.050 444.900 ;
        RECT 380.400 444.600 381.600 448.950 ;
        RECT 404.400 445.050 405.600 449.100 ;
        RECT 412.950 447.600 415.050 451.050 ;
        RECT 427.950 450.750 430.050 451.200 ;
        RECT 433.950 450.750 436.050 451.200 ;
        RECT 427.950 449.550 436.050 450.750 ;
        RECT 427.950 449.100 430.050 449.550 ;
        RECT 433.950 449.100 436.050 449.550 ;
        RECT 439.950 450.600 442.050 451.050 ;
        RECT 445.950 450.600 448.050 451.200 ;
        RECT 439.950 449.400 448.050 450.600 ;
        RECT 439.950 448.950 442.050 449.400 ;
        RECT 445.950 449.100 448.050 449.400 ;
        RECT 505.950 450.600 508.050 451.200 ;
        RECT 523.950 450.600 526.050 451.200 ;
        RECT 505.950 449.400 526.050 450.600 ;
        RECT 505.950 449.100 508.050 449.400 ;
        RECT 523.950 449.100 526.050 449.400 ;
        RECT 472.950 447.600 475.050 448.050 ;
        RECT 412.950 447.000 420.600 447.600 ;
        RECT 413.400 446.400 420.600 447.000 ;
        RECT 382.950 444.600 385.050 444.900 ;
        RECT 355.950 443.400 366.600 444.600 ;
        RECT 380.400 443.400 385.050 444.600 ;
        RECT 404.400 443.400 409.050 445.050 ;
        RECT 419.400 444.900 420.600 446.400 ;
        RECT 464.400 446.400 475.050 447.600 ;
        RECT 464.400 444.900 465.600 446.400 ;
        RECT 472.950 445.950 475.050 446.400 ;
        RECT 478.950 447.600 481.050 448.050 ;
        RECT 496.950 447.600 499.050 448.050 ;
        RECT 478.950 446.400 499.050 447.600 ;
        RECT 478.950 445.950 481.050 446.400 ;
        RECT 496.950 445.950 499.050 446.400 ;
        RECT 524.400 445.050 525.600 449.100 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 571.950 450.600 574.050 451.200 ;
        RECT 595.950 450.600 598.050 451.200 ;
        RECT 571.950 449.400 598.050 450.600 ;
        RECT 571.950 449.100 574.050 449.400 ;
        RECT 595.950 449.100 598.050 449.400 ;
        RECT 601.950 449.100 604.050 451.200 ;
        RECT 355.950 442.950 358.050 443.400 ;
        RECT 361.950 442.800 364.050 443.400 ;
        RECT 103.950 440.400 117.600 441.600 ;
        RECT 139.950 441.600 142.050 442.050 ;
        RECT 145.950 441.600 148.050 442.050 ;
        RECT 139.950 440.400 148.050 441.600 ;
        RECT 103.950 439.950 106.050 440.400 ;
        RECT 139.950 439.950 142.050 440.400 ;
        RECT 145.950 439.950 148.050 440.400 ;
        RECT 214.950 440.400 219.600 442.050 ;
        RECT 265.950 441.600 268.050 442.050 ;
        RECT 277.950 441.600 280.050 442.050 ;
        RECT 265.950 440.400 280.050 441.600 ;
        RECT 214.950 439.950 219.000 440.400 ;
        RECT 265.950 439.950 268.050 440.400 ;
        RECT 277.950 439.950 280.050 440.400 ;
        RECT 292.950 441.600 295.050 442.050 ;
        RECT 301.950 441.600 304.050 441.750 ;
        RECT 319.950 441.600 322.050 442.050 ;
        RECT 292.950 440.400 322.050 441.600 ;
        RECT 365.400 441.600 366.600 443.400 ;
        RECT 382.950 442.800 385.050 443.400 ;
        RECT 405.000 442.950 409.050 443.400 ;
        RECT 418.950 442.800 421.050 444.900 ;
        RECT 436.950 444.450 439.050 444.900 ;
        RECT 442.950 444.450 445.050 444.900 ;
        RECT 436.950 443.250 445.050 444.450 ;
        RECT 436.950 442.800 439.050 443.250 ;
        RECT 442.950 442.800 445.050 443.250 ;
        RECT 463.950 442.800 466.050 444.900 ;
        RECT 520.950 443.400 525.600 445.050 ;
        RECT 526.950 444.600 529.050 444.900 ;
        RECT 536.400 444.600 537.600 448.950 ;
        RECT 550.950 444.600 553.050 444.900 ;
        RECT 526.950 443.400 553.050 444.600 ;
        RECT 520.950 442.950 525.000 443.400 ;
        RECT 526.950 442.800 529.050 443.400 ;
        RECT 550.950 442.800 553.050 443.400 ;
        RECT 565.950 444.450 568.050 444.900 ;
        RECT 574.950 444.450 577.050 444.900 ;
        RECT 565.950 443.250 577.050 444.450 ;
        RECT 565.950 442.800 568.050 443.250 ;
        RECT 574.950 442.800 577.050 443.250 ;
        RECT 580.950 444.600 583.050 444.900 ;
        RECT 602.400 444.600 603.600 449.100 ;
        RECT 623.400 444.900 624.600 451.950 ;
        RECT 625.950 450.600 628.050 451.200 ;
        RECT 652.950 450.600 655.050 451.200 ;
        RECT 667.950 450.600 670.050 451.200 ;
        RECT 625.950 449.400 651.600 450.600 ;
        RECT 625.950 449.100 628.050 449.400 ;
        RECT 650.400 447.600 651.600 449.400 ;
        RECT 652.950 449.400 670.050 450.600 ;
        RECT 652.950 449.100 655.050 449.400 ;
        RECT 667.950 449.100 670.050 449.400 ;
        RECT 676.950 450.600 681.000 451.050 ;
        RECT 682.950 450.600 685.050 451.200 ;
        RECT 709.950 450.600 712.050 451.050 ;
        RECT 718.950 450.600 721.050 451.200 ;
        RECT 676.950 448.950 681.600 450.600 ;
        RECT 682.950 449.400 721.050 450.600 ;
        RECT 682.950 449.100 685.050 449.400 ;
        RECT 709.950 448.950 712.050 449.400 ;
        RECT 718.950 449.100 721.050 449.400 ;
        RECT 754.950 450.750 757.050 451.200 ;
        RECT 784.950 450.750 787.050 451.200 ;
        RECT 754.950 449.550 787.050 450.750 ;
        RECT 817.950 450.600 820.050 451.050 ;
        RECT 754.950 449.100 757.050 449.550 ;
        RECT 784.950 449.100 787.050 449.550 ;
        RECT 809.400 449.400 820.050 450.600 ;
        RECT 680.400 447.600 681.600 448.950 ;
        RECT 809.400 447.600 810.600 449.400 ;
        RECT 817.950 448.950 820.050 449.400 ;
        RECT 826.950 449.100 829.050 451.200 ;
        RECT 841.950 450.750 844.050 451.200 ;
        RECT 853.950 450.750 856.050 451.200 ;
        RECT 841.950 449.550 856.050 450.750 ;
        RECT 841.950 449.100 844.050 449.550 ;
        RECT 853.950 449.100 856.050 449.550 ;
        RECT 859.950 449.100 862.050 451.200 ;
        RECT 629.400 446.400 648.600 447.600 ;
        RECT 650.400 446.400 666.600 447.600 ;
        RECT 680.400 446.400 687.600 447.600 ;
        RECT 629.400 444.900 630.600 446.400 ;
        RECT 616.950 444.600 619.050 444.900 ;
        RECT 580.950 443.400 603.600 444.600 ;
        RECT 608.400 443.400 619.050 444.600 ;
        RECT 580.950 442.800 583.050 443.400 ;
        RECT 379.950 441.600 382.050 442.050 ;
        RECT 365.400 440.400 382.050 441.600 ;
        RECT 292.950 439.950 295.050 440.400 ;
        RECT 301.950 439.650 304.050 440.400 ;
        RECT 319.950 439.950 322.050 440.400 ;
        RECT 379.950 439.950 382.050 440.400 ;
        RECT 394.950 441.600 397.050 442.050 ;
        RECT 418.950 441.600 421.050 442.050 ;
        RECT 394.950 440.400 421.050 441.600 ;
        RECT 394.950 439.950 397.050 440.400 ;
        RECT 418.950 439.950 421.050 440.400 ;
        RECT 469.950 441.600 472.050 442.050 ;
        RECT 475.950 441.600 478.050 442.050 ;
        RECT 469.950 440.400 478.050 441.600 ;
        RECT 469.950 439.950 472.050 440.400 ;
        RECT 475.950 439.950 478.050 440.400 ;
        RECT 598.950 441.600 601.050 442.050 ;
        RECT 608.400 441.600 609.600 443.400 ;
        RECT 616.950 442.800 619.050 443.400 ;
        RECT 622.950 442.800 625.050 444.900 ;
        RECT 628.950 442.800 631.050 444.900 ;
        RECT 643.950 444.600 646.050 444.900 ;
        RECT 638.400 443.400 646.050 444.600 ;
        RECT 598.950 440.400 609.600 441.600 ;
        RECT 616.950 441.600 619.050 442.050 ;
        RECT 638.400 441.600 639.600 443.400 ;
        RECT 643.950 442.800 646.050 443.400 ;
        RECT 647.400 442.050 648.600 446.400 ;
        RECT 665.400 444.900 666.600 446.400 ;
        RECT 686.400 444.900 687.600 446.400 ;
        RECT 806.400 446.400 810.600 447.600 ;
        RECT 664.950 442.800 667.050 444.900 ;
        RECT 685.950 442.800 688.050 444.900 ;
        RECT 697.950 444.450 700.050 444.900 ;
        RECT 709.950 444.450 712.050 444.900 ;
        RECT 697.950 443.250 712.050 444.450 ;
        RECT 697.950 442.800 700.050 443.250 ;
        RECT 709.950 442.800 712.050 443.250 ;
        RECT 721.950 444.600 724.050 444.900 ;
        RECT 733.950 444.600 736.050 445.050 ;
        RECT 742.950 444.600 745.050 444.900 ;
        RECT 721.950 443.400 745.050 444.600 ;
        RECT 721.950 442.800 724.050 443.400 ;
        RECT 733.950 442.950 736.050 443.400 ;
        RECT 742.950 442.800 745.050 443.400 ;
        RECT 793.950 444.600 796.050 445.050 ;
        RECT 806.400 444.600 807.600 446.400 ;
        RECT 827.400 444.600 828.600 449.100 ;
        RECT 793.950 443.400 807.600 444.600 ;
        RECT 815.400 444.000 828.600 444.600 ;
        RECT 814.950 443.400 828.600 444.000 ;
        RECT 860.400 445.050 861.600 449.100 ;
        RECT 871.950 448.950 874.050 451.050 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 860.400 443.400 865.050 445.050 ;
        RECT 793.950 442.950 796.050 443.400 ;
        RECT 616.950 440.400 639.600 441.600 ;
        RECT 598.950 439.950 601.050 440.400 ;
        RECT 616.950 439.950 619.050 440.400 ;
        RECT 646.950 439.950 649.050 442.050 ;
        RECT 658.950 441.600 661.050 442.050 ;
        RECT 658.950 440.400 684.600 441.600 ;
        RECT 658.950 439.950 661.050 440.400 ;
        RECT 178.950 438.600 181.050 439.050 ;
        RECT 211.950 438.600 214.050 439.050 ;
        RECT 178.950 437.400 214.050 438.600 ;
        RECT 178.950 436.950 181.050 437.400 ;
        RECT 211.950 436.950 214.050 437.400 ;
        RECT 226.950 438.600 229.050 439.050 ;
        RECT 247.950 438.600 250.050 439.050 ;
        RECT 226.950 437.400 250.050 438.600 ;
        RECT 226.950 436.950 229.050 437.400 ;
        RECT 247.950 436.950 250.050 437.400 ;
        RECT 256.950 438.600 259.050 439.050 ;
        RECT 286.950 438.600 289.050 439.050 ;
        RECT 256.950 437.400 289.050 438.600 ;
        RECT 256.950 436.950 259.050 437.400 ;
        RECT 286.950 436.950 289.050 437.400 ;
        RECT 400.950 438.600 403.050 439.050 ;
        RECT 475.950 438.600 478.050 438.900 ;
        RECT 520.950 438.600 523.050 439.050 ;
        RECT 400.950 437.400 523.050 438.600 ;
        RECT 400.950 436.950 403.050 437.400 ;
        RECT 475.950 436.800 478.050 437.400 ;
        RECT 520.950 436.950 523.050 437.400 ;
        RECT 541.950 438.600 544.050 439.050 ;
        RECT 547.950 438.600 550.050 439.050 ;
        RECT 541.950 437.400 550.050 438.600 ;
        RECT 541.950 436.950 544.050 437.400 ;
        RECT 547.950 436.950 550.050 437.400 ;
        RECT 574.950 438.600 577.050 439.050 ;
        RECT 580.950 438.600 583.050 439.050 ;
        RECT 574.950 437.400 583.050 438.600 ;
        RECT 574.950 436.950 577.050 437.400 ;
        RECT 580.950 436.950 583.050 437.400 ;
        RECT 592.950 438.600 595.050 439.050 ;
        RECT 610.950 438.600 613.050 439.050 ;
        RECT 592.950 437.400 613.050 438.600 ;
        RECT 683.400 438.600 684.600 440.400 ;
        RECT 814.950 439.950 817.050 443.400 ;
        RECT 861.000 442.950 865.050 443.400 ;
        RECT 820.950 441.600 823.050 442.050 ;
        RECT 835.950 441.600 838.050 442.050 ;
        RECT 820.950 440.400 838.050 441.600 ;
        RECT 820.950 439.950 823.050 440.400 ;
        RECT 835.950 439.950 838.050 440.400 ;
        RECT 844.950 441.600 847.050 442.050 ;
        RECT 856.950 441.600 859.050 442.050 ;
        RECT 844.950 440.400 859.050 441.600 ;
        RECT 872.400 441.600 873.600 448.950 ;
        RECT 883.950 444.600 886.050 444.900 ;
        RECT 889.950 444.600 892.050 445.050 ;
        RECT 883.950 443.400 892.050 444.600 ;
        RECT 893.400 444.600 894.600 448.950 ;
        RECT 907.950 447.600 910.050 451.050 ;
        RECT 907.950 447.000 915.600 447.600 ;
        RECT 908.400 446.400 915.600 447.000 ;
        RECT 901.950 444.600 904.050 444.900 ;
        RECT 893.400 443.400 904.050 444.600 ;
        RECT 914.400 444.600 915.600 446.400 ;
        RECT 923.400 444.900 924.600 452.400 ;
        RECT 925.950 449.100 928.050 451.200 ;
        RECT 916.950 444.600 919.050 444.900 ;
        RECT 914.400 443.400 919.050 444.600 ;
        RECT 883.950 442.800 886.050 443.400 ;
        RECT 889.950 442.950 892.050 443.400 ;
        RECT 901.950 442.800 904.050 443.400 ;
        RECT 916.950 442.800 919.050 443.400 ;
        RECT 922.950 442.800 925.050 444.900 ;
        RECT 880.950 441.600 883.050 442.050 ;
        RECT 872.400 440.400 883.050 441.600 ;
        RECT 844.950 439.950 847.050 440.400 ;
        RECT 856.950 439.950 859.050 440.400 ;
        RECT 880.950 439.950 883.050 440.400 ;
        RECT 919.950 441.600 922.050 442.050 ;
        RECT 926.400 441.600 927.600 449.100 ;
        RECT 934.950 448.950 937.050 451.050 ;
        RECT 919.950 440.400 927.600 441.600 ;
        RECT 935.400 442.050 936.600 448.950 ;
        RECT 935.400 440.400 940.050 442.050 ;
        RECT 919.950 439.950 922.050 440.400 ;
        RECT 936.000 439.950 940.050 440.400 ;
        RECT 703.950 438.600 706.050 439.050 ;
        RECT 727.800 438.600 729.900 439.050 ;
        RECT 683.400 437.400 729.900 438.600 ;
        RECT 592.950 436.950 595.050 437.400 ;
        RECT 610.950 436.950 613.050 437.400 ;
        RECT 703.950 436.950 706.050 437.400 ;
        RECT 727.800 436.950 729.900 437.400 ;
        RECT 730.950 438.600 733.050 439.050 ;
        RECT 748.950 438.600 751.050 439.050 ;
        RECT 730.950 437.400 751.050 438.600 ;
        RECT 730.950 436.950 733.050 437.400 ;
        RECT 748.950 436.950 751.050 437.400 ;
        RECT 778.950 438.600 781.050 439.050 ;
        RECT 787.950 438.600 790.050 439.050 ;
        RECT 778.950 437.400 790.050 438.600 ;
        RECT 778.950 436.950 781.050 437.400 ;
        RECT 787.950 436.950 790.050 437.400 ;
        RECT 925.950 438.600 928.050 439.050 ;
        RECT 946.950 438.600 949.050 439.050 ;
        RECT 925.950 437.400 949.050 438.600 ;
        RECT 925.950 436.950 928.050 437.400 ;
        RECT 946.950 436.950 949.050 437.400 ;
        RECT 49.950 435.600 52.050 436.050 ;
        RECT 58.950 435.600 61.050 436.050 ;
        RECT 49.950 434.400 61.050 435.600 ;
        RECT 49.950 433.950 52.050 434.400 ;
        RECT 58.950 433.950 61.050 434.400 ;
        RECT 217.950 435.600 220.050 436.050 ;
        RECT 283.950 435.600 286.050 436.050 ;
        RECT 217.950 434.400 286.050 435.600 ;
        RECT 217.950 433.950 220.050 434.400 ;
        RECT 283.950 433.950 286.050 434.400 ;
        RECT 310.950 435.600 313.050 436.050 ;
        RECT 334.950 435.600 337.050 436.050 ;
        RECT 310.950 434.400 337.050 435.600 ;
        RECT 310.950 433.950 313.050 434.400 ;
        RECT 334.950 433.950 337.050 434.400 ;
        RECT 412.950 435.600 415.050 436.050 ;
        RECT 451.950 435.600 454.050 436.050 ;
        RECT 412.950 434.400 454.050 435.600 ;
        RECT 412.950 433.950 415.050 434.400 ;
        RECT 451.950 433.950 454.050 434.400 ;
        RECT 457.950 435.600 460.050 436.050 ;
        RECT 469.950 435.600 472.050 436.050 ;
        RECT 457.950 434.400 472.050 435.600 ;
        RECT 457.950 433.950 460.050 434.400 ;
        RECT 469.950 433.950 472.050 434.400 ;
        RECT 487.950 435.600 490.050 436.050 ;
        RECT 517.950 435.600 520.050 436.050 ;
        RECT 487.950 434.400 520.050 435.600 ;
        RECT 487.950 433.950 490.050 434.400 ;
        RECT 517.950 433.950 520.050 434.400 ;
        RECT 562.950 435.600 565.050 436.050 ;
        RECT 571.950 435.600 574.050 436.050 ;
        RECT 562.950 434.400 574.050 435.600 ;
        RECT 562.950 433.950 565.050 434.400 ;
        RECT 571.950 433.950 574.050 434.400 ;
        RECT 634.950 435.600 637.050 436.050 ;
        RECT 679.950 435.600 682.050 436.050 ;
        RECT 634.950 434.400 682.050 435.600 ;
        RECT 634.950 433.950 637.050 434.400 ;
        RECT 679.950 433.950 682.050 434.400 ;
        RECT 742.950 435.600 745.050 436.050 ;
        RECT 754.950 435.600 757.050 436.050 ;
        RECT 742.950 434.400 757.050 435.600 ;
        RECT 742.950 433.950 745.050 434.400 ;
        RECT 754.950 433.950 757.050 434.400 ;
        RECT 838.950 435.600 841.050 436.050 ;
        RECT 874.950 435.600 877.050 436.050 ;
        RECT 838.950 434.400 877.050 435.600 ;
        RECT 838.950 433.950 841.050 434.400 ;
        RECT 874.950 433.950 877.050 434.400 ;
        RECT 883.950 435.600 886.050 436.050 ;
        RECT 940.950 435.600 943.050 436.050 ;
        RECT 883.950 434.400 943.050 435.600 ;
        RECT 883.950 433.950 886.050 434.400 ;
        RECT 940.950 433.950 943.050 434.400 ;
        RECT 37.950 432.600 40.050 433.050 ;
        RECT 85.950 432.600 88.050 433.050 ;
        RECT 37.950 431.400 88.050 432.600 ;
        RECT 37.950 430.950 40.050 431.400 ;
        RECT 85.950 430.950 88.050 431.400 ;
        RECT 94.950 432.600 97.050 433.050 ;
        RECT 121.950 432.600 124.050 433.050 ;
        RECT 94.950 431.400 124.050 432.600 ;
        RECT 94.950 430.950 97.050 431.400 ;
        RECT 121.950 430.950 124.050 431.400 ;
        RECT 160.950 432.600 163.050 433.050 ;
        RECT 181.950 432.600 184.050 433.050 ;
        RECT 160.950 431.400 184.050 432.600 ;
        RECT 160.950 430.950 163.050 431.400 ;
        RECT 181.950 430.950 184.050 431.400 ;
        RECT 193.950 432.600 196.050 433.050 ;
        RECT 229.950 432.600 232.050 433.050 ;
        RECT 193.950 431.400 232.050 432.600 ;
        RECT 193.950 430.950 196.050 431.400 ;
        RECT 229.950 430.950 232.050 431.400 ;
        RECT 268.950 432.600 271.050 433.050 ;
        RECT 292.950 432.600 295.050 433.050 ;
        RECT 349.950 432.600 352.050 433.050 ;
        RECT 376.950 432.600 379.050 433.050 ;
        RECT 268.950 431.400 352.050 432.600 ;
        RECT 268.950 430.950 271.050 431.400 ;
        RECT 292.950 430.950 295.050 431.400 ;
        RECT 349.950 430.950 352.050 431.400 ;
        RECT 356.400 431.400 379.050 432.600 ;
        RECT 88.950 429.600 91.050 430.050 ;
        RECT 127.950 429.600 130.050 430.050 ;
        RECT 88.950 428.400 130.050 429.600 ;
        RECT 88.950 427.950 91.050 428.400 ;
        RECT 127.950 427.950 130.050 428.400 ;
        RECT 295.950 429.600 298.050 430.050 ;
        RECT 356.400 429.600 357.600 431.400 ;
        RECT 376.950 430.950 379.050 431.400 ;
        RECT 442.950 432.600 445.050 433.050 ;
        RECT 478.950 432.600 481.050 433.050 ;
        RECT 442.950 431.400 481.050 432.600 ;
        RECT 442.950 430.950 445.050 431.400 ;
        RECT 478.950 430.950 481.050 431.400 ;
        RECT 490.950 432.600 493.050 433.050 ;
        RECT 502.950 432.600 505.050 433.050 ;
        RECT 490.950 431.400 505.050 432.600 ;
        RECT 490.950 430.950 493.050 431.400 ;
        RECT 502.950 430.950 505.050 431.400 ;
        RECT 508.950 432.600 511.050 433.050 ;
        RECT 538.950 432.600 541.050 433.050 ;
        RECT 508.950 431.400 541.050 432.600 ;
        RECT 508.950 430.950 511.050 431.400 ;
        RECT 538.950 430.950 541.050 431.400 ;
        RECT 562.950 432.600 565.050 432.900 ;
        RECT 604.950 432.600 607.050 433.050 ;
        RECT 562.950 431.400 607.050 432.600 ;
        RECT 562.950 430.800 565.050 431.400 ;
        RECT 604.950 430.950 607.050 431.400 ;
        RECT 790.950 432.600 793.050 433.050 ;
        RECT 829.950 432.600 832.050 433.050 ;
        RECT 790.950 431.400 832.050 432.600 ;
        RECT 790.950 430.950 793.050 431.400 ;
        RECT 829.950 430.950 832.050 431.400 ;
        RECT 865.950 432.600 868.050 433.050 ;
        RECT 884.400 432.600 885.600 433.950 ;
        RECT 865.950 431.400 885.600 432.600 ;
        RECT 865.950 430.950 868.050 431.400 ;
        RECT 295.950 428.400 357.600 429.600 ;
        RECT 436.950 429.600 439.050 430.050 ;
        RECT 460.950 429.600 463.050 430.050 ;
        RECT 436.950 428.400 463.050 429.600 ;
        RECT 295.950 427.950 298.050 428.400 ;
        RECT 436.950 427.950 439.050 428.400 ;
        RECT 460.950 427.950 463.050 428.400 ;
        RECT 556.950 429.600 559.050 430.050 ;
        RECT 607.950 429.600 610.050 430.050 ;
        RECT 556.950 428.400 610.050 429.600 ;
        RECT 556.950 427.950 559.050 428.400 ;
        RECT 607.950 427.950 610.050 428.400 ;
        RECT 679.950 429.600 682.050 430.050 ;
        RECT 691.950 429.600 694.050 430.050 ;
        RECT 679.950 428.400 694.050 429.600 ;
        RECT 679.950 427.950 682.050 428.400 ;
        RECT 691.950 427.950 694.050 428.400 ;
        RECT 712.950 429.600 715.050 430.050 ;
        RECT 763.950 429.600 766.050 430.050 ;
        RECT 712.950 428.400 766.050 429.600 ;
        RECT 712.950 427.950 715.050 428.400 ;
        RECT 763.950 427.950 766.050 428.400 ;
        RECT 109.950 426.600 112.050 427.050 ;
        RECT 211.950 426.600 214.050 427.050 ;
        RECT 109.950 425.400 214.050 426.600 ;
        RECT 109.950 424.950 112.050 425.400 ;
        RECT 211.950 424.950 214.050 425.400 ;
        RECT 229.950 426.600 232.050 427.050 ;
        RECT 289.950 426.600 292.050 427.050 ;
        RECT 367.950 426.600 370.050 427.050 ;
        RECT 229.950 425.400 370.050 426.600 ;
        RECT 229.950 424.950 232.050 425.400 ;
        RECT 289.950 424.950 292.050 425.400 ;
        RECT 367.950 424.950 370.050 425.400 ;
        RECT 376.950 426.600 379.050 427.050 ;
        RECT 382.950 426.600 385.050 427.050 ;
        RECT 376.950 425.400 385.050 426.600 ;
        RECT 376.950 424.950 379.050 425.400 ;
        RECT 382.950 424.950 385.050 425.400 ;
        RECT 418.950 426.600 421.050 427.050 ;
        RECT 490.950 426.600 493.050 427.050 ;
        RECT 418.950 425.400 493.050 426.600 ;
        RECT 418.950 424.950 421.050 425.400 ;
        RECT 490.950 424.950 493.050 425.400 ;
        RECT 496.950 426.600 499.050 427.050 ;
        RECT 505.950 426.600 508.050 427.050 ;
        RECT 496.950 425.400 508.050 426.600 ;
        RECT 496.950 424.950 499.050 425.400 ;
        RECT 505.950 424.950 508.050 425.400 ;
        RECT 532.950 426.600 535.050 427.050 ;
        RECT 550.950 426.600 553.050 427.050 ;
        RECT 532.950 425.400 553.050 426.600 ;
        RECT 532.950 424.950 535.050 425.400 ;
        RECT 550.950 424.950 553.050 425.400 ;
        RECT 580.950 426.600 583.050 427.050 ;
        RECT 631.950 426.600 634.050 427.050 ;
        RECT 580.950 425.400 634.050 426.600 ;
        RECT 580.950 424.950 583.050 425.400 ;
        RECT 631.950 424.950 634.050 425.400 ;
        RECT 649.950 426.600 652.050 427.050 ;
        RECT 655.950 426.600 658.050 427.050 ;
        RECT 649.950 425.400 658.050 426.600 ;
        RECT 649.950 424.950 652.050 425.400 ;
        RECT 655.950 424.950 658.050 425.400 ;
        RECT 685.950 426.600 688.050 427.050 ;
        RECT 700.950 426.600 703.050 427.050 ;
        RECT 685.950 425.400 703.050 426.600 ;
        RECT 685.950 424.950 688.050 425.400 ;
        RECT 700.950 424.950 703.050 425.400 ;
        RECT 829.950 426.600 832.050 427.050 ;
        RECT 841.950 426.600 844.050 427.050 ;
        RECT 829.950 425.400 844.050 426.600 ;
        RECT 829.950 424.950 832.050 425.400 ;
        RECT 841.950 424.950 844.050 425.400 ;
        RECT 856.950 426.600 859.050 427.050 ;
        RECT 871.950 426.600 874.050 427.050 ;
        RECT 856.950 425.400 874.050 426.600 ;
        RECT 856.950 424.950 859.050 425.400 ;
        RECT 871.950 424.950 874.050 425.400 ;
        RECT 910.950 426.600 913.050 427.050 ;
        RECT 922.950 426.600 925.050 427.050 ;
        RECT 910.950 425.400 925.050 426.600 ;
        RECT 910.950 424.950 913.050 425.400 ;
        RECT 922.950 424.950 925.050 425.400 ;
        RECT 40.950 423.600 43.050 424.050 ;
        RECT 133.950 423.600 136.050 424.050 ;
        RECT 40.950 422.400 136.050 423.600 ;
        RECT 40.950 421.950 43.050 422.400 ;
        RECT 133.950 421.950 136.050 422.400 ;
        RECT 157.950 423.600 160.050 424.050 ;
        RECT 175.950 423.600 178.050 424.050 ;
        RECT 301.950 423.600 304.050 424.050 ;
        RECT 157.950 422.400 178.050 423.600 ;
        RECT 157.950 421.950 160.050 422.400 ;
        RECT 175.950 421.950 178.050 422.400 ;
        RECT 293.400 422.400 304.050 423.600 ;
        RECT 142.950 420.600 145.050 421.050 ;
        RECT 154.950 420.600 157.050 421.050 ;
        RECT 163.950 420.600 166.050 421.050 ;
        RECT 142.950 419.400 166.050 420.600 ;
        RECT 142.950 418.950 145.050 419.400 ;
        RECT 154.950 418.950 157.050 419.400 ;
        RECT 163.950 418.950 166.050 419.400 ;
        RECT 274.950 420.600 277.050 421.050 ;
        RECT 293.400 420.600 294.600 422.400 ;
        RECT 301.950 421.950 304.050 422.400 ;
        RECT 424.950 423.600 427.050 424.050 ;
        RECT 463.950 423.600 466.050 424.050 ;
        RECT 424.950 422.400 466.050 423.600 ;
        RECT 424.950 421.950 427.050 422.400 ;
        RECT 463.950 421.950 466.050 422.400 ;
        RECT 469.950 423.600 472.050 424.050 ;
        RECT 481.950 423.600 484.050 424.050 ;
        RECT 469.950 422.400 484.050 423.600 ;
        RECT 469.950 421.950 472.050 422.400 ;
        RECT 481.950 421.950 484.050 422.400 ;
        RECT 496.950 423.600 499.050 423.900 ;
        RECT 511.950 423.600 514.050 424.050 ;
        RECT 496.950 422.400 514.050 423.600 ;
        RECT 496.950 421.800 499.050 422.400 ;
        RECT 511.950 421.950 514.050 422.400 ;
        RECT 523.950 423.600 526.050 424.050 ;
        RECT 553.950 423.600 556.050 424.050 ;
        RECT 523.950 422.400 556.050 423.600 ;
        RECT 523.950 421.950 526.050 422.400 ;
        RECT 553.950 421.950 556.050 422.400 ;
        RECT 604.950 423.600 607.050 424.050 ;
        RECT 634.950 423.600 637.050 424.050 ;
        RECT 643.950 423.600 646.050 424.050 ;
        RECT 604.950 422.400 633.600 423.600 ;
        RECT 604.950 421.950 607.050 422.400 ;
        RECT 274.950 419.400 294.600 420.600 ;
        RECT 316.950 420.600 319.050 421.050 ;
        RECT 325.950 420.600 328.050 421.050 ;
        RECT 316.950 419.400 328.050 420.600 ;
        RECT 274.950 418.950 277.050 419.400 ;
        RECT 316.950 418.950 319.050 419.400 ;
        RECT 325.950 418.950 328.050 419.400 ;
        RECT 406.950 420.600 409.050 421.050 ;
        RECT 472.950 420.600 475.050 421.050 ;
        RECT 406.950 419.400 475.050 420.600 ;
        RECT 406.950 418.950 409.050 419.400 ;
        RECT 16.950 417.750 19.050 418.200 ;
        RECT 31.950 417.750 34.050 418.200 ;
        RECT 16.950 416.550 34.050 417.750 ;
        RECT 16.950 416.100 19.050 416.550 ;
        RECT 31.950 416.100 34.050 416.550 ;
        RECT 46.950 417.600 49.050 418.050 ;
        RECT 64.950 417.600 67.050 418.050 ;
        RECT 76.950 417.600 79.050 418.200 ;
        RECT 46.950 416.400 67.050 417.600 ;
        RECT 46.950 415.950 49.050 416.400 ;
        RECT 64.950 415.950 67.050 416.400 ;
        RECT 71.400 416.400 79.050 417.600 ;
        RECT 71.400 414.600 72.600 416.400 ;
        RECT 76.950 416.100 79.050 416.400 ;
        RECT 85.950 417.600 88.050 418.050 ;
        RECT 94.950 417.600 97.050 418.200 ;
        RECT 85.950 416.400 97.050 417.600 ;
        RECT 85.950 415.950 88.050 416.400 ;
        RECT 94.950 416.100 97.050 416.400 ;
        RECT 106.950 417.750 109.050 418.200 ;
        RECT 115.950 417.750 118.050 418.200 ;
        RECT 106.950 416.550 118.050 417.750 ;
        RECT 106.950 416.100 109.050 416.550 ;
        RECT 115.950 416.100 118.050 416.550 ;
        RECT 121.950 417.600 124.050 418.200 ;
        RECT 151.950 417.600 154.050 418.050 ;
        RECT 121.950 416.400 154.050 417.600 ;
        RECT 121.950 416.100 124.050 416.400 ;
        RECT 151.950 415.950 154.050 416.400 ;
        RECT 199.950 416.100 202.050 418.200 ;
        RECT 211.950 417.750 214.050 418.200 ;
        RECT 220.950 417.750 223.050 418.200 ;
        RECT 211.950 417.600 223.050 417.750 ;
        RECT 238.950 417.600 241.050 418.050 ;
        RECT 265.950 417.750 268.050 418.200 ;
        RECT 271.950 417.750 274.050 418.200 ;
        RECT 211.950 416.550 252.600 417.600 ;
        RECT 211.950 416.100 214.050 416.550 ;
        RECT 220.950 416.400 252.600 416.550 ;
        RECT 220.950 416.100 223.050 416.400 ;
        RECT 62.400 413.400 72.600 414.600 ;
        RECT 62.400 411.900 63.600 413.400 ;
        RECT 22.950 411.600 25.050 411.900 ;
        RECT 55.950 411.600 58.050 411.900 ;
        RECT 22.950 410.400 58.050 411.600 ;
        RECT 22.950 409.800 25.050 410.400 ;
        RECT 55.950 409.800 58.050 410.400 ;
        RECT 61.950 409.800 64.050 411.900 ;
        RECT 187.950 411.600 190.050 412.050 ;
        RECT 200.400 411.600 201.600 416.100 ;
        RECT 238.950 415.950 241.050 416.400 ;
        RECT 251.400 414.600 252.600 416.400 ;
        RECT 265.950 416.550 274.050 417.750 ;
        RECT 265.950 416.100 268.050 416.550 ;
        RECT 271.950 416.100 274.050 416.550 ;
        RECT 295.950 414.600 298.050 418.050 ;
        RECT 328.950 417.750 331.050 418.200 ;
        RECT 334.950 417.750 337.050 418.200 ;
        RECT 328.950 416.550 337.050 417.750 ;
        RECT 328.950 416.100 331.050 416.550 ;
        RECT 334.950 416.100 337.050 416.550 ;
        RECT 349.950 417.750 352.050 418.200 ;
        RECT 355.950 417.750 358.050 418.200 ;
        RECT 349.950 416.550 358.050 417.750 ;
        RECT 379.950 417.600 382.050 418.200 ;
        RECT 349.950 416.100 352.050 416.550 ;
        RECT 355.950 416.100 358.050 416.550 ;
        RECT 359.400 416.400 382.050 417.600 ;
        RECT 359.400 414.600 360.600 416.400 ;
        RECT 379.950 416.100 382.050 416.400 ;
        RECT 424.950 417.600 427.050 418.200 ;
        RECT 439.950 417.750 442.050 418.200 ;
        RECT 445.950 417.750 448.050 418.200 ;
        RECT 439.950 417.600 448.050 417.750 ;
        RECT 424.950 416.550 448.050 417.600 ;
        RECT 424.950 416.400 442.050 416.550 ;
        RECT 424.950 416.100 427.050 416.400 ;
        RECT 439.950 416.100 442.050 416.400 ;
        RECT 445.950 416.100 448.050 416.550 ;
        RECT 451.950 417.600 454.050 418.200 ;
        RECT 460.950 417.600 463.050 418.050 ;
        RECT 451.950 416.400 463.050 417.600 ;
        RECT 464.400 417.600 465.600 419.400 ;
        RECT 472.950 418.950 475.050 419.400 ;
        RECT 532.950 420.600 535.050 421.050 ;
        RECT 544.950 420.600 547.050 421.050 ;
        RECT 532.950 419.400 547.050 420.600 ;
        RECT 532.950 418.950 535.050 419.400 ;
        RECT 544.950 418.950 547.050 419.400 ;
        RECT 586.950 420.600 589.050 421.050 ;
        RECT 610.950 420.600 613.050 421.050 ;
        RECT 586.950 419.400 613.050 420.600 ;
        RECT 632.400 420.600 633.600 422.400 ;
        RECT 634.950 422.400 646.050 423.600 ;
        RECT 634.950 421.950 637.050 422.400 ;
        RECT 643.950 421.950 646.050 422.400 ;
        RECT 697.950 423.600 700.050 424.050 ;
        RECT 709.950 423.600 712.050 424.050 ;
        RECT 697.950 422.400 712.050 423.600 ;
        RECT 697.950 421.950 700.050 422.400 ;
        RECT 709.950 421.950 712.050 422.400 ;
        RECT 760.950 423.600 763.050 424.050 ;
        RECT 808.950 423.600 811.050 424.050 ;
        RECT 760.950 422.400 811.050 423.600 ;
        RECT 760.950 421.950 763.050 422.400 ;
        RECT 808.950 421.950 811.050 422.400 ;
        RECT 859.950 423.600 862.050 424.050 ;
        RECT 868.950 423.600 871.050 424.050 ;
        RECT 859.950 422.400 871.050 423.600 ;
        RECT 859.950 421.950 862.050 422.400 ;
        RECT 868.950 421.950 871.050 422.400 ;
        RECT 646.950 420.600 649.050 421.050 ;
        RECT 632.400 419.400 649.050 420.600 ;
        RECT 586.950 418.950 589.050 419.400 ;
        RECT 610.950 418.950 613.050 419.400 ;
        RECT 638.400 418.200 639.600 419.400 ;
        RECT 646.950 418.950 649.050 419.400 ;
        RECT 796.950 420.600 799.050 421.050 ;
        RECT 805.950 420.600 808.050 421.050 ;
        RECT 796.950 419.400 808.050 420.600 ;
        RECT 796.950 418.950 799.050 419.400 ;
        RECT 805.950 418.950 808.050 419.400 ;
        RECT 874.950 420.600 877.050 421.050 ;
        RECT 895.950 420.600 898.050 421.050 ;
        RECT 874.950 419.400 898.050 420.600 ;
        RECT 874.950 418.950 877.050 419.400 ;
        RECT 895.950 418.950 898.050 419.400 ;
        RECT 484.950 417.600 487.050 418.050 ;
        RECT 502.950 417.600 505.050 418.200 ;
        RECT 523.950 417.600 526.050 418.200 ;
        RECT 464.400 416.400 477.600 417.600 ;
        RECT 451.950 416.100 454.050 416.400 ;
        RECT 460.950 415.950 463.050 416.400 ;
        RECT 251.400 414.000 298.050 414.600 ;
        RECT 353.400 414.000 360.600 414.600 ;
        RECT 251.400 413.400 297.600 414.000 ;
        RECT 208.800 411.600 210.900 412.050 ;
        RECT 187.950 410.400 210.900 411.600 ;
        RECT 187.950 409.950 190.050 410.400 ;
        RECT 208.800 409.950 210.900 410.400 ;
        RECT 211.950 411.600 214.050 412.050 ;
        RECT 217.950 411.600 220.050 412.050 ;
        RECT 211.950 410.400 220.050 411.600 ;
        RECT 211.950 409.950 214.050 410.400 ;
        RECT 217.950 409.950 220.050 410.400 ;
        RECT 223.950 411.600 226.050 411.900 ;
        RECT 244.950 411.600 247.050 411.900 ;
        RECT 223.950 410.400 247.050 411.600 ;
        RECT 223.950 409.800 226.050 410.400 ;
        RECT 244.950 409.800 247.050 410.400 ;
        RECT 253.950 411.600 256.050 412.050 ;
        RECT 262.950 411.600 265.050 411.900 ;
        RECT 253.950 410.400 265.050 411.600 ;
        RECT 253.950 409.950 256.050 410.400 ;
        RECT 262.950 409.800 265.050 410.400 ;
        RECT 271.950 411.600 274.050 412.050 ;
        RECT 280.950 411.600 283.050 411.900 ;
        RECT 271.950 410.400 283.050 411.600 ;
        RECT 296.400 411.600 297.600 413.400 ;
        RECT 352.950 413.400 360.600 414.000 ;
        RECT 298.950 411.600 301.050 411.900 ;
        RECT 296.400 410.400 301.050 411.600 ;
        RECT 271.950 409.950 274.050 410.400 ;
        RECT 280.950 409.800 283.050 410.400 ;
        RECT 298.950 409.800 301.050 410.400 ;
        RECT 304.950 411.450 307.050 411.900 ;
        RECT 310.950 411.450 313.050 411.900 ;
        RECT 304.950 410.250 313.050 411.450 ;
        RECT 304.950 409.800 307.050 410.250 ;
        RECT 310.950 409.800 313.050 410.250 ;
        RECT 352.950 409.950 355.050 413.400 ;
        RECT 476.400 412.050 477.600 416.400 ;
        RECT 484.950 416.400 501.600 417.600 ;
        RECT 484.950 415.950 487.050 416.400 ;
        RECT 403.950 411.600 406.050 411.900 ;
        RECT 421.950 411.600 424.050 411.900 ;
        RECT 403.950 410.400 424.050 411.600 ;
        RECT 403.950 409.800 406.050 410.400 ;
        RECT 421.950 409.800 424.050 410.400 ;
        RECT 439.950 411.600 442.050 412.050 ;
        RECT 457.950 411.600 460.050 412.050 ;
        RECT 439.950 410.400 460.050 411.600 ;
        RECT 476.400 410.400 481.050 412.050 ;
        RECT 500.400 411.900 501.600 416.400 ;
        RECT 502.950 416.400 526.050 417.600 ;
        RECT 502.950 416.100 505.050 416.400 ;
        RECT 523.950 416.100 526.050 416.400 ;
        RECT 529.950 417.750 532.050 418.200 ;
        RECT 538.950 417.750 541.050 418.200 ;
        RECT 529.950 416.550 541.050 417.750 ;
        RECT 529.950 416.100 532.050 416.550 ;
        RECT 538.950 416.100 541.050 416.550 ;
        RECT 574.950 414.600 577.050 418.050 ;
        RECT 601.950 417.600 604.050 418.200 ;
        RECT 613.950 417.600 616.050 418.050 ;
        RECT 601.950 416.400 616.050 417.600 ;
        RECT 601.950 416.100 604.050 416.400 ;
        RECT 613.950 415.950 616.050 416.400 ;
        RECT 619.950 416.100 622.050 418.200 ;
        RECT 637.950 416.100 640.050 418.200 ;
        RECT 664.950 417.600 667.050 418.200 ;
        RECT 688.950 417.600 691.050 418.200 ;
        RECT 664.950 416.400 691.050 417.600 ;
        RECT 664.950 416.100 667.050 416.400 ;
        RECT 688.950 416.100 691.050 416.400 ;
        RECT 715.950 417.600 718.050 418.200 ;
        RECT 721.950 417.600 724.050 418.050 ;
        RECT 715.950 416.400 724.050 417.600 ;
        RECT 715.950 416.100 718.050 416.400 ;
        RECT 563.400 414.000 577.050 414.600 ;
        RECT 563.400 413.400 576.600 414.000 ;
        RECT 439.950 409.950 442.050 410.400 ;
        RECT 457.950 409.950 460.050 410.400 ;
        RECT 477.000 409.950 481.050 410.400 ;
        RECT 484.950 411.450 487.050 411.900 ;
        RECT 493.950 411.450 496.050 411.900 ;
        RECT 484.950 410.250 496.050 411.450 ;
        RECT 484.950 409.800 487.050 410.250 ;
        RECT 493.950 409.800 496.050 410.250 ;
        RECT 499.950 409.800 502.050 411.900 ;
        RECT 541.950 411.450 544.050 411.900 ;
        RECT 550.950 411.450 553.050 412.050 ;
        RECT 541.950 410.250 553.050 411.450 ;
        RECT 541.950 409.800 544.050 410.250 ;
        RECT 550.950 409.950 553.050 410.250 ;
        RECT 31.950 408.600 34.050 409.050 ;
        RECT 37.950 408.600 40.050 409.050 ;
        RECT 31.950 407.400 40.050 408.600 ;
        RECT 31.950 406.950 34.050 407.400 ;
        RECT 37.950 406.950 40.050 407.400 ;
        RECT 145.950 408.600 148.050 409.050 ;
        RECT 154.950 408.600 157.050 409.050 ;
        RECT 145.950 407.400 157.050 408.600 ;
        RECT 145.950 406.950 148.050 407.400 ;
        RECT 154.950 406.950 157.050 407.400 ;
        RECT 286.950 408.600 289.050 409.050 ;
        RECT 292.950 408.600 295.050 409.050 ;
        RECT 286.950 407.400 295.050 408.600 ;
        RECT 286.950 406.950 289.050 407.400 ;
        RECT 292.950 406.950 295.050 407.400 ;
        RECT 391.950 408.600 394.050 409.050 ;
        RECT 457.950 408.600 460.050 408.900 ;
        RECT 391.950 407.400 460.050 408.600 ;
        RECT 391.950 406.950 394.050 407.400 ;
        RECT 457.950 406.800 460.050 407.400 ;
        RECT 550.950 408.600 553.050 408.900 ;
        RECT 563.400 408.600 564.600 413.400 ;
        RECT 583.950 411.450 586.050 411.900 ;
        RECT 595.950 411.450 598.050 411.900 ;
        RECT 583.950 410.250 598.050 411.450 ;
        RECT 583.950 409.800 586.050 410.250 ;
        RECT 595.950 409.800 598.050 410.250 ;
        RECT 604.950 411.600 607.050 411.900 ;
        RECT 620.400 411.600 621.600 416.100 ;
        RECT 631.950 414.600 634.050 415.050 ;
        RECT 665.400 414.600 666.600 416.100 ;
        RECT 721.950 415.950 724.050 416.400 ;
        RECT 730.950 417.600 733.050 418.200 ;
        RECT 739.950 417.600 742.050 418.050 ;
        RECT 730.950 416.400 742.050 417.600 ;
        RECT 730.950 416.100 733.050 416.400 ;
        RECT 739.950 415.950 742.050 416.400 ;
        RECT 748.950 417.750 751.050 418.200 ;
        RECT 757.950 417.750 760.050 418.200 ;
        RECT 748.950 417.600 760.050 417.750 ;
        RECT 781.950 417.600 784.050 418.200 ;
        RECT 748.950 416.550 784.050 417.600 ;
        RECT 748.950 416.100 751.050 416.550 ;
        RECT 757.950 416.400 784.050 416.550 ;
        RECT 757.950 416.100 760.050 416.400 ;
        RECT 781.950 416.100 784.050 416.400 ;
        RECT 823.950 416.100 826.050 418.200 ;
        RECT 862.950 417.750 865.050 418.200 ;
        RECT 871.950 417.750 874.050 418.200 ;
        RECT 862.950 416.550 874.050 417.750 ;
        RECT 862.950 416.100 865.050 416.550 ;
        RECT 871.950 416.100 874.050 416.550 ;
        RECT 904.950 417.750 907.050 418.200 ;
        RECT 913.950 417.750 916.050 418.200 ;
        RECT 904.950 416.550 916.050 417.750 ;
        RECT 921.000 417.600 925.050 418.050 ;
        RECT 904.950 416.100 907.050 416.550 ;
        RECT 913.950 416.100 916.050 416.550 ;
        RECT 631.950 413.400 666.600 414.600 ;
        RECT 631.950 412.950 634.050 413.400 ;
        RECT 824.400 412.050 825.600 416.100 ;
        RECT 920.400 415.950 925.050 417.600 ;
        RECT 937.950 417.600 940.050 418.200 ;
        RECT 946.950 417.600 949.050 418.050 ;
        RECT 937.950 416.400 949.050 417.600 ;
        RECT 937.950 416.100 940.050 416.400 ;
        RECT 946.950 415.950 949.050 416.400 ;
        RECT 920.400 414.600 921.600 415.950 ;
        RECT 917.400 413.400 921.600 414.600 ;
        RECT 604.950 410.400 621.600 411.600 ;
        RECT 673.950 411.600 676.050 411.900 ;
        RECT 697.950 411.600 700.050 412.050 ;
        RECT 673.950 410.400 700.050 411.600 ;
        RECT 604.950 409.800 607.050 410.400 ;
        RECT 673.950 409.800 676.050 410.400 ;
        RECT 697.950 409.950 700.050 410.400 ;
        RECT 757.950 411.600 760.050 412.050 ;
        RECT 772.950 411.600 775.050 412.050 ;
        RECT 757.950 410.400 775.050 411.600 ;
        RECT 757.950 409.950 760.050 410.400 ;
        RECT 772.950 409.950 775.050 410.400 ;
        RECT 790.950 411.450 793.050 411.900 ;
        RECT 802.950 411.450 805.050 411.900 ;
        RECT 790.950 410.250 805.050 411.450 ;
        RECT 790.950 409.800 793.050 410.250 ;
        RECT 802.950 409.800 805.050 410.250 ;
        RECT 808.950 411.600 811.050 411.900 ;
        RECT 814.950 411.600 817.050 412.050 ;
        RECT 808.950 410.400 817.050 411.600 ;
        RECT 808.950 409.800 811.050 410.400 ;
        RECT 814.950 409.950 817.050 410.400 ;
        RECT 820.950 410.400 825.600 412.050 ;
        RECT 850.950 411.450 853.050 411.900 ;
        RECT 862.950 411.450 865.050 411.900 ;
        RECT 820.950 409.950 825.000 410.400 ;
        RECT 850.950 410.250 865.050 411.450 ;
        RECT 850.950 409.800 853.050 410.250 ;
        RECT 862.950 409.800 865.050 410.250 ;
        RECT 874.950 411.600 877.050 411.900 ;
        RECT 880.950 411.600 883.050 412.050 ;
        RECT 889.950 411.600 892.050 411.900 ;
        RECT 907.950 411.600 910.050 412.050 ;
        RECT 917.400 411.900 918.600 413.400 ;
        RECT 874.950 410.400 910.050 411.600 ;
        RECT 874.950 409.800 877.050 410.400 ;
        RECT 880.950 409.950 883.050 410.400 ;
        RECT 889.950 409.800 892.050 410.400 ;
        RECT 907.950 409.950 910.050 410.400 ;
        RECT 916.950 409.800 919.050 411.900 ;
        RECT 550.950 407.400 564.600 408.600 ;
        RECT 565.950 408.600 568.050 409.050 ;
        RECT 580.950 408.600 583.050 409.050 ;
        RECT 565.950 407.400 583.050 408.600 ;
        RECT 550.950 406.800 553.050 407.400 ;
        RECT 565.950 406.950 568.050 407.400 ;
        RECT 580.950 406.950 583.050 407.400 ;
        RECT 598.950 408.600 601.050 409.050 ;
        RECT 616.950 408.600 619.050 409.050 ;
        RECT 598.950 407.400 619.050 408.600 ;
        RECT 598.950 406.950 601.050 407.400 ;
        RECT 616.950 406.950 619.050 407.400 ;
        RECT 721.950 408.600 724.050 409.050 ;
        RECT 733.950 408.600 736.050 409.050 ;
        RECT 721.950 407.400 736.050 408.600 ;
        RECT 721.950 406.950 724.050 407.400 ;
        RECT 733.950 406.950 736.050 407.400 ;
        RECT 751.950 408.600 754.050 409.050 ;
        RECT 775.950 408.600 778.050 409.050 ;
        RECT 751.950 407.400 778.050 408.600 ;
        RECT 751.950 406.950 754.050 407.400 ;
        RECT 775.950 406.950 778.050 407.400 ;
        RECT 925.950 408.600 928.050 409.050 ;
        RECT 943.950 408.600 946.050 409.050 ;
        RECT 925.950 407.400 946.050 408.600 ;
        RECT 925.950 406.950 928.050 407.400 ;
        RECT 943.950 406.950 946.050 407.400 ;
        RECT 73.950 405.600 76.050 406.050 ;
        RECT 160.950 405.600 163.050 406.050 ;
        RECT 73.950 404.400 163.050 405.600 ;
        RECT 73.950 403.950 76.050 404.400 ;
        RECT 160.950 403.950 163.050 404.400 ;
        RECT 208.950 405.600 211.050 406.050 ;
        RECT 274.950 405.600 277.050 406.050 ;
        RECT 208.950 404.400 277.050 405.600 ;
        RECT 208.950 403.950 211.050 404.400 ;
        RECT 274.950 403.950 277.050 404.400 ;
        RECT 319.950 405.600 322.050 406.050 ;
        RECT 334.950 405.600 337.050 406.050 ;
        RECT 346.950 405.600 349.050 406.050 ;
        RECT 358.950 405.600 361.050 406.050 ;
        RECT 319.950 404.400 361.050 405.600 ;
        RECT 319.950 403.950 322.050 404.400 ;
        RECT 334.950 403.950 337.050 404.400 ;
        RECT 346.950 403.950 349.050 404.400 ;
        RECT 358.950 403.950 361.050 404.400 ;
        RECT 400.950 405.600 403.050 406.050 ;
        RECT 409.950 405.600 412.050 406.050 ;
        RECT 400.950 404.400 412.050 405.600 ;
        RECT 400.950 403.950 403.050 404.400 ;
        RECT 409.950 403.950 412.050 404.400 ;
        RECT 427.950 405.600 430.050 406.050 ;
        RECT 433.950 405.600 436.050 406.050 ;
        RECT 448.950 405.600 451.050 406.050 ;
        RECT 466.950 405.600 469.050 406.050 ;
        RECT 427.950 404.400 469.050 405.600 ;
        RECT 427.950 403.950 430.050 404.400 ;
        RECT 433.950 403.950 436.050 404.400 ;
        RECT 448.950 403.950 451.050 404.400 ;
        RECT 466.950 403.950 469.050 404.400 ;
        RECT 478.950 405.600 481.050 406.050 ;
        RECT 487.950 405.600 490.050 406.050 ;
        RECT 517.950 405.600 520.050 406.050 ;
        RECT 478.950 404.400 520.050 405.600 ;
        RECT 478.950 403.950 481.050 404.400 ;
        RECT 487.950 403.950 490.050 404.400 ;
        RECT 517.950 403.950 520.050 404.400 ;
        RECT 526.950 405.600 529.050 406.050 ;
        RECT 577.950 405.600 580.050 406.050 ;
        RECT 526.950 404.400 580.050 405.600 ;
        RECT 526.950 403.950 529.050 404.400 ;
        RECT 577.950 403.950 580.050 404.400 ;
        RECT 604.950 405.600 607.050 406.050 ;
        RECT 616.950 405.600 619.050 405.900 ;
        RECT 604.950 404.400 619.050 405.600 ;
        RECT 604.950 403.950 607.050 404.400 ;
        RECT 616.950 403.800 619.050 404.400 ;
        RECT 625.950 405.600 628.050 406.050 ;
        RECT 712.950 405.600 715.050 406.050 ;
        RECT 625.950 404.400 715.050 405.600 ;
        RECT 625.950 403.950 628.050 404.400 ;
        RECT 712.950 403.950 715.050 404.400 ;
        RECT 844.950 405.600 847.050 406.050 ;
        RECT 859.950 405.600 862.050 406.050 ;
        RECT 844.950 404.400 862.050 405.600 ;
        RECT 844.950 403.950 847.050 404.400 ;
        RECT 859.950 403.950 862.050 404.400 ;
        RECT 877.950 405.600 880.050 406.050 ;
        RECT 910.950 405.600 913.050 406.050 ;
        RECT 877.950 404.400 913.050 405.600 ;
        RECT 877.950 403.950 880.050 404.400 ;
        RECT 910.950 403.950 913.050 404.400 ;
        RECT 931.950 405.600 934.050 406.050 ;
        RECT 940.950 405.600 943.050 406.050 ;
        RECT 931.950 404.400 943.050 405.600 ;
        RECT 931.950 403.950 934.050 404.400 ;
        RECT 940.950 403.950 943.050 404.400 ;
        RECT 127.950 402.600 130.050 403.050 ;
        RECT 178.950 402.600 181.050 403.050 ;
        RECT 127.950 401.400 181.050 402.600 ;
        RECT 127.950 400.950 130.050 401.400 ;
        RECT 178.950 400.950 181.050 401.400 ;
        RECT 298.950 402.600 301.050 403.050 ;
        RECT 373.950 402.600 376.050 403.050 ;
        RECT 298.950 401.400 376.050 402.600 ;
        RECT 298.950 400.950 301.050 401.400 ;
        RECT 373.950 400.950 376.050 401.400 ;
        RECT 472.950 402.600 475.050 403.050 ;
        RECT 529.950 402.600 532.050 403.050 ;
        RECT 472.950 401.400 532.050 402.600 ;
        RECT 472.950 400.950 475.050 401.400 ;
        RECT 529.950 400.950 532.050 401.400 ;
        RECT 586.950 402.600 589.050 403.050 ;
        RECT 691.950 402.600 694.050 403.050 ;
        RECT 586.950 401.400 694.050 402.600 ;
        RECT 586.950 400.950 589.050 401.400 ;
        RECT 691.950 400.950 694.050 401.400 ;
        RECT 742.950 402.600 745.050 403.050 ;
        RECT 766.950 402.600 769.050 403.050 ;
        RECT 742.950 401.400 769.050 402.600 ;
        RECT 742.950 400.950 745.050 401.400 ;
        RECT 766.950 400.950 769.050 401.400 ;
        RECT 856.950 402.600 859.050 403.050 ;
        RECT 907.950 402.600 910.050 403.050 ;
        RECT 856.950 401.400 910.050 402.600 ;
        RECT 856.950 400.950 859.050 401.400 ;
        RECT 907.950 400.950 910.050 401.400 ;
        RECT 106.950 399.600 109.050 400.050 ;
        RECT 115.950 399.600 118.050 400.050 ;
        RECT 106.950 398.400 118.050 399.600 ;
        RECT 106.950 397.950 109.050 398.400 ;
        RECT 115.950 397.950 118.050 398.400 ;
        RECT 163.950 399.600 166.050 400.050 ;
        RECT 205.950 399.600 208.050 400.050 ;
        RECT 163.950 398.400 208.050 399.600 ;
        RECT 163.950 397.950 166.050 398.400 ;
        RECT 205.950 397.950 208.050 398.400 ;
        RECT 268.950 399.600 271.050 400.050 ;
        RECT 379.950 399.600 382.050 400.050 ;
        RECT 268.950 398.400 382.050 399.600 ;
        RECT 268.950 397.950 271.050 398.400 ;
        RECT 379.950 397.950 382.050 398.400 ;
        RECT 460.950 399.600 463.050 400.050 ;
        RECT 469.950 399.600 472.050 400.050 ;
        RECT 460.950 398.400 472.050 399.600 ;
        RECT 460.950 397.950 463.050 398.400 ;
        RECT 469.950 397.950 472.050 398.400 ;
        RECT 514.950 399.600 517.050 400.050 ;
        RECT 559.950 399.600 562.050 400.050 ;
        RECT 514.950 398.400 562.050 399.600 ;
        RECT 514.950 397.950 517.050 398.400 ;
        RECT 559.950 397.950 562.050 398.400 ;
        RECT 610.950 399.600 613.050 400.050 ;
        RECT 622.950 399.600 625.050 400.050 ;
        RECT 610.950 398.400 625.050 399.600 ;
        RECT 610.950 397.950 613.050 398.400 ;
        RECT 622.950 397.950 625.050 398.400 ;
        RECT 634.950 399.600 637.050 400.050 ;
        RECT 637.950 399.600 640.050 400.050 ;
        RECT 646.950 399.600 649.050 400.050 ;
        RECT 634.950 398.400 649.050 399.600 ;
        RECT 634.950 397.950 637.050 398.400 ;
        RECT 637.950 397.950 640.050 398.400 ;
        RECT 646.950 397.950 649.050 398.400 ;
        RECT 694.950 399.600 697.050 400.050 ;
        RECT 739.950 399.600 742.050 400.050 ;
        RECT 754.950 399.600 757.050 400.050 ;
        RECT 694.950 398.400 757.050 399.600 ;
        RECT 694.950 397.950 697.050 398.400 ;
        RECT 739.950 397.950 742.050 398.400 ;
        RECT 754.950 397.950 757.050 398.400 ;
        RECT 841.950 399.600 844.050 400.050 ;
        RECT 865.950 399.600 868.050 400.050 ;
        RECT 841.950 398.400 868.050 399.600 ;
        RECT 841.950 397.950 844.050 398.400 ;
        RECT 865.950 397.950 868.050 398.400 ;
        RECT 307.950 396.600 310.050 397.050 ;
        RECT 349.950 396.600 352.050 397.050 ;
        RECT 307.950 395.400 352.050 396.600 ;
        RECT 307.950 394.950 310.050 395.400 ;
        RECT 349.950 394.950 352.050 395.400 ;
        RECT 358.950 396.600 361.050 397.050 ;
        RECT 571.950 396.600 574.050 397.050 ;
        RECT 589.950 396.600 592.050 397.050 ;
        RECT 358.950 395.400 393.600 396.600 ;
        RECT 358.950 394.950 361.050 395.400 ;
        RECT 52.950 393.600 55.050 394.050 ;
        RECT 97.950 393.600 100.050 394.050 ;
        RECT 52.950 392.400 100.050 393.600 ;
        RECT 52.950 391.950 55.050 392.400 ;
        RECT 97.950 391.950 100.050 392.400 ;
        RECT 112.950 393.600 115.050 394.050 ;
        RECT 118.950 393.600 121.050 394.050 ;
        RECT 202.950 393.600 205.050 394.050 ;
        RECT 112.950 392.400 205.050 393.600 ;
        RECT 112.950 391.950 115.050 392.400 ;
        RECT 118.950 391.950 121.050 392.400 ;
        RECT 202.950 391.950 205.050 392.400 ;
        RECT 316.950 393.600 319.050 394.050 ;
        RECT 337.950 393.600 340.050 394.050 ;
        RECT 316.950 392.400 340.050 393.600 ;
        RECT 392.400 393.600 393.600 395.400 ;
        RECT 473.400 395.400 592.050 396.600 ;
        RECT 473.400 393.600 474.600 395.400 ;
        RECT 571.950 394.950 574.050 395.400 ;
        RECT 589.950 394.950 592.050 395.400 ;
        RECT 691.950 396.600 694.050 397.050 ;
        RECT 838.950 396.600 841.050 397.050 ;
        RECT 691.950 395.400 841.050 396.600 ;
        RECT 691.950 394.950 694.050 395.400 ;
        RECT 838.950 394.950 841.050 395.400 ;
        RECT 392.400 392.400 474.600 393.600 ;
        RECT 490.950 393.600 493.050 394.050 ;
        RECT 538.950 393.600 541.050 394.050 ;
        RECT 490.950 392.400 541.050 393.600 ;
        RECT 316.950 391.950 319.050 392.400 ;
        RECT 337.950 391.950 340.050 392.400 ;
        RECT 490.950 391.950 493.050 392.400 ;
        RECT 538.950 391.950 541.050 392.400 ;
        RECT 547.950 393.600 550.050 394.050 ;
        RECT 583.950 393.600 586.050 394.050 ;
        RECT 547.950 392.400 586.050 393.600 ;
        RECT 547.950 391.950 550.050 392.400 ;
        RECT 583.950 391.950 586.050 392.400 ;
        RECT 595.950 393.600 598.050 394.050 ;
        RECT 628.950 393.600 631.050 394.050 ;
        RECT 595.950 392.400 631.050 393.600 ;
        RECT 595.950 391.950 598.050 392.400 ;
        RECT 628.950 391.950 631.050 392.400 ;
        RECT 640.950 393.600 643.050 394.050 ;
        RECT 667.950 393.600 670.050 394.050 ;
        RECT 640.950 392.400 670.050 393.600 ;
        RECT 640.950 391.950 643.050 392.400 ;
        RECT 667.950 391.950 670.050 392.400 ;
        RECT 4.950 390.600 7.050 391.050 ;
        RECT 199.950 390.600 202.050 391.050 ;
        RECT 4.950 389.400 202.050 390.600 ;
        RECT 4.950 388.950 7.050 389.400 ;
        RECT 199.950 388.950 202.050 389.400 ;
        RECT 205.950 390.600 208.050 391.050 ;
        RECT 256.950 390.600 259.050 391.050 ;
        RECT 289.950 390.600 292.050 391.050 ;
        RECT 205.950 389.400 292.050 390.600 ;
        RECT 205.950 388.950 208.050 389.400 ;
        RECT 256.950 388.950 259.050 389.400 ;
        RECT 289.950 388.950 292.050 389.400 ;
        RECT 352.950 390.600 355.050 391.050 ;
        RECT 370.950 390.600 373.050 391.050 ;
        RECT 352.950 389.400 373.050 390.600 ;
        RECT 352.950 388.950 355.050 389.400 ;
        RECT 370.950 388.950 373.050 389.400 ;
        RECT 379.950 390.600 382.050 391.050 ;
        RECT 430.950 390.600 433.050 391.050 ;
        RECT 469.950 390.600 472.050 391.050 ;
        RECT 586.950 390.600 589.050 391.050 ;
        RECT 379.950 389.400 433.050 390.600 ;
        RECT 379.950 388.950 382.050 389.400 ;
        RECT 430.950 388.950 433.050 389.400 ;
        RECT 461.400 389.400 472.050 390.600 ;
        RECT 461.400 388.050 462.600 389.400 ;
        RECT 469.950 388.950 472.050 389.400 ;
        RECT 479.400 389.400 589.050 390.600 ;
        RECT 28.950 387.600 31.050 388.050 ;
        RECT 61.950 387.600 64.050 388.050 ;
        RECT 187.950 387.600 190.050 388.050 ;
        RECT 28.950 386.400 190.050 387.600 ;
        RECT 28.950 385.950 31.050 386.400 ;
        RECT 61.950 385.950 64.050 386.400 ;
        RECT 187.950 385.950 190.050 386.400 ;
        RECT 292.950 387.600 295.050 388.050 ;
        RECT 358.950 387.600 361.050 388.050 ;
        RECT 292.950 386.400 361.050 387.600 ;
        RECT 292.950 385.950 295.050 386.400 ;
        RECT 358.950 385.950 361.050 386.400 ;
        RECT 385.950 387.600 388.050 388.050 ;
        RECT 460.950 387.600 463.050 388.050 ;
        RECT 479.400 387.600 480.600 389.400 ;
        RECT 586.950 388.950 589.050 389.400 ;
        RECT 634.950 390.600 637.050 391.050 ;
        RECT 727.950 390.600 730.050 391.050 ;
        RECT 634.950 389.400 730.050 390.600 ;
        RECT 634.950 388.950 637.050 389.400 ;
        RECT 727.950 388.950 730.050 389.400 ;
        RECT 742.950 390.600 745.050 391.050 ;
        RECT 805.950 390.600 808.050 391.050 ;
        RECT 742.950 389.400 808.050 390.600 ;
        RECT 742.950 388.950 745.050 389.400 ;
        RECT 805.950 388.950 808.050 389.400 ;
        RECT 385.950 386.400 463.050 387.600 ;
        RECT 385.950 385.950 388.050 386.400 ;
        RECT 460.950 385.950 463.050 386.400 ;
        RECT 473.400 386.400 480.600 387.600 ;
        RECT 481.950 387.600 484.050 388.050 ;
        RECT 547.950 387.600 550.050 388.050 ;
        RECT 481.950 386.400 550.050 387.600 ;
        RECT 202.950 384.600 205.050 385.050 ;
        RECT 223.950 384.600 226.050 385.050 ;
        RECT 280.950 384.600 283.050 385.050 ;
        RECT 202.950 383.400 283.050 384.600 ;
        RECT 202.950 382.950 205.050 383.400 ;
        RECT 223.950 382.950 226.050 383.400 ;
        RECT 280.950 382.950 283.050 383.400 ;
        RECT 373.950 384.600 376.050 385.050 ;
        RECT 473.400 384.600 474.600 386.400 ;
        RECT 481.950 385.950 484.050 386.400 ;
        RECT 547.950 385.950 550.050 386.400 ;
        RECT 559.950 387.600 562.050 388.050 ;
        RECT 568.950 387.600 571.050 388.050 ;
        RECT 580.950 387.600 583.050 388.050 ;
        RECT 559.950 386.400 583.050 387.600 ;
        RECT 559.950 385.950 562.050 386.400 ;
        RECT 568.950 385.950 571.050 386.400 ;
        RECT 580.950 385.950 583.050 386.400 ;
        RECT 613.950 387.600 616.050 388.050 ;
        RECT 673.950 387.600 676.050 388.050 ;
        RECT 613.950 386.400 676.050 387.600 ;
        RECT 613.950 385.950 616.050 386.400 ;
        RECT 673.950 385.950 676.050 386.400 ;
        RECT 373.950 383.400 474.600 384.600 ;
        RECT 478.950 384.600 481.050 385.050 ;
        RECT 502.950 384.600 505.050 385.050 ;
        RECT 550.950 384.600 553.050 385.050 ;
        RECT 478.950 383.400 553.050 384.600 ;
        RECT 373.950 382.950 376.050 383.400 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 502.950 382.950 505.050 383.400 ;
        RECT 550.950 382.950 553.050 383.400 ;
        RECT 199.950 381.600 202.050 382.050 ;
        RECT 226.950 381.600 229.050 382.050 ;
        RECT 199.950 380.400 229.050 381.600 ;
        RECT 199.950 379.950 202.050 380.400 ;
        RECT 226.950 379.950 229.050 380.400 ;
        RECT 247.950 381.600 250.050 382.050 ;
        RECT 259.950 381.600 262.050 382.050 ;
        RECT 304.950 381.600 307.050 382.050 ;
        RECT 247.950 380.400 307.050 381.600 ;
        RECT 247.950 379.950 250.050 380.400 ;
        RECT 259.950 379.950 262.050 380.400 ;
        RECT 304.950 379.950 307.050 380.400 ;
        RECT 364.950 381.600 367.050 382.050 ;
        RECT 418.950 381.600 421.050 382.050 ;
        RECT 469.950 381.600 472.050 382.050 ;
        RECT 364.950 380.400 472.050 381.600 ;
        RECT 364.950 379.950 367.050 380.400 ;
        RECT 418.950 379.950 421.050 380.400 ;
        RECT 469.950 379.950 472.050 380.400 ;
        RECT 475.950 381.600 478.050 382.050 ;
        RECT 544.950 381.600 547.050 382.050 ;
        RECT 553.950 381.600 556.050 382.050 ;
        RECT 475.950 380.400 556.050 381.600 ;
        RECT 475.950 379.950 478.050 380.400 ;
        RECT 544.950 379.950 547.050 380.400 ;
        RECT 553.950 379.950 556.050 380.400 ;
        RECT 583.950 381.600 586.050 382.050 ;
        RECT 589.950 381.600 592.050 382.050 ;
        RECT 598.950 381.600 601.050 382.050 ;
        RECT 583.950 380.400 601.050 381.600 ;
        RECT 583.950 379.950 586.050 380.400 ;
        RECT 589.950 379.950 592.050 380.400 ;
        RECT 598.950 379.950 601.050 380.400 ;
        RECT 721.950 381.600 724.050 382.050 ;
        RECT 769.950 381.600 772.050 382.050 ;
        RECT 787.950 381.600 790.050 382.050 ;
        RECT 721.950 380.400 790.050 381.600 ;
        RECT 721.950 379.950 724.050 380.400 ;
        RECT 769.950 379.950 772.050 380.400 ;
        RECT 787.950 379.950 790.050 380.400 ;
        RECT 820.950 381.600 823.050 382.050 ;
        RECT 853.950 381.600 856.050 382.050 ;
        RECT 895.950 381.600 898.050 382.050 ;
        RECT 820.950 380.400 898.050 381.600 ;
        RECT 820.950 379.950 823.050 380.400 ;
        RECT 853.950 379.950 856.050 380.400 ;
        RECT 895.950 379.950 898.050 380.400 ;
        RECT 4.950 378.600 7.050 379.050 ;
        RECT 46.950 378.600 49.050 379.050 ;
        RECT 97.950 378.600 100.050 379.050 ;
        RECT 4.950 377.400 100.050 378.600 ;
        RECT 4.950 376.950 7.050 377.400 ;
        RECT 46.950 376.950 49.050 377.400 ;
        RECT 97.950 376.950 100.050 377.400 ;
        RECT 196.950 378.600 199.050 379.050 ;
        RECT 229.950 378.600 232.050 379.050 ;
        RECT 196.950 377.400 232.050 378.600 ;
        RECT 196.950 376.950 199.050 377.400 ;
        RECT 229.950 376.950 232.050 377.400 ;
        RECT 481.950 378.600 484.050 379.050 ;
        RECT 505.950 378.600 508.050 379.050 ;
        RECT 481.950 377.400 508.050 378.600 ;
        RECT 481.950 376.950 484.050 377.400 ;
        RECT 505.950 376.950 508.050 377.400 ;
        RECT 580.950 378.600 583.050 379.050 ;
        RECT 610.950 378.600 613.050 379.050 ;
        RECT 580.950 377.400 613.050 378.600 ;
        RECT 580.950 376.950 583.050 377.400 ;
        RECT 610.950 376.950 613.050 377.400 ;
        RECT 781.950 378.600 784.050 379.050 ;
        RECT 811.950 378.600 814.050 379.050 ;
        RECT 832.950 378.600 835.050 379.050 ;
        RECT 781.950 377.400 835.050 378.600 ;
        RECT 781.950 376.950 784.050 377.400 ;
        RECT 811.950 376.950 814.050 377.400 ;
        RECT 832.950 376.950 835.050 377.400 ;
        RECT 922.950 378.600 925.050 379.050 ;
        RECT 940.950 378.600 943.050 379.050 ;
        RECT 922.950 377.400 943.050 378.600 ;
        RECT 922.950 376.950 925.050 377.400 ;
        RECT 940.950 376.950 943.050 377.400 ;
        RECT 241.950 375.600 244.050 376.050 ;
        RECT 292.950 375.600 295.050 376.050 ;
        RECT 241.950 374.400 295.050 375.600 ;
        RECT 241.950 373.950 244.050 374.400 ;
        RECT 292.950 373.950 295.050 374.400 ;
        RECT 388.950 375.600 391.050 376.050 ;
        RECT 436.950 375.600 439.050 375.900 ;
        RECT 388.950 374.400 439.050 375.600 ;
        RECT 388.950 373.950 391.050 374.400 ;
        RECT 436.950 373.800 439.050 374.400 ;
        RECT 463.950 375.600 466.050 376.050 ;
        RECT 508.950 375.600 511.050 376.050 ;
        RECT 463.950 374.400 511.050 375.600 ;
        RECT 463.950 373.950 466.050 374.400 ;
        RECT 508.950 373.950 511.050 374.400 ;
        RECT 604.950 375.600 607.050 376.050 ;
        RECT 613.950 375.600 616.050 376.050 ;
        RECT 604.950 374.400 616.050 375.600 ;
        RECT 604.950 373.950 607.050 374.400 ;
        RECT 613.950 373.950 616.050 374.400 ;
        RECT 622.950 373.950 625.050 376.050 ;
        RECT 796.950 375.600 801.000 376.050 ;
        RECT 877.950 375.600 880.050 376.050 ;
        RECT 889.950 375.600 892.050 376.050 ;
        RECT 796.950 373.950 801.600 375.600 ;
        RECT 877.950 374.400 892.050 375.600 ;
        RECT 877.950 373.950 880.050 374.400 ;
        RECT 889.950 373.950 892.050 374.400 ;
        RECT 913.950 375.600 916.050 376.050 ;
        RECT 928.950 375.600 931.050 376.050 ;
        RECT 913.950 374.400 931.050 375.600 ;
        RECT 913.950 373.950 916.050 374.400 ;
        RECT 928.950 373.950 931.050 374.400 ;
        RECT 37.950 372.750 40.050 373.200 ;
        RECT 52.950 372.750 55.050 373.200 ;
        RECT 37.950 371.550 55.050 372.750 ;
        RECT 37.950 371.100 40.050 371.550 ;
        RECT 52.950 371.100 55.050 371.550 ;
        RECT 67.950 371.100 70.050 373.200 ;
        RECT 88.950 372.600 91.050 373.200 ;
        RECT 106.950 372.600 109.050 373.200 ;
        RECT 88.950 371.400 109.050 372.600 ;
        RECT 88.950 371.100 91.050 371.400 ;
        RECT 106.950 371.100 109.050 371.400 ;
        RECT 28.950 369.600 31.050 370.050 ;
        RECT 17.400 368.400 31.050 369.600 ;
        RECT 17.400 366.900 18.600 368.400 ;
        RECT 28.950 367.950 31.050 368.400 ;
        RECT 68.400 367.050 69.600 371.100 ;
        RECT 115.950 370.950 118.050 373.050 ;
        RECT 139.950 371.100 142.050 373.200 ;
        RECT 160.950 371.100 163.050 373.200 ;
        RECT 181.950 372.600 184.050 373.200 ;
        RECT 202.950 372.600 205.050 373.200 ;
        RECT 181.950 371.400 205.050 372.600 ;
        RECT 181.950 371.100 184.050 371.400 ;
        RECT 202.950 371.100 205.050 371.400 ;
        RECT 208.950 371.100 211.050 373.200 ;
        RECT 265.950 372.600 268.050 373.050 ;
        RECT 271.950 372.600 274.050 373.200 ;
        RECT 265.950 371.400 274.050 372.600 ;
        RECT 16.950 364.800 19.050 366.900 ;
        RECT 68.400 365.400 73.050 367.050 ;
        RECT 116.400 366.900 117.600 370.950 ;
        RECT 69.000 364.950 73.050 365.400 ;
        RECT 109.950 366.450 112.050 366.900 ;
        RECT 115.950 366.450 118.050 366.900 ;
        RECT 109.950 365.250 118.050 366.450 ;
        RECT 109.950 364.800 112.050 365.250 ;
        RECT 115.950 364.800 118.050 365.250 ;
        RECT 124.950 366.600 127.050 366.900 ;
        RECT 140.400 366.600 141.600 371.100 ;
        RECT 161.400 369.600 162.600 371.100 ;
        RECT 152.400 368.400 162.600 369.600 ;
        RECT 124.950 365.400 141.600 366.600 ;
        RECT 142.950 366.600 145.050 366.900 ;
        RECT 152.400 366.600 153.600 368.400 ;
        RECT 142.950 365.400 153.600 366.600 ;
        RECT 154.950 366.600 157.050 367.050 ;
        RECT 163.950 366.600 166.050 366.900 ;
        RECT 154.950 365.400 166.050 366.600 ;
        RECT 209.400 366.600 210.600 371.100 ;
        RECT 265.950 370.950 268.050 371.400 ;
        RECT 271.950 371.100 274.050 371.400 ;
        RECT 298.950 372.600 301.050 373.200 ;
        RECT 364.950 372.600 367.050 373.200 ;
        RECT 298.950 371.400 367.050 372.600 ;
        RECT 298.950 371.100 301.050 371.400 ;
        RECT 364.950 371.100 367.050 371.400 ;
        RECT 409.950 372.600 412.050 373.200 ;
        RECT 424.950 372.600 427.050 373.200 ;
        RECT 409.950 371.400 427.050 372.600 ;
        RECT 409.950 371.100 412.050 371.400 ;
        RECT 424.950 371.100 427.050 371.400 ;
        RECT 283.950 369.600 286.050 370.050 ;
        RECT 325.950 369.600 328.050 370.050 ;
        RECT 433.950 369.600 436.050 373.050 ;
        RECT 451.950 371.100 454.050 373.200 ;
        RECT 283.950 368.400 328.050 369.600 ;
        RECT 283.950 367.950 286.050 368.400 ;
        RECT 314.400 366.900 315.600 368.400 ;
        RECT 325.950 367.950 328.050 368.400 ;
        RECT 431.400 369.000 436.050 369.600 ;
        RECT 431.400 368.400 435.600 369.000 ;
        RECT 232.950 366.600 235.050 366.900 ;
        RECT 253.950 366.600 256.050 366.900 ;
        RECT 209.400 366.450 256.050 366.600 ;
        RECT 268.950 366.450 271.050 366.900 ;
        RECT 209.400 365.400 271.050 366.450 ;
        RECT 124.950 364.800 127.050 365.400 ;
        RECT 142.950 364.800 145.050 365.400 ;
        RECT 154.950 364.950 157.050 365.400 ;
        RECT 163.950 364.800 166.050 365.400 ;
        RECT 232.950 364.800 235.050 365.400 ;
        RECT 253.950 365.250 271.050 365.400 ;
        RECT 253.950 364.800 256.050 365.250 ;
        RECT 268.950 364.800 271.050 365.250 ;
        RECT 292.950 366.450 295.050 366.900 ;
        RECT 301.950 366.450 304.050 366.900 ;
        RECT 292.950 365.250 304.050 366.450 ;
        RECT 292.950 364.800 295.050 365.250 ;
        RECT 301.950 364.800 304.050 365.250 ;
        RECT 313.950 364.800 316.050 366.900 ;
        RECT 394.950 366.450 397.050 366.900 ;
        RECT 406.950 366.450 409.050 366.900 ;
        RECT 394.950 365.250 409.050 366.450 ;
        RECT 394.950 364.800 397.050 365.250 ;
        RECT 406.950 364.800 409.050 365.250 ;
        RECT 427.950 366.600 430.050 366.900 ;
        RECT 431.400 366.600 432.600 368.400 ;
        RECT 427.950 365.400 432.600 366.600 ;
        RECT 433.950 366.600 436.050 367.050 ;
        RECT 439.950 366.600 442.050 367.050 ;
        RECT 433.950 365.400 442.050 366.600 ;
        RECT 452.400 366.600 453.600 371.100 ;
        RECT 457.950 369.600 460.050 373.050 ;
        RECT 469.950 372.600 472.050 373.200 ;
        RECT 496.950 372.600 499.050 373.200 ;
        RECT 469.950 371.400 499.050 372.600 ;
        RECT 469.950 371.100 472.050 371.400 ;
        RECT 496.950 371.100 499.050 371.400 ;
        RECT 565.950 372.600 568.050 373.200 ;
        RECT 577.950 372.600 580.050 373.050 ;
        RECT 565.950 371.400 580.050 372.600 ;
        RECT 565.950 371.100 568.050 371.400 ;
        RECT 577.950 370.950 580.050 371.400 ;
        RECT 589.950 372.600 592.050 373.200 ;
        RECT 589.950 371.400 600.600 372.600 ;
        RECT 589.950 371.100 592.050 371.400 ;
        RECT 592.950 369.600 595.050 370.050 ;
        RECT 457.950 369.000 595.050 369.600 ;
        RECT 458.400 368.400 595.050 369.000 ;
        RECT 592.950 367.950 595.050 368.400 ;
        RECT 599.400 367.050 600.600 371.400 ;
        RECT 466.950 366.600 469.050 367.050 ;
        RECT 452.400 365.400 469.050 366.600 ;
        RECT 427.950 364.800 430.050 365.400 ;
        RECT 433.950 364.950 436.050 365.400 ;
        RECT 439.950 364.950 442.050 365.400 ;
        RECT 466.950 364.950 469.050 365.400 ;
        RECT 490.950 366.600 493.050 367.050 ;
        RECT 499.950 366.600 502.050 366.900 ;
        RECT 490.950 365.400 502.050 366.600 ;
        RECT 490.950 364.950 493.050 365.400 ;
        RECT 499.950 364.800 502.050 365.400 ;
        RECT 517.950 366.600 520.050 366.900 ;
        RECT 535.950 366.600 538.050 366.900 ;
        RECT 517.950 365.400 538.050 366.600 ;
        RECT 517.950 364.800 520.050 365.400 ;
        RECT 535.950 364.800 538.050 365.400 ;
        RECT 553.950 366.450 556.050 366.900 ;
        RECT 562.950 366.450 565.050 366.900 ;
        RECT 553.950 365.250 565.050 366.450 ;
        RECT 553.950 364.800 556.050 365.250 ;
        RECT 562.950 364.800 565.050 365.250 ;
        RECT 598.950 364.950 601.050 367.050 ;
        RECT 623.400 366.600 624.600 373.950 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 652.950 372.750 655.050 373.200 ;
        RECT 658.950 372.750 661.050 373.200 ;
        RECT 652.950 371.550 661.050 372.750 ;
        RECT 652.950 371.100 655.050 371.550 ;
        RECT 658.950 371.100 661.050 371.550 ;
        RECT 673.950 372.600 676.050 373.200 ;
        RECT 688.950 372.600 691.050 373.200 ;
        RECT 673.950 371.400 691.050 372.600 ;
        RECT 673.950 371.100 676.050 371.400 ;
        RECT 688.950 371.100 691.050 371.400 ;
        RECT 712.950 372.600 715.050 373.200 ;
        RECT 736.950 372.600 739.050 373.200 ;
        RECT 712.950 371.400 739.050 372.600 ;
        RECT 712.950 371.100 715.050 371.400 ;
        RECT 736.950 371.100 739.050 371.400 ;
        RECT 748.950 372.600 751.050 373.200 ;
        RECT 763.950 372.600 766.050 373.200 ;
        RECT 748.950 371.400 766.050 372.600 ;
        RECT 748.950 371.100 751.050 371.400 ;
        RECT 763.950 371.100 766.050 371.400 ;
        RECT 778.950 372.750 781.050 373.200 ;
        RECT 793.950 372.750 796.050 373.200 ;
        RECT 778.950 371.550 796.050 372.750 ;
        RECT 778.950 371.100 781.050 371.550 ;
        RECT 793.950 371.100 796.050 371.550 ;
        RECT 628.950 366.600 631.050 366.900 ;
        RECT 635.400 366.600 636.600 370.950 ;
        RECT 764.400 367.050 765.600 371.100 ;
        RECT 800.400 369.600 801.600 373.950 ;
        RECT 805.950 372.600 810.000 373.050 ;
        RECT 805.950 370.950 810.600 372.600 ;
        RECT 817.950 371.100 820.050 373.200 ;
        RECT 623.400 366.000 627.600 366.600 ;
        RECT 623.400 365.400 628.050 366.000 ;
        RECT 64.950 363.600 67.050 364.050 ;
        RECT 76.950 363.600 79.050 364.050 ;
        RECT 64.950 362.400 79.050 363.600 ;
        RECT 64.950 361.950 67.050 362.400 ;
        RECT 76.950 361.950 79.050 362.400 ;
        RECT 226.950 363.600 229.050 364.050 ;
        RECT 232.950 363.600 235.050 363.750 ;
        RECT 226.950 362.400 235.050 363.600 ;
        RECT 226.950 361.950 229.050 362.400 ;
        RECT 232.950 361.650 235.050 362.400 ;
        RECT 319.950 363.600 322.050 364.050 ;
        RECT 325.950 363.600 328.050 364.050 ;
        RECT 319.950 362.400 328.050 363.600 ;
        RECT 319.950 361.950 322.050 362.400 ;
        RECT 325.950 361.950 328.050 362.400 ;
        RECT 337.950 363.600 340.050 364.050 ;
        RECT 355.950 363.600 358.050 364.050 ;
        RECT 337.950 362.400 358.050 363.600 ;
        RECT 337.950 361.950 340.050 362.400 ;
        RECT 355.950 361.950 358.050 362.400 ;
        RECT 385.950 363.600 388.050 364.050 ;
        RECT 395.400 363.600 396.600 364.800 ;
        RECT 385.950 362.400 396.600 363.600 ;
        RECT 448.950 363.600 451.050 364.050 ;
        RECT 463.950 363.600 466.050 364.050 ;
        RECT 574.950 363.600 577.050 364.050 ;
        RECT 448.950 362.400 466.050 363.600 ;
        RECT 385.950 361.950 388.050 362.400 ;
        RECT 448.950 361.950 451.050 362.400 ;
        RECT 463.950 361.950 466.050 362.400 ;
        RECT 527.400 362.400 577.050 363.600 ;
        RECT 527.400 361.050 528.600 362.400 ;
        RECT 574.950 361.950 577.050 362.400 ;
        RECT 583.950 363.600 586.050 364.050 ;
        RECT 607.950 363.600 610.050 364.050 ;
        RECT 616.950 363.600 619.050 364.050 ;
        RECT 583.950 362.400 619.050 363.600 ;
        RECT 583.950 361.950 586.050 362.400 ;
        RECT 607.950 361.950 610.050 362.400 ;
        RECT 616.950 361.950 619.050 362.400 ;
        RECT 625.950 361.950 628.050 365.400 ;
        RECT 628.950 365.400 636.600 366.600 ;
        RECT 637.950 366.450 640.050 366.900 ;
        RECT 667.950 366.450 670.050 366.900 ;
        RECT 628.950 364.800 631.050 365.400 ;
        RECT 637.950 365.250 670.050 366.450 ;
        RECT 637.950 364.800 640.050 365.250 ;
        RECT 667.950 364.800 670.050 365.250 ;
        RECT 718.950 366.450 721.050 366.900 ;
        RECT 727.950 366.600 730.050 366.900 ;
        RECT 739.950 366.600 742.050 366.900 ;
        RECT 727.950 366.450 742.050 366.600 ;
        RECT 718.950 365.400 742.050 366.450 ;
        RECT 718.950 365.250 730.050 365.400 ;
        RECT 718.950 364.800 721.050 365.250 ;
        RECT 727.950 364.800 730.050 365.250 ;
        RECT 739.950 364.800 742.050 365.400 ;
        RECT 760.950 365.400 765.600 367.050 ;
        RECT 797.400 368.400 801.600 369.600 ;
        RECT 797.400 366.600 798.600 368.400 ;
        RECT 809.400 366.900 810.600 370.950 ;
        RECT 794.400 366.000 798.600 366.600 ;
        RECT 793.950 365.400 798.600 366.000 ;
        RECT 760.950 364.950 765.000 365.400 ;
        RECT 781.950 363.600 784.050 364.050 ;
        RECT 752.400 362.400 784.050 363.600 ;
        RECT 10.950 360.600 13.050 361.050 ;
        RECT 58.950 360.600 61.050 361.050 ;
        RECT 10.950 359.400 61.050 360.600 ;
        RECT 10.950 358.950 13.050 359.400 ;
        RECT 58.950 358.950 61.050 359.400 ;
        RECT 103.950 360.600 106.050 361.050 ;
        RECT 124.950 360.600 127.050 361.050 ;
        RECT 103.950 359.400 127.050 360.600 ;
        RECT 103.950 358.950 106.050 359.400 ;
        RECT 124.950 358.950 127.050 359.400 ;
        RECT 139.950 360.600 142.050 361.050 ;
        RECT 151.950 360.600 154.050 361.050 ;
        RECT 139.950 359.400 154.050 360.600 ;
        RECT 139.950 358.950 142.050 359.400 ;
        RECT 151.950 358.950 154.050 359.400 ;
        RECT 214.950 360.600 217.050 361.050 ;
        RECT 238.950 360.600 241.050 361.050 ;
        RECT 214.950 359.400 241.050 360.600 ;
        RECT 214.950 358.950 217.050 359.400 ;
        RECT 238.950 358.950 241.050 359.400 ;
        RECT 289.950 360.600 292.050 361.050 ;
        RECT 301.950 360.600 304.050 361.050 ;
        RECT 289.950 359.400 304.050 360.600 ;
        RECT 289.950 358.950 292.050 359.400 ;
        RECT 301.950 358.950 304.050 359.400 ;
        RECT 472.950 360.600 475.050 361.050 ;
        RECT 481.950 360.600 484.050 361.050 ;
        RECT 472.950 359.400 484.050 360.600 ;
        RECT 472.950 358.950 475.050 359.400 ;
        RECT 481.950 358.950 484.050 359.400 ;
        RECT 493.950 360.600 496.050 361.050 ;
        RECT 523.950 360.600 528.600 361.050 ;
        RECT 493.950 359.400 528.600 360.600 ;
        RECT 595.950 360.600 598.050 361.050 ;
        RECT 604.950 360.600 607.050 361.050 ;
        RECT 595.950 359.400 607.050 360.600 ;
        RECT 493.950 358.950 496.050 359.400 ;
        RECT 523.950 358.950 528.000 359.400 ;
        RECT 595.950 358.950 598.050 359.400 ;
        RECT 604.950 358.950 607.050 359.400 ;
        RECT 613.950 360.600 616.050 361.050 ;
        RECT 622.950 360.600 625.050 361.050 ;
        RECT 640.950 360.600 643.050 361.050 ;
        RECT 613.950 359.400 643.050 360.600 ;
        RECT 613.950 358.950 616.050 359.400 ;
        RECT 622.950 358.950 625.050 359.400 ;
        RECT 640.950 358.950 643.050 359.400 ;
        RECT 649.950 360.600 652.050 361.050 ;
        RECT 691.950 360.600 694.050 361.050 ;
        RECT 649.950 359.400 694.050 360.600 ;
        RECT 649.950 358.950 652.050 359.400 ;
        RECT 691.950 358.950 694.050 359.400 ;
        RECT 697.950 360.600 700.050 361.050 ;
        RECT 752.400 360.600 753.600 362.400 ;
        RECT 781.950 361.950 784.050 362.400 ;
        RECT 793.950 361.950 796.050 365.400 ;
        RECT 808.950 364.800 811.050 366.900 ;
        RECT 818.400 366.600 819.600 371.100 ;
        RECT 841.950 370.950 844.050 373.050 ;
        RECT 865.950 372.750 868.050 373.200 ;
        RECT 901.950 372.750 904.050 373.200 ;
        RECT 865.950 371.550 904.050 372.750 ;
        RECT 865.950 371.100 868.050 371.550 ;
        RECT 901.950 371.100 904.050 371.550 ;
        RECT 931.950 370.950 934.050 373.050 ;
        RECT 842.400 367.050 843.600 370.950 ;
        RECT 812.400 366.000 819.600 366.600 ;
        RECT 811.950 365.400 819.600 366.000 ;
        RECT 811.950 361.950 814.050 365.400 ;
        RECT 841.950 364.950 844.050 367.050 ;
        RECT 919.950 366.600 922.050 366.900 ;
        RECT 932.400 366.600 933.600 370.950 ;
        RECT 919.950 365.400 933.600 366.600 ;
        RECT 919.950 364.800 922.050 365.400 ;
        RECT 844.950 363.600 847.050 364.050 ;
        RECT 874.950 363.600 877.050 364.050 ;
        RECT 844.950 362.400 877.050 363.600 ;
        RECT 844.950 361.950 847.050 362.400 ;
        RECT 874.950 361.950 877.050 362.400 ;
        RECT 880.950 363.600 883.050 364.050 ;
        RECT 910.950 363.600 913.050 364.050 ;
        RECT 925.800 363.600 927.900 364.050 ;
        RECT 880.950 362.400 927.900 363.600 ;
        RECT 880.950 361.950 883.050 362.400 ;
        RECT 910.950 361.950 913.050 362.400 ;
        RECT 925.800 361.950 927.900 362.400 ;
        RECT 928.950 363.600 931.050 364.050 ;
        RECT 943.950 363.600 946.050 364.050 ;
        RECT 928.950 362.400 946.050 363.600 ;
        RECT 928.950 361.950 931.050 362.400 ;
        RECT 943.950 361.950 946.050 362.400 ;
        RECT 697.950 359.400 753.600 360.600 ;
        RECT 754.950 360.600 757.050 361.050 ;
        RECT 787.950 360.600 790.050 361.050 ;
        RECT 754.950 359.400 790.050 360.600 ;
        RECT 697.950 358.950 700.050 359.400 ;
        RECT 754.950 358.950 757.050 359.400 ;
        RECT 787.950 358.950 790.050 359.400 ;
        RECT 817.950 360.600 820.050 361.050 ;
        RECT 829.950 360.600 832.050 361.050 ;
        RECT 817.950 359.400 832.050 360.600 ;
        RECT 817.950 358.950 820.050 359.400 ;
        RECT 829.950 358.950 832.050 359.400 ;
        RECT 853.950 360.600 856.050 361.050 ;
        RECT 865.950 360.600 868.050 361.050 ;
        RECT 853.950 359.400 868.050 360.600 ;
        RECT 853.950 358.950 856.050 359.400 ;
        RECT 865.950 358.950 868.050 359.400 ;
        RECT 877.950 360.600 880.050 361.050 ;
        RECT 886.950 360.600 889.050 361.050 ;
        RECT 877.950 359.400 889.050 360.600 ;
        RECT 877.950 358.950 880.050 359.400 ;
        RECT 886.950 358.950 889.050 359.400 ;
        RECT 244.950 357.600 247.050 358.050 ;
        RECT 286.950 357.600 289.050 358.050 ;
        RECT 367.950 357.600 370.050 358.050 ;
        RECT 391.950 357.600 394.050 358.050 ;
        RECT 244.950 356.400 318.600 357.600 ;
        RECT 244.950 355.950 247.050 356.400 ;
        RECT 286.950 355.950 289.050 356.400 ;
        RECT 40.950 354.600 43.050 355.050 ;
        RECT 82.950 354.600 85.050 355.050 ;
        RECT 40.950 353.400 85.050 354.600 ;
        RECT 40.950 352.950 43.050 353.400 ;
        RECT 82.950 352.950 85.050 353.400 ;
        RECT 205.950 354.600 208.050 355.050 ;
        RECT 265.950 354.600 268.050 355.050 ;
        RECT 205.950 353.400 268.050 354.600 ;
        RECT 317.400 354.600 318.600 356.400 ;
        RECT 367.950 356.400 394.050 357.600 ;
        RECT 367.950 355.950 370.050 356.400 ;
        RECT 391.950 355.950 394.050 356.400 ;
        RECT 418.950 357.600 421.050 358.050 ;
        RECT 424.950 357.600 427.050 358.050 ;
        RECT 418.950 356.400 427.050 357.600 ;
        RECT 418.950 355.950 421.050 356.400 ;
        RECT 424.950 355.950 427.050 356.400 ;
        RECT 544.950 357.600 547.050 358.050 ;
        RECT 586.950 357.600 589.050 358.050 ;
        RECT 544.950 356.400 589.050 357.600 ;
        RECT 544.950 355.950 547.050 356.400 ;
        RECT 586.950 355.950 589.050 356.400 ;
        RECT 745.950 357.600 748.050 358.050 ;
        RECT 766.950 357.600 769.050 358.050 ;
        RECT 745.950 356.400 769.050 357.600 ;
        RECT 745.950 355.950 748.050 356.400 ;
        RECT 766.950 355.950 769.050 356.400 ;
        RECT 835.950 357.600 838.050 358.050 ;
        RECT 847.950 357.600 850.050 358.050 ;
        RECT 835.950 356.400 850.050 357.600 ;
        RECT 835.950 355.950 838.050 356.400 ;
        RECT 847.950 355.950 850.050 356.400 ;
        RECT 904.950 357.600 907.050 358.050 ;
        RECT 913.950 357.600 916.050 358.050 ;
        RECT 904.950 356.400 916.050 357.600 ;
        RECT 904.950 355.950 907.050 356.400 ;
        RECT 913.950 355.950 916.050 356.400 ;
        RECT 364.950 354.600 367.050 355.050 ;
        RECT 317.400 353.400 367.050 354.600 ;
        RECT 205.950 352.950 208.050 353.400 ;
        RECT 265.950 352.950 268.050 353.400 ;
        RECT 364.950 352.950 367.050 353.400 ;
        RECT 541.950 354.600 544.050 355.050 ;
        RECT 571.950 354.600 574.050 355.050 ;
        RECT 580.950 354.600 583.050 355.050 ;
        RECT 541.950 353.400 570.600 354.600 ;
        RECT 541.950 352.950 544.050 353.400 ;
        RECT 193.950 351.600 196.050 352.050 ;
        RECT 110.400 350.400 196.050 351.600 ;
        RECT 19.950 348.600 22.050 349.050 ;
        RECT 79.950 348.600 82.050 349.050 ;
        RECT 19.950 347.400 82.050 348.600 ;
        RECT 19.950 346.950 22.050 347.400 ;
        RECT 79.950 346.950 82.050 347.400 ;
        RECT 103.950 348.600 106.050 349.050 ;
        RECT 110.400 348.600 111.600 350.400 ;
        RECT 193.950 349.950 196.050 350.400 ;
        RECT 211.950 351.600 214.050 352.050 ;
        RECT 226.950 351.600 229.050 352.050 ;
        RECT 211.950 350.400 229.050 351.600 ;
        RECT 211.950 349.950 214.050 350.400 ;
        RECT 226.950 349.950 229.050 350.400 ;
        RECT 280.950 351.600 283.050 352.050 ;
        RECT 292.950 351.600 295.050 352.050 ;
        RECT 280.950 350.400 295.050 351.600 ;
        RECT 280.950 349.950 283.050 350.400 ;
        RECT 292.950 349.950 295.050 350.400 ;
        RECT 298.950 351.600 301.050 352.050 ;
        RECT 313.950 351.600 316.050 352.050 ;
        RECT 298.950 350.400 316.050 351.600 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 313.950 349.950 316.050 350.400 ;
        RECT 352.950 351.600 355.050 352.050 ;
        RECT 442.950 351.600 445.050 352.050 ;
        RECT 352.950 350.400 445.050 351.600 ;
        RECT 352.950 349.950 355.050 350.400 ;
        RECT 442.950 349.950 445.050 350.400 ;
        RECT 463.950 351.600 466.050 352.050 ;
        RECT 478.950 351.600 481.050 352.050 ;
        RECT 463.950 350.400 481.050 351.600 ;
        RECT 463.950 349.950 466.050 350.400 ;
        RECT 478.950 349.950 481.050 350.400 ;
        RECT 499.950 351.600 502.050 352.050 ;
        RECT 538.950 351.600 541.050 352.050 ;
        RECT 499.950 350.400 541.050 351.600 ;
        RECT 499.950 349.950 502.050 350.400 ;
        RECT 538.950 349.950 541.050 350.400 ;
        RECT 550.950 351.600 553.050 352.050 ;
        RECT 556.950 351.600 559.050 352.050 ;
        RECT 550.950 350.400 559.050 351.600 ;
        RECT 569.400 351.600 570.600 353.400 ;
        RECT 571.950 353.400 583.050 354.600 ;
        RECT 571.950 352.950 574.050 353.400 ;
        RECT 580.950 352.950 583.050 353.400 ;
        RECT 589.950 354.600 592.050 355.050 ;
        RECT 616.950 354.600 619.050 355.050 ;
        RECT 589.950 353.400 619.050 354.600 ;
        RECT 589.950 352.950 592.050 353.400 ;
        RECT 616.950 352.950 619.050 353.400 ;
        RECT 667.950 354.600 670.050 355.050 ;
        RECT 682.950 354.600 685.050 355.050 ;
        RECT 667.950 353.400 685.050 354.600 ;
        RECT 767.400 354.600 768.600 355.950 ;
        RECT 790.950 354.600 793.050 355.050 ;
        RECT 767.400 353.400 793.050 354.600 ;
        RECT 667.950 352.950 670.050 353.400 ;
        RECT 682.950 352.950 685.050 353.400 ;
        RECT 790.950 352.950 793.050 353.400 ;
        RECT 814.950 354.600 817.050 355.050 ;
        RECT 898.950 354.600 901.050 355.050 ;
        RECT 814.950 353.400 901.050 354.600 ;
        RECT 814.950 352.950 817.050 353.400 ;
        RECT 898.950 352.950 901.050 353.400 ;
        RECT 628.950 351.600 631.050 352.050 ;
        RECT 569.400 350.400 631.050 351.600 ;
        RECT 550.950 349.950 553.050 350.400 ;
        RECT 556.950 349.950 559.050 350.400 ;
        RECT 628.950 349.950 631.050 350.400 ;
        RECT 805.950 351.600 808.050 352.050 ;
        RECT 823.950 351.600 826.050 352.050 ;
        RECT 805.950 350.400 826.050 351.600 ;
        RECT 805.950 349.950 808.050 350.400 ;
        RECT 823.950 349.950 826.050 350.400 ;
        RECT 838.950 351.600 841.050 352.050 ;
        RECT 889.950 351.600 892.050 352.050 ;
        RECT 838.950 350.400 892.050 351.600 ;
        RECT 838.950 349.950 841.050 350.400 ;
        RECT 889.950 349.950 892.050 350.400 ;
        RECT 103.950 347.400 111.600 348.600 ;
        RECT 148.950 348.600 151.050 349.050 ;
        RECT 178.950 348.600 181.050 349.050 ;
        RECT 148.950 347.400 181.050 348.600 ;
        RECT 103.950 346.950 106.050 347.400 ;
        RECT 148.950 346.950 151.050 347.400 ;
        RECT 178.950 346.950 181.050 347.400 ;
        RECT 187.950 348.600 190.050 349.050 ;
        RECT 214.950 348.600 217.050 349.050 ;
        RECT 244.950 348.600 247.050 349.050 ;
        RECT 187.950 347.400 247.050 348.600 ;
        RECT 187.950 346.950 190.050 347.400 ;
        RECT 214.950 346.950 217.050 347.400 ;
        RECT 244.950 346.950 247.050 347.400 ;
        RECT 250.950 348.600 253.050 349.050 ;
        RECT 277.950 348.600 280.050 349.050 ;
        RECT 250.950 347.400 280.050 348.600 ;
        RECT 250.950 346.950 253.050 347.400 ;
        RECT 277.950 346.950 280.050 347.400 ;
        RECT 364.950 348.600 367.050 349.050 ;
        RECT 382.950 348.600 385.050 349.050 ;
        RECT 364.950 347.400 385.050 348.600 ;
        RECT 364.950 346.950 367.050 347.400 ;
        RECT 382.950 346.950 385.050 347.400 ;
        RECT 397.950 348.600 400.050 349.050 ;
        RECT 445.950 348.600 448.050 349.050 ;
        RECT 451.950 348.600 454.050 349.050 ;
        RECT 397.950 347.400 454.050 348.600 ;
        RECT 397.950 346.950 400.050 347.400 ;
        RECT 445.950 346.950 448.050 347.400 ;
        RECT 451.950 346.950 454.050 347.400 ;
        RECT 544.950 348.600 547.050 349.050 ;
        RECT 565.950 348.600 568.050 349.050 ;
        RECT 544.950 347.400 568.050 348.600 ;
        RECT 544.950 346.950 547.050 347.400 ;
        RECT 565.950 346.950 568.050 347.400 ;
        RECT 577.950 348.600 580.050 349.050 ;
        RECT 613.950 348.600 616.050 349.050 ;
        RECT 577.950 347.400 616.050 348.600 ;
        RECT 577.950 346.950 580.050 347.400 ;
        RECT 613.950 346.950 616.050 347.400 ;
        RECT 652.950 348.600 655.050 349.050 ;
        RECT 748.950 348.600 751.050 349.050 ;
        RECT 760.950 348.600 763.050 349.050 ;
        RECT 652.950 347.400 763.050 348.600 ;
        RECT 652.950 346.950 655.050 347.400 ;
        RECT 748.950 346.950 751.050 347.400 ;
        RECT 760.950 346.950 763.050 347.400 ;
        RECT 808.950 348.600 811.050 349.050 ;
        RECT 817.950 348.600 820.050 349.050 ;
        RECT 808.950 347.400 820.050 348.600 ;
        RECT 808.950 346.950 811.050 347.400 ;
        RECT 817.950 346.950 820.050 347.400 ;
        RECT 40.950 345.600 43.050 346.050 ;
        RECT 46.950 345.600 49.050 346.050 ;
        RECT 40.950 344.400 49.050 345.600 ;
        RECT 40.950 343.950 43.050 344.400 ;
        RECT 46.950 343.950 49.050 344.400 ;
        RECT 55.950 345.600 58.050 346.050 ;
        RECT 67.950 345.600 70.050 346.050 ;
        RECT 55.950 344.400 70.050 345.600 ;
        RECT 55.950 343.950 58.050 344.400 ;
        RECT 67.950 343.950 70.050 344.400 ;
        RECT 229.950 345.600 232.050 346.050 ;
        RECT 241.950 345.600 244.050 346.050 ;
        RECT 229.950 344.400 244.050 345.600 ;
        RECT 229.950 343.950 232.050 344.400 ;
        RECT 241.950 343.950 244.050 344.400 ;
        RECT 268.950 345.600 271.050 346.050 ;
        RECT 283.950 345.600 286.050 346.050 ;
        RECT 268.950 344.400 286.050 345.600 ;
        RECT 268.950 343.950 271.050 344.400 ;
        RECT 283.950 343.950 286.050 344.400 ;
        RECT 352.950 345.600 355.050 346.050 ;
        RECT 361.950 345.600 364.050 346.050 ;
        RECT 352.950 344.400 364.050 345.600 ;
        RECT 352.950 343.950 355.050 344.400 ;
        RECT 361.950 343.950 364.050 344.400 ;
        RECT 454.950 345.600 457.050 346.050 ;
        RECT 463.950 345.600 466.050 346.050 ;
        RECT 454.950 344.400 466.050 345.600 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 463.950 343.950 466.050 344.400 ;
        RECT 481.950 345.600 484.050 346.050 ;
        RECT 490.950 345.600 493.050 346.050 ;
        RECT 481.950 344.400 493.050 345.600 ;
        RECT 481.950 343.950 484.050 344.400 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 547.950 345.600 550.050 346.050 ;
        RECT 559.950 345.600 562.050 346.050 ;
        RECT 547.950 344.400 562.050 345.600 ;
        RECT 547.950 343.950 550.050 344.400 ;
        RECT 559.950 343.950 562.050 344.400 ;
        RECT 661.950 345.600 664.050 346.050 ;
        RECT 679.950 345.600 682.050 346.050 ;
        RECT 661.950 344.400 682.050 345.600 ;
        RECT 661.950 343.950 664.050 344.400 ;
        RECT 679.950 343.950 682.050 344.400 ;
        RECT 697.950 345.600 700.050 346.050 ;
        RECT 733.950 345.600 736.050 346.050 ;
        RECT 745.950 345.600 748.050 346.050 ;
        RECT 697.950 344.400 748.050 345.600 ;
        RECT 697.950 343.950 700.050 344.400 ;
        RECT 733.950 343.950 736.050 344.400 ;
        RECT 745.950 343.950 748.050 344.400 ;
        RECT 781.950 345.600 784.050 346.050 ;
        RECT 790.950 345.600 793.050 346.050 ;
        RECT 823.950 345.600 826.050 346.050 ;
        RECT 781.950 344.400 826.050 345.600 ;
        RECT 781.950 343.950 784.050 344.400 ;
        RECT 790.950 343.950 793.050 344.400 ;
        RECT 823.950 343.950 826.050 344.400 ;
        RECT 829.950 345.600 832.050 346.050 ;
        RECT 844.950 345.600 847.050 346.050 ;
        RECT 829.950 344.400 847.050 345.600 ;
        RECT 829.950 343.950 832.050 344.400 ;
        RECT 844.950 343.950 847.050 344.400 ;
        RECT 886.950 345.600 889.050 346.050 ;
        RECT 892.950 345.600 895.050 346.050 ;
        RECT 886.950 344.400 895.050 345.600 ;
        RECT 886.950 343.950 889.050 344.400 ;
        RECT 892.950 343.950 895.050 344.400 ;
        RECT 76.950 342.600 79.050 343.050 ;
        RECT 88.950 342.600 91.050 343.050 ;
        RECT 76.950 341.400 91.050 342.600 ;
        RECT 76.950 340.950 79.050 341.400 ;
        RECT 88.950 340.950 91.050 341.400 ;
        RECT 166.950 342.600 169.050 343.050 ;
        RECT 172.950 342.600 175.050 343.050 ;
        RECT 193.950 342.600 196.050 343.050 ;
        RECT 166.950 341.400 196.050 342.600 ;
        RECT 166.950 340.950 169.050 341.400 ;
        RECT 172.950 340.950 175.050 341.400 ;
        RECT 193.950 340.950 196.050 341.400 ;
        RECT 214.950 340.950 217.050 343.050 ;
        RECT 220.950 342.600 223.050 343.050 ;
        RECT 256.950 342.600 259.050 343.050 ;
        RECT 289.950 342.600 292.050 343.050 ;
        RECT 298.950 342.600 301.050 343.050 ;
        RECT 220.950 341.400 301.050 342.600 ;
        RECT 220.950 340.950 223.050 341.400 ;
        RECT 256.950 340.950 259.050 341.400 ;
        RECT 289.950 340.950 292.050 341.400 ;
        RECT 298.950 340.950 301.050 341.400 ;
        RECT 304.950 342.600 307.050 343.050 ;
        RECT 364.950 342.600 367.050 343.050 ;
        RECT 304.950 341.400 367.050 342.600 ;
        RECT 304.950 340.950 307.050 341.400 ;
        RECT 364.950 340.950 367.050 341.400 ;
        RECT 370.950 342.600 373.050 343.050 ;
        RECT 379.950 342.600 382.050 343.050 ;
        RECT 370.950 341.400 382.050 342.600 ;
        RECT 370.950 340.950 373.050 341.400 ;
        RECT 379.950 340.950 382.050 341.400 ;
        RECT 436.950 342.600 439.050 343.050 ;
        RECT 448.950 342.600 451.050 343.050 ;
        RECT 436.950 341.400 451.050 342.600 ;
        RECT 436.950 340.950 439.050 341.400 ;
        RECT 448.950 340.950 451.050 341.400 ;
        RECT 469.950 342.600 472.050 343.050 ;
        RECT 475.950 342.600 478.050 343.050 ;
        RECT 469.950 341.400 478.050 342.600 ;
        RECT 560.400 342.600 561.600 343.950 ;
        RECT 571.950 342.600 574.050 343.050 ;
        RECT 589.950 342.600 592.050 343.050 ;
        RECT 560.400 341.400 574.050 342.600 ;
        RECT 469.950 340.950 472.050 341.400 ;
        RECT 475.950 340.950 478.050 341.400 ;
        RECT 571.950 340.950 574.050 341.400 ;
        RECT 581.400 341.400 592.050 342.600 ;
        RECT 19.950 339.750 22.050 340.200 ;
        RECT 25.950 339.750 28.050 340.200 ;
        RECT 19.950 338.550 28.050 339.750 ;
        RECT 19.950 338.100 22.050 338.550 ;
        RECT 25.950 338.100 28.050 338.550 ;
        RECT 40.950 339.600 43.050 340.200 ;
        RECT 55.800 339.600 57.900 340.050 ;
        RECT 40.950 338.400 57.900 339.600 ;
        RECT 40.950 338.100 43.050 338.400 ;
        RECT 55.800 337.950 57.900 338.400 ;
        RECT 58.950 338.100 61.050 340.200 ;
        RECT 28.950 333.450 31.050 333.900 ;
        RECT 37.950 333.450 40.050 333.900 ;
        RECT 28.950 332.250 40.050 333.450 ;
        RECT 28.950 331.800 31.050 332.250 ;
        RECT 37.950 331.800 40.050 332.250 ;
        RECT 43.950 333.600 46.050 333.900 ;
        RECT 59.400 333.600 60.600 338.100 ;
        RECT 73.950 336.600 76.050 340.050 ;
        RECT 121.950 339.750 124.050 340.200 ;
        RECT 127.950 339.750 130.050 340.200 ;
        RECT 121.950 338.550 130.050 339.750 ;
        RECT 121.950 338.100 124.050 338.550 ;
        RECT 127.950 338.100 130.050 338.550 ;
        RECT 151.950 339.750 154.050 340.200 ;
        RECT 160.950 339.750 163.050 340.200 ;
        RECT 151.950 338.550 163.050 339.750 ;
        RECT 151.950 338.100 154.050 338.550 ;
        RECT 160.950 338.100 163.050 338.550 ;
        RECT 172.950 339.750 175.050 339.900 ;
        RECT 178.950 339.750 181.050 340.200 ;
        RECT 172.950 338.550 181.050 339.750 ;
        RECT 172.950 337.800 175.050 338.550 ;
        RECT 178.950 338.100 181.050 338.550 ;
        RECT 184.950 339.600 187.050 340.200 ;
        RECT 184.950 338.400 207.600 339.600 ;
        RECT 184.950 338.100 187.050 338.400 ;
        RECT 73.950 336.000 78.600 336.600 ;
        RECT 74.400 335.400 78.600 336.000 ;
        RECT 43.950 332.400 60.600 333.600 ;
        RECT 61.950 333.600 64.050 333.900 ;
        RECT 70.950 333.600 73.050 334.050 ;
        RECT 77.400 333.900 78.600 335.400 ;
        RECT 206.400 334.050 207.600 338.400 ;
        RECT 61.950 332.400 73.050 333.600 ;
        RECT 43.950 331.800 46.050 332.400 ;
        RECT 61.950 331.800 64.050 332.400 ;
        RECT 70.950 331.950 73.050 332.400 ;
        RECT 76.950 331.800 79.050 333.900 ;
        RECT 88.950 333.450 91.050 333.900 ;
        RECT 112.950 333.450 115.050 333.900 ;
        RECT 88.950 332.250 115.050 333.450 ;
        RECT 88.950 331.800 91.050 332.250 ;
        RECT 112.950 331.800 115.050 332.250 ;
        RECT 148.950 333.450 151.050 333.900 ;
        RECT 157.950 333.450 160.050 333.900 ;
        RECT 148.950 332.250 160.050 333.450 ;
        RECT 148.950 331.800 151.050 332.250 ;
        RECT 157.950 331.800 160.050 332.250 ;
        RECT 187.950 333.450 190.050 333.900 ;
        RECT 193.950 333.450 196.050 333.900 ;
        RECT 187.950 332.250 196.050 333.450 ;
        RECT 187.950 331.800 190.050 332.250 ;
        RECT 193.950 331.800 196.050 332.250 ;
        RECT 205.950 331.950 208.050 334.050 ;
        RECT 22.950 330.600 25.050 331.050 ;
        RECT 37.950 330.600 40.050 330.750 ;
        RECT 22.950 329.400 40.050 330.600 ;
        RECT 22.950 328.950 25.050 329.400 ;
        RECT 37.950 328.650 40.050 329.400 ;
        RECT 127.950 330.600 130.050 331.050 ;
        RECT 145.950 330.600 148.050 331.050 ;
        RECT 127.950 329.400 148.050 330.600 ;
        RECT 194.400 330.600 195.600 331.800 ;
        RECT 215.400 331.050 216.600 340.950 ;
        RECT 581.400 340.200 582.600 341.400 ;
        RECT 589.950 340.950 592.050 341.400 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 616.950 342.600 619.050 343.050 ;
        RECT 643.950 342.600 646.050 343.050 ;
        RECT 616.950 341.400 646.050 342.600 ;
        RECT 616.950 340.950 619.050 341.400 ;
        RECT 643.950 340.950 646.050 341.400 ;
        RECT 799.950 342.600 802.050 343.050 ;
        RECT 814.950 342.600 817.050 343.050 ;
        RECT 820.950 342.600 823.050 343.050 ;
        RECT 799.950 341.400 823.050 342.600 ;
        RECT 799.950 340.950 802.050 341.400 ;
        RECT 814.950 340.950 817.050 341.400 ;
        RECT 820.950 340.950 823.050 341.400 ;
        RECT 826.950 342.600 829.050 343.050 ;
        RECT 844.950 342.600 847.050 342.900 ;
        RECT 826.950 341.400 847.050 342.600 ;
        RECT 826.950 340.950 829.050 341.400 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 262.950 337.950 265.050 340.050 ;
        RECT 277.950 339.600 280.050 340.200 ;
        RECT 301.950 339.600 304.050 340.200 ;
        RECT 277.950 338.400 304.050 339.600 ;
        RECT 277.950 338.100 280.050 338.400 ;
        RECT 301.950 338.100 304.050 338.400 ;
        RECT 316.950 339.600 319.050 340.050 ;
        RECT 346.950 339.600 349.050 340.050 ;
        RECT 355.950 339.600 358.050 340.050 ;
        RECT 316.950 338.400 358.050 339.600 ;
        RECT 316.950 337.950 319.050 338.400 ;
        RECT 346.950 337.950 349.050 338.400 ;
        RECT 355.950 337.950 358.050 338.400 ;
        RECT 361.950 339.750 364.050 340.200 ;
        RECT 418.950 339.750 421.050 340.200 ;
        RECT 361.950 338.550 421.050 339.750 ;
        RECT 361.950 338.100 364.050 338.550 ;
        RECT 418.950 338.100 421.050 338.550 ;
        RECT 439.950 338.100 442.050 340.200 ;
        RECT 463.950 339.600 466.050 340.050 ;
        RECT 487.950 339.600 490.050 340.050 ;
        RECT 463.950 338.400 490.050 339.600 ;
        RECT 233.400 334.050 234.600 337.950 ;
        RECT 263.400 334.050 264.600 337.950 ;
        RECT 440.400 334.050 441.600 338.100 ;
        RECT 463.950 337.950 466.050 338.400 ;
        RECT 487.950 337.950 490.050 338.400 ;
        RECT 511.950 337.950 514.050 340.050 ;
        RECT 517.950 339.600 520.050 340.200 ;
        RECT 538.950 339.600 541.050 340.200 ;
        RECT 547.950 339.600 550.050 340.050 ;
        RECT 517.950 338.400 541.050 339.600 ;
        RECT 517.950 338.100 520.050 338.400 ;
        RECT 538.950 338.100 541.050 338.400 ;
        RECT 542.400 338.400 550.050 339.600 ;
        RECT 448.950 336.600 451.050 337.050 ;
        RECT 448.950 335.400 474.600 336.600 ;
        RECT 448.950 334.950 451.050 335.400 ;
        RECT 232.950 331.950 235.050 334.050 ;
        RECT 241.950 333.600 244.050 333.900 ;
        RECT 259.800 333.600 261.900 333.900 ;
        RECT 241.950 332.400 261.900 333.600 ;
        RECT 241.950 331.800 244.050 332.400 ;
        RECT 259.800 331.800 261.900 332.400 ;
        RECT 262.950 331.950 265.050 334.050 ;
        RECT 280.950 333.450 283.050 333.900 ;
        RECT 289.950 333.450 292.050 333.900 ;
        RECT 280.950 332.250 292.050 333.450 ;
        RECT 280.950 331.800 283.050 332.250 ;
        RECT 289.950 331.800 292.050 332.250 ;
        RECT 304.950 333.450 307.050 333.900 ;
        RECT 313.950 333.450 316.050 333.900 ;
        RECT 304.950 332.250 316.050 333.450 ;
        RECT 304.950 331.800 307.050 332.250 ;
        RECT 313.950 331.800 316.050 332.250 ;
        RECT 337.950 333.450 340.050 333.900 ;
        RECT 343.950 333.450 346.050 333.900 ;
        RECT 337.950 332.250 346.050 333.450 ;
        RECT 337.950 331.800 340.050 332.250 ;
        RECT 343.950 331.800 346.050 332.250 ;
        RECT 421.950 333.450 424.050 333.900 ;
        RECT 436.950 333.450 439.050 333.900 ;
        RECT 421.950 332.250 439.050 333.450 ;
        RECT 440.400 332.400 445.050 334.050 ;
        RECT 473.400 333.600 474.600 335.400 ;
        RECT 512.400 334.050 513.600 337.950 ;
        RECT 542.400 336.600 543.600 338.400 ;
        RECT 547.950 337.950 550.050 338.400 ;
        RECT 565.950 339.600 570.000 340.050 ;
        RECT 565.950 337.950 570.600 339.600 ;
        RECT 574.950 337.950 577.050 340.050 ;
        RECT 580.800 338.100 582.900 340.200 ;
        RECT 583.950 339.600 586.050 340.050 ;
        RECT 589.950 339.600 592.050 339.900 ;
        RECT 583.950 338.400 592.050 339.600 ;
        RECT 583.950 337.950 586.050 338.400 ;
        RECT 539.400 335.400 543.600 336.600 ;
        RECT 484.950 333.600 487.050 333.900 ;
        RECT 496.950 333.600 499.050 333.900 ;
        RECT 473.400 332.400 499.050 333.600 ;
        RECT 421.950 331.800 424.050 332.250 ;
        RECT 436.950 331.800 439.050 332.250 ;
        RECT 441.000 331.950 445.050 332.400 ;
        RECT 484.950 331.800 487.050 332.400 ;
        RECT 496.950 331.800 499.050 332.400 ;
        RECT 511.950 331.950 514.050 334.050 ;
        RECT 535.950 333.600 538.050 333.900 ;
        RECT 539.400 333.600 540.600 335.400 ;
        RECT 535.950 332.400 540.600 333.600 ;
        RECT 535.950 331.800 538.050 332.400 ;
        RECT 569.400 331.050 570.600 337.950 ;
        RECT 575.400 331.050 576.600 337.950 ;
        RECT 589.950 337.800 592.050 338.400 ;
        RECT 577.950 333.600 580.050 333.900 ;
        RECT 589.950 333.600 592.050 334.050 ;
        RECT 577.950 332.400 592.050 333.600 ;
        RECT 577.950 331.800 580.050 332.400 ;
        RECT 589.950 331.950 592.050 332.400 ;
        RECT 208.950 330.600 211.050 331.050 ;
        RECT 194.400 329.400 211.050 330.600 ;
        RECT 127.950 328.950 130.050 329.400 ;
        RECT 145.950 328.950 148.050 329.400 ;
        RECT 208.950 328.950 211.050 329.400 ;
        RECT 214.950 328.950 217.050 331.050 ;
        RECT 298.950 330.600 301.050 331.050 ;
        RECT 307.950 330.600 310.050 331.050 ;
        RECT 298.950 329.400 310.050 330.600 ;
        RECT 298.950 328.950 301.050 329.400 ;
        RECT 307.950 328.950 310.050 329.400 ;
        RECT 448.950 330.600 451.050 331.050 ;
        RECT 502.950 330.600 505.050 331.050 ;
        RECT 448.950 329.400 505.050 330.600 ;
        RECT 448.950 328.950 451.050 329.400 ;
        RECT 502.950 328.950 505.050 329.400 ;
        RECT 520.950 330.600 523.050 331.050 ;
        RECT 532.950 330.600 535.050 331.050 ;
        RECT 520.950 329.400 535.050 330.600 ;
        RECT 520.950 328.950 523.050 329.400 ;
        RECT 532.950 328.950 535.050 329.400 ;
        RECT 559.950 330.600 562.050 331.050 ;
        RECT 565.800 330.600 567.900 331.050 ;
        RECT 559.950 329.400 567.900 330.600 ;
        RECT 559.950 328.950 562.050 329.400 ;
        RECT 565.800 328.950 567.900 329.400 ;
        RECT 568.950 328.950 571.050 331.050 ;
        RECT 574.950 328.950 577.050 331.050 ;
        RECT 583.950 330.600 586.050 331.050 ;
        RECT 596.400 330.600 597.600 340.950 ;
        RECT 844.950 340.800 847.050 341.400 ;
        RECT 913.950 342.600 916.050 343.050 ;
        RECT 925.950 342.600 928.050 343.050 ;
        RECT 913.950 341.400 928.050 342.600 ;
        RECT 913.950 340.950 916.050 341.400 ;
        RECT 925.950 340.950 928.050 341.400 ;
        RECT 940.950 340.950 943.050 343.050 ;
        RECT 619.950 339.600 622.050 340.200 ;
        RECT 658.950 339.600 661.050 340.050 ;
        RECT 670.950 339.600 673.050 340.200 ;
        RECT 619.950 338.400 624.600 339.600 ;
        RECT 619.950 338.100 622.050 338.400 ;
        RECT 623.400 334.050 624.600 338.400 ;
        RECT 656.400 338.400 673.050 339.600 ;
        RECT 598.950 333.600 601.050 333.900 ;
        RECT 610.950 333.600 613.050 333.900 ;
        RECT 598.950 332.400 613.050 333.600 ;
        RECT 598.950 331.800 601.050 332.400 ;
        RECT 610.950 331.800 613.050 332.400 ;
        RECT 622.950 331.950 625.050 334.050 ;
        RECT 656.400 333.900 657.600 338.400 ;
        RECT 658.950 337.950 661.050 338.400 ;
        RECT 670.950 338.100 673.050 338.400 ;
        RECT 679.950 339.750 682.050 340.200 ;
        RECT 691.950 339.750 694.050 340.200 ;
        RECT 679.950 339.600 694.050 339.750 ;
        RECT 715.950 339.600 718.050 340.200 ;
        RECT 679.950 338.550 718.050 339.600 ;
        RECT 679.950 338.100 682.050 338.550 ;
        RECT 691.950 338.400 718.050 338.550 ;
        RECT 691.950 338.100 694.050 338.400 ;
        RECT 715.950 338.100 718.050 338.400 ;
        RECT 721.950 339.600 724.050 340.200 ;
        RECT 742.950 339.600 745.050 340.050 ;
        RECT 721.950 338.400 745.050 339.600 ;
        RECT 721.950 338.100 724.050 338.400 ;
        RECT 742.950 337.950 745.050 338.400 ;
        RECT 748.950 339.600 751.050 340.050 ;
        RECT 766.950 339.750 769.050 340.200 ;
        RECT 775.950 339.750 778.050 340.200 ;
        RECT 748.950 338.400 762.600 339.600 ;
        RECT 748.950 337.950 751.050 338.400 ;
        RECT 761.400 333.900 762.600 338.400 ;
        RECT 766.950 338.550 778.050 339.750 ;
        RECT 786.000 339.600 790.050 340.050 ;
        RECT 766.950 338.100 769.050 338.550 ;
        RECT 775.950 338.100 778.050 338.550 ;
        RECT 785.400 337.950 790.050 339.600 ;
        RECT 823.950 339.600 826.050 340.200 ;
        RECT 871.950 339.600 874.050 340.200 ;
        RECT 883.950 339.600 886.050 340.050 ;
        RECT 892.950 339.600 895.050 340.200 ;
        RECT 823.950 338.400 846.600 339.600 ;
        RECT 823.950 338.100 826.050 338.400 ;
        RECT 785.400 333.900 786.600 337.950 ;
        RECT 845.400 333.900 846.600 338.400 ;
        RECT 871.950 338.400 895.050 339.600 ;
        RECT 871.950 338.100 874.050 338.400 ;
        RECT 883.950 337.950 886.050 338.400 ;
        RECT 892.950 338.100 895.050 338.400 ;
        RECT 898.950 339.750 901.050 340.200 ;
        RECT 907.950 339.750 910.050 340.200 ;
        RECT 898.950 338.550 910.050 339.750 ;
        RECT 898.950 338.100 901.050 338.550 ;
        RECT 907.950 338.100 910.050 338.550 ;
        RECT 937.950 338.100 940.050 340.200 ;
        RECT 938.400 336.600 939.600 338.100 ;
        RECT 932.400 335.400 939.600 336.600 ;
        RECT 634.950 333.600 637.050 333.900 ;
        RECT 649.950 333.600 652.050 333.900 ;
        RECT 634.950 332.400 652.050 333.600 ;
        RECT 634.950 331.800 637.050 332.400 ;
        RECT 649.950 331.800 652.050 332.400 ;
        RECT 655.950 331.800 658.050 333.900 ;
        RECT 664.950 333.450 667.050 333.900 ;
        RECT 673.950 333.450 676.050 333.900 ;
        RECT 664.950 332.250 676.050 333.450 ;
        RECT 664.950 331.800 667.050 332.250 ;
        RECT 673.950 331.800 676.050 332.250 ;
        RECT 682.950 333.450 685.050 333.900 ;
        RECT 694.950 333.450 697.050 333.900 ;
        RECT 682.950 332.250 697.050 333.450 ;
        RECT 682.950 331.800 685.050 332.250 ;
        RECT 694.950 331.800 697.050 332.250 ;
        RECT 736.950 333.600 739.050 333.900 ;
        RECT 754.950 333.600 757.050 333.900 ;
        RECT 736.950 332.400 757.050 333.600 ;
        RECT 736.950 331.800 739.050 332.400 ;
        RECT 754.950 331.800 757.050 332.400 ;
        RECT 760.950 331.800 763.050 333.900 ;
        RECT 784.950 331.800 787.050 333.900 ;
        RECT 790.950 333.450 793.050 333.900 ;
        RECT 796.950 333.450 799.050 333.900 ;
        RECT 790.950 332.250 799.050 333.450 ;
        RECT 790.950 331.800 793.050 332.250 ;
        RECT 796.950 331.800 799.050 332.250 ;
        RECT 802.950 333.450 805.050 333.900 ;
        RECT 808.950 333.450 811.050 333.900 ;
        RECT 802.950 332.250 811.050 333.450 ;
        RECT 802.950 331.800 805.050 332.250 ;
        RECT 808.950 331.800 811.050 332.250 ;
        RECT 844.950 331.800 847.050 333.900 ;
        RECT 904.950 333.600 907.050 334.050 ;
        RECT 932.400 333.600 933.600 335.400 ;
        RECT 941.400 333.600 942.600 340.950 ;
        RECT 946.950 337.950 949.050 340.050 ;
        RECT 947.400 334.050 948.600 337.950 ;
        RECT 904.950 332.400 933.600 333.600 ;
        RECT 938.400 333.000 942.600 333.600 ;
        RECT 937.950 332.400 942.600 333.000 ;
        RECT 904.950 331.950 907.050 332.400 ;
        RECT 583.950 329.400 597.600 330.600 ;
        RECT 694.950 330.600 697.050 331.050 ;
        RECT 718.950 330.600 721.050 331.050 ;
        RECT 694.950 329.400 721.050 330.600 ;
        RECT 583.950 328.950 586.050 329.400 ;
        RECT 694.950 328.950 697.050 329.400 ;
        RECT 718.950 328.950 721.050 329.400 ;
        RECT 883.950 330.600 886.050 331.050 ;
        RECT 898.950 330.600 901.050 331.050 ;
        RECT 883.950 329.400 901.050 330.600 ;
        RECT 883.950 328.950 886.050 329.400 ;
        RECT 898.950 328.950 901.050 329.400 ;
        RECT 916.950 330.600 919.050 331.050 ;
        RECT 922.950 330.600 925.050 331.050 ;
        RECT 916.950 329.400 925.050 330.600 ;
        RECT 916.950 328.950 919.050 329.400 ;
        RECT 922.950 328.950 925.050 329.400 ;
        RECT 937.950 328.950 940.050 332.400 ;
        RECT 946.950 331.950 949.050 334.050 ;
        RECT 94.950 327.600 97.050 328.050 ;
        RECT 118.950 327.600 121.050 328.050 ;
        RECT 94.950 326.400 121.050 327.600 ;
        RECT 94.950 325.950 97.050 326.400 ;
        RECT 118.950 325.950 121.050 326.400 ;
        RECT 205.950 327.600 208.050 328.050 ;
        RECT 235.950 327.600 238.050 328.050 ;
        RECT 205.950 326.400 238.050 327.600 ;
        RECT 205.950 325.950 208.050 326.400 ;
        RECT 235.950 325.950 238.050 326.400 ;
        RECT 274.950 327.600 277.050 328.050 ;
        RECT 299.400 327.600 300.600 328.950 ;
        RECT 274.950 326.400 300.600 327.600 ;
        RECT 409.950 327.600 412.050 328.050 ;
        RECT 442.950 327.600 445.050 328.050 ;
        RECT 409.950 326.400 445.050 327.600 ;
        RECT 274.950 325.950 277.050 326.400 ;
        RECT 409.950 325.950 412.050 326.400 ;
        RECT 442.950 325.950 445.050 326.400 ;
        RECT 448.950 327.600 451.050 327.900 ;
        RECT 466.950 327.600 469.050 328.050 ;
        RECT 448.950 326.400 469.050 327.600 ;
        RECT 448.950 325.800 451.050 326.400 ;
        RECT 466.950 325.950 469.050 326.400 ;
        RECT 490.950 327.600 493.050 328.050 ;
        RECT 541.950 327.600 544.050 328.050 ;
        RECT 490.950 326.400 544.050 327.600 ;
        RECT 490.950 325.950 493.050 326.400 ;
        RECT 541.950 325.950 544.050 326.400 ;
        RECT 601.950 327.600 604.050 328.050 ;
        RECT 625.950 327.600 628.050 328.050 ;
        RECT 601.950 326.400 628.050 327.600 ;
        RECT 601.950 325.950 604.050 326.400 ;
        RECT 625.950 325.950 628.050 326.400 ;
        RECT 649.950 327.600 652.050 328.050 ;
        RECT 661.950 327.600 664.050 328.050 ;
        RECT 649.950 326.400 664.050 327.600 ;
        RECT 649.950 325.950 652.050 326.400 ;
        RECT 661.950 325.950 664.050 326.400 ;
        RECT 742.950 327.600 745.050 328.050 ;
        RECT 763.950 327.600 766.050 328.050 ;
        RECT 742.950 326.400 766.050 327.600 ;
        RECT 742.950 325.950 745.050 326.400 ;
        RECT 763.950 325.950 766.050 326.400 ;
        RECT 769.950 327.600 772.050 328.050 ;
        RECT 814.950 327.600 817.050 328.050 ;
        RECT 820.950 327.600 823.050 328.050 ;
        RECT 769.950 326.400 823.050 327.600 ;
        RECT 769.950 325.950 772.050 326.400 ;
        RECT 814.950 325.950 817.050 326.400 ;
        RECT 820.950 325.950 823.050 326.400 ;
        RECT 136.950 324.600 139.050 325.050 ;
        RECT 154.950 324.600 157.050 325.050 ;
        RECT 136.950 323.400 157.050 324.600 ;
        RECT 136.950 322.950 139.050 323.400 ;
        RECT 154.950 322.950 157.050 323.400 ;
        RECT 181.950 324.600 184.050 325.050 ;
        RECT 193.950 324.600 196.050 325.050 ;
        RECT 226.950 324.600 229.050 325.050 ;
        RECT 181.950 323.400 229.050 324.600 ;
        RECT 181.950 322.950 184.050 323.400 ;
        RECT 193.950 322.950 196.050 323.400 ;
        RECT 226.950 322.950 229.050 323.400 ;
        RECT 265.950 324.600 268.050 325.050 ;
        RECT 298.950 324.600 301.050 324.900 ;
        RECT 265.950 323.400 301.050 324.600 ;
        RECT 265.950 322.950 268.050 323.400 ;
        RECT 298.950 322.800 301.050 323.400 ;
        RECT 403.950 324.600 406.050 325.050 ;
        RECT 430.950 324.600 433.050 325.050 ;
        RECT 403.950 323.400 433.050 324.600 ;
        RECT 403.950 322.950 406.050 323.400 ;
        RECT 430.950 322.950 433.050 323.400 ;
        RECT 439.950 324.600 442.050 325.050 ;
        RECT 445.950 324.600 448.050 325.050 ;
        RECT 496.950 324.600 499.050 325.050 ;
        RECT 439.950 323.400 499.050 324.600 ;
        RECT 439.950 322.950 442.050 323.400 ;
        RECT 445.950 322.950 448.050 323.400 ;
        RECT 496.950 322.950 499.050 323.400 ;
        RECT 520.950 324.600 523.050 325.050 ;
        RECT 550.950 324.600 553.050 325.050 ;
        RECT 520.950 323.400 553.050 324.600 ;
        RECT 520.950 322.950 523.050 323.400 ;
        RECT 550.950 322.950 553.050 323.400 ;
        RECT 556.950 324.600 559.050 325.050 ;
        RECT 565.950 324.600 568.050 325.050 ;
        RECT 583.800 324.600 585.900 325.050 ;
        RECT 556.950 323.400 585.900 324.600 ;
        RECT 556.950 322.950 559.050 323.400 ;
        RECT 565.950 322.950 568.050 323.400 ;
        RECT 583.800 322.950 585.900 323.400 ;
        RECT 586.950 324.600 589.050 325.050 ;
        RECT 616.950 324.600 619.050 325.050 ;
        RECT 586.950 323.400 619.050 324.600 ;
        RECT 586.950 322.950 589.050 323.400 ;
        RECT 616.950 322.950 619.050 323.400 ;
        RECT 232.950 321.600 235.050 322.050 ;
        RECT 253.950 321.600 256.050 322.050 ;
        RECT 232.950 320.400 256.050 321.600 ;
        RECT 232.950 319.950 235.050 320.400 ;
        RECT 253.950 319.950 256.050 320.400 ;
        RECT 460.950 321.600 463.050 322.050 ;
        RECT 493.950 321.600 496.050 322.050 ;
        RECT 460.950 320.400 496.050 321.600 ;
        RECT 460.950 319.950 463.050 320.400 ;
        RECT 493.950 319.950 496.050 320.400 ;
        RECT 595.950 321.600 598.050 322.050 ;
        RECT 637.950 321.600 640.050 322.050 ;
        RECT 595.950 320.400 640.050 321.600 ;
        RECT 595.950 319.950 598.050 320.400 ;
        RECT 637.950 319.950 640.050 320.400 ;
        RECT 688.950 321.600 691.050 322.050 ;
        RECT 712.950 321.600 715.050 322.050 ;
        RECT 688.950 320.400 715.050 321.600 ;
        RECT 688.950 319.950 691.050 320.400 ;
        RECT 712.950 319.950 715.050 320.400 ;
        RECT 43.950 318.600 46.050 319.050 ;
        RECT 124.950 318.600 127.050 319.050 ;
        RECT 43.950 317.400 127.050 318.600 ;
        RECT 43.950 316.950 46.050 317.400 ;
        RECT 124.950 316.950 127.050 317.400 ;
        RECT 145.950 318.600 148.050 319.050 ;
        RECT 211.950 318.600 214.050 319.050 ;
        RECT 145.950 317.400 214.050 318.600 ;
        RECT 145.950 316.950 148.050 317.400 ;
        RECT 211.950 316.950 214.050 317.400 ;
        RECT 277.950 318.600 280.050 319.050 ;
        RECT 295.950 318.600 298.050 319.050 ;
        RECT 277.950 317.400 298.050 318.600 ;
        RECT 277.950 316.950 280.050 317.400 ;
        RECT 295.950 316.950 298.050 317.400 ;
        RECT 301.950 318.600 304.050 319.050 ;
        RECT 358.950 318.600 361.050 319.050 ;
        RECT 430.950 318.600 433.050 319.050 ;
        RECT 301.950 317.400 433.050 318.600 ;
        RECT 301.950 316.950 304.050 317.400 ;
        RECT 358.950 316.950 361.050 317.400 ;
        RECT 430.950 316.950 433.050 317.400 ;
        RECT 538.950 318.600 541.050 319.050 ;
        RECT 571.950 318.600 574.050 319.050 ;
        RECT 580.950 318.600 583.050 319.050 ;
        RECT 640.950 318.600 643.050 319.050 ;
        RECT 538.950 317.400 570.600 318.600 ;
        RECT 538.950 316.950 541.050 317.400 ;
        RECT 136.950 315.600 139.050 316.050 ;
        RECT 223.950 315.600 226.050 316.050 ;
        RECT 136.950 314.400 226.050 315.600 ;
        RECT 136.950 313.950 139.050 314.400 ;
        RECT 223.950 313.950 226.050 314.400 ;
        RECT 280.950 315.600 283.050 316.050 ;
        RECT 325.950 315.600 328.050 316.050 ;
        RECT 280.950 314.400 328.050 315.600 ;
        RECT 280.950 313.950 283.050 314.400 ;
        RECT 325.950 313.950 328.050 314.400 ;
        RECT 361.950 315.600 364.050 316.050 ;
        RECT 394.950 315.600 397.050 316.050 ;
        RECT 361.950 314.400 397.050 315.600 ;
        RECT 361.950 313.950 364.050 314.400 ;
        RECT 394.950 313.950 397.050 314.400 ;
        RECT 451.950 315.600 454.050 316.050 ;
        RECT 520.950 315.600 523.050 316.050 ;
        RECT 451.950 314.400 523.050 315.600 ;
        RECT 451.950 313.950 454.050 314.400 ;
        RECT 520.950 313.950 523.050 314.400 ;
        RECT 556.950 315.600 559.050 316.050 ;
        RECT 562.950 315.600 565.050 316.050 ;
        RECT 556.950 314.400 565.050 315.600 ;
        RECT 569.400 315.600 570.600 317.400 ;
        RECT 571.950 317.400 643.050 318.600 ;
        RECT 571.950 316.950 574.050 317.400 ;
        RECT 580.950 316.950 583.050 317.400 ;
        RECT 640.950 316.950 643.050 317.400 ;
        RECT 886.950 318.600 889.050 319.050 ;
        RECT 898.950 318.600 901.050 319.050 ;
        RECT 886.950 317.400 901.050 318.600 ;
        RECT 886.950 316.950 889.050 317.400 ;
        RECT 898.950 316.950 901.050 317.400 ;
        RECT 595.800 315.600 597.900 316.050 ;
        RECT 569.400 314.400 597.900 315.600 ;
        RECT 556.950 313.950 559.050 314.400 ;
        RECT 562.950 313.950 565.050 314.400 ;
        RECT 595.800 313.950 597.900 314.400 ;
        RECT 598.950 315.600 601.050 316.050 ;
        RECT 604.950 315.600 607.050 316.050 ;
        RECT 598.950 314.400 607.050 315.600 ;
        RECT 598.950 313.950 601.050 314.400 ;
        RECT 604.950 313.950 607.050 314.400 ;
        RECT 637.950 315.600 640.050 316.050 ;
        RECT 667.950 315.600 670.050 316.050 ;
        RECT 679.950 315.600 682.050 316.050 ;
        RECT 637.950 314.400 682.050 315.600 ;
        RECT 637.950 313.950 640.050 314.400 ;
        RECT 667.950 313.950 670.050 314.400 ;
        RECT 679.950 313.950 682.050 314.400 ;
        RECT 691.950 315.600 694.050 316.050 ;
        RECT 703.950 315.600 706.050 316.050 ;
        RECT 691.950 314.400 706.050 315.600 ;
        RECT 691.950 313.950 694.050 314.400 ;
        RECT 703.950 313.950 706.050 314.400 ;
        RECT 241.950 312.600 244.050 313.050 ;
        RECT 247.950 312.600 250.050 313.050 ;
        RECT 418.950 312.600 421.050 313.050 ;
        RECT 241.950 311.400 421.050 312.600 ;
        RECT 241.950 310.950 244.050 311.400 ;
        RECT 247.950 310.950 250.050 311.400 ;
        RECT 418.950 310.950 421.050 311.400 ;
        RECT 445.950 312.600 448.050 313.050 ;
        RECT 505.950 312.600 508.050 313.050 ;
        RECT 526.950 312.600 529.050 313.050 ;
        RECT 541.800 312.600 543.900 313.050 ;
        RECT 445.950 311.400 543.900 312.600 ;
        RECT 445.950 310.950 448.050 311.400 ;
        RECT 505.950 310.950 508.050 311.400 ;
        RECT 526.950 310.950 529.050 311.400 ;
        RECT 541.800 310.950 543.900 311.400 ;
        RECT 544.950 312.600 547.050 313.050 ;
        RECT 574.950 312.600 577.050 313.050 ;
        RECT 601.950 312.600 604.050 313.050 ;
        RECT 544.950 311.400 604.050 312.600 ;
        RECT 544.950 310.950 547.050 311.400 ;
        RECT 574.950 310.950 577.050 311.400 ;
        RECT 601.950 310.950 604.050 311.400 ;
        RECT 628.950 312.600 631.050 313.050 ;
        RECT 745.950 312.600 748.050 313.050 ;
        RECT 754.950 312.600 757.050 313.050 ;
        RECT 628.950 311.400 757.050 312.600 ;
        RECT 628.950 310.950 631.050 311.400 ;
        RECT 745.950 310.950 748.050 311.400 ;
        RECT 754.950 310.950 757.050 311.400 ;
        RECT 805.950 312.600 808.050 313.050 ;
        RECT 859.950 312.600 862.050 313.050 ;
        RECT 805.950 311.400 862.050 312.600 ;
        RECT 805.950 310.950 808.050 311.400 ;
        RECT 859.950 310.950 862.050 311.400 ;
        RECT 913.950 312.600 916.050 313.050 ;
        RECT 934.950 312.600 937.050 313.050 ;
        RECT 913.950 311.400 937.050 312.600 ;
        RECT 913.950 310.950 916.050 311.400 ;
        RECT 934.950 310.950 937.050 311.400 ;
        RECT 82.950 309.600 85.050 310.050 ;
        RECT 133.950 309.600 136.050 310.050 ;
        RECT 205.950 309.600 208.050 310.050 ;
        RECT 82.950 308.400 208.050 309.600 ;
        RECT 82.950 307.950 85.050 308.400 ;
        RECT 133.950 307.950 136.050 308.400 ;
        RECT 205.950 307.950 208.050 308.400 ;
        RECT 289.950 309.600 292.050 310.050 ;
        RECT 349.950 309.600 352.050 310.050 ;
        RECT 289.950 308.400 352.050 309.600 ;
        RECT 289.950 307.950 292.050 308.400 ;
        RECT 349.950 307.950 352.050 308.400 ;
        RECT 388.950 309.600 391.050 310.050 ;
        RECT 412.950 309.600 415.050 310.050 ;
        RECT 388.950 308.400 415.050 309.600 ;
        RECT 388.950 307.950 391.050 308.400 ;
        RECT 412.950 307.950 415.050 308.400 ;
        RECT 430.950 309.600 433.050 310.050 ;
        RECT 442.950 309.600 445.050 310.050 ;
        RECT 430.950 308.400 445.050 309.600 ;
        RECT 430.950 307.950 433.050 308.400 ;
        RECT 442.950 307.950 445.050 308.400 ;
        RECT 493.950 309.600 496.050 310.050 ;
        RECT 553.950 309.600 556.050 310.050 ;
        RECT 493.950 308.400 556.050 309.600 ;
        RECT 493.950 307.950 496.050 308.400 ;
        RECT 553.950 307.950 556.050 308.400 ;
        RECT 568.950 309.600 571.050 310.050 ;
        RECT 700.950 309.600 703.050 310.050 ;
        RECT 568.950 308.400 703.050 309.600 ;
        RECT 568.950 307.950 571.050 308.400 ;
        RECT 700.950 307.950 703.050 308.400 ;
        RECT 910.950 309.600 913.050 310.050 ;
        RECT 940.950 309.600 943.050 310.050 ;
        RECT 910.950 308.400 943.050 309.600 ;
        RECT 910.950 307.950 913.050 308.400 ;
        RECT 940.950 307.950 943.050 308.400 ;
        RECT 52.950 306.600 55.050 307.050 ;
        RECT 148.950 306.600 151.050 307.050 ;
        RECT 229.950 306.600 232.050 307.050 ;
        RECT 52.950 305.400 232.050 306.600 ;
        RECT 52.950 304.950 55.050 305.400 ;
        RECT 148.950 304.950 151.050 305.400 ;
        RECT 229.950 304.950 232.050 305.400 ;
        RECT 370.950 306.600 373.050 307.050 ;
        RECT 445.950 306.600 448.050 307.050 ;
        RECT 370.950 305.400 448.050 306.600 ;
        RECT 370.950 304.950 373.050 305.400 ;
        RECT 445.950 304.950 448.050 305.400 ;
        RECT 451.950 306.600 454.050 307.050 ;
        RECT 478.950 306.600 481.050 307.050 ;
        RECT 571.950 306.600 574.050 307.050 ;
        RECT 451.950 305.400 574.050 306.600 ;
        RECT 451.950 304.950 454.050 305.400 ;
        RECT 478.950 304.950 481.050 305.400 ;
        RECT 571.950 304.950 574.050 305.400 ;
        RECT 643.950 306.600 646.050 307.050 ;
        RECT 691.950 306.600 694.050 307.050 ;
        RECT 643.950 305.400 694.050 306.600 ;
        RECT 643.950 304.950 646.050 305.400 ;
        RECT 691.950 304.950 694.050 305.400 ;
        RECT 757.950 306.600 760.050 307.050 ;
        RECT 790.950 306.600 793.050 307.050 ;
        RECT 757.950 305.400 793.050 306.600 ;
        RECT 757.950 304.950 760.050 305.400 ;
        RECT 790.950 304.950 793.050 305.400 ;
        RECT 868.950 306.600 871.050 307.050 ;
        RECT 922.950 306.600 925.050 307.050 ;
        RECT 868.950 305.400 925.050 306.600 ;
        RECT 868.950 304.950 871.050 305.400 ;
        RECT 922.950 304.950 925.050 305.400 ;
        RECT 76.950 303.600 79.050 304.050 ;
        RECT 115.950 303.600 118.050 304.050 ;
        RECT 130.950 303.600 133.050 304.050 ;
        RECT 76.950 302.400 133.050 303.600 ;
        RECT 76.950 301.950 79.050 302.400 ;
        RECT 115.950 301.950 118.050 302.400 ;
        RECT 130.950 301.950 133.050 302.400 ;
        RECT 172.950 303.600 175.050 304.050 ;
        RECT 295.950 303.600 298.050 304.050 ;
        RECT 172.950 302.400 298.050 303.600 ;
        RECT 172.950 301.950 175.050 302.400 ;
        RECT 295.950 301.950 298.050 302.400 ;
        RECT 328.950 303.600 331.050 304.050 ;
        RECT 361.950 303.600 364.050 304.050 ;
        RECT 328.950 302.400 364.050 303.600 ;
        RECT 328.950 301.950 331.050 302.400 ;
        RECT 361.950 301.950 364.050 302.400 ;
        RECT 496.950 303.600 499.050 304.050 ;
        RECT 562.950 303.600 565.050 304.050 ;
        RECT 583.950 303.600 586.050 304.050 ;
        RECT 496.950 302.400 586.050 303.600 ;
        RECT 496.950 301.950 499.050 302.400 ;
        RECT 562.950 301.950 565.050 302.400 ;
        RECT 583.950 301.950 586.050 302.400 ;
        RECT 700.950 303.600 703.050 304.050 ;
        RECT 730.950 303.600 733.050 304.050 ;
        RECT 700.950 302.400 733.050 303.600 ;
        RECT 700.950 301.950 703.050 302.400 ;
        RECT 730.950 301.950 733.050 302.400 ;
        RECT 13.950 300.600 16.050 301.050 ;
        RECT 28.950 300.600 31.050 301.050 ;
        RECT 13.950 299.400 31.050 300.600 ;
        RECT 13.950 298.950 16.050 299.400 ;
        RECT 28.950 298.950 31.050 299.400 ;
        RECT 103.950 300.600 106.050 301.050 ;
        RECT 112.950 300.600 115.050 301.050 ;
        RECT 292.950 300.600 295.050 301.050 ;
        RECT 103.950 299.400 115.050 300.600 ;
        RECT 103.950 298.950 106.050 299.400 ;
        RECT 112.950 298.950 115.050 299.400 ;
        RECT 218.400 299.400 295.050 300.600 ;
        RECT 205.950 297.600 208.050 298.050 ;
        RECT 218.400 297.600 219.600 299.400 ;
        RECT 292.950 298.950 295.050 299.400 ;
        RECT 382.950 300.600 385.050 301.050 ;
        RECT 403.950 300.600 406.050 301.050 ;
        RECT 382.950 299.400 406.050 300.600 ;
        RECT 382.950 298.950 385.050 299.400 ;
        RECT 403.950 298.950 406.050 299.400 ;
        RECT 424.950 300.600 427.050 300.900 ;
        RECT 448.950 300.600 451.050 301.050 ;
        RECT 424.950 299.400 451.050 300.600 ;
        RECT 424.950 298.800 427.050 299.400 ;
        RECT 448.950 298.950 451.050 299.400 ;
        RECT 487.950 300.600 490.050 301.050 ;
        RECT 511.950 300.600 514.050 301.050 ;
        RECT 487.950 299.400 514.050 300.600 ;
        RECT 487.950 298.950 490.050 299.400 ;
        RECT 511.950 298.950 514.050 299.400 ;
        RECT 529.950 300.600 532.050 301.050 ;
        RECT 535.950 300.600 538.050 301.050 ;
        RECT 556.950 300.600 559.050 301.050 ;
        RECT 529.950 299.400 559.050 300.600 ;
        RECT 529.950 298.950 532.050 299.400 ;
        RECT 535.950 298.950 538.050 299.400 ;
        RECT 556.950 298.950 559.050 299.400 ;
        RECT 604.950 300.600 607.050 301.050 ;
        RECT 655.950 300.600 658.050 301.050 ;
        RECT 604.950 299.400 658.050 300.600 ;
        RECT 604.950 298.950 607.050 299.400 ;
        RECT 655.950 298.950 658.050 299.400 ;
        RECT 679.950 300.600 682.050 301.050 ;
        RECT 760.950 300.600 763.050 301.050 ;
        RECT 679.950 299.400 763.050 300.600 ;
        RECT 679.950 298.950 682.050 299.400 ;
        RECT 760.950 298.950 763.050 299.400 ;
        RECT 910.950 300.600 913.050 301.050 ;
        RECT 916.950 300.600 919.050 301.050 ;
        RECT 910.950 299.400 919.050 300.600 ;
        RECT 910.950 298.950 913.050 299.400 ;
        RECT 916.950 298.950 919.050 299.400 ;
        RECT 205.950 296.400 219.600 297.600 ;
        RECT 301.950 297.600 304.050 298.050 ;
        RECT 310.950 297.600 313.050 298.050 ;
        RECT 301.950 296.400 313.050 297.600 ;
        RECT 205.950 295.950 208.050 296.400 ;
        RECT 301.950 295.950 304.050 296.400 ;
        RECT 310.950 295.950 313.050 296.400 ;
        RECT 322.950 297.600 325.050 298.050 ;
        RECT 334.950 297.600 337.050 298.050 ;
        RECT 322.950 296.400 337.050 297.600 ;
        RECT 322.950 295.950 325.050 296.400 ;
        RECT 334.950 295.950 337.050 296.400 ;
        RECT 400.950 295.950 403.050 298.050 ;
        RECT 496.950 295.950 499.050 298.050 ;
        RECT 544.800 297.000 546.900 298.050 ;
        RECT 547.950 297.600 550.050 298.050 ;
        RECT 601.950 297.600 604.050 298.050 ;
        RECT 544.800 295.950 547.050 297.000 ;
        RECT 547.950 296.400 604.050 297.600 ;
        RECT 547.950 295.950 550.050 296.400 ;
        RECT 601.950 295.950 604.050 296.400 ;
        RECT 622.950 297.600 625.050 298.050 ;
        RECT 706.950 297.600 709.050 298.050 ;
        RECT 712.950 297.600 715.050 298.050 ;
        RECT 754.950 297.600 757.050 298.050 ;
        RECT 921.000 297.600 925.050 298.050 ;
        RECT 622.950 296.400 715.050 297.600 ;
        RECT 622.950 295.950 625.050 296.400 ;
        RECT 706.950 295.950 709.050 296.400 ;
        RECT 712.950 295.950 715.050 296.400 ;
        RECT 734.400 296.400 750.600 297.600 ;
        RECT 16.950 294.600 19.050 295.200 ;
        RECT 16.950 293.400 24.600 294.600 ;
        RECT 16.950 293.100 19.050 293.400 ;
        RECT 23.400 289.050 24.600 293.400 ;
        RECT 43.950 293.100 46.050 295.200 ;
        RECT 49.950 294.750 52.050 295.200 ;
        RECT 55.950 294.750 58.050 295.200 ;
        RECT 49.950 293.550 58.050 294.750 ;
        RECT 49.950 293.100 52.050 293.550 ;
        RECT 55.950 293.100 58.050 293.550 ;
        RECT 61.950 294.600 64.050 295.200 ;
        RECT 70.950 294.750 73.050 295.200 ;
        RECT 79.950 294.750 82.050 295.200 ;
        RECT 70.950 294.600 82.050 294.750 ;
        RECT 61.950 293.550 82.050 294.600 ;
        RECT 61.950 293.400 73.050 293.550 ;
        RECT 61.950 293.100 64.050 293.400 ;
        RECT 70.950 293.100 73.050 293.400 ;
        RECT 79.950 293.100 82.050 293.550 ;
        RECT 94.950 294.750 97.050 295.200 ;
        RECT 106.950 294.750 109.050 295.200 ;
        RECT 94.950 294.600 109.050 294.750 ;
        RECT 118.950 294.600 121.050 295.200 ;
        RECT 147.000 294.600 151.050 295.050 ;
        RECT 94.950 293.550 121.050 294.600 ;
        RECT 94.950 293.100 97.050 293.550 ;
        RECT 106.950 293.400 121.050 293.550 ;
        RECT 106.950 293.100 109.050 293.400 ;
        RECT 118.950 293.100 121.050 293.400 ;
        RECT 22.950 286.950 25.050 289.050 ;
        RECT 31.950 288.600 34.050 289.050 ;
        RECT 44.400 288.600 45.600 293.100 ;
        RECT 146.400 292.950 151.050 294.600 ;
        RECT 163.950 294.600 166.050 295.200 ;
        RECT 181.950 294.600 184.050 295.200 ;
        RECT 163.950 293.400 184.050 294.600 ;
        RECT 163.950 293.100 166.050 293.400 ;
        RECT 181.950 293.100 184.050 293.400 ;
        RECT 187.950 294.600 190.050 295.200 ;
        RECT 223.950 294.600 226.050 295.200 ;
        RECT 235.950 294.600 238.050 295.200 ;
        RECT 253.950 294.600 256.050 295.050 ;
        RECT 277.950 294.600 280.050 295.050 ;
        RECT 187.950 293.400 192.600 294.600 ;
        RECT 187.950 293.100 190.050 293.400 ;
        RECT 31.950 287.400 45.600 288.600 ;
        RECT 58.950 288.450 61.050 288.900 ;
        RECT 73.950 288.450 76.050 288.900 ;
        RECT 31.950 286.950 34.050 287.400 ;
        RECT 58.950 287.250 76.050 288.450 ;
        RECT 58.950 286.800 61.050 287.250 ;
        RECT 73.950 286.800 76.050 287.250 ;
        RECT 94.950 288.450 97.050 288.900 ;
        RECT 121.950 288.600 124.050 288.900 ;
        RECT 136.950 288.600 139.050 289.050 ;
        RECT 121.950 288.450 139.050 288.600 ;
        RECT 94.950 287.400 139.050 288.450 ;
        RECT 94.950 287.250 124.050 287.400 ;
        RECT 94.950 286.800 97.050 287.250 ;
        RECT 121.950 286.800 124.050 287.250 ;
        RECT 136.950 286.950 139.050 287.400 ;
        RECT 142.950 288.600 145.050 288.900 ;
        RECT 146.400 288.600 147.600 292.950 ;
        RECT 191.400 289.050 192.600 293.400 ;
        RECT 223.950 293.400 238.050 294.600 ;
        RECT 223.950 293.100 226.050 293.400 ;
        RECT 235.950 293.100 238.050 293.400 ;
        RECT 242.400 293.400 280.050 294.600 ;
        RECT 242.400 291.600 243.600 293.400 ;
        RECT 253.950 292.950 256.050 293.400 ;
        RECT 277.950 292.950 280.050 293.400 ;
        RECT 307.950 293.100 310.050 295.200 ;
        RECT 308.400 291.600 309.600 293.100 ;
        RECT 319.950 292.950 322.050 295.050 ;
        RECT 340.950 294.750 343.050 295.200 ;
        RECT 346.950 294.750 349.050 295.200 ;
        RECT 340.950 293.550 349.050 294.750 ;
        RECT 340.950 293.100 343.050 293.550 ;
        RECT 346.950 293.100 349.050 293.550 ;
        RECT 361.950 294.600 364.050 295.200 ;
        RECT 388.950 294.750 391.050 295.200 ;
        RECT 397.950 294.750 400.050 295.200 ;
        RECT 361.950 293.400 369.600 294.600 ;
        RECT 361.950 293.100 364.050 293.400 ;
        RECT 239.400 290.400 243.600 291.600 ;
        RECT 281.400 290.400 309.600 291.600 ;
        RECT 142.950 287.400 147.600 288.600 ;
        RECT 154.950 288.600 157.050 289.050 ;
        RECT 178.950 288.600 181.050 288.900 ;
        RECT 154.950 287.400 181.050 288.600 ;
        RECT 142.950 286.800 145.050 287.400 ;
        RECT 154.950 286.950 157.050 287.400 ;
        RECT 178.950 286.800 181.050 287.400 ;
        RECT 190.950 286.950 193.050 289.050 ;
        RECT 239.400 288.900 240.600 290.400 ;
        RECT 281.400 289.050 282.600 290.400 ;
        RECT 238.950 288.600 241.050 288.900 ;
        RECT 197.400 287.400 241.050 288.600 ;
        RECT 197.400 286.050 198.600 287.400 ;
        RECT 238.950 286.800 241.050 287.400 ;
        RECT 277.950 287.400 282.600 289.050 ;
        RECT 283.950 288.450 286.050 288.900 ;
        RECT 301.950 288.450 304.050 288.900 ;
        RECT 277.950 286.950 282.000 287.400 ;
        RECT 283.950 287.250 304.050 288.450 ;
        RECT 283.950 286.800 286.050 287.250 ;
        RECT 301.950 286.800 304.050 287.250 ;
        RECT 310.950 288.600 313.050 288.900 ;
        RECT 320.400 288.600 321.600 292.950 ;
        RECT 368.400 291.600 369.600 293.400 ;
        RECT 388.950 293.550 400.050 294.750 ;
        RECT 388.950 293.100 391.050 293.550 ;
        RECT 397.950 293.100 400.050 293.550 ;
        RECT 368.400 290.400 375.600 291.600 ;
        RECT 310.950 287.400 321.600 288.600 ;
        RECT 337.950 288.600 340.050 288.900 ;
        RECT 349.950 288.600 352.050 289.050 ;
        RECT 337.950 287.400 352.050 288.600 ;
        RECT 310.950 286.800 313.050 287.400 ;
        RECT 337.950 286.800 340.050 287.400 ;
        RECT 349.950 286.950 352.050 287.400 ;
        RECT 364.950 288.600 367.050 288.900 ;
        RECT 370.950 288.600 373.050 289.050 ;
        RECT 364.950 287.400 373.050 288.600 ;
        RECT 374.400 288.600 375.600 290.400 ;
        RECT 401.400 288.900 402.600 295.950 ;
        RECT 457.950 294.600 460.050 295.200 ;
        RECT 446.400 293.400 460.050 294.600 ;
        RECT 446.400 291.600 447.600 293.400 ;
        RECT 457.950 293.100 460.050 293.400 ;
        RECT 469.800 294.000 471.900 295.050 ;
        RECT 472.950 294.600 475.050 295.050 ;
        RECT 478.950 294.600 481.050 295.200 ;
        RECT 469.800 292.950 472.050 294.000 ;
        RECT 472.950 293.400 481.050 294.600 ;
        RECT 472.950 292.950 475.050 293.400 ;
        RECT 478.950 293.100 481.050 293.400 ;
        RECT 493.950 293.100 496.050 295.200 ;
        RECT 469.950 291.600 472.050 292.950 ;
        RECT 443.400 290.400 447.600 291.600 ;
        RECT 464.400 291.000 472.050 291.600 ;
        RECT 464.400 290.400 471.450 291.000 ;
        RECT 443.400 288.900 444.600 290.400 ;
        RECT 379.950 288.600 382.050 288.900 ;
        RECT 374.400 287.400 382.050 288.600 ;
        RECT 364.950 286.800 367.050 287.400 ;
        RECT 370.950 286.950 373.050 287.400 ;
        RECT 379.950 286.800 382.050 287.400 ;
        RECT 400.950 286.800 403.050 288.900 ;
        RECT 442.950 286.800 445.050 288.900 ;
        RECT 448.950 288.600 451.050 289.050 ;
        RECT 464.400 288.600 465.600 290.400 ;
        RECT 448.950 287.400 465.600 288.600 ;
        RECT 466.950 288.450 469.050 288.900 ;
        RECT 472.950 288.450 475.050 288.900 ;
        RECT 448.950 286.950 451.050 287.400 ;
        RECT 466.950 287.250 475.050 288.450 ;
        RECT 466.950 286.800 469.050 287.250 ;
        RECT 472.950 286.800 475.050 287.250 ;
        RECT 481.950 288.600 484.050 288.900 ;
        RECT 494.400 288.600 495.600 293.100 ;
        RECT 497.400 291.600 498.600 295.950 ;
        RECT 499.950 294.600 502.050 295.200 ;
        RECT 544.950 294.600 547.050 295.950 ;
        RECT 499.950 293.400 510.600 294.600 ;
        RECT 499.950 293.100 502.050 293.400 ;
        RECT 497.400 290.400 504.600 291.600 ;
        RECT 503.400 288.900 504.600 290.400 ;
        RECT 509.400 289.050 510.600 293.400 ;
        RECT 542.400 294.000 547.050 294.600 ;
        RECT 553.950 294.600 556.050 295.200 ;
        RECT 568.950 294.600 571.050 295.200 ;
        RECT 542.400 293.400 546.450 294.000 ;
        RECT 553.950 293.400 571.050 294.600 ;
        RECT 481.950 287.400 495.600 288.600 ;
        RECT 481.950 286.800 484.050 287.400 ;
        RECT 502.950 286.800 505.050 288.900 ;
        RECT 508.950 286.950 511.050 289.050 ;
        RECT 523.950 288.600 526.050 288.900 ;
        RECT 542.400 288.600 543.600 293.400 ;
        RECT 553.950 293.100 556.050 293.400 ;
        RECT 568.950 293.100 571.050 293.400 ;
        RECT 592.950 294.750 595.050 295.200 ;
        RECT 598.950 294.750 601.050 295.200 ;
        RECT 592.950 293.550 601.050 294.750 ;
        RECT 592.950 293.100 595.050 293.550 ;
        RECT 598.950 293.100 601.050 293.550 ;
        RECT 634.950 294.750 637.050 295.200 ;
        RECT 649.950 294.750 652.050 295.200 ;
        RECT 634.950 293.550 652.050 294.750 ;
        RECT 634.950 293.100 637.050 293.550 ;
        RECT 649.950 293.100 652.050 293.550 ;
        RECT 682.950 294.600 685.050 295.200 ;
        RECT 734.400 294.600 735.600 296.400 ;
        RECT 682.950 293.400 735.600 294.600 ;
        RECT 749.400 294.600 750.600 296.400 ;
        RECT 754.950 296.400 765.600 297.600 ;
        RECT 754.950 295.950 757.050 296.400 ;
        RECT 764.400 295.200 765.600 296.400 ;
        RECT 920.400 295.950 925.050 297.600 ;
        RECT 937.950 297.600 940.050 298.050 ;
        RECT 937.950 296.400 948.600 297.600 ;
        RECT 937.950 295.950 940.050 296.400 ;
        RECT 751.950 294.600 754.050 295.200 ;
        RECT 749.400 293.400 762.600 294.600 ;
        RECT 682.950 293.100 685.050 293.400 ;
        RECT 751.950 293.100 754.050 293.400 ;
        RECT 761.400 291.600 762.600 293.400 ;
        RECT 763.950 293.100 766.050 295.200 ;
        RECT 781.950 294.750 784.050 295.200 ;
        RECT 796.950 294.750 799.050 295.200 ;
        RECT 781.950 293.550 799.050 294.750 ;
        RECT 781.950 293.100 784.050 293.550 ;
        RECT 796.950 293.100 799.050 293.550 ;
        RECT 814.950 294.600 817.050 295.200 ;
        RECT 859.950 294.600 862.050 295.200 ;
        RECT 814.950 293.400 862.050 294.600 ;
        RECT 814.950 293.100 817.050 293.400 ;
        RECT 859.950 293.100 862.050 293.400 ;
        RECT 871.950 292.950 874.050 295.050 ;
        RECT 883.950 294.600 886.050 295.200 ;
        RECT 920.400 295.050 921.600 295.950 ;
        RECT 904.950 294.600 907.050 295.050 ;
        RECT 883.950 293.400 907.050 294.600 ;
        RECT 883.950 293.100 886.050 293.400 ;
        RECT 761.400 290.400 780.600 291.600 ;
        RECT 544.950 288.600 547.050 288.900 ;
        RECT 523.950 287.400 547.050 288.600 ;
        RECT 523.950 286.800 526.050 287.400 ;
        RECT 544.950 286.800 547.050 287.400 ;
        RECT 571.950 288.600 574.050 288.900 ;
        RECT 604.950 288.600 607.050 289.050 ;
        RECT 679.950 288.600 682.050 288.900 ;
        RECT 571.950 287.400 607.050 288.600 ;
        RECT 571.950 286.800 574.050 287.400 ;
        RECT 604.950 286.950 607.050 287.400 ;
        RECT 635.400 287.400 682.050 288.600 ;
        RECT 19.950 285.600 22.050 286.050 ;
        RECT 25.950 285.600 28.050 286.050 ;
        RECT 55.950 285.600 58.050 286.050 ;
        RECT 19.950 284.400 58.050 285.600 ;
        RECT 19.950 283.950 22.050 284.400 ;
        RECT 25.950 283.950 28.050 284.400 ;
        RECT 55.950 283.950 58.050 284.400 ;
        RECT 76.950 285.600 79.050 286.050 ;
        RECT 97.950 285.600 100.050 286.050 ;
        RECT 76.950 284.400 100.050 285.600 ;
        RECT 76.950 283.950 79.050 284.400 ;
        RECT 97.950 283.950 100.050 284.400 ;
        RECT 151.950 285.600 154.050 286.050 ;
        RECT 166.950 285.600 169.050 286.050 ;
        RECT 195.000 285.900 198.600 286.050 ;
        RECT 151.950 284.400 169.050 285.600 ;
        RECT 151.950 283.950 154.050 284.400 ;
        RECT 166.950 283.950 169.050 284.400 ;
        RECT 193.950 284.400 198.600 285.900 ;
        RECT 217.950 285.600 220.050 286.050 ;
        RECT 244.950 285.600 247.050 286.050 ;
        RECT 217.950 284.400 247.050 285.600 ;
        RECT 193.950 283.950 198.000 284.400 ;
        RECT 217.950 283.950 220.050 284.400 ;
        RECT 244.950 283.950 247.050 284.400 ;
        RECT 316.950 285.600 319.050 286.050 ;
        RECT 325.950 285.600 328.050 286.050 ;
        RECT 361.950 285.600 364.050 286.050 ;
        RECT 316.950 284.400 364.050 285.600 ;
        RECT 316.950 283.950 319.050 284.400 ;
        RECT 325.950 283.950 328.050 284.400 ;
        RECT 361.950 283.950 364.050 284.400 ;
        RECT 382.950 285.600 385.050 286.050 ;
        RECT 391.950 285.600 394.050 286.050 ;
        RECT 382.950 284.400 394.050 285.600 ;
        RECT 382.950 283.950 385.050 284.400 ;
        RECT 391.950 283.950 394.050 284.400 ;
        RECT 487.950 285.600 490.050 286.050 ;
        RECT 496.950 285.600 499.050 286.050 ;
        RECT 514.950 285.600 517.050 286.050 ;
        RECT 487.950 284.400 517.050 285.600 ;
        RECT 487.950 283.950 490.050 284.400 ;
        RECT 496.950 283.950 499.050 284.400 ;
        RECT 514.950 283.950 517.050 284.400 ;
        RECT 550.950 285.600 553.050 286.050 ;
        RECT 562.950 285.600 565.050 286.050 ;
        RECT 550.950 284.400 565.050 285.600 ;
        RECT 550.950 283.950 553.050 284.400 ;
        RECT 562.950 283.950 565.050 284.400 ;
        RECT 595.950 285.600 598.050 286.050 ;
        RECT 635.400 285.600 636.600 287.400 ;
        RECT 679.950 286.800 682.050 287.400 ;
        RECT 712.950 288.450 715.050 288.900 ;
        RECT 724.950 288.450 727.050 288.900 ;
        RECT 712.950 287.250 727.050 288.450 ;
        RECT 712.950 286.800 715.050 287.250 ;
        RECT 724.950 286.800 727.050 287.250 ;
        RECT 748.950 288.600 751.050 288.900 ;
        RECT 757.950 288.600 760.050 289.050 ;
        RECT 779.400 288.900 780.600 290.400 ;
        RECT 748.950 287.400 760.050 288.600 ;
        RECT 748.950 286.800 751.050 287.400 ;
        RECT 757.950 286.950 760.050 287.400 ;
        RECT 778.950 286.800 781.050 288.900 ;
        RECT 799.950 288.600 802.050 288.900 ;
        RECT 829.950 288.600 832.050 288.900 ;
        RECT 844.950 288.600 847.050 288.900 ;
        RECT 799.950 287.400 847.050 288.600 ;
        RECT 872.400 288.600 873.600 292.950 ;
        RECT 893.400 291.600 894.600 293.400 ;
        RECT 904.950 292.950 907.050 293.400 ;
        RECT 910.950 294.600 915.000 295.050 ;
        RECT 910.950 292.950 915.600 294.600 ;
        RECT 919.950 292.950 922.050 295.050 ;
        RECT 925.950 294.750 928.050 295.200 ;
        RECT 934.950 294.750 937.050 295.200 ;
        RECT 925.950 293.550 937.050 294.750 ;
        RECT 925.950 293.100 928.050 293.550 ;
        RECT 934.950 293.100 937.050 293.550 ;
        RECT 943.950 292.950 946.050 295.050 ;
        RECT 893.400 290.400 897.600 291.600 ;
        RECT 874.950 288.600 877.050 288.900 ;
        RECT 872.400 287.400 877.050 288.600 ;
        RECT 896.400 288.600 897.600 290.400 ;
        RECT 910.950 288.600 913.050 289.050 ;
        RECT 896.400 287.400 913.050 288.600 ;
        RECT 914.400 288.600 915.600 292.950 ;
        RECT 916.950 288.600 919.050 288.900 ;
        RECT 914.400 287.400 919.050 288.600 ;
        RECT 799.950 286.800 802.050 287.400 ;
        RECT 829.950 286.800 832.050 287.400 ;
        RECT 844.950 286.800 847.050 287.400 ;
        RECT 874.950 286.800 877.050 287.400 ;
        RECT 910.950 286.950 913.050 287.400 ;
        RECT 916.950 286.800 919.050 287.400 ;
        RECT 922.950 288.450 925.050 288.900 ;
        RECT 931.950 288.450 934.050 288.900 ;
        RECT 922.950 287.250 934.050 288.450 ;
        RECT 922.950 286.800 925.050 287.250 ;
        RECT 931.950 286.800 934.050 287.250 ;
        RECT 937.950 288.600 940.050 288.900 ;
        RECT 944.400 288.600 945.600 292.950 ;
        RECT 937.950 287.400 945.600 288.600 ;
        RECT 937.950 286.800 940.050 287.400 ;
        RECT 947.400 286.050 948.600 296.400 ;
        RECT 595.950 284.400 636.600 285.600 ;
        RECT 637.950 285.600 640.050 286.050 ;
        RECT 874.950 285.600 877.050 286.050 ;
        RECT 895.950 285.600 898.050 286.050 ;
        RECT 637.950 284.400 723.600 285.600 ;
        RECT 595.950 283.950 598.050 284.400 ;
        RECT 637.950 283.950 640.050 284.400 ;
        RECT 193.950 283.800 196.050 283.950 ;
        RECT 13.950 282.600 16.050 283.050 ;
        RECT 28.950 282.600 31.050 283.050 ;
        RECT 103.950 282.600 106.050 283.050 ;
        RECT 13.950 281.400 106.050 282.600 ;
        RECT 13.950 280.950 16.050 281.400 ;
        RECT 28.950 280.950 31.050 281.400 ;
        RECT 103.950 280.950 106.050 281.400 ;
        RECT 112.950 282.600 115.050 283.050 ;
        RECT 127.950 282.600 130.050 283.050 ;
        RECT 112.950 281.400 130.050 282.600 ;
        RECT 112.950 280.950 115.050 281.400 ;
        RECT 127.950 280.950 130.050 281.400 ;
        RECT 139.950 282.600 142.050 283.050 ;
        RECT 202.950 282.600 205.050 283.050 ;
        RECT 139.950 281.400 205.050 282.600 ;
        RECT 139.950 280.950 142.050 281.400 ;
        RECT 202.950 280.950 205.050 281.400 ;
        RECT 256.950 282.600 259.050 283.050 ;
        RECT 283.950 282.600 286.050 283.050 ;
        RECT 256.950 281.400 286.050 282.600 ;
        RECT 256.950 280.950 259.050 281.400 ;
        RECT 283.950 280.950 286.050 281.400 ;
        RECT 295.950 282.600 298.050 283.050 ;
        RECT 367.950 282.600 370.050 283.050 ;
        RECT 295.950 281.400 370.050 282.600 ;
        RECT 295.950 280.950 298.050 281.400 ;
        RECT 367.950 280.950 370.050 281.400 ;
        RECT 376.950 282.600 379.050 283.050 ;
        RECT 415.950 282.600 418.050 283.050 ;
        RECT 376.950 281.400 418.050 282.600 ;
        RECT 376.950 280.950 379.050 281.400 ;
        RECT 415.950 280.950 418.050 281.400 ;
        RECT 589.950 282.600 592.050 283.050 ;
        RECT 625.950 282.600 628.050 283.050 ;
        RECT 589.950 281.400 628.050 282.600 ;
        RECT 722.400 282.600 723.600 284.400 ;
        RECT 874.950 284.400 898.050 285.600 ;
        RECT 874.950 283.950 877.050 284.400 ;
        RECT 895.950 283.950 898.050 284.400 ;
        RECT 943.950 284.400 948.600 286.050 ;
        RECT 943.950 283.950 948.000 284.400 ;
        RECT 799.950 282.600 802.050 283.050 ;
        RECT 722.400 281.400 802.050 282.600 ;
        RECT 589.950 280.950 592.050 281.400 ;
        RECT 625.950 280.950 628.050 281.400 ;
        RECT 799.950 280.950 802.050 281.400 ;
        RECT 22.950 279.600 25.050 280.050 ;
        RECT 34.950 279.600 37.050 280.050 ;
        RECT 22.950 278.400 37.050 279.600 ;
        RECT 22.950 277.950 25.050 278.400 ;
        RECT 34.950 277.950 37.050 278.400 ;
        RECT 40.950 279.600 43.050 280.050 ;
        RECT 49.950 279.600 52.050 280.050 ;
        RECT 82.950 279.600 85.050 280.050 ;
        RECT 40.950 278.400 85.050 279.600 ;
        RECT 40.950 277.950 43.050 278.400 ;
        RECT 49.950 277.950 52.050 278.400 ;
        RECT 82.950 277.950 85.050 278.400 ;
        RECT 88.950 279.600 91.050 280.050 ;
        RECT 160.950 279.600 163.050 280.050 ;
        RECT 187.950 279.600 190.050 280.050 ;
        RECT 88.950 278.400 190.050 279.600 ;
        RECT 88.950 277.950 91.050 278.400 ;
        RECT 160.950 277.950 163.050 278.400 ;
        RECT 187.950 277.950 190.050 278.400 ;
        RECT 220.950 279.600 223.050 280.050 ;
        RECT 229.950 279.600 232.050 280.050 ;
        RECT 220.950 278.400 232.050 279.600 ;
        RECT 220.950 277.950 223.050 278.400 ;
        RECT 229.950 277.950 232.050 278.400 ;
        RECT 292.950 279.600 295.050 280.050 ;
        RECT 364.950 279.600 367.050 280.050 ;
        RECT 373.950 279.600 376.050 280.050 ;
        RECT 292.950 278.400 312.600 279.600 ;
        RECT 292.950 277.950 295.050 278.400 ;
        RECT 97.950 276.600 100.050 277.050 ;
        RECT 112.950 276.600 115.050 277.050 ;
        RECT 97.950 275.400 115.050 276.600 ;
        RECT 97.950 274.950 100.050 275.400 ;
        RECT 112.950 274.950 115.050 275.400 ;
        RECT 211.950 276.600 214.050 277.050 ;
        RECT 235.950 276.600 238.050 277.050 ;
        RECT 241.950 276.600 244.050 277.050 ;
        RECT 271.950 276.600 274.050 277.050 ;
        RECT 211.950 275.400 274.050 276.600 ;
        RECT 211.950 274.950 214.050 275.400 ;
        RECT 235.950 274.950 238.050 275.400 ;
        RECT 241.950 274.950 244.050 275.400 ;
        RECT 271.950 274.950 274.050 275.400 ;
        RECT 277.950 276.600 280.050 277.050 ;
        RECT 307.950 276.600 310.050 277.050 ;
        RECT 277.950 275.400 310.050 276.600 ;
        RECT 311.400 276.600 312.600 278.400 ;
        RECT 364.950 278.400 376.050 279.600 ;
        RECT 364.950 277.950 367.050 278.400 ;
        RECT 373.950 277.950 376.050 278.400 ;
        RECT 433.950 279.600 436.050 280.050 ;
        RECT 445.950 279.600 448.050 280.050 ;
        RECT 433.950 278.400 448.050 279.600 ;
        RECT 433.950 277.950 436.050 278.400 ;
        RECT 445.950 277.950 448.050 278.400 ;
        RECT 460.950 279.600 463.050 280.050 ;
        RECT 469.950 279.600 472.050 280.050 ;
        RECT 460.950 278.400 472.050 279.600 ;
        RECT 460.950 277.950 463.050 278.400 ;
        RECT 469.950 277.950 472.050 278.400 ;
        RECT 517.950 279.600 520.050 280.050 ;
        RECT 574.950 279.600 577.050 280.050 ;
        RECT 517.950 278.400 577.050 279.600 ;
        RECT 626.400 279.600 627.600 280.950 ;
        RECT 643.950 279.600 646.050 280.050 ;
        RECT 658.950 279.600 661.050 280.050 ;
        RECT 626.400 278.400 661.050 279.600 ;
        RECT 517.950 277.950 520.050 278.400 ;
        RECT 574.950 277.950 577.050 278.400 ;
        RECT 643.950 277.950 646.050 278.400 ;
        RECT 658.950 277.950 661.050 278.400 ;
        RECT 772.950 279.600 775.050 280.050 ;
        RECT 781.950 279.600 784.050 280.050 ;
        RECT 811.950 279.600 814.050 280.050 ;
        RECT 772.950 278.400 814.050 279.600 ;
        RECT 772.950 277.950 775.050 278.400 ;
        RECT 781.950 277.950 784.050 278.400 ;
        RECT 811.950 277.950 814.050 278.400 ;
        RECT 838.950 279.600 841.050 280.050 ;
        RECT 847.950 279.600 850.050 280.050 ;
        RECT 838.950 278.400 850.050 279.600 ;
        RECT 838.950 277.950 841.050 278.400 ;
        RECT 847.950 277.950 850.050 278.400 ;
        RECT 868.950 279.600 871.050 280.050 ;
        RECT 880.950 279.600 883.050 280.050 ;
        RECT 868.950 278.400 883.050 279.600 ;
        RECT 868.950 277.950 871.050 278.400 ;
        RECT 880.950 277.950 883.050 278.400 ;
        RECT 889.950 279.600 892.050 280.050 ;
        RECT 901.950 279.600 904.050 280.050 ;
        RECT 889.950 278.400 904.050 279.600 ;
        RECT 889.950 277.950 892.050 278.400 ;
        RECT 901.950 277.950 904.050 278.400 ;
        RECT 916.950 279.600 919.050 280.050 ;
        RECT 928.950 279.600 931.050 280.050 ;
        RECT 916.950 278.400 931.050 279.600 ;
        RECT 916.950 277.950 919.050 278.400 ;
        RECT 928.950 277.950 931.050 278.400 ;
        RECT 394.950 276.600 397.050 277.050 ;
        RECT 311.400 275.400 397.050 276.600 ;
        RECT 277.950 274.950 280.050 275.400 ;
        RECT 307.950 274.950 310.050 275.400 ;
        RECT 394.950 274.950 397.050 275.400 ;
        RECT 412.950 276.600 415.050 277.050 ;
        RECT 481.950 276.600 484.050 277.050 ;
        RECT 412.950 275.400 484.050 276.600 ;
        RECT 412.950 274.950 415.050 275.400 ;
        RECT 481.950 274.950 484.050 275.400 ;
        RECT 532.950 276.600 535.050 277.050 ;
        RECT 556.950 276.600 559.050 277.050 ;
        RECT 532.950 275.400 559.050 276.600 ;
        RECT 532.950 274.950 535.050 275.400 ;
        RECT 556.950 274.950 559.050 275.400 ;
        RECT 718.950 276.600 721.050 277.050 ;
        RECT 727.950 276.600 730.050 277.050 ;
        RECT 718.950 275.400 730.050 276.600 ;
        RECT 718.950 274.950 721.050 275.400 ;
        RECT 727.950 274.950 730.050 275.400 ;
        RECT 793.950 276.600 796.050 277.050 ;
        RECT 805.950 276.600 808.050 277.050 ;
        RECT 793.950 275.400 808.050 276.600 ;
        RECT 793.950 274.950 796.050 275.400 ;
        RECT 805.950 274.950 808.050 275.400 ;
        RECT 64.950 273.600 67.050 274.050 ;
        RECT 145.950 273.600 148.050 274.050 ;
        RECT 178.950 273.600 181.050 274.050 ;
        RECT 184.950 273.600 187.050 274.050 ;
        RECT 64.950 272.400 187.050 273.600 ;
        RECT 64.950 271.950 67.050 272.400 ;
        RECT 145.950 271.950 148.050 272.400 ;
        RECT 178.950 271.950 181.050 272.400 ;
        RECT 184.950 271.950 187.050 272.400 ;
        RECT 268.950 273.600 271.050 274.050 ;
        RECT 331.950 273.600 334.050 274.050 ;
        RECT 268.950 272.400 334.050 273.600 ;
        RECT 268.950 271.950 271.050 272.400 ;
        RECT 331.950 271.950 334.050 272.400 ;
        RECT 415.950 273.600 418.050 274.050 ;
        RECT 457.950 273.600 460.050 274.050 ;
        RECT 415.950 272.400 460.050 273.600 ;
        RECT 415.950 271.950 418.050 272.400 ;
        RECT 457.950 271.950 460.050 272.400 ;
        RECT 493.950 273.600 496.050 274.050 ;
        RECT 508.950 273.600 511.050 274.050 ;
        RECT 493.950 272.400 511.050 273.600 ;
        RECT 493.950 271.950 496.050 272.400 ;
        RECT 508.950 271.950 511.050 272.400 ;
        RECT 550.950 273.600 553.050 274.050 ;
        RECT 559.950 273.600 562.050 274.050 ;
        RECT 550.950 272.400 562.050 273.600 ;
        RECT 550.950 271.950 553.050 272.400 ;
        RECT 559.950 271.950 562.050 272.400 ;
        RECT 616.950 273.600 619.050 274.050 ;
        RECT 646.950 273.600 649.050 274.050 ;
        RECT 616.950 272.400 649.050 273.600 ;
        RECT 616.950 271.950 619.050 272.400 ;
        RECT 646.950 271.950 649.050 272.400 ;
        RECT 925.950 273.600 928.050 274.050 ;
        RECT 934.950 273.600 937.050 274.050 ;
        RECT 925.950 272.400 937.050 273.600 ;
        RECT 925.950 271.950 928.050 272.400 ;
        RECT 934.950 271.950 937.050 272.400 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 118.950 270.600 121.050 271.050 ;
        RECT 106.950 269.400 121.050 270.600 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 118.950 268.950 121.050 269.400 ;
        RECT 154.950 270.600 157.050 271.050 ;
        RECT 169.950 270.600 172.050 271.050 ;
        RECT 154.950 269.400 172.050 270.600 ;
        RECT 154.950 268.950 157.050 269.400 ;
        RECT 169.950 268.950 172.050 269.400 ;
        RECT 190.950 270.600 193.050 271.050 ;
        RECT 205.950 270.600 208.050 271.050 ;
        RECT 238.950 270.600 241.050 271.050 ;
        RECT 190.950 269.400 241.050 270.600 ;
        RECT 190.950 268.950 193.050 269.400 ;
        RECT 205.950 268.950 208.050 269.400 ;
        RECT 238.950 268.950 241.050 269.400 ;
        RECT 271.950 270.600 274.050 271.050 ;
        RECT 280.950 270.600 283.050 271.050 ;
        RECT 271.950 269.400 283.050 270.600 ;
        RECT 271.950 268.950 274.050 269.400 ;
        RECT 280.950 268.950 283.050 269.400 ;
        RECT 298.950 270.600 301.050 271.050 ;
        RECT 376.950 270.600 379.050 271.050 ;
        RECT 298.950 269.400 379.050 270.600 ;
        RECT 298.950 268.950 301.050 269.400 ;
        RECT 376.950 268.950 379.050 269.400 ;
        RECT 430.950 270.600 433.050 271.050 ;
        RECT 454.950 270.600 457.050 271.050 ;
        RECT 580.950 270.600 583.050 271.050 ;
        RECT 430.950 269.400 457.050 270.600 ;
        RECT 430.950 268.950 433.050 269.400 ;
        RECT 454.950 268.950 457.050 269.400 ;
        RECT 464.400 269.400 583.050 270.600 ;
        RECT 464.400 268.050 465.600 269.400 ;
        RECT 580.950 268.950 583.050 269.400 ;
        RECT 598.950 270.600 601.050 271.050 ;
        RECT 616.950 270.600 619.050 270.900 ;
        RECT 598.950 269.400 619.050 270.600 ;
        RECT 598.950 268.950 601.050 269.400 ;
        RECT 616.950 268.800 619.050 269.400 ;
        RECT 718.950 270.600 721.050 271.050 ;
        RECT 751.950 270.600 754.050 271.050 ;
        RECT 718.950 269.400 754.050 270.600 ;
        RECT 718.950 268.950 721.050 269.400 ;
        RECT 751.950 268.950 754.050 269.400 ;
        RECT 883.950 270.600 886.050 271.050 ;
        RECT 907.950 270.600 910.050 271.050 ;
        RECT 919.950 270.600 922.050 271.050 ;
        RECT 883.950 269.400 922.050 270.600 ;
        RECT 883.950 268.950 886.050 269.400 ;
        RECT 907.950 268.950 910.050 269.400 ;
        RECT 919.950 268.950 922.050 269.400 ;
        RECT 49.950 267.600 52.050 268.050 ;
        RECT 73.950 267.600 76.050 268.050 ;
        RECT 49.950 266.400 76.050 267.600 ;
        RECT 49.950 265.950 52.050 266.400 ;
        RECT 73.950 265.950 76.050 266.400 ;
        RECT 91.950 267.600 94.050 268.050 ;
        RECT 226.950 267.600 229.050 268.050 ;
        RECT 91.950 266.400 229.050 267.600 ;
        RECT 91.950 265.950 94.050 266.400 ;
        RECT 226.950 265.950 229.050 266.400 ;
        RECT 283.950 267.600 286.050 268.050 ;
        RECT 295.950 267.600 298.050 268.050 ;
        RECT 283.950 266.400 298.050 267.600 ;
        RECT 283.950 265.950 286.050 266.400 ;
        RECT 295.950 265.950 298.050 266.400 ;
        RECT 358.950 267.600 361.050 268.050 ;
        RECT 388.950 267.600 391.050 268.050 ;
        RECT 358.950 266.400 391.050 267.600 ;
        RECT 358.950 265.950 361.050 266.400 ;
        RECT 388.950 265.950 391.050 266.400 ;
        RECT 394.950 267.600 397.050 268.050 ;
        RECT 436.950 267.600 439.050 268.050 ;
        RECT 394.950 266.400 439.050 267.600 ;
        RECT 394.950 265.950 397.050 266.400 ;
        RECT 436.950 265.950 439.050 266.400 ;
        RECT 442.950 267.600 445.050 268.050 ;
        RECT 463.950 267.600 466.050 268.050 ;
        RECT 442.950 266.400 466.050 267.600 ;
        RECT 442.950 265.950 445.050 266.400 ;
        RECT 463.950 265.950 466.050 266.400 ;
        RECT 484.950 267.600 487.050 268.050 ;
        RECT 535.950 267.600 538.050 268.050 ;
        RECT 484.950 266.400 538.050 267.600 ;
        RECT 484.950 265.950 487.050 266.400 ;
        RECT 535.950 265.950 538.050 266.400 ;
        RECT 634.950 267.600 637.050 268.050 ;
        RECT 664.950 267.600 667.050 268.050 ;
        RECT 634.950 266.400 667.050 267.600 ;
        RECT 634.950 265.950 637.050 266.400 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 784.950 267.600 787.050 268.050 ;
        RECT 793.950 267.600 796.050 268.050 ;
        RECT 784.950 266.400 796.050 267.600 ;
        RECT 784.950 265.950 787.050 266.400 ;
        RECT 793.950 265.950 796.050 266.400 ;
        RECT 937.950 267.600 940.050 268.050 ;
        RECT 946.950 267.600 949.050 268.050 ;
        RECT 937.950 266.400 949.050 267.600 ;
        RECT 937.950 265.950 940.050 266.400 ;
        RECT 946.950 265.950 949.050 266.400 ;
        RECT 21.000 264.600 25.050 265.050 ;
        RECT 20.400 262.950 25.050 264.600 ;
        RECT 28.950 264.600 31.050 265.050 ;
        RECT 55.950 264.600 58.050 265.050 ;
        RECT 85.950 264.600 88.050 265.050 ;
        RECT 28.950 263.400 39.600 264.600 ;
        RECT 28.950 262.950 31.050 263.400 ;
        RECT 7.950 261.750 10.050 262.200 ;
        RECT 16.950 261.750 19.050 262.200 ;
        RECT 7.950 260.550 19.050 261.750 ;
        RECT 7.950 260.100 10.050 260.550 ;
        RECT 16.950 260.100 19.050 260.550 ;
        RECT 20.400 255.900 21.600 262.950 ;
        RECT 28.950 261.750 31.050 261.900 ;
        RECT 34.950 261.750 37.050 262.200 ;
        RECT 28.950 260.550 37.050 261.750 ;
        RECT 28.950 259.800 31.050 260.550 ;
        RECT 34.950 260.100 37.050 260.550 ;
        RECT 38.400 255.900 39.600 263.400 ;
        RECT 55.950 263.400 88.050 264.600 ;
        RECT 55.950 262.950 58.050 263.400 ;
        RECT 85.950 262.950 88.050 263.400 ;
        RECT 97.950 264.600 100.050 265.050 ;
        RECT 103.950 264.600 106.050 265.050 ;
        RECT 97.950 263.400 106.050 264.600 ;
        RECT 97.950 262.950 100.050 263.400 ;
        RECT 103.950 262.950 106.050 263.400 ;
        RECT 136.950 264.600 139.050 265.050 ;
        RECT 184.800 264.600 186.900 265.050 ;
        RECT 136.950 263.400 186.900 264.600 ;
        RECT 136.950 262.950 139.050 263.400 ;
        RECT 184.800 262.950 186.900 263.400 ;
        RECT 187.950 262.950 190.050 265.050 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 478.950 264.600 481.050 265.050 ;
        RECT 529.950 264.600 532.050 265.050 ;
        RECT 454.950 263.400 481.050 264.600 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 478.950 262.950 481.050 263.400 ;
        RECT 497.400 263.400 532.050 264.600 ;
        RECT 40.950 261.600 43.050 262.200 ;
        RECT 52.950 261.600 55.050 262.050 ;
        RECT 40.950 260.400 55.050 261.600 ;
        RECT 40.950 260.100 43.050 260.400 ;
        RECT 52.950 259.950 55.050 260.400 ;
        RECT 61.950 260.100 64.050 262.200 ;
        RECT 112.800 260.100 115.050 262.200 ;
        RECT 115.950 261.750 118.050 262.200 ;
        RECT 121.950 261.750 124.050 262.050 ;
        RECT 130.800 261.750 132.900 262.200 ;
        RECT 115.950 260.550 132.900 261.750 ;
        RECT 115.950 260.100 118.050 260.550 ;
        RECT 19.950 253.800 22.050 255.900 ;
        RECT 37.950 253.800 40.050 255.900 ;
        RECT 43.950 255.450 46.050 255.900 ;
        RECT 49.950 255.450 52.050 255.900 ;
        RECT 43.950 254.250 52.050 255.450 ;
        RECT 43.950 253.800 46.050 254.250 ;
        RECT 49.950 253.800 52.050 254.250 ;
        RECT 55.950 255.600 58.050 256.050 ;
        RECT 62.400 255.600 63.600 260.100 ;
        RECT 113.400 258.600 114.600 260.100 ;
        RECT 121.950 259.950 124.050 260.550 ;
        RECT 130.800 260.100 132.900 260.550 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 178.950 261.600 183.000 262.050 ;
        RECT 178.950 259.950 183.600 261.600 ;
        RECT 113.400 257.400 120.600 258.600 ;
        RECT 55.950 254.400 63.600 255.600 ;
        RECT 64.950 255.600 67.050 255.900 ;
        RECT 73.950 255.600 76.050 256.050 ;
        RECT 79.950 255.600 82.050 255.900 ;
        RECT 64.950 254.400 82.050 255.600 ;
        RECT 55.950 253.950 58.050 254.400 ;
        RECT 64.950 253.800 67.050 254.400 ;
        RECT 73.950 253.950 76.050 254.400 ;
        RECT 79.950 253.800 82.050 254.400 ;
        RECT 88.950 255.600 91.050 255.900 ;
        RECT 97.950 255.600 100.050 255.900 ;
        RECT 88.950 255.450 100.050 255.600 ;
        RECT 103.950 255.450 106.050 255.900 ;
        RECT 88.950 254.400 106.050 255.450 ;
        RECT 119.400 255.600 120.600 257.400 ;
        RECT 134.400 256.050 135.600 259.950 ;
        RECT 124.950 255.600 127.050 256.050 ;
        RECT 119.400 254.400 127.050 255.600 ;
        RECT 88.950 253.800 91.050 254.400 ;
        RECT 97.950 254.250 106.050 254.400 ;
        RECT 97.950 253.800 100.050 254.250 ;
        RECT 103.950 253.800 106.050 254.250 ;
        RECT 124.950 253.950 127.050 254.400 ;
        RECT 133.950 253.950 136.050 256.050 ;
        RECT 182.400 255.900 183.600 259.950 ;
        RECT 188.400 255.900 189.600 262.950 ;
        RECT 190.950 261.600 193.050 262.200 ;
        RECT 214.950 261.750 217.050 262.200 ;
        RECT 226.950 261.750 229.050 262.200 ;
        RECT 190.950 260.400 201.600 261.600 ;
        RECT 190.950 260.100 193.050 260.400 ;
        RECT 148.950 255.600 151.050 255.900 ;
        RECT 163.950 255.600 166.050 255.900 ;
        RECT 148.950 254.400 166.050 255.600 ;
        RECT 148.950 253.800 151.050 254.400 ;
        RECT 163.950 253.800 166.050 254.400 ;
        RECT 181.950 253.800 184.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 193.950 255.600 196.050 256.050 ;
        RECT 200.400 255.600 201.600 260.400 ;
        RECT 214.950 260.550 229.050 261.750 ;
        RECT 214.950 260.100 217.050 260.550 ;
        RECT 226.950 260.100 229.050 260.550 ;
        RECT 238.950 258.600 241.050 262.050 ;
        RECT 265.950 261.750 268.050 262.200 ;
        RECT 274.950 261.750 277.050 262.200 ;
        RECT 265.950 260.550 277.050 261.750 ;
        RECT 265.950 260.100 268.050 260.550 ;
        RECT 274.950 260.100 277.050 260.550 ;
        RECT 286.950 260.100 289.050 262.200 ;
        RECT 328.950 261.750 331.050 262.200 ;
        RECT 337.800 261.750 339.900 262.200 ;
        RECT 328.950 260.550 339.900 261.750 ;
        RECT 328.950 260.100 331.050 260.550 ;
        RECT 337.800 260.100 339.900 260.550 ;
        RECT 340.950 261.750 343.050 262.200 ;
        RECT 352.950 261.750 355.050 262.200 ;
        RECT 340.950 260.550 355.050 261.750 ;
        RECT 340.950 260.100 343.050 260.550 ;
        RECT 352.950 260.100 355.050 260.550 ;
        RECT 367.950 261.600 370.050 262.050 ;
        RECT 406.950 261.600 409.050 262.050 ;
        RECT 367.950 260.400 409.050 261.600 ;
        RECT 238.950 258.000 246.600 258.600 ;
        RECT 239.400 257.400 246.600 258.000 ;
        RECT 245.400 255.900 246.600 257.400 ;
        RECT 208.950 255.600 211.050 255.900 ;
        RECT 193.950 254.400 211.050 255.600 ;
        RECT 193.950 253.950 196.050 254.400 ;
        RECT 208.950 253.800 211.050 254.400 ;
        RECT 244.950 255.600 247.050 255.900 ;
        RECT 262.950 255.600 265.050 255.900 ;
        RECT 287.400 255.600 288.600 260.100 ;
        RECT 367.950 259.950 370.050 260.400 ;
        RECT 406.950 259.950 409.050 260.400 ;
        RECT 418.950 261.750 421.050 262.200 ;
        RECT 430.950 261.750 433.050 262.200 ;
        RECT 418.950 260.550 433.050 261.750 ;
        RECT 418.950 260.100 421.050 260.550 ;
        RECT 430.950 260.100 433.050 260.550 ;
        RECT 436.950 261.600 439.050 262.200 ;
        RECT 484.950 261.600 487.050 262.200 ;
        RECT 436.950 260.400 487.050 261.600 ;
        RECT 436.950 260.100 439.050 260.400 ;
        RECT 484.950 260.100 487.050 260.400 ;
        RECT 361.950 258.600 364.050 259.050 ;
        RECT 427.950 258.600 430.050 259.050 ;
        RECT 361.950 257.400 430.050 258.600 ;
        RECT 361.950 256.950 364.050 257.400 ;
        RECT 427.950 256.950 430.050 257.400 ;
        RECT 497.400 256.050 498.600 263.400 ;
        RECT 529.950 262.950 532.050 263.400 ;
        RECT 553.950 264.600 556.050 265.050 ;
        RECT 562.950 264.600 565.050 265.050 ;
        RECT 553.950 263.400 565.050 264.600 ;
        RECT 553.950 262.950 556.050 263.400 ;
        RECT 562.950 262.950 565.050 263.400 ;
        RECT 586.950 264.600 589.050 265.050 ;
        RECT 622.950 264.600 625.050 265.050 ;
        RECT 586.950 263.400 625.050 264.600 ;
        RECT 586.950 262.950 589.050 263.400 ;
        RECT 622.950 262.950 625.050 263.400 ;
        RECT 667.950 264.600 670.050 265.050 ;
        RECT 679.950 264.600 682.050 265.050 ;
        RECT 685.950 264.600 688.050 265.050 ;
        RECT 667.950 263.400 688.050 264.600 ;
        RECT 667.950 262.950 670.050 263.400 ;
        RECT 679.950 262.950 682.050 263.400 ;
        RECT 685.950 262.950 688.050 263.400 ;
        RECT 691.950 264.600 694.050 265.050 ;
        RECT 706.950 264.600 709.050 265.050 ;
        RECT 691.950 263.400 709.050 264.600 ;
        RECT 691.950 262.950 694.050 263.400 ;
        RECT 706.950 262.950 709.050 263.400 ;
        RECT 733.950 262.950 736.050 265.050 ;
        RECT 760.950 264.600 763.050 265.050 ;
        RECT 772.950 264.600 775.050 265.050 ;
        RECT 781.950 264.600 784.050 265.050 ;
        RECT 760.950 263.400 784.050 264.600 ;
        RECT 760.950 262.950 763.050 263.400 ;
        RECT 772.950 262.950 775.050 263.400 ;
        RECT 781.950 262.950 784.050 263.400 ;
        RECT 808.950 264.600 811.050 265.050 ;
        RECT 817.950 264.600 820.050 265.050 ;
        RECT 823.950 264.600 826.050 265.050 ;
        RECT 808.950 263.400 826.050 264.600 ;
        RECT 808.950 262.950 811.050 263.400 ;
        RECT 817.950 262.950 820.050 263.400 ;
        RECT 823.950 262.950 826.050 263.400 ;
        RECT 850.950 264.600 853.050 265.050 ;
        RECT 904.950 264.600 907.050 265.050 ;
        RECT 913.950 264.600 916.050 265.050 ;
        RECT 850.950 263.400 861.600 264.600 ;
        RECT 850.950 262.950 853.050 263.400 ;
        RECT 502.950 261.600 505.050 262.200 ;
        RECT 523.950 261.600 526.050 262.200 ;
        RECT 502.950 260.400 507.600 261.600 ;
        RECT 502.950 260.100 505.050 260.400 ;
        RECT 244.950 254.400 265.050 255.600 ;
        RECT 244.950 253.800 247.050 254.400 ;
        RECT 262.950 253.800 265.050 254.400 ;
        RECT 284.400 254.400 288.600 255.600 ;
        RECT 295.950 255.600 298.050 256.050 ;
        RECT 319.950 255.600 322.050 256.050 ;
        RECT 295.950 254.400 322.050 255.600 ;
        RECT 247.950 252.600 250.050 253.050 ;
        RECT 284.400 252.600 285.600 254.400 ;
        RECT 295.950 253.950 298.050 254.400 ;
        RECT 319.950 253.950 322.050 254.400 ;
        RECT 334.950 255.600 337.050 256.050 ;
        RECT 364.950 255.600 367.050 256.050 ;
        RECT 421.950 255.600 424.050 256.050 ;
        RECT 334.950 254.400 424.050 255.600 ;
        RECT 334.950 253.950 337.050 254.400 ;
        RECT 364.950 253.950 367.050 254.400 ;
        RECT 421.950 253.950 424.050 254.400 ;
        RECT 445.950 255.450 448.050 255.900 ;
        RECT 487.950 255.450 490.050 255.900 ;
        RECT 445.950 254.250 490.050 255.450 ;
        RECT 445.950 253.800 448.050 254.250 ;
        RECT 487.950 253.800 490.050 254.250 ;
        RECT 496.950 253.950 499.050 256.050 ;
        RECT 506.400 253.050 507.600 260.400 ;
        RECT 521.250 260.400 526.050 261.600 ;
        RECT 508.950 255.600 511.050 256.050 ;
        RECT 514.950 255.600 517.050 256.050 ;
        RECT 508.950 254.400 517.050 255.600 ;
        RECT 508.950 253.950 511.050 254.400 ;
        RECT 514.950 253.950 517.050 254.400 ;
        RECT 521.250 253.050 522.450 260.400 ;
        RECT 523.950 260.100 526.050 260.400 ;
        RECT 535.950 261.750 538.050 262.200 ;
        RECT 541.950 261.750 544.050 262.200 ;
        RECT 535.950 260.550 544.050 261.750 ;
        RECT 535.950 260.100 538.050 260.550 ;
        RECT 541.950 260.100 544.050 260.550 ;
        RECT 571.950 261.750 574.050 262.050 ;
        RECT 586.950 261.750 589.050 262.200 ;
        RECT 571.950 260.550 589.050 261.750 ;
        RECT 571.950 259.950 574.050 260.550 ;
        RECT 586.950 260.100 589.050 260.550 ;
        RECT 592.950 261.600 595.050 262.050 ;
        RECT 601.950 261.600 604.050 262.200 ;
        RECT 592.950 260.400 604.050 261.600 ;
        RECT 592.950 259.950 595.050 260.400 ;
        RECT 601.950 260.100 604.050 260.400 ;
        RECT 607.950 261.600 610.050 262.200 ;
        RECT 619.950 261.600 622.050 262.050 ;
        RECT 649.950 261.600 652.050 262.050 ;
        RECT 607.950 260.400 622.050 261.600 ;
        RECT 644.400 261.000 652.050 261.600 ;
        RECT 607.950 260.100 610.050 260.400 ;
        RECT 619.950 259.950 622.050 260.400 ;
        RECT 643.950 260.400 652.050 261.000 ;
        RECT 643.950 256.950 646.050 260.400 ;
        RECT 649.950 259.950 652.050 260.400 ;
        RECT 655.950 261.600 658.050 262.200 ;
        RECT 664.950 261.600 667.050 261.900 ;
        RECT 655.950 260.400 667.050 261.600 ;
        RECT 655.950 260.100 658.050 260.400 ;
        RECT 664.950 259.800 667.050 260.400 ;
        RECT 673.950 261.600 676.050 262.200 ;
        RECT 694.950 261.600 697.050 262.200 ;
        RECT 703.950 261.750 706.050 262.200 ;
        RECT 712.950 261.750 715.050 262.200 ;
        RECT 673.950 260.400 678.600 261.600 ;
        RECT 673.950 260.100 676.050 260.400 ;
        RECT 677.400 258.600 678.600 260.400 ;
        RECT 694.950 260.400 702.600 261.600 ;
        RECT 694.950 260.100 697.050 260.400 ;
        RECT 701.400 258.600 702.600 260.400 ;
        RECT 703.950 260.550 715.050 261.750 ;
        RECT 703.950 260.100 706.050 260.550 ;
        RECT 712.950 260.100 715.050 260.550 ;
        RECT 671.400 258.000 693.600 258.600 ;
        RECT 670.950 257.400 693.600 258.000 ;
        RECT 701.400 258.000 726.600 258.600 ;
        RECT 701.400 257.400 727.050 258.000 ;
        RECT 529.950 255.600 532.050 256.050 ;
        RECT 547.950 255.600 550.050 256.050 ;
        RECT 529.950 254.400 550.050 255.600 ;
        RECT 529.950 253.950 532.050 254.400 ;
        RECT 547.950 253.950 550.050 254.400 ;
        RECT 559.950 255.600 562.050 255.900 ;
        RECT 571.950 255.600 574.050 256.050 ;
        RECT 559.950 254.400 574.050 255.600 ;
        RECT 559.950 253.800 562.050 254.400 ;
        RECT 571.950 253.950 574.050 254.400 ;
        RECT 646.950 255.450 649.050 255.900 ;
        RECT 652.950 255.450 655.050 255.900 ;
        RECT 646.950 254.250 655.050 255.450 ;
        RECT 646.950 253.800 649.050 254.250 ;
        RECT 652.950 253.800 655.050 254.250 ;
        RECT 670.950 253.950 673.050 257.400 ;
        RECT 692.400 255.600 693.600 257.400 ;
        RECT 697.950 255.600 700.050 255.900 ;
        RECT 692.400 254.400 700.050 255.600 ;
        RECT 697.950 253.800 700.050 254.400 ;
        RECT 724.950 253.950 727.050 257.400 ;
        RECT 734.400 255.900 735.600 262.950 ;
        RECT 742.950 260.100 745.050 262.200 ;
        RECT 766.950 261.600 769.050 262.200 ;
        RECT 787.950 261.600 790.050 262.200 ;
        RECT 811.950 261.600 814.050 262.050 ;
        RECT 766.950 260.400 786.600 261.600 ;
        RECT 766.950 260.100 769.050 260.400 ;
        RECT 733.950 253.800 736.050 255.900 ;
        RECT 247.950 251.400 285.600 252.600 ;
        RECT 286.950 252.600 289.050 253.050 ;
        RECT 301.950 252.600 304.050 253.050 ;
        RECT 286.950 251.400 304.050 252.600 ;
        RECT 247.950 250.950 250.050 251.400 ;
        RECT 286.950 250.950 289.050 251.400 ;
        RECT 301.950 250.950 304.050 251.400 ;
        RECT 310.950 252.600 313.050 253.050 ;
        RECT 325.950 252.600 328.050 253.050 ;
        RECT 310.950 251.400 328.050 252.600 ;
        RECT 310.950 250.950 313.050 251.400 ;
        RECT 325.950 250.950 328.050 251.400 ;
        RECT 331.950 252.600 334.050 253.050 ;
        RECT 349.950 252.600 352.050 253.050 ;
        RECT 331.950 251.400 352.050 252.600 ;
        RECT 331.950 250.950 334.050 251.400 ;
        RECT 349.950 250.950 352.050 251.400 ;
        RECT 370.950 252.600 373.050 253.050 ;
        RECT 376.950 252.600 379.050 253.050 ;
        RECT 400.950 252.600 403.050 253.050 ;
        RECT 370.950 251.400 403.050 252.600 ;
        RECT 370.950 250.950 373.050 251.400 ;
        RECT 376.950 250.950 379.050 251.400 ;
        RECT 400.950 250.950 403.050 251.400 ;
        RECT 409.950 252.600 412.050 253.050 ;
        RECT 418.950 252.600 421.050 253.050 ;
        RECT 409.950 251.400 421.050 252.600 ;
        RECT 409.950 250.950 412.050 251.400 ;
        RECT 418.950 250.950 421.050 251.400 ;
        RECT 427.950 252.600 430.050 253.050 ;
        RECT 457.950 252.600 460.050 253.050 ;
        RECT 427.950 251.400 460.050 252.600 ;
        RECT 427.950 250.950 430.050 251.400 ;
        RECT 457.950 250.950 460.050 251.400 ;
        RECT 493.950 252.600 496.050 253.050 ;
        RECT 502.800 252.600 504.900 253.050 ;
        RECT 493.950 251.400 504.900 252.600 ;
        RECT 493.950 250.950 496.050 251.400 ;
        RECT 502.800 250.950 504.900 251.400 ;
        RECT 505.950 250.950 508.050 253.050 ;
        RECT 520.800 250.950 522.900 253.050 ;
        RECT 523.950 252.600 526.050 253.050 ;
        RECT 532.950 252.600 535.050 253.050 ;
        RECT 523.950 251.400 535.050 252.600 ;
        RECT 523.950 250.950 526.050 251.400 ;
        RECT 532.950 250.950 535.050 251.400 ;
        RECT 574.950 252.600 577.050 253.050 ;
        RECT 580.950 252.600 583.050 253.050 ;
        RECT 610.950 252.600 613.050 253.050 ;
        RECT 574.950 251.400 613.050 252.600 ;
        RECT 574.950 250.950 577.050 251.400 ;
        RECT 580.950 250.950 583.050 251.400 ;
        RECT 610.950 250.950 613.050 251.400 ;
        RECT 619.950 252.600 622.050 253.050 ;
        RECT 658.950 252.600 661.050 253.050 ;
        RECT 667.950 252.600 670.050 253.050 ;
        RECT 619.950 251.400 670.050 252.600 ;
        RECT 619.950 250.950 622.050 251.400 ;
        RECT 658.950 250.950 661.050 251.400 ;
        RECT 667.950 250.950 670.050 251.400 ;
        RECT 676.950 252.600 679.050 253.050 ;
        RECT 715.950 252.600 718.050 253.050 ;
        RECT 676.950 251.400 718.050 252.600 ;
        RECT 676.950 250.950 679.050 251.400 ;
        RECT 715.950 250.950 718.050 251.400 ;
        RECT 7.950 249.600 10.050 250.050 ;
        RECT 58.950 249.600 61.050 250.050 ;
        RECT 7.950 248.400 61.050 249.600 ;
        RECT 7.950 247.950 10.050 248.400 ;
        RECT 58.950 247.950 61.050 248.400 ;
        RECT 64.950 249.600 67.050 250.050 ;
        RECT 118.950 249.600 121.050 250.050 ;
        RECT 64.950 248.400 121.050 249.600 ;
        RECT 64.950 247.950 67.050 248.400 ;
        RECT 118.950 247.950 121.050 248.400 ;
        RECT 148.950 249.600 151.050 250.050 ;
        RECT 154.950 249.600 157.050 250.050 ;
        RECT 148.950 248.400 157.050 249.600 ;
        RECT 148.950 247.950 151.050 248.400 ;
        RECT 154.950 247.950 157.050 248.400 ;
        RECT 169.950 249.600 172.050 250.050 ;
        RECT 184.950 249.600 187.050 250.050 ;
        RECT 193.950 249.600 196.050 250.050 ;
        RECT 169.950 248.400 196.050 249.600 ;
        RECT 169.950 247.950 172.050 248.400 ;
        RECT 184.950 247.950 187.050 248.400 ;
        RECT 193.950 247.950 196.050 248.400 ;
        RECT 244.950 249.600 247.050 250.050 ;
        RECT 253.800 249.600 255.900 250.050 ;
        RECT 244.950 248.400 255.900 249.600 ;
        RECT 244.950 247.950 247.050 248.400 ;
        RECT 253.800 247.950 255.900 248.400 ;
        RECT 256.950 249.600 259.050 250.050 ;
        RECT 271.950 249.600 274.050 250.050 ;
        RECT 256.950 248.400 274.050 249.600 ;
        RECT 256.950 247.950 259.050 248.400 ;
        RECT 271.950 247.950 274.050 248.400 ;
        RECT 280.950 249.600 283.050 250.050 ;
        RECT 379.950 249.600 382.050 250.050 ;
        RECT 397.950 249.600 400.050 250.050 ;
        RECT 280.950 248.400 288.600 249.600 ;
        RECT 280.950 247.950 283.050 248.400 ;
        RECT 10.950 246.600 13.050 247.050 ;
        RECT 55.950 246.600 58.050 247.050 ;
        RECT 10.950 245.400 58.050 246.600 ;
        RECT 10.950 244.950 13.050 245.400 ;
        RECT 55.950 244.950 58.050 245.400 ;
        RECT 196.950 246.600 199.050 247.050 ;
        RECT 208.950 246.600 211.050 247.050 ;
        RECT 196.950 245.400 211.050 246.600 ;
        RECT 196.950 244.950 199.050 245.400 ;
        RECT 208.950 244.950 211.050 245.400 ;
        RECT 268.950 246.600 271.050 247.050 ;
        RECT 283.950 246.600 286.050 247.050 ;
        RECT 268.950 245.400 286.050 246.600 ;
        RECT 287.400 246.600 288.600 248.400 ;
        RECT 379.950 248.400 400.050 249.600 ;
        RECT 379.950 247.950 382.050 248.400 ;
        RECT 397.950 247.950 400.050 248.400 ;
        RECT 406.950 249.600 409.050 250.050 ;
        RECT 415.950 249.600 418.050 250.050 ;
        RECT 451.950 249.600 454.050 250.050 ;
        RECT 493.950 249.600 496.050 249.900 ;
        RECT 406.950 248.400 496.050 249.600 ;
        RECT 406.950 247.950 409.050 248.400 ;
        RECT 415.950 247.950 418.050 248.400 ;
        RECT 451.950 247.950 454.050 248.400 ;
        RECT 493.950 247.800 496.050 248.400 ;
        RECT 550.950 249.600 553.050 250.050 ;
        RECT 565.950 249.600 568.050 250.050 ;
        RECT 550.950 248.400 568.050 249.600 ;
        RECT 550.950 247.950 553.050 248.400 ;
        RECT 565.950 247.950 568.050 248.400 ;
        RECT 724.950 249.600 727.050 250.050 ;
        RECT 743.400 249.600 744.600 260.100 ;
        RECT 785.400 258.600 786.600 260.400 ;
        RECT 787.950 260.400 814.050 261.600 ;
        RECT 787.950 260.100 790.050 260.400 ;
        RECT 785.400 257.400 789.600 258.600 ;
        RECT 788.400 255.600 789.600 257.400 ;
        RECT 806.400 255.900 807.600 260.400 ;
        RECT 811.950 259.950 814.050 260.400 ;
        RECT 829.950 261.600 832.050 262.200 ;
        RECT 838.950 261.600 841.050 262.050 ;
        RECT 829.950 260.400 841.050 261.600 ;
        RECT 829.950 260.100 832.050 260.400 ;
        RECT 838.950 259.950 841.050 260.400 ;
        RECT 860.400 256.050 861.600 263.400 ;
        RECT 904.950 263.400 916.050 264.600 ;
        RECT 904.950 262.950 907.050 263.400 ;
        RECT 913.950 262.950 916.050 263.400 ;
        RECT 943.950 262.950 946.050 265.050 ;
        RECT 874.950 261.750 877.050 262.200 ;
        RECT 886.950 261.750 889.050 262.200 ;
        RECT 874.950 260.550 889.050 261.750 ;
        RECT 874.950 260.100 877.050 260.550 ;
        RECT 886.950 260.100 889.050 260.550 ;
        RECT 892.950 258.600 895.050 262.050 ;
        RECT 898.950 260.100 901.050 262.200 ;
        RECT 925.950 260.100 928.050 262.200 ;
        RECT 890.400 258.000 895.050 258.600 ;
        RECT 890.400 257.400 894.600 258.000 ;
        RECT 799.950 255.600 802.050 255.900 ;
        RECT 788.400 254.400 802.050 255.600 ;
        RECT 799.950 253.800 802.050 254.400 ;
        RECT 805.950 253.800 808.050 255.900 ;
        RECT 817.950 255.450 820.050 255.900 ;
        RECT 832.950 255.450 835.050 255.900 ;
        RECT 817.950 254.250 835.050 255.450 ;
        RECT 817.950 253.800 820.050 254.250 ;
        RECT 832.950 253.800 835.050 254.250 ;
        RECT 859.950 253.950 862.050 256.050 ;
        RECT 751.950 252.600 754.050 253.050 ;
        RECT 763.950 252.600 766.050 253.050 ;
        RECT 751.950 251.400 766.050 252.600 ;
        RECT 751.950 250.950 754.050 251.400 ;
        RECT 763.950 250.950 766.050 251.400 ;
        RECT 856.950 252.600 859.050 253.050 ;
        RECT 865.950 252.600 868.050 253.050 ;
        RECT 856.950 251.400 868.050 252.600 ;
        RECT 856.950 250.950 859.050 251.400 ;
        RECT 865.950 250.950 868.050 251.400 ;
        RECT 880.950 252.600 883.050 253.050 ;
        RECT 890.400 252.600 891.600 257.400 ;
        RECT 892.950 255.600 895.050 256.050 ;
        RECT 899.400 255.600 900.600 260.100 ;
        RECT 910.950 258.600 913.050 258.900 ;
        RECT 926.400 258.600 927.600 260.100 ;
        RECT 931.950 259.950 934.050 262.050 ;
        RECT 910.950 257.400 927.600 258.600 ;
        RECT 910.950 256.800 913.050 257.400 ;
        RECT 932.400 256.050 933.600 259.950 ;
        RECT 944.400 258.600 945.600 262.950 ;
        RECT 946.950 261.600 951.000 262.050 ;
        RECT 946.950 259.950 951.600 261.600 ;
        RECT 944.400 258.000 948.600 258.600 ;
        RECT 944.400 257.400 949.050 258.000 ;
        RECT 892.950 254.400 900.600 255.600 ;
        RECT 928.950 255.600 931.050 255.900 ;
        RECT 931.950 255.600 934.050 256.050 ;
        RECT 940.950 255.600 943.050 255.900 ;
        RECT 928.950 254.400 943.050 255.600 ;
        RECT 892.950 253.950 895.050 254.400 ;
        RECT 928.950 253.800 931.050 254.400 ;
        RECT 931.950 253.950 934.050 254.400 ;
        RECT 940.950 253.800 943.050 254.400 ;
        RECT 946.950 253.950 949.050 257.400 ;
        RECT 880.950 251.400 891.600 252.600 ;
        RECT 916.950 252.600 919.050 253.050 ;
        RECT 925.950 252.600 928.050 253.050 ;
        RECT 916.950 251.400 928.050 252.600 ;
        RECT 880.950 250.950 883.050 251.400 ;
        RECT 916.950 250.950 919.050 251.400 ;
        RECT 925.950 250.950 928.050 251.400 ;
        RECT 724.950 248.400 744.600 249.600 ;
        RECT 847.950 249.600 850.050 250.050 ;
        RECT 859.950 249.600 862.050 250.050 ;
        RECT 847.950 248.400 862.050 249.600 ;
        RECT 724.950 247.950 727.050 248.400 ;
        RECT 847.950 247.950 850.050 248.400 ;
        RECT 859.950 247.950 862.050 248.400 ;
        RECT 877.950 249.600 880.050 250.050 ;
        RECT 886.950 249.600 889.050 250.050 ;
        RECT 895.950 249.600 898.050 250.050 ;
        RECT 877.950 248.400 898.050 249.600 ;
        RECT 877.950 247.950 880.050 248.400 ;
        RECT 886.950 247.950 889.050 248.400 ;
        RECT 895.950 247.950 898.050 248.400 ;
        RECT 910.950 249.600 913.050 250.050 ;
        RECT 928.950 249.600 931.050 250.050 ;
        RECT 910.950 248.400 931.050 249.600 ;
        RECT 910.950 247.950 913.050 248.400 ;
        RECT 928.950 247.950 931.050 248.400 ;
        RECT 943.950 249.600 946.050 250.050 ;
        RECT 950.400 249.600 951.600 259.950 ;
        RECT 943.950 248.400 951.600 249.600 ;
        RECT 943.950 247.950 946.050 248.400 ;
        RECT 349.950 246.600 352.050 247.050 ;
        RECT 287.400 245.400 352.050 246.600 ;
        RECT 268.950 244.950 271.050 245.400 ;
        RECT 283.950 244.950 286.050 245.400 ;
        RECT 349.950 244.950 352.050 245.400 ;
        RECT 373.950 246.600 376.050 247.050 ;
        RECT 388.950 246.600 391.050 247.050 ;
        RECT 373.950 245.400 391.050 246.600 ;
        RECT 373.950 244.950 376.050 245.400 ;
        RECT 388.950 244.950 391.050 245.400 ;
        RECT 553.950 246.600 556.050 247.050 ;
        RECT 838.950 246.600 841.050 247.050 ;
        RECT 871.950 246.600 874.050 247.050 ;
        RECT 886.950 246.600 889.050 246.900 ;
        RECT 892.950 246.600 895.050 247.050 ;
        RECT 553.950 245.400 609.600 246.600 ;
        RECT 553.950 244.950 556.050 245.400 ;
        RECT 28.950 243.600 31.050 244.050 ;
        RECT 40.950 243.600 43.050 244.050 ;
        RECT 28.950 242.400 43.050 243.600 ;
        RECT 28.950 241.950 31.050 242.400 ;
        RECT 40.950 241.950 43.050 242.400 ;
        RECT 64.950 243.600 67.050 244.050 ;
        RECT 124.950 243.600 127.050 244.050 ;
        RECT 64.950 242.400 127.050 243.600 ;
        RECT 64.950 241.950 67.050 242.400 ;
        RECT 124.950 241.950 127.050 242.400 ;
        RECT 172.950 243.600 175.050 244.050 ;
        RECT 199.950 243.600 202.050 244.050 ;
        RECT 205.950 243.600 208.050 244.050 ;
        RECT 172.950 242.400 208.050 243.600 ;
        RECT 172.950 241.950 175.050 242.400 ;
        RECT 199.950 241.950 202.050 242.400 ;
        RECT 205.950 241.950 208.050 242.400 ;
        RECT 232.950 243.600 235.050 244.050 ;
        RECT 256.950 243.600 259.050 244.050 ;
        RECT 232.950 242.400 259.050 243.600 ;
        RECT 232.950 241.950 235.050 242.400 ;
        RECT 256.950 241.950 259.050 242.400 ;
        RECT 262.950 243.600 265.050 244.050 ;
        RECT 277.950 243.600 280.050 244.050 ;
        RECT 262.950 242.400 280.050 243.600 ;
        RECT 262.950 241.950 265.050 242.400 ;
        RECT 277.950 241.950 280.050 242.400 ;
        RECT 298.950 243.600 301.050 244.050 ;
        RECT 310.950 243.600 313.050 244.050 ;
        RECT 298.950 242.400 313.050 243.600 ;
        RECT 298.950 241.950 301.050 242.400 ;
        RECT 310.950 241.950 313.050 242.400 ;
        RECT 421.950 243.600 424.050 244.050 ;
        RECT 478.950 243.600 481.050 244.050 ;
        RECT 496.950 243.600 499.050 244.050 ;
        RECT 595.950 243.600 598.050 244.050 ;
        RECT 421.950 242.400 499.050 243.600 ;
        RECT 421.950 241.950 424.050 242.400 ;
        RECT 478.950 241.950 481.050 242.400 ;
        RECT 496.950 241.950 499.050 242.400 ;
        RECT 515.400 242.400 598.050 243.600 ;
        RECT 608.400 243.600 609.600 245.400 ;
        RECT 838.950 245.400 895.050 246.600 ;
        RECT 838.950 244.950 841.050 245.400 ;
        RECT 871.950 244.950 874.050 245.400 ;
        RECT 886.950 244.800 889.050 245.400 ;
        RECT 892.950 244.950 895.050 245.400 ;
        RECT 901.950 246.600 904.050 246.900 ;
        RECT 934.950 246.600 937.050 247.050 ;
        RECT 901.950 245.400 937.050 246.600 ;
        RECT 901.950 244.800 904.050 245.400 ;
        RECT 934.950 244.950 937.050 245.400 ;
        RECT 676.950 243.600 679.050 244.050 ;
        RECT 608.400 242.400 679.050 243.600 ;
        RECT 4.950 240.600 7.050 241.050 ;
        RECT 70.950 240.600 73.050 241.050 ;
        RECT 175.950 240.600 178.050 241.050 ;
        RECT 4.950 239.400 33.600 240.600 ;
        RECT 4.950 238.950 7.050 239.400 ;
        RECT 32.400 238.050 33.600 239.400 ;
        RECT 70.950 239.400 178.050 240.600 ;
        RECT 70.950 238.950 73.050 239.400 ;
        RECT 175.950 238.950 178.050 239.400 ;
        RECT 181.950 240.600 184.050 241.050 ;
        RECT 217.950 240.600 220.050 241.050 ;
        RECT 181.950 239.400 220.050 240.600 ;
        RECT 181.950 238.950 184.050 239.400 ;
        RECT 217.950 238.950 220.050 239.400 ;
        RECT 229.950 240.600 232.050 241.050 ;
        RECT 295.950 240.600 298.050 241.050 ;
        RECT 229.950 239.400 298.050 240.600 ;
        RECT 229.950 238.950 232.050 239.400 ;
        RECT 295.950 238.950 298.050 239.400 ;
        RECT 301.950 240.600 304.050 241.050 ;
        RECT 334.950 240.600 337.050 241.050 ;
        RECT 301.950 239.400 337.050 240.600 ;
        RECT 301.950 238.950 304.050 239.400 ;
        RECT 334.950 238.950 337.050 239.400 ;
        RECT 343.950 240.600 346.050 241.050 ;
        RECT 379.950 240.600 382.050 241.050 ;
        RECT 515.400 240.600 516.600 242.400 ;
        RECT 595.950 241.950 598.050 242.400 ;
        RECT 676.950 241.950 679.050 242.400 ;
        RECT 763.950 243.600 766.050 244.050 ;
        RECT 784.950 243.600 787.050 244.050 ;
        RECT 763.950 242.400 787.050 243.600 ;
        RECT 763.950 241.950 766.050 242.400 ;
        RECT 784.950 241.950 787.050 242.400 ;
        RECT 343.950 239.400 382.050 240.600 ;
        RECT 343.950 238.950 346.050 239.400 ;
        RECT 379.950 238.950 382.050 239.400 ;
        RECT 443.400 239.400 516.600 240.600 ;
        RECT 517.950 240.600 520.050 241.050 ;
        RECT 616.950 240.600 619.050 241.050 ;
        RECT 517.950 239.400 619.050 240.600 ;
        RECT 32.400 237.600 37.050 238.050 ;
        RECT 88.950 237.600 91.050 238.050 ;
        RECT 32.400 236.400 91.050 237.600 ;
        RECT 33.000 235.950 37.050 236.400 ;
        RECT 88.950 235.950 91.050 236.400 ;
        RECT 109.950 237.600 112.050 238.050 ;
        RECT 139.950 237.600 142.050 238.050 ;
        RECT 286.950 237.600 289.050 238.050 ;
        RECT 355.950 237.600 358.050 238.050 ;
        RECT 443.400 237.600 444.600 239.400 ;
        RECT 517.950 238.950 520.050 239.400 ;
        RECT 616.950 238.950 619.050 239.400 ;
        RECT 625.950 240.600 628.050 241.050 ;
        RECT 745.950 240.600 748.050 241.050 ;
        RECT 625.950 239.400 748.050 240.600 ;
        RECT 625.950 238.950 628.050 239.400 ;
        RECT 745.950 238.950 748.050 239.400 ;
        RECT 874.950 240.600 877.050 241.050 ;
        RECT 898.950 240.600 901.050 241.050 ;
        RECT 874.950 239.400 901.050 240.600 ;
        RECT 874.950 238.950 877.050 239.400 ;
        RECT 898.950 238.950 901.050 239.400 ;
        RECT 109.950 236.400 444.600 237.600 ;
        RECT 445.950 237.600 448.050 238.050 ;
        RECT 475.950 237.600 478.050 238.050 ;
        RECT 445.950 236.400 478.050 237.600 ;
        RECT 109.950 235.950 112.050 236.400 ;
        RECT 139.950 235.950 142.050 236.400 ;
        RECT 286.950 235.950 289.050 236.400 ;
        RECT 355.950 235.950 358.050 236.400 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 475.950 235.950 478.050 236.400 ;
        RECT 511.950 237.600 514.050 238.050 ;
        RECT 757.950 237.600 760.050 238.050 ;
        RECT 778.950 237.600 781.050 238.050 ;
        RECT 511.950 236.400 781.050 237.600 ;
        RECT 511.950 235.950 514.050 236.400 ;
        RECT 757.950 235.950 760.050 236.400 ;
        RECT 778.950 235.950 781.050 236.400 ;
        RECT 823.950 237.600 826.050 238.050 ;
        RECT 850.950 237.600 853.050 238.050 ;
        RECT 823.950 236.400 853.050 237.600 ;
        RECT 823.950 235.950 826.050 236.400 ;
        RECT 850.950 235.950 853.050 236.400 ;
        RECT 904.950 237.600 907.050 238.050 ;
        RECT 910.950 237.600 913.050 238.050 ;
        RECT 934.950 237.600 937.050 238.050 ;
        RECT 904.950 236.400 937.050 237.600 ;
        RECT 904.950 235.950 907.050 236.400 ;
        RECT 910.950 235.950 913.050 236.400 ;
        RECT 934.950 235.950 937.050 236.400 ;
        RECT 193.950 234.600 196.050 235.050 ;
        RECT 214.950 234.600 217.050 235.050 ;
        RECT 226.950 234.600 229.050 235.050 ;
        RECT 193.950 233.400 229.050 234.600 ;
        RECT 193.950 232.950 196.050 233.400 ;
        RECT 214.950 232.950 217.050 233.400 ;
        RECT 226.950 232.950 229.050 233.400 ;
        RECT 259.950 234.600 262.050 235.050 ;
        RECT 292.950 234.600 295.050 235.050 ;
        RECT 259.950 233.400 295.050 234.600 ;
        RECT 259.950 232.950 262.050 233.400 ;
        RECT 292.950 232.950 295.050 233.400 ;
        RECT 298.950 234.600 301.050 235.050 ;
        RECT 322.950 234.600 325.050 235.050 ;
        RECT 298.950 233.400 325.050 234.600 ;
        RECT 298.950 232.950 301.050 233.400 ;
        RECT 322.950 232.950 325.050 233.400 ;
        RECT 337.950 234.600 340.050 235.050 ;
        RECT 358.800 234.600 360.900 235.050 ;
        RECT 337.950 233.400 360.900 234.600 ;
        RECT 337.950 232.950 340.050 233.400 ;
        RECT 358.800 232.950 360.900 233.400 ;
        RECT 361.950 234.600 364.050 235.050 ;
        RECT 472.950 234.600 475.050 235.050 ;
        RECT 361.950 233.400 475.050 234.600 ;
        RECT 361.950 232.950 364.050 233.400 ;
        RECT 472.950 232.950 475.050 233.400 ;
        RECT 619.950 234.600 622.050 235.050 ;
        RECT 643.950 234.600 646.050 235.050 ;
        RECT 619.950 233.400 646.050 234.600 ;
        RECT 619.950 232.950 622.050 233.400 ;
        RECT 643.950 232.950 646.050 233.400 ;
        RECT 874.950 234.600 877.050 235.050 ;
        RECT 883.950 234.600 886.050 235.050 ;
        RECT 874.950 233.400 886.050 234.600 ;
        RECT 874.950 232.950 877.050 233.400 ;
        RECT 883.950 232.950 886.050 233.400 ;
        RECT 28.950 231.600 31.050 232.050 ;
        RECT 94.950 231.600 97.050 232.050 ;
        RECT 100.950 231.600 103.050 232.050 ;
        RECT 28.950 230.400 103.050 231.600 ;
        RECT 28.950 229.950 31.050 230.400 ;
        RECT 94.950 229.950 97.050 230.400 ;
        RECT 100.950 229.950 103.050 230.400 ;
        RECT 160.950 231.600 163.050 232.050 ;
        RECT 190.950 231.600 193.050 232.050 ;
        RECT 160.950 230.400 193.050 231.600 ;
        RECT 160.950 229.950 163.050 230.400 ;
        RECT 190.950 229.950 193.050 230.400 ;
        RECT 196.950 231.600 199.050 232.050 ;
        RECT 307.950 231.600 310.050 232.050 ;
        RECT 196.950 230.400 310.050 231.600 ;
        RECT 196.950 229.950 199.050 230.400 ;
        RECT 307.950 229.950 310.050 230.400 ;
        RECT 379.950 231.600 382.050 232.050 ;
        RECT 391.950 231.600 394.050 232.050 ;
        RECT 379.950 230.400 394.050 231.600 ;
        RECT 379.950 229.950 382.050 230.400 ;
        RECT 391.950 229.950 394.050 230.400 ;
        RECT 403.950 231.600 406.050 232.050 ;
        RECT 433.950 231.600 436.050 232.050 ;
        RECT 442.950 231.600 445.050 232.050 ;
        RECT 475.950 231.600 478.050 232.050 ;
        RECT 403.950 230.400 432.600 231.600 ;
        RECT 403.950 229.950 406.050 230.400 ;
        RECT 214.950 228.600 217.050 229.050 ;
        RECT 268.950 228.600 271.050 229.050 ;
        RECT 331.950 228.600 334.050 229.050 ;
        RECT 214.950 227.400 271.050 228.600 ;
        RECT 214.950 226.950 217.050 227.400 ;
        RECT 268.950 226.950 271.050 227.400 ;
        RECT 317.400 227.400 334.050 228.600 ;
        RECT 317.400 226.050 318.600 227.400 ;
        RECT 331.950 226.950 334.050 227.400 ;
        RECT 337.950 228.600 340.050 229.050 ;
        RECT 364.950 228.600 367.050 229.050 ;
        RECT 337.950 227.400 367.050 228.600 ;
        RECT 337.950 226.950 340.050 227.400 ;
        RECT 364.950 226.950 367.050 227.400 ;
        RECT 391.950 228.600 394.050 228.900 ;
        RECT 427.950 228.600 430.050 229.050 ;
        RECT 391.950 227.400 430.050 228.600 ;
        RECT 431.400 228.600 432.600 230.400 ;
        RECT 433.950 230.400 478.050 231.600 ;
        RECT 433.950 229.950 436.050 230.400 ;
        RECT 442.950 229.950 445.050 230.400 ;
        RECT 475.950 229.950 478.050 230.400 ;
        RECT 499.950 231.600 502.050 232.050 ;
        RECT 517.950 231.600 520.050 232.050 ;
        RECT 499.950 230.400 520.050 231.600 ;
        RECT 499.950 229.950 502.050 230.400 ;
        RECT 517.950 229.950 520.050 230.400 ;
        RECT 583.950 231.600 586.050 232.050 ;
        RECT 595.950 231.600 598.050 232.050 ;
        RECT 610.950 231.600 613.050 232.050 ;
        RECT 583.950 230.400 613.050 231.600 ;
        RECT 583.950 229.950 586.050 230.400 ;
        RECT 595.950 229.950 598.050 230.400 ;
        RECT 610.950 229.950 613.050 230.400 ;
        RECT 898.950 231.600 901.050 232.050 ;
        RECT 916.950 231.600 919.050 232.050 ;
        RECT 943.950 231.600 946.050 232.050 ;
        RECT 898.950 230.400 946.050 231.600 ;
        RECT 898.950 229.950 901.050 230.400 ;
        RECT 916.950 229.950 919.050 230.400 ;
        RECT 943.950 229.950 946.050 230.400 ;
        RECT 445.950 228.600 448.050 229.050 ;
        RECT 431.400 227.400 448.050 228.600 ;
        RECT 391.950 226.800 394.050 227.400 ;
        RECT 427.950 226.950 430.050 227.400 ;
        RECT 445.950 226.950 448.050 227.400 ;
        RECT 481.950 228.600 484.050 229.050 ;
        RECT 529.950 228.600 532.050 229.050 ;
        RECT 535.950 228.600 538.050 229.050 ;
        RECT 481.950 227.400 538.050 228.600 ;
        RECT 481.950 226.950 484.050 227.400 ;
        RECT 529.950 226.950 532.050 227.400 ;
        RECT 535.950 226.950 538.050 227.400 ;
        RECT 883.950 228.600 886.050 229.050 ;
        RECT 895.950 228.600 898.050 229.050 ;
        RECT 883.950 227.400 898.050 228.600 ;
        RECT 883.950 226.950 886.050 227.400 ;
        RECT 895.950 226.950 898.050 227.400 ;
        RECT 49.950 225.600 52.050 226.050 ;
        RECT 76.950 225.600 79.050 226.050 ;
        RECT 49.950 224.400 79.050 225.600 ;
        RECT 49.950 223.950 52.050 224.400 ;
        RECT 76.950 223.950 79.050 224.400 ;
        RECT 211.950 225.600 214.050 226.050 ;
        RECT 250.950 225.600 253.050 226.050 ;
        RECT 211.950 224.400 253.050 225.600 ;
        RECT 211.950 223.950 214.050 224.400 ;
        RECT 250.950 223.950 253.050 224.400 ;
        RECT 256.950 225.600 259.050 226.050 ;
        RECT 265.950 225.600 268.050 226.050 ;
        RECT 256.950 224.400 268.050 225.600 ;
        RECT 256.950 223.950 259.050 224.400 ;
        RECT 265.950 223.950 268.050 224.400 ;
        RECT 271.950 225.600 274.050 226.050 ;
        RECT 292.950 225.600 295.050 226.050 ;
        RECT 316.950 225.600 319.050 226.050 ;
        RECT 271.950 224.400 291.600 225.600 ;
        RECT 271.950 223.950 274.050 224.400 ;
        RECT 52.950 222.600 55.050 223.050 ;
        RECT 61.950 222.600 64.050 223.050 ;
        RECT 52.950 221.400 64.050 222.600 ;
        RECT 52.950 220.950 55.050 221.400 ;
        RECT 61.950 220.950 64.050 221.400 ;
        RECT 88.950 222.600 91.050 223.050 ;
        RECT 109.950 222.600 112.050 223.050 ;
        RECT 88.950 221.400 112.050 222.600 ;
        RECT 88.950 220.950 91.050 221.400 ;
        RECT 109.950 220.950 112.050 221.400 ;
        RECT 166.950 222.600 169.050 223.050 ;
        RECT 247.950 222.600 250.050 223.050 ;
        RECT 166.950 221.400 250.050 222.600 ;
        RECT 290.400 222.600 291.600 224.400 ;
        RECT 292.950 224.400 319.050 225.600 ;
        RECT 292.950 223.950 295.050 224.400 ;
        RECT 316.950 223.950 319.050 224.400 ;
        RECT 322.950 225.600 325.050 226.050 ;
        RECT 361.950 225.600 364.050 226.050 ;
        RECT 322.950 224.400 364.050 225.600 ;
        RECT 322.950 223.950 325.050 224.400 ;
        RECT 361.950 223.950 364.050 224.400 ;
        RECT 505.950 225.600 508.050 226.050 ;
        RECT 562.950 225.600 565.050 226.050 ;
        RECT 604.950 225.600 607.050 226.050 ;
        RECT 640.950 225.600 643.050 226.050 ;
        RECT 505.950 224.400 643.050 225.600 ;
        RECT 505.950 223.950 508.050 224.400 ;
        RECT 562.950 223.950 565.050 224.400 ;
        RECT 604.950 223.950 607.050 224.400 ;
        RECT 640.950 223.950 643.050 224.400 ;
        RECT 664.950 225.600 667.050 226.050 ;
        RECT 682.950 225.600 685.050 226.050 ;
        RECT 709.950 225.600 712.050 226.050 ;
        RECT 664.950 224.400 712.050 225.600 ;
        RECT 664.950 223.950 667.050 224.400 ;
        RECT 682.950 223.950 685.050 224.400 ;
        RECT 709.950 223.950 712.050 224.400 ;
        RECT 772.950 225.600 775.050 226.050 ;
        RECT 784.950 225.600 787.050 226.050 ;
        RECT 793.950 225.600 796.050 226.050 ;
        RECT 772.950 224.400 796.050 225.600 ;
        RECT 772.950 223.950 775.050 224.400 ;
        RECT 784.950 223.950 787.050 224.400 ;
        RECT 793.950 223.950 796.050 224.400 ;
        RECT 898.950 225.600 901.050 226.050 ;
        RECT 907.950 225.600 910.050 226.050 ;
        RECT 898.950 224.400 910.050 225.600 ;
        RECT 898.950 223.950 901.050 224.400 ;
        RECT 907.950 223.950 910.050 224.400 ;
        RECT 304.950 222.600 307.050 223.050 ;
        RECT 290.400 221.400 307.050 222.600 ;
        RECT 166.950 220.950 169.050 221.400 ;
        RECT 247.950 220.950 250.050 221.400 ;
        RECT 304.950 220.950 307.050 221.400 ;
        RECT 325.950 222.600 328.050 223.050 ;
        RECT 352.950 222.600 355.050 223.050 ;
        RECT 325.950 221.400 355.050 222.600 ;
        RECT 325.950 220.950 328.050 221.400 ;
        RECT 352.950 220.950 355.050 221.400 ;
        RECT 358.950 222.600 361.050 223.050 ;
        RECT 400.950 222.600 403.050 223.050 ;
        RECT 358.950 221.400 403.050 222.600 ;
        RECT 358.950 220.950 361.050 221.400 ;
        RECT 400.950 220.950 403.050 221.400 ;
        RECT 427.950 222.600 430.050 223.050 ;
        RECT 439.950 222.600 442.050 223.050 ;
        RECT 448.950 222.600 451.050 223.050 ;
        RECT 499.950 222.600 502.050 223.050 ;
        RECT 427.950 221.400 451.050 222.600 ;
        RECT 427.950 220.950 430.050 221.400 ;
        RECT 439.950 220.950 442.050 221.400 ;
        RECT 448.950 220.950 451.050 221.400 ;
        RECT 461.400 221.400 502.050 222.600 ;
        RECT 121.950 219.600 124.050 220.050 ;
        RECT 154.950 219.600 157.050 220.050 ;
        RECT 121.950 218.400 157.050 219.600 ;
        RECT 121.950 217.950 124.050 218.400 ;
        RECT 154.950 217.950 157.050 218.400 ;
        RECT 229.950 219.600 232.050 220.050 ;
        RECT 235.950 219.600 238.050 220.050 ;
        RECT 229.950 218.400 238.050 219.600 ;
        RECT 229.950 217.950 232.050 218.400 ;
        RECT 235.950 217.950 238.050 218.400 ;
        RECT 265.950 219.600 268.050 219.900 ;
        RECT 274.950 219.600 277.050 220.050 ;
        RECT 265.950 218.400 277.050 219.600 ;
        RECT 265.950 217.800 268.050 218.400 ;
        RECT 274.950 217.950 277.050 218.400 ;
        RECT 313.950 219.600 316.050 220.050 ;
        RECT 322.950 219.600 325.050 220.050 ;
        RECT 313.950 218.400 325.050 219.600 ;
        RECT 313.950 217.950 316.050 218.400 ;
        RECT 322.950 217.950 325.050 218.400 ;
        RECT 382.950 219.600 385.050 220.050 ;
        RECT 427.950 219.600 430.050 219.900 ;
        RECT 461.400 219.600 462.600 221.400 ;
        RECT 499.950 220.950 502.050 221.400 ;
        RECT 505.950 222.600 508.050 222.900 ;
        RECT 511.950 222.600 514.050 223.050 ;
        RECT 541.950 222.600 544.050 223.050 ;
        RECT 505.950 221.400 544.050 222.600 ;
        RECT 505.950 220.800 508.050 221.400 ;
        RECT 511.950 220.950 514.050 221.400 ;
        RECT 541.950 220.950 544.050 221.400 ;
        RECT 577.950 222.600 580.050 223.050 ;
        RECT 592.950 222.600 595.050 223.050 ;
        RECT 577.950 221.400 595.050 222.600 ;
        RECT 577.950 220.950 580.050 221.400 ;
        RECT 592.950 220.950 595.050 221.400 ;
        RECT 799.950 222.600 802.050 223.050 ;
        RECT 841.950 222.600 844.050 223.050 ;
        RECT 868.950 222.600 871.050 223.050 ;
        RECT 799.950 221.400 871.050 222.600 ;
        RECT 799.950 220.950 802.050 221.400 ;
        RECT 841.950 220.950 844.050 221.400 ;
        RECT 868.950 220.950 871.050 221.400 ;
        RECT 937.950 222.600 940.050 223.050 ;
        RECT 943.950 222.600 946.050 223.050 ;
        RECT 937.950 221.400 946.050 222.600 ;
        RECT 937.950 220.950 940.050 221.400 ;
        RECT 943.950 220.950 946.050 221.400 ;
        RECT 382.950 218.400 399.600 219.600 ;
        RECT 382.950 217.950 385.050 218.400 ;
        RECT 34.950 216.600 37.050 217.200 ;
        RECT 55.950 216.600 58.050 217.200 ;
        RECT 34.950 215.400 58.050 216.600 ;
        RECT 34.950 215.100 37.050 215.400 ;
        RECT 55.950 215.100 58.050 215.400 ;
        RECT 64.950 216.600 69.000 217.050 ;
        RECT 76.950 216.750 79.050 217.200 ;
        RECT 82.950 216.750 85.050 217.200 ;
        RECT 64.950 214.950 69.600 216.600 ;
        RECT 76.950 215.550 85.050 216.750 ;
        RECT 76.950 215.100 79.050 215.550 ;
        RECT 82.950 215.100 85.050 215.550 ;
        RECT 94.950 216.600 97.050 217.200 ;
        RECT 115.950 216.600 118.050 217.200 ;
        RECT 94.950 215.400 118.050 216.600 ;
        RECT 94.950 215.100 97.050 215.400 ;
        RECT 115.950 215.100 118.050 215.400 ;
        RECT 124.950 216.750 127.050 217.200 ;
        RECT 130.950 216.750 133.050 217.200 ;
        RECT 124.950 215.550 133.050 216.750 ;
        RECT 124.950 215.100 127.050 215.550 ;
        RECT 130.950 215.100 133.050 215.550 ;
        RECT 136.950 216.600 139.050 217.200 ;
        RECT 145.950 216.600 148.050 217.050 ;
        RECT 136.950 215.400 148.050 216.600 ;
        RECT 136.950 215.100 139.050 215.400 ;
        RECT 145.950 214.950 148.050 215.400 ;
        RECT 220.950 215.100 223.050 217.200 ;
        RECT 13.950 210.600 16.050 210.900 ;
        RECT 31.950 210.600 34.050 210.900 ;
        RECT 40.950 210.600 43.050 211.050 ;
        RECT 68.400 210.900 69.600 214.950 ;
        RECT 13.950 209.400 43.050 210.600 ;
        RECT 13.950 208.800 16.050 209.400 ;
        RECT 31.950 208.800 34.050 209.400 ;
        RECT 40.950 208.950 43.050 209.400 ;
        RECT 67.950 208.800 70.050 210.900 ;
        RECT 82.950 210.600 85.050 211.050 ;
        RECT 91.950 210.600 94.050 210.900 ;
        RECT 82.950 209.400 94.050 210.600 ;
        RECT 82.950 208.950 85.050 209.400 ;
        RECT 91.950 208.800 94.050 209.400 ;
        RECT 139.950 210.600 142.050 210.900 ;
        RECT 148.950 210.600 151.050 211.050 ;
        RECT 139.950 209.400 151.050 210.600 ;
        RECT 139.950 208.800 142.050 209.400 ;
        RECT 148.950 208.950 151.050 209.400 ;
        RECT 193.950 210.600 196.050 210.900 ;
        RECT 217.950 210.600 220.050 210.900 ;
        RECT 193.950 209.400 220.050 210.600 ;
        RECT 193.950 208.800 196.050 209.400 ;
        RECT 217.950 208.800 220.050 209.400 ;
        RECT 221.400 208.050 222.600 215.100 ;
        RECT 226.950 214.950 229.050 217.050 ;
        RECT 238.950 216.600 241.050 217.200 ;
        RECT 238.950 215.400 255.600 216.600 ;
        RECT 238.950 215.100 241.050 215.400 ;
        RECT 227.400 210.600 228.600 214.950 ;
        RECT 254.400 210.900 255.600 215.400 ;
        RECT 262.950 214.950 265.050 217.050 ;
        RECT 268.950 214.950 271.050 217.050 ;
        RECT 292.950 215.100 295.050 217.200 ;
        RECT 325.950 216.600 328.050 217.200 ;
        RECT 337.950 216.600 340.050 217.200 ;
        RECT 325.950 215.400 340.050 216.600 ;
        RECT 325.950 215.100 328.050 215.400 ;
        RECT 337.950 215.100 340.050 215.400 ;
        RECT 352.950 216.600 355.050 217.050 ;
        RECT 390.000 216.600 394.050 217.050 ;
        RECT 352.950 215.400 394.050 216.600 ;
        RECT 235.950 210.600 238.050 210.900 ;
        RECT 227.400 209.400 238.050 210.600 ;
        RECT 235.950 208.800 238.050 209.400 ;
        RECT 253.950 208.800 256.050 210.900 ;
        RECT 100.950 207.600 103.050 208.050 ;
        RECT 169.950 207.600 172.050 208.050 ;
        RECT 100.950 206.400 172.050 207.600 ;
        RECT 221.400 206.400 226.050 208.050 ;
        RECT 100.950 205.950 103.050 206.400 ;
        RECT 169.950 205.950 172.050 206.400 ;
        RECT 222.000 205.950 226.050 206.400 ;
        RECT 256.950 207.600 259.050 208.050 ;
        RECT 263.400 207.600 264.600 214.950 ;
        RECT 269.400 210.600 270.600 214.950 ;
        RECT 293.400 213.600 294.600 215.100 ;
        RECT 352.950 214.950 355.050 215.400 ;
        RECT 389.400 214.950 394.050 215.400 ;
        RECT 290.400 213.000 294.600 213.600 ;
        RECT 289.950 212.400 294.600 213.000 ;
        RECT 274.950 210.600 277.050 210.900 ;
        RECT 269.400 209.400 277.050 210.600 ;
        RECT 274.950 208.800 277.050 209.400 ;
        RECT 289.950 208.950 292.050 212.400 ;
        RECT 301.950 210.600 304.050 210.900 ;
        RECT 313.950 210.600 316.050 214.050 ;
        RECT 322.950 210.600 325.050 210.900 ;
        RECT 293.400 210.000 316.050 210.600 ;
        RECT 292.950 209.400 315.600 210.000 ;
        RECT 320.400 209.400 325.050 210.600 ;
        RECT 256.950 206.400 264.600 207.600 ;
        RECT 256.950 205.950 259.050 206.400 ;
        RECT 292.950 205.950 295.050 209.400 ;
        RECT 301.950 208.800 304.050 209.400 ;
        RECT 310.950 207.600 313.050 208.050 ;
        RECT 320.400 207.600 321.600 209.400 ;
        RECT 322.950 208.800 325.050 209.400 ;
        RECT 340.950 210.600 343.050 210.900 ;
        RECT 346.950 210.600 349.050 211.050 ;
        RECT 340.950 209.400 349.050 210.600 ;
        RECT 340.950 208.800 343.050 209.400 ;
        RECT 346.950 208.950 349.050 209.400 ;
        RECT 352.950 210.600 355.050 211.050 ;
        RECT 370.950 210.600 373.050 211.050 ;
        RECT 389.400 210.900 390.600 214.950 ;
        RECT 398.400 213.600 399.600 218.400 ;
        RECT 427.950 218.400 462.600 219.600 ;
        RECT 463.950 219.600 466.050 220.050 ;
        RECT 469.800 219.600 471.900 220.050 ;
        RECT 463.950 218.400 471.900 219.600 ;
        RECT 427.950 217.800 430.050 218.400 ;
        RECT 463.950 217.950 466.050 218.400 ;
        RECT 469.800 217.950 471.900 218.400 ;
        RECT 472.950 219.600 475.050 220.050 ;
        RECT 634.950 219.600 637.050 220.050 ;
        RECT 646.950 219.600 649.050 220.050 ;
        RECT 472.950 218.400 492.600 219.600 ;
        RECT 472.950 217.950 475.050 218.400 ;
        RECT 433.950 216.600 436.050 217.200 ;
        RECT 454.950 216.600 457.050 217.200 ;
        RECT 466.950 216.600 469.050 217.050 ;
        RECT 433.950 215.400 444.600 216.600 ;
        RECT 433.950 215.100 436.050 215.400 ;
        RECT 398.400 212.400 408.600 213.600 ;
        RECT 352.950 209.400 373.050 210.600 ;
        RECT 352.950 208.950 355.050 209.400 ;
        RECT 370.950 208.950 373.050 209.400 ;
        RECT 388.950 208.800 391.050 210.900 ;
        RECT 407.400 210.600 408.600 212.400 ;
        RECT 409.950 210.600 412.050 210.900 ;
        RECT 407.400 209.400 412.050 210.600 ;
        RECT 409.950 208.800 412.050 209.400 ;
        RECT 418.950 210.600 421.050 211.050 ;
        RECT 424.950 210.600 427.050 211.050 ;
        RECT 418.950 209.400 427.050 210.600 ;
        RECT 443.400 210.600 444.600 215.400 ;
        RECT 454.950 215.400 469.050 216.600 ;
        RECT 454.950 215.100 457.050 215.400 ;
        RECT 466.950 214.950 469.050 215.400 ;
        RECT 475.950 216.600 478.050 217.200 ;
        RECT 487.950 216.600 490.050 217.200 ;
        RECT 475.950 215.400 490.050 216.600 ;
        RECT 491.400 216.600 492.600 218.400 ;
        RECT 634.950 218.400 649.050 219.600 ;
        RECT 634.950 217.950 637.050 218.400 ;
        RECT 646.950 217.950 649.050 218.400 ;
        RECT 691.950 219.600 694.050 220.050 ;
        RECT 703.950 219.600 706.050 220.050 ;
        RECT 691.950 218.400 706.050 219.600 ;
        RECT 691.950 217.950 694.050 218.400 ;
        RECT 703.950 217.950 706.050 218.400 ;
        RECT 739.950 219.600 742.050 220.050 ;
        RECT 772.950 219.600 775.050 220.050 ;
        RECT 739.950 218.400 775.050 219.600 ;
        RECT 739.950 217.950 742.050 218.400 ;
        RECT 772.950 217.950 775.050 218.400 ;
        RECT 505.950 216.600 508.050 217.050 ;
        RECT 491.400 215.400 508.050 216.600 ;
        RECT 475.950 215.100 478.050 215.400 ;
        RECT 487.950 215.100 490.050 215.400 ;
        RECT 505.950 214.950 508.050 215.400 ;
        RECT 514.800 216.000 516.900 217.050 ;
        RECT 517.950 216.750 520.050 217.200 ;
        RECT 535.950 216.750 538.050 217.200 ;
        RECT 514.800 214.950 517.050 216.000 ;
        RECT 517.950 215.550 538.050 216.750 ;
        RECT 517.950 215.100 520.050 215.550 ;
        RECT 535.950 215.100 538.050 215.550 ;
        RECT 553.950 216.600 556.050 217.200 ;
        RECT 559.950 216.600 562.050 217.050 ;
        RECT 553.950 215.400 562.050 216.600 ;
        RECT 553.950 215.100 556.050 215.400 ;
        RECT 559.950 214.950 562.050 215.400 ;
        RECT 568.950 216.600 571.050 217.200 ;
        RECT 589.950 216.600 592.050 217.200 ;
        RECT 598.950 216.600 601.050 217.050 ;
        RECT 568.950 215.400 576.600 216.600 ;
        RECT 568.950 215.100 571.050 215.400 ;
        RECT 467.400 211.050 468.600 214.950 ;
        RECT 514.950 213.600 517.050 214.950 ;
        RECT 509.400 213.000 517.050 213.600 ;
        RECT 509.400 212.400 516.450 213.000 ;
        RECT 451.950 210.600 454.050 210.900 ;
        RECT 443.400 209.400 454.050 210.600 ;
        RECT 418.950 208.950 421.050 209.400 ;
        RECT 424.950 208.950 427.050 209.400 ;
        RECT 451.950 208.800 454.050 209.400 ;
        RECT 466.950 208.950 469.050 211.050 ;
        RECT 509.400 210.900 510.600 212.400 ;
        RECT 481.950 210.450 484.050 210.900 ;
        RECT 496.950 210.450 499.050 210.900 ;
        RECT 481.950 209.250 499.050 210.450 ;
        RECT 481.950 208.800 484.050 209.250 ;
        RECT 496.950 208.800 499.050 209.250 ;
        RECT 508.950 208.800 511.050 210.900 ;
        RECT 523.950 210.450 526.050 210.900 ;
        RECT 550.950 210.450 553.050 210.900 ;
        RECT 523.950 209.250 553.050 210.450 ;
        RECT 575.400 210.600 576.600 215.400 ;
        RECT 589.950 215.400 601.050 216.600 ;
        RECT 589.950 215.100 592.050 215.400 ;
        RECT 598.950 214.950 601.050 215.400 ;
        RECT 604.950 215.100 607.050 217.200 ;
        RECT 622.950 216.750 625.050 217.200 ;
        RECT 628.950 216.750 631.050 217.200 ;
        RECT 622.950 215.550 631.050 216.750 ;
        RECT 622.950 215.100 625.050 215.550 ;
        RECT 628.950 215.100 631.050 215.550 ;
        RECT 649.950 216.600 652.050 217.200 ;
        RECT 658.950 216.600 661.050 217.050 ;
        RECT 649.950 215.400 661.050 216.600 ;
        RECT 649.950 215.100 652.050 215.400 ;
        RECT 605.400 210.600 606.600 215.100 ;
        RECT 623.400 213.600 624.600 215.100 ;
        RECT 658.950 214.950 661.050 215.400 ;
        RECT 664.950 215.100 667.050 217.200 ;
        RECT 679.950 216.750 682.050 217.200 ;
        RECT 685.950 216.750 688.050 217.200 ;
        RECT 679.950 216.600 688.050 216.750 ;
        RECT 697.950 216.600 700.050 217.050 ;
        RECT 679.950 215.550 700.050 216.600 ;
        RECT 679.950 215.100 682.050 215.550 ;
        RECT 685.950 215.400 700.050 215.550 ;
        RECT 685.950 215.100 688.050 215.400 ;
        RECT 665.400 213.600 666.600 215.100 ;
        RECT 697.950 214.950 700.050 215.400 ;
        RECT 727.950 216.750 730.050 217.200 ;
        RECT 736.950 216.750 739.050 217.200 ;
        RECT 727.950 216.600 739.050 216.750 ;
        RECT 754.950 216.600 757.050 217.200 ;
        RECT 727.950 215.550 757.050 216.600 ;
        RECT 727.950 215.100 730.050 215.550 ;
        RECT 736.950 215.400 757.050 215.550 ;
        RECT 736.950 215.100 739.050 215.400 ;
        RECT 754.950 215.100 757.050 215.400 ;
        RECT 778.950 216.600 781.050 217.200 ;
        RECT 799.950 216.600 802.050 217.200 ;
        RECT 778.950 215.400 802.050 216.600 ;
        RECT 778.950 215.100 781.050 215.400 ;
        RECT 799.950 215.100 802.050 215.400 ;
        RECT 805.950 216.750 808.050 217.200 ;
        RECT 814.950 216.750 817.050 217.200 ;
        RECT 805.950 215.550 817.050 216.750 ;
        RECT 805.950 215.100 808.050 215.550 ;
        RECT 814.950 215.100 817.050 215.550 ;
        RECT 847.950 216.600 850.050 217.200 ;
        RECT 862.950 216.600 865.050 217.200 ;
        RECT 847.950 215.400 865.050 216.600 ;
        RECT 871.950 216.600 874.050 220.050 ;
        RECT 889.950 219.600 892.050 220.050 ;
        RECT 901.950 219.600 904.050 220.050 ;
        RECT 889.950 218.400 904.050 219.600 ;
        RECT 889.950 217.950 892.050 218.400 ;
        RECT 901.950 217.950 904.050 218.400 ;
        RECT 913.950 219.600 916.050 220.050 ;
        RECT 922.950 219.600 925.050 219.900 ;
        RECT 913.950 218.400 925.050 219.600 ;
        RECT 913.950 217.950 916.050 218.400 ;
        RECT 922.950 217.800 925.050 218.400 ;
        RECT 871.950 216.000 882.600 216.600 ;
        RECT 872.400 215.400 882.600 216.000 ;
        RECT 847.950 215.100 850.050 215.400 ;
        RECT 862.950 215.100 865.050 215.400 ;
        RECT 623.400 212.400 666.600 213.600 ;
        RECT 631.950 210.600 634.050 210.900 ;
        RECT 575.400 210.000 606.600 210.600 ;
        RECT 626.400 210.000 634.050 210.600 ;
        RECT 575.400 209.400 607.050 210.000 ;
        RECT 523.950 208.800 526.050 209.250 ;
        RECT 550.950 208.800 553.050 209.250 ;
        RECT 310.950 206.400 321.600 207.600 ;
        RECT 328.950 207.600 331.050 208.050 ;
        RECT 337.950 207.600 340.050 208.050 ;
        RECT 328.950 206.400 340.050 207.600 ;
        RECT 310.950 205.950 313.050 206.400 ;
        RECT 328.950 205.950 331.050 206.400 ;
        RECT 337.950 205.950 340.050 206.400 ;
        RECT 373.950 207.600 376.050 208.050 ;
        RECT 403.950 207.600 406.050 208.050 ;
        RECT 373.950 206.400 406.050 207.600 ;
        RECT 373.950 205.950 376.050 206.400 ;
        RECT 403.950 205.950 406.050 206.400 ;
        RECT 430.950 207.600 433.050 208.050 ;
        RECT 448.950 207.600 451.050 208.050 ;
        RECT 430.950 206.400 451.050 207.600 ;
        RECT 430.950 205.950 433.050 206.400 ;
        RECT 448.950 205.950 451.050 206.400 ;
        RECT 604.950 205.950 607.050 209.400 ;
        RECT 625.950 209.400 634.050 210.000 ;
        RECT 625.950 205.950 628.050 209.400 ;
        RECT 631.950 208.800 634.050 209.400 ;
        RECT 643.950 210.450 646.050 210.900 ;
        RECT 652.950 210.450 655.050 210.900 ;
        RECT 643.950 209.250 655.050 210.450 ;
        RECT 643.950 208.800 646.050 209.250 ;
        RECT 652.950 208.800 655.050 209.250 ;
        RECT 667.950 210.600 670.050 210.900 ;
        RECT 679.950 210.600 682.050 211.050 ;
        RECT 667.950 209.400 682.050 210.600 ;
        RECT 667.950 208.800 670.050 209.400 ;
        RECT 679.950 208.950 682.050 209.400 ;
        RECT 703.950 210.450 706.050 210.900 ;
        RECT 712.950 210.450 715.050 210.900 ;
        RECT 703.950 209.250 715.050 210.450 ;
        RECT 703.950 208.800 706.050 209.250 ;
        RECT 712.950 208.800 715.050 209.250 ;
        RECT 745.950 210.450 748.050 210.900 ;
        RECT 757.950 210.450 760.050 210.900 ;
        RECT 745.950 209.250 760.050 210.450 ;
        RECT 745.950 208.800 748.050 209.250 ;
        RECT 757.950 208.800 760.050 209.250 ;
        RECT 793.950 210.450 796.050 210.900 ;
        RECT 802.950 210.450 805.050 210.900 ;
        RECT 793.950 209.250 805.050 210.450 ;
        RECT 793.950 208.800 796.050 209.250 ;
        RECT 802.950 208.800 805.050 209.250 ;
        RECT 832.950 210.600 835.050 211.050 ;
        RECT 838.950 210.600 841.050 211.050 ;
        RECT 832.950 209.400 841.050 210.600 ;
        RECT 832.950 208.950 835.050 209.400 ;
        RECT 838.950 208.950 841.050 209.400 ;
        RECT 844.950 210.600 847.050 210.900 ;
        RECT 865.950 210.600 868.050 210.900 ;
        RECT 844.950 209.400 868.050 210.600 ;
        RECT 844.950 208.800 847.050 209.400 ;
        RECT 736.950 207.600 739.050 208.050 ;
        RECT 746.400 207.600 747.600 208.800 ;
        RECT 736.950 206.400 747.600 207.600 ;
        RECT 817.950 207.600 820.050 208.050 ;
        RECT 817.950 206.400 831.600 207.600 ;
        RECT 736.950 205.950 739.050 206.400 ;
        RECT 817.950 205.950 820.050 206.400 ;
        RECT 193.950 204.600 196.050 205.050 ;
        RECT 229.950 204.600 232.050 205.050 ;
        RECT 193.950 203.400 232.050 204.600 ;
        RECT 193.950 202.950 196.050 203.400 ;
        RECT 229.950 202.950 232.050 203.400 ;
        RECT 265.950 204.600 268.050 205.050 ;
        RECT 274.950 204.600 277.050 205.050 ;
        RECT 265.950 203.400 277.050 204.600 ;
        RECT 265.950 202.950 268.050 203.400 ;
        RECT 274.950 202.950 277.050 203.400 ;
        RECT 298.950 204.600 301.050 205.050 ;
        RECT 307.950 204.600 310.050 205.050 ;
        RECT 298.950 203.400 310.050 204.600 ;
        RECT 298.950 202.950 301.050 203.400 ;
        RECT 307.950 202.950 310.050 203.400 ;
        RECT 340.950 204.600 343.050 205.050 ;
        RECT 349.950 204.600 352.050 205.050 ;
        RECT 340.950 203.400 352.050 204.600 ;
        RECT 340.950 202.950 343.050 203.400 ;
        RECT 349.950 202.950 352.050 203.400 ;
        RECT 385.950 204.600 388.050 205.050 ;
        RECT 397.950 204.600 400.050 205.050 ;
        RECT 385.950 203.400 400.050 204.600 ;
        RECT 385.950 202.950 388.050 203.400 ;
        RECT 397.950 202.950 400.050 203.400 ;
        RECT 409.950 204.600 412.050 205.050 ;
        RECT 418.950 204.600 421.050 205.050 ;
        RECT 472.950 204.600 475.050 205.050 ;
        RECT 517.950 204.600 520.050 205.050 ;
        RECT 409.950 203.400 471.600 204.600 ;
        RECT 409.950 202.950 412.050 203.400 ;
        RECT 418.950 202.950 421.050 203.400 ;
        RECT 88.950 201.600 91.050 202.050 ;
        RECT 124.950 201.600 127.050 202.050 ;
        RECT 142.950 201.600 145.050 202.050 ;
        RECT 88.950 200.400 145.050 201.600 ;
        RECT 88.950 199.950 91.050 200.400 ;
        RECT 124.950 199.950 127.050 200.400 ;
        RECT 142.950 199.950 145.050 200.400 ;
        RECT 166.950 201.600 169.050 202.050 ;
        RECT 199.950 201.600 202.050 202.050 ;
        RECT 166.950 200.400 202.050 201.600 ;
        RECT 166.950 199.950 169.050 200.400 ;
        RECT 199.950 199.950 202.050 200.400 ;
        RECT 211.950 201.600 214.050 202.050 ;
        RECT 220.950 201.600 223.050 202.050 ;
        RECT 211.950 200.400 223.050 201.600 ;
        RECT 211.950 199.950 214.050 200.400 ;
        RECT 220.950 199.950 223.050 200.400 ;
        RECT 283.950 201.600 286.050 202.050 ;
        RECT 295.950 201.600 298.050 202.050 ;
        RECT 283.950 200.400 298.050 201.600 ;
        RECT 283.950 199.950 286.050 200.400 ;
        RECT 295.950 199.950 298.050 200.400 ;
        RECT 301.950 201.600 304.050 202.050 ;
        RECT 352.950 201.600 355.050 202.050 ;
        RECT 301.950 200.400 355.050 201.600 ;
        RECT 470.400 201.600 471.600 203.400 ;
        RECT 472.950 203.400 520.050 204.600 ;
        RECT 472.950 202.950 475.050 203.400 ;
        RECT 517.950 202.950 520.050 203.400 ;
        RECT 562.950 204.600 565.050 205.050 ;
        RECT 605.400 204.600 606.600 205.950 ;
        RECT 562.950 203.400 606.600 204.600 ;
        RECT 613.950 204.600 616.050 205.050 ;
        RECT 622.950 204.600 625.050 205.050 ;
        RECT 646.950 204.600 649.050 205.050 ;
        RECT 613.950 203.400 649.050 204.600 ;
        RECT 562.950 202.950 565.050 203.400 ;
        RECT 613.950 202.950 616.050 203.400 ;
        RECT 622.950 202.950 625.050 203.400 ;
        RECT 646.950 202.950 649.050 203.400 ;
        RECT 763.950 204.600 766.050 205.050 ;
        RECT 814.950 204.600 817.050 205.050 ;
        RECT 820.950 204.600 823.050 205.050 ;
        RECT 763.950 203.400 823.050 204.600 ;
        RECT 830.400 204.600 831.600 206.400 ;
        RECT 859.950 205.950 862.050 209.400 ;
        RECT 865.950 208.800 868.050 209.400 ;
        RECT 871.950 210.600 874.050 210.900 ;
        RECT 877.950 210.600 880.050 211.050 ;
        RECT 871.950 209.400 880.050 210.600 ;
        RECT 871.950 208.800 874.050 209.400 ;
        RECT 877.950 208.950 880.050 209.400 ;
        RECT 881.400 207.600 882.600 215.400 ;
        RECT 892.950 215.100 895.050 217.200 ;
        RECT 893.400 208.050 894.600 215.100 ;
        RECT 898.950 214.950 901.050 217.050 ;
        RECT 928.950 214.950 931.050 217.050 ;
        RECT 943.950 214.950 946.050 217.050 ;
        RECT 899.400 210.600 900.600 214.950 ;
        RECT 929.400 211.050 930.600 214.950 ;
        RECT 944.400 211.050 945.600 214.950 ;
        RECT 907.950 210.600 910.050 210.900 ;
        RECT 899.400 209.400 910.050 210.600 ;
        RECT 907.950 208.800 910.050 209.400 ;
        RECT 913.950 210.450 916.050 210.900 ;
        RECT 922.950 210.450 925.050 210.900 ;
        RECT 913.950 209.250 925.050 210.450 ;
        RECT 913.950 208.800 916.050 209.250 ;
        RECT 922.950 208.800 925.050 209.250 ;
        RECT 928.950 208.950 931.050 211.050 ;
        RECT 943.950 208.950 946.050 211.050 ;
        RECT 886.950 207.600 889.050 208.050 ;
        RECT 881.400 206.400 889.050 207.600 ;
        RECT 886.950 205.950 889.050 206.400 ;
        RECT 892.950 205.950 895.050 208.050 ;
        RECT 844.950 204.600 847.050 205.050 ;
        RECT 830.400 203.400 847.050 204.600 ;
        RECT 763.950 202.950 766.050 203.400 ;
        RECT 814.950 202.950 817.050 203.400 ;
        RECT 820.950 202.950 823.050 203.400 ;
        RECT 844.950 202.950 847.050 203.400 ;
        RECT 895.950 204.600 898.050 205.050 ;
        RECT 907.950 204.600 910.050 205.050 ;
        RECT 895.950 203.400 910.050 204.600 ;
        RECT 895.950 202.950 898.050 203.400 ;
        RECT 907.950 202.950 910.050 203.400 ;
        RECT 919.950 204.600 922.050 204.900 ;
        RECT 928.950 204.600 931.050 205.050 ;
        RECT 937.950 204.600 940.050 205.050 ;
        RECT 919.950 203.400 940.050 204.600 ;
        RECT 919.950 202.800 922.050 203.400 ;
        RECT 928.950 202.950 931.050 203.400 ;
        RECT 937.950 202.950 940.050 203.400 ;
        RECT 550.950 201.600 553.050 202.050 ;
        RECT 559.950 201.600 562.050 202.050 ;
        RECT 470.400 200.400 492.600 201.600 ;
        RECT 301.950 199.950 304.050 200.400 ;
        RECT 352.950 199.950 355.050 200.400 ;
        RECT 112.950 198.600 115.050 199.050 ;
        RECT 121.950 198.600 124.050 199.050 ;
        RECT 112.950 197.400 124.050 198.600 ;
        RECT 112.950 196.950 115.050 197.400 ;
        RECT 121.950 196.950 124.050 197.400 ;
        RECT 136.950 198.600 139.050 199.050 ;
        RECT 175.950 198.600 178.050 199.050 ;
        RECT 229.950 198.600 232.050 199.050 ;
        RECT 136.950 197.400 232.050 198.600 ;
        RECT 136.950 196.950 139.050 197.400 ;
        RECT 175.950 196.950 178.050 197.400 ;
        RECT 229.950 196.950 232.050 197.400 ;
        RECT 298.950 198.600 301.050 199.050 ;
        RECT 331.950 198.600 334.050 199.050 ;
        RECT 298.950 197.400 334.050 198.600 ;
        RECT 298.950 196.950 301.050 197.400 ;
        RECT 331.950 196.950 334.050 197.400 ;
        RECT 343.950 198.600 346.050 199.050 ;
        RECT 355.950 198.600 358.050 199.050 ;
        RECT 343.950 197.400 358.050 198.600 ;
        RECT 343.950 196.950 346.050 197.400 ;
        RECT 355.950 196.950 358.050 197.400 ;
        RECT 361.950 198.600 364.050 199.050 ;
        RECT 373.950 198.600 376.050 199.050 ;
        RECT 361.950 197.400 376.050 198.600 ;
        RECT 361.950 196.950 364.050 197.400 ;
        RECT 373.950 196.950 376.050 197.400 ;
        RECT 466.950 198.600 469.050 199.050 ;
        RECT 472.950 198.600 475.050 199.050 ;
        RECT 466.950 197.400 475.050 198.600 ;
        RECT 491.400 198.600 492.600 200.400 ;
        RECT 550.950 200.400 562.050 201.600 ;
        RECT 550.950 199.950 553.050 200.400 ;
        RECT 559.950 199.950 562.050 200.400 ;
        RECT 565.950 201.600 568.050 202.050 ;
        RECT 586.950 201.600 589.050 202.050 ;
        RECT 565.950 200.400 589.050 201.600 ;
        RECT 565.950 199.950 568.050 200.400 ;
        RECT 586.950 199.950 589.050 200.400 ;
        RECT 661.950 201.600 664.050 202.050 ;
        RECT 685.950 201.600 688.050 202.050 ;
        RECT 700.950 201.600 703.050 202.050 ;
        RECT 808.950 201.600 811.050 202.050 ;
        RECT 862.950 201.600 865.050 202.050 ;
        RECT 877.950 201.600 880.050 202.050 ;
        RECT 661.950 200.400 703.050 201.600 ;
        RECT 661.950 199.950 664.050 200.400 ;
        RECT 685.950 199.950 688.050 200.400 ;
        RECT 700.950 199.950 703.050 200.400 ;
        RECT 749.400 200.400 807.600 201.600 ;
        RECT 749.400 199.050 750.600 200.400 ;
        RECT 493.950 198.600 496.050 199.050 ;
        RECT 523.950 198.600 526.050 199.050 ;
        RECT 491.400 197.400 526.050 198.600 ;
        RECT 466.950 196.950 469.050 197.400 ;
        RECT 472.950 196.950 475.050 197.400 ;
        RECT 493.950 196.950 496.050 197.400 ;
        RECT 523.950 196.950 526.050 197.400 ;
        RECT 532.950 198.600 535.050 199.050 ;
        RECT 646.950 198.600 649.050 199.050 ;
        RECT 532.950 197.400 649.050 198.600 ;
        RECT 532.950 196.950 535.050 197.400 ;
        RECT 646.950 196.950 649.050 197.400 ;
        RECT 658.950 198.600 661.050 199.050 ;
        RECT 748.950 198.600 751.050 199.050 ;
        RECT 658.950 197.400 751.050 198.600 ;
        RECT 806.400 198.600 807.600 200.400 ;
        RECT 808.950 200.400 880.050 201.600 ;
        RECT 808.950 199.950 811.050 200.400 ;
        RECT 862.950 199.950 865.050 200.400 ;
        RECT 877.950 199.950 880.050 200.400 ;
        RECT 922.950 201.600 925.050 202.050 ;
        RECT 934.950 201.600 937.050 202.050 ;
        RECT 922.950 200.400 937.050 201.600 ;
        RECT 922.950 199.950 925.050 200.400 ;
        RECT 934.950 199.950 937.050 200.400 ;
        RECT 817.950 198.600 820.050 199.050 ;
        RECT 806.400 197.400 820.050 198.600 ;
        RECT 658.950 196.950 661.050 197.400 ;
        RECT 748.950 196.950 751.050 197.400 ;
        RECT 817.950 196.950 820.050 197.400 ;
        RECT 874.950 198.600 877.050 199.050 ;
        RECT 895.950 198.600 898.050 199.050 ;
        RECT 874.950 197.400 898.050 198.600 ;
        RECT 874.950 196.950 877.050 197.400 ;
        RECT 895.950 196.950 898.050 197.400 ;
        RECT 910.950 198.600 913.050 199.050 ;
        RECT 916.950 198.600 919.050 199.050 ;
        RECT 910.950 197.400 919.050 198.600 ;
        RECT 910.950 196.950 913.050 197.400 ;
        RECT 916.950 196.950 919.050 197.400 ;
        RECT 232.950 195.600 235.050 196.050 ;
        RECT 268.950 195.600 271.050 196.050 ;
        RECT 232.950 194.400 271.050 195.600 ;
        RECT 232.950 193.950 235.050 194.400 ;
        RECT 268.950 193.950 271.050 194.400 ;
        RECT 289.950 195.600 292.050 196.050 ;
        RECT 334.950 195.600 337.050 196.050 ;
        RECT 289.950 194.400 337.050 195.600 ;
        RECT 289.950 193.950 292.050 194.400 ;
        RECT 334.950 193.950 337.050 194.400 ;
        RECT 361.950 195.600 364.050 195.900 ;
        RECT 382.950 195.600 385.050 196.050 ;
        RECT 361.950 194.400 385.050 195.600 ;
        RECT 361.950 193.800 364.050 194.400 ;
        RECT 382.950 193.950 385.050 194.400 ;
        RECT 406.950 195.600 409.050 196.050 ;
        RECT 433.950 195.600 436.050 196.050 ;
        RECT 406.950 194.400 436.050 195.600 ;
        RECT 406.950 193.950 409.050 194.400 ;
        RECT 433.950 193.950 436.050 194.400 ;
        RECT 460.950 195.600 463.050 196.050 ;
        RECT 475.950 195.600 478.050 196.050 ;
        RECT 460.950 194.400 478.050 195.600 ;
        RECT 460.950 193.950 463.050 194.400 ;
        RECT 475.950 193.950 478.050 194.400 ;
        RECT 499.950 195.600 502.050 196.050 ;
        RECT 508.950 195.600 511.050 196.050 ;
        RECT 499.950 194.400 511.050 195.600 ;
        RECT 499.950 193.950 502.050 194.400 ;
        RECT 508.950 193.950 511.050 194.400 ;
        RECT 520.950 195.600 523.050 196.050 ;
        RECT 529.950 195.600 532.050 196.050 ;
        RECT 520.950 194.400 532.050 195.600 ;
        RECT 520.950 193.950 523.050 194.400 ;
        RECT 529.950 193.950 532.050 194.400 ;
        RECT 559.950 195.600 562.050 196.050 ;
        RECT 619.950 195.600 622.050 196.050 ;
        RECT 559.950 194.400 622.050 195.600 ;
        RECT 559.950 193.950 562.050 194.400 ;
        RECT 619.950 193.950 622.050 194.400 ;
        RECT 712.950 195.600 715.050 196.050 ;
        RECT 718.950 195.600 721.050 196.050 ;
        RECT 712.950 194.400 721.050 195.600 ;
        RECT 712.950 193.950 715.050 194.400 ;
        RECT 718.950 193.950 721.050 194.400 ;
        RECT 781.950 195.600 784.050 196.050 ;
        RECT 826.950 195.600 829.050 196.050 ;
        RECT 781.950 194.400 829.050 195.600 ;
        RECT 781.950 193.950 784.050 194.400 ;
        RECT 826.950 193.950 829.050 194.400 ;
        RECT 850.950 195.600 853.050 196.050 ;
        RECT 898.950 195.600 901.050 196.050 ;
        RECT 850.950 194.400 901.050 195.600 ;
        RECT 850.950 193.950 853.050 194.400 ;
        RECT 898.950 193.950 901.050 194.400 ;
        RECT 103.950 192.600 106.050 193.050 ;
        RECT 151.950 192.600 154.050 193.050 ;
        RECT 103.950 191.400 154.050 192.600 ;
        RECT 103.950 190.950 106.050 191.400 ;
        RECT 151.950 190.950 154.050 191.400 ;
        RECT 223.950 192.600 226.050 193.050 ;
        RECT 394.950 192.600 397.050 193.050 ;
        RECT 556.950 192.600 559.050 193.050 ;
        RECT 652.950 192.600 655.050 193.050 ;
        RECT 223.950 191.400 655.050 192.600 ;
        RECT 223.950 190.950 226.050 191.400 ;
        RECT 394.950 190.950 397.050 191.400 ;
        RECT 556.950 190.950 559.050 191.400 ;
        RECT 652.950 190.950 655.050 191.400 ;
        RECT 694.950 192.600 697.050 193.050 ;
        RECT 754.950 192.600 757.050 193.050 ;
        RECT 694.950 191.400 757.050 192.600 ;
        RECT 694.950 190.950 697.050 191.400 ;
        RECT 754.950 190.950 757.050 191.400 ;
        RECT 829.950 192.600 832.050 193.050 ;
        RECT 865.950 192.600 868.050 193.050 ;
        RECT 829.950 191.400 868.050 192.600 ;
        RECT 829.950 190.950 832.050 191.400 ;
        RECT 865.950 190.950 868.050 191.400 ;
        RECT 871.950 192.600 874.050 193.050 ;
        RECT 889.950 192.600 892.050 193.050 ;
        RECT 871.950 191.400 892.050 192.600 ;
        RECT 871.950 190.950 874.050 191.400 ;
        RECT 889.950 190.950 892.050 191.400 ;
        RECT 916.950 192.600 919.050 193.050 ;
        RECT 931.950 192.600 934.050 193.050 ;
        RECT 940.950 192.600 943.050 193.050 ;
        RECT 916.950 192.000 927.450 192.600 ;
        RECT 916.950 191.400 928.050 192.000 ;
        RECT 916.950 190.950 919.050 191.400 ;
        RECT 925.950 190.050 928.050 191.400 ;
        RECT 931.950 191.400 943.050 192.600 ;
        RECT 931.950 190.950 934.050 191.400 ;
        RECT 940.950 190.950 943.050 191.400 ;
        RECT 67.950 189.600 70.050 190.050 ;
        RECT 97.950 189.600 100.050 190.050 ;
        RECT 67.950 188.400 100.050 189.600 ;
        RECT 67.950 187.950 70.050 188.400 ;
        RECT 97.950 187.950 100.050 188.400 ;
        RECT 109.950 189.600 112.050 190.050 ;
        RECT 118.950 189.600 121.050 190.050 ;
        RECT 109.950 188.400 121.050 189.600 ;
        RECT 109.950 187.950 112.050 188.400 ;
        RECT 118.950 187.950 121.050 188.400 ;
        RECT 160.950 189.600 163.050 190.050 ;
        RECT 175.950 189.600 178.050 190.050 ;
        RECT 160.950 188.400 178.050 189.600 ;
        RECT 160.950 187.950 163.050 188.400 ;
        RECT 175.950 187.950 178.050 188.400 ;
        RECT 277.950 189.600 280.050 190.050 ;
        RECT 286.950 189.600 289.050 190.050 ;
        RECT 277.950 188.400 289.050 189.600 ;
        RECT 277.950 187.950 280.050 188.400 ;
        RECT 286.950 187.950 289.050 188.400 ;
        RECT 304.950 189.600 307.050 190.050 ;
        RECT 331.950 189.600 334.050 190.050 ;
        RECT 304.950 188.400 334.050 189.600 ;
        RECT 304.950 187.950 307.050 188.400 ;
        RECT 331.950 187.950 334.050 188.400 ;
        RECT 349.950 189.600 352.050 190.050 ;
        RECT 358.950 189.600 361.050 190.050 ;
        RECT 349.950 188.400 361.050 189.600 ;
        RECT 349.950 187.950 352.050 188.400 ;
        RECT 358.950 187.950 361.050 188.400 ;
        RECT 364.950 189.600 367.050 190.050 ;
        RECT 391.950 189.600 394.050 190.050 ;
        RECT 364.950 188.400 394.050 189.600 ;
        RECT 364.950 187.950 367.050 188.400 ;
        RECT 391.950 187.950 394.050 188.400 ;
        RECT 439.950 189.600 442.050 190.050 ;
        RECT 457.950 189.600 460.050 190.050 ;
        RECT 439.950 188.400 460.050 189.600 ;
        RECT 439.950 187.950 442.050 188.400 ;
        RECT 457.950 187.950 460.050 188.400 ;
        RECT 463.950 189.600 466.050 190.050 ;
        RECT 469.950 189.600 472.050 190.050 ;
        RECT 463.950 188.400 472.050 189.600 ;
        RECT 463.950 187.950 466.050 188.400 ;
        RECT 469.950 187.950 472.050 188.400 ;
        RECT 496.950 189.600 499.050 190.050 ;
        RECT 505.950 189.600 508.050 190.050 ;
        RECT 523.950 189.600 526.050 190.050 ;
        RECT 496.950 188.400 526.050 189.600 ;
        RECT 496.950 187.950 499.050 188.400 ;
        RECT 505.950 187.950 508.050 188.400 ;
        RECT 523.950 187.950 526.050 188.400 ;
        RECT 583.950 189.600 586.050 190.050 ;
        RECT 592.950 189.600 595.050 190.050 ;
        RECT 583.950 188.400 595.050 189.600 ;
        RECT 583.950 187.950 586.050 188.400 ;
        RECT 592.950 187.950 595.050 188.400 ;
        RECT 598.950 189.600 601.050 190.050 ;
        RECT 625.950 189.600 628.050 190.050 ;
        RECT 598.950 188.400 628.050 189.600 ;
        RECT 598.950 187.950 601.050 188.400 ;
        RECT 625.950 187.950 628.050 188.400 ;
        RECT 691.950 189.600 694.050 190.050 ;
        RECT 718.950 189.600 721.050 190.050 ;
        RECT 691.950 188.400 721.050 189.600 ;
        RECT 691.950 187.950 694.050 188.400 ;
        RECT 718.950 187.950 721.050 188.400 ;
        RECT 739.950 189.600 742.050 190.050 ;
        RECT 769.950 189.600 772.050 190.050 ;
        RECT 739.950 188.400 772.050 189.600 ;
        RECT 739.950 187.950 742.050 188.400 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 784.950 189.600 787.050 190.050 ;
        RECT 820.950 189.600 823.050 190.050 ;
        RECT 784.950 188.400 823.050 189.600 ;
        RECT 784.950 187.950 787.050 188.400 ;
        RECT 820.950 187.950 823.050 188.400 ;
        RECT 850.950 189.600 853.050 190.050 ;
        RECT 874.950 189.600 877.050 190.050 ;
        RECT 850.950 188.400 877.050 189.600 ;
        RECT 850.950 187.950 853.050 188.400 ;
        RECT 874.950 187.950 877.050 188.400 ;
        RECT 892.950 187.950 895.050 190.050 ;
        RECT 925.800 189.000 928.050 190.050 ;
        RECT 928.950 189.600 931.050 190.050 ;
        RECT 943.950 189.600 946.050 190.050 ;
        RECT 925.800 187.950 927.900 189.000 ;
        RECT 928.950 188.400 946.050 189.600 ;
        RECT 928.950 187.950 931.050 188.400 ;
        RECT 943.950 187.950 946.050 188.400 ;
        RECT 22.950 186.600 25.050 187.050 ;
        RECT 31.950 186.600 34.050 187.050 ;
        RECT 61.950 186.600 64.050 187.050 ;
        RECT 22.950 185.400 34.050 186.600 ;
        RECT 22.950 184.950 25.050 185.400 ;
        RECT 31.950 184.950 34.050 185.400 ;
        RECT 44.400 185.400 64.050 186.600 ;
        RECT 4.950 183.750 7.050 184.200 ;
        RECT 16.950 183.750 19.050 184.200 ;
        RECT 4.950 182.550 19.050 183.750 ;
        RECT 4.950 182.100 7.050 182.550 ;
        RECT 16.950 182.100 19.050 182.550 ;
        RECT 25.950 183.600 28.050 184.050 ;
        RECT 25.950 182.400 33.600 183.600 ;
        RECT 25.950 181.950 28.050 182.400 ;
        RECT 32.400 177.600 33.600 182.400 ;
        RECT 44.400 177.900 45.600 185.400 ;
        RECT 61.950 184.950 64.050 185.400 ;
        RECT 91.950 184.950 94.050 187.050 ;
        RECT 133.950 186.600 136.050 187.050 ;
        RECT 128.400 185.400 136.050 186.600 ;
        RECT 46.950 183.750 49.050 184.200 ;
        RECT 52.950 183.750 55.050 184.200 ;
        RECT 46.950 182.550 55.050 183.750 ;
        RECT 46.950 182.100 49.050 182.550 ;
        RECT 52.950 182.100 55.050 182.550 ;
        RECT 76.950 183.750 79.050 184.200 ;
        RECT 82.950 183.750 85.050 184.200 ;
        RECT 76.950 182.550 85.050 183.750 ;
        RECT 76.950 182.100 79.050 182.550 ;
        RECT 82.950 182.100 85.050 182.550 ;
        RECT 37.950 177.600 40.050 177.900 ;
        RECT 32.400 176.400 40.050 177.600 ;
        RECT 37.950 175.800 40.050 176.400 ;
        RECT 43.950 175.800 46.050 177.900 ;
        RECT 52.950 177.600 55.050 178.050 ;
        RECT 85.950 177.600 88.050 177.900 ;
        RECT 52.950 176.400 88.050 177.600 ;
        RECT 52.950 175.950 55.050 176.400 ;
        RECT 85.950 175.800 88.050 176.400 ;
        RECT 92.400 175.050 93.600 184.950 ;
        RECT 103.950 182.100 106.050 184.200 ;
        RECT 94.950 177.600 97.050 178.050 ;
        RECT 104.400 177.600 105.600 182.100 ;
        RECT 128.400 177.900 129.600 185.400 ;
        RECT 133.950 184.950 136.050 185.400 ;
        RECT 157.950 186.600 160.050 187.050 ;
        RECT 163.950 186.600 166.050 187.050 ;
        RECT 157.950 185.400 166.050 186.600 ;
        RECT 157.950 184.950 160.050 185.400 ;
        RECT 163.950 184.950 166.050 185.400 ;
        RECT 223.950 184.950 226.050 187.050 ;
        RECT 241.950 186.600 244.050 187.050 ;
        RECT 253.950 186.600 256.050 187.050 ;
        RECT 241.950 185.400 256.050 186.600 ;
        RECT 241.950 184.950 244.050 185.400 ;
        RECT 253.950 184.950 256.050 185.400 ;
        RECT 259.950 184.950 262.050 187.050 ;
        RECT 301.950 186.600 304.050 187.050 ;
        RECT 290.400 185.400 304.050 186.600 ;
        RECT 130.950 183.750 133.050 184.200 ;
        RECT 145.950 183.750 148.050 184.200 ;
        RECT 130.950 182.550 148.050 183.750 ;
        RECT 130.950 182.100 133.050 182.550 ;
        RECT 145.950 182.100 148.050 182.550 ;
        RECT 169.950 181.950 172.050 184.050 ;
        RECT 175.950 183.750 178.050 184.200 ;
        RECT 187.950 183.750 190.050 184.200 ;
        RECT 175.950 182.550 190.050 183.750 ;
        RECT 175.950 182.100 178.050 182.550 ;
        RECT 187.950 182.100 190.050 182.550 ;
        RECT 199.950 182.100 202.050 184.200 ;
        RECT 94.950 176.400 105.600 177.600 ;
        RECT 94.950 175.950 97.050 176.400 ;
        RECT 127.950 175.800 130.050 177.900 ;
        RECT 133.950 177.450 136.050 177.900 ;
        RECT 142.950 177.450 145.050 177.900 ;
        RECT 133.950 176.250 145.050 177.450 ;
        RECT 133.950 175.800 136.050 176.250 ;
        RECT 142.950 175.800 145.050 176.250 ;
        RECT 91.950 172.950 94.050 175.050 ;
        RECT 97.950 174.600 100.050 175.050 ;
        RECT 112.950 174.600 115.050 175.050 ;
        RECT 97.950 173.400 115.050 174.600 ;
        RECT 97.950 172.950 100.050 173.400 ;
        RECT 112.950 172.950 115.050 173.400 ;
        RECT 148.950 174.600 151.050 175.050 ;
        RECT 157.950 174.600 160.050 175.050 ;
        RECT 148.950 173.400 160.050 174.600 ;
        RECT 170.400 174.600 171.600 181.950 ;
        RECT 181.950 177.600 184.050 178.050 ;
        RECT 200.400 177.600 201.600 182.100 ;
        RECT 224.400 177.900 225.600 184.950 ;
        RECT 229.950 183.600 232.050 184.050 ;
        RECT 229.950 182.400 240.600 183.600 ;
        RECT 229.950 181.950 232.050 182.400 ;
        RECT 239.400 177.900 240.600 182.400 ;
        RECT 256.950 181.950 259.050 184.050 ;
        RECT 257.400 178.050 258.600 181.950 ;
        RECT 181.950 176.400 201.600 177.600 ;
        RECT 181.950 175.950 184.050 176.400 ;
        RECT 223.950 175.800 226.050 177.900 ;
        RECT 238.950 175.800 241.050 177.900 ;
        RECT 256.800 175.950 258.900 178.050 ;
        RECT 260.400 177.900 261.600 184.950 ;
        RECT 262.950 183.600 265.050 184.200 ;
        RECT 268.950 183.600 271.050 184.200 ;
        RECT 286.950 183.600 289.050 184.200 ;
        RECT 262.950 182.400 267.600 183.600 ;
        RECT 262.950 182.100 265.050 182.400 ;
        RECT 266.400 180.600 267.600 182.400 ;
        RECT 268.950 182.400 289.050 183.600 ;
        RECT 268.950 182.100 271.050 182.400 ;
        RECT 286.950 182.100 289.050 182.400 ;
        RECT 266.400 180.000 273.600 180.600 ;
        RECT 266.400 179.400 274.050 180.000 ;
        RECT 259.950 175.800 262.050 177.900 ;
        RECT 271.950 175.950 274.050 179.400 ;
        RECT 290.400 177.900 291.600 185.400 ;
        RECT 301.950 184.950 304.050 185.400 ;
        RECT 334.950 186.600 337.050 187.050 ;
        RECT 415.950 186.600 418.050 187.050 ;
        RECT 334.950 185.400 418.050 186.600 ;
        RECT 334.950 184.950 337.050 185.400 ;
        RECT 415.950 184.950 418.050 185.400 ;
        RECT 502.950 186.600 505.050 187.050 ;
        RECT 514.950 186.600 517.050 187.050 ;
        RECT 502.950 185.400 517.050 186.600 ;
        RECT 502.950 184.950 505.050 185.400 ;
        RECT 514.950 184.950 517.050 185.400 ;
        RECT 535.950 186.600 538.050 187.050 ;
        RECT 541.950 186.600 544.050 187.050 ;
        RECT 535.950 185.400 544.050 186.600 ;
        RECT 535.950 184.950 538.050 185.400 ;
        RECT 541.950 184.950 544.050 185.400 ;
        RECT 559.950 186.600 562.050 187.050 ;
        RECT 574.950 186.600 577.050 187.050 ;
        RECT 559.950 185.400 577.050 186.600 ;
        RECT 559.950 184.950 562.050 185.400 ;
        RECT 574.950 184.950 577.050 185.400 ;
        RECT 586.950 186.600 589.050 187.050 ;
        RECT 628.950 186.600 631.050 187.050 ;
        RECT 586.950 185.400 631.050 186.600 ;
        RECT 586.950 184.950 589.050 185.400 ;
        RECT 628.950 184.950 631.050 185.400 ;
        RECT 634.950 186.600 637.050 187.050 ;
        RECT 643.950 186.600 646.050 187.050 ;
        RECT 634.950 185.400 646.050 186.600 ;
        RECT 634.950 184.950 637.050 185.400 ;
        RECT 643.950 184.950 646.050 185.400 ;
        RECT 670.950 186.600 673.050 187.050 ;
        RECT 676.950 186.600 679.050 187.050 ;
        RECT 724.950 186.600 727.050 187.050 ;
        RECT 748.950 186.600 751.050 187.050 ;
        RECT 811.950 186.600 814.050 187.050 ;
        RECT 817.950 186.600 820.050 187.050 ;
        RECT 670.950 185.400 679.050 186.600 ;
        RECT 670.950 184.950 673.050 185.400 ;
        RECT 676.950 184.950 679.050 185.400 ;
        RECT 716.400 185.400 762.600 186.600 ;
        RECT 298.950 180.600 301.050 184.050 ;
        RECT 304.950 182.100 307.050 184.200 ;
        RECT 298.950 180.000 303.600 180.600 ;
        RECT 299.400 179.400 303.600 180.000 ;
        RECT 302.400 177.900 303.600 179.400 ;
        RECT 289.950 175.800 292.050 177.900 ;
        RECT 301.950 175.800 304.050 177.900 ;
        RECT 305.400 175.050 306.600 182.100 ;
        RECT 310.950 181.950 313.050 184.050 ;
        RECT 316.950 183.600 319.050 184.050 ;
        RECT 325.950 183.600 328.050 184.200 ;
        RECT 316.950 182.400 328.050 183.600 ;
        RECT 316.950 181.950 319.050 182.400 ;
        RECT 325.950 182.100 328.050 182.400 ;
        RECT 343.950 183.600 346.050 184.050 ;
        RECT 355.950 183.600 358.050 184.200 ;
        RECT 367.950 183.600 370.050 184.050 ;
        RECT 391.950 183.600 394.050 184.200 ;
        RECT 412.950 183.600 415.050 184.200 ;
        RECT 343.950 182.400 354.600 183.600 ;
        RECT 343.950 181.950 346.050 182.400 ;
        RECT 307.950 177.450 310.050 177.900 ;
        RECT 311.400 177.450 312.600 181.950 ;
        RECT 319.950 177.450 322.050 177.900 ;
        RECT 307.950 176.250 322.050 177.450 ;
        RECT 307.950 175.800 310.050 176.250 ;
        RECT 319.950 175.800 322.050 176.250 ;
        RECT 337.950 177.600 340.050 178.050 ;
        RECT 343.950 177.600 346.050 178.050 ;
        RECT 353.400 177.900 354.600 182.400 ;
        RECT 355.950 182.400 360.600 183.600 ;
        RECT 355.950 182.100 358.050 182.400 ;
        RECT 359.400 178.050 360.600 182.400 ;
        RECT 367.950 182.400 381.600 183.600 ;
        RECT 367.950 181.950 370.050 182.400 ;
        RECT 361.950 180.600 364.050 181.050 ;
        RECT 361.950 179.400 378.600 180.600 ;
        RECT 361.950 178.950 364.050 179.400 ;
        RECT 337.950 176.400 346.050 177.600 ;
        RECT 337.950 175.950 340.050 176.400 ;
        RECT 343.950 175.950 346.050 176.400 ;
        RECT 352.950 175.800 355.050 177.900 ;
        RECT 358.950 175.950 361.050 178.050 ;
        RECT 377.400 177.900 378.600 179.400 ;
        RECT 364.950 177.450 367.050 177.900 ;
        RECT 370.950 177.450 373.050 177.900 ;
        RECT 364.950 176.250 373.050 177.450 ;
        RECT 364.950 175.800 367.050 176.250 ;
        RECT 370.950 175.800 373.050 176.250 ;
        RECT 376.950 175.800 379.050 177.900 ;
        RECT 380.400 177.600 381.600 182.400 ;
        RECT 391.950 182.400 415.050 183.600 ;
        RECT 391.950 182.100 394.050 182.400 ;
        RECT 412.950 182.100 415.050 182.400 ;
        RECT 418.950 181.950 421.050 184.050 ;
        RECT 427.950 183.600 430.050 184.050 ;
        RECT 451.950 183.600 454.050 184.050 ;
        RECT 463.950 183.600 466.050 184.200 ;
        RECT 427.950 182.400 444.600 183.600 ;
        RECT 427.950 181.950 430.050 182.400 ;
        RECT 419.400 178.050 420.600 181.950 ;
        RECT 394.950 177.600 397.050 177.900 ;
        RECT 380.400 176.400 397.050 177.600 ;
        RECT 394.950 175.800 397.050 176.400 ;
        RECT 403.950 175.950 406.050 178.050 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 443.400 177.900 444.600 182.400 ;
        RECT 451.950 182.400 466.050 183.600 ;
        RECT 451.950 181.950 454.050 182.400 ;
        RECT 463.950 182.100 466.050 182.400 ;
        RECT 469.950 181.950 472.050 184.050 ;
        RECT 481.950 183.600 484.050 184.200 ;
        RECT 479.400 182.400 484.050 183.600 ;
        RECT 470.400 178.050 471.600 181.950 ;
        RECT 479.400 178.050 480.600 182.400 ;
        RECT 481.950 182.100 484.050 182.400 ;
        RECT 493.950 183.600 496.050 184.050 ;
        RECT 493.950 182.400 504.600 183.600 ;
        RECT 493.950 181.950 496.050 182.400 ;
        RECT 172.950 174.600 175.050 175.050 ;
        RECT 199.800 174.600 201.900 175.050 ;
        RECT 170.400 173.400 201.900 174.600 ;
        RECT 148.950 172.950 151.050 173.400 ;
        RECT 157.950 172.950 160.050 173.400 ;
        RECT 172.950 172.950 175.050 173.400 ;
        RECT 199.800 172.950 201.900 173.400 ;
        RECT 202.950 174.600 205.050 175.050 ;
        RECT 232.950 174.600 235.050 175.050 ;
        RECT 202.950 173.400 235.050 174.600 ;
        RECT 202.950 172.950 205.050 173.400 ;
        RECT 232.950 172.950 235.050 173.400 ;
        RECT 247.950 174.600 250.050 175.050 ;
        RECT 274.950 174.600 277.050 175.050 ;
        RECT 247.950 173.400 277.050 174.600 ;
        RECT 247.950 172.950 250.050 173.400 ;
        RECT 274.950 172.950 277.050 173.400 ;
        RECT 304.950 172.950 307.050 175.050 ;
        RECT 127.950 171.600 130.050 172.050 ;
        RECT 139.950 171.600 142.050 172.050 ;
        RECT 127.950 170.400 142.050 171.600 ;
        RECT 127.950 169.950 130.050 170.400 ;
        RECT 139.950 169.950 142.050 170.400 ;
        RECT 154.950 171.600 157.050 172.050 ;
        RECT 184.950 171.600 187.050 172.050 ;
        RECT 154.950 170.400 187.050 171.600 ;
        RECT 154.950 169.950 157.050 170.400 ;
        RECT 184.950 169.950 187.050 170.400 ;
        RECT 196.950 171.600 199.050 172.050 ;
        RECT 289.950 171.600 292.050 172.050 ;
        RECT 196.950 170.400 292.050 171.600 ;
        RECT 196.950 169.950 199.050 170.400 ;
        RECT 289.950 169.950 292.050 170.400 ;
        RECT 295.950 171.600 298.050 172.050 ;
        RECT 370.950 171.600 373.050 172.050 ;
        RECT 295.950 170.400 373.050 171.600 ;
        RECT 295.950 169.950 298.050 170.400 ;
        RECT 370.950 169.950 373.050 170.400 ;
        RECT 388.950 171.600 391.050 172.050 ;
        RECT 404.400 171.600 405.600 175.950 ;
        RECT 442.950 175.800 445.050 177.900 ;
        RECT 469.950 175.950 472.050 178.050 ;
        RECT 478.950 175.950 481.050 178.050 ;
        RECT 503.400 177.900 504.600 182.400 ;
        RECT 511.950 181.950 514.050 184.050 ;
        RECT 550.950 183.600 553.050 184.200 ;
        RECT 556.950 183.600 559.050 184.050 ;
        RECT 550.950 182.400 559.050 183.600 ;
        RECT 550.950 182.100 553.050 182.400 ;
        RECT 556.950 181.950 559.050 182.400 ;
        RECT 562.950 183.600 567.000 184.050 ;
        RECT 577.950 183.750 580.050 184.200 ;
        RECT 586.950 183.750 589.050 184.200 ;
        RECT 562.950 181.950 567.600 183.600 ;
        RECT 577.950 182.550 589.050 183.750 ;
        RECT 598.950 183.600 601.050 184.050 ;
        RECT 577.950 182.100 580.050 182.550 ;
        RECT 586.950 182.100 589.050 182.550 ;
        RECT 593.400 182.400 601.050 183.600 ;
        RECT 490.950 177.450 493.050 177.900 ;
        RECT 496.950 177.450 499.050 177.900 ;
        RECT 490.950 176.250 499.050 177.450 ;
        RECT 490.950 175.800 493.050 176.250 ;
        RECT 496.950 175.800 499.050 176.250 ;
        RECT 502.950 175.800 505.050 177.900 ;
        RECT 508.950 177.600 511.050 177.900 ;
        RECT 512.400 177.600 513.600 181.950 ;
        RECT 566.400 177.900 567.600 181.950 ;
        RECT 593.400 180.600 594.600 182.400 ;
        RECT 598.950 181.950 601.050 182.400 ;
        RECT 604.950 183.600 609.000 184.050 ;
        RECT 625.950 183.600 628.050 184.050 ;
        RECT 639.000 183.600 643.050 184.050 ;
        RECT 604.950 181.950 609.600 183.600 ;
        RECT 625.950 182.400 633.600 183.600 ;
        RECT 625.950 181.950 628.050 182.400 ;
        RECT 590.400 179.400 594.600 180.600 ;
        RECT 590.400 177.900 591.600 179.400 ;
        RECT 608.400 177.900 609.600 181.950 ;
        RECT 632.400 177.900 633.600 182.400 ;
        RECT 638.400 181.950 643.050 183.600 ;
        RECT 667.950 183.750 670.050 184.200 ;
        RECT 679.950 183.750 682.050 184.200 ;
        RECT 667.950 183.600 682.050 183.750 ;
        RECT 716.400 183.600 717.600 185.400 ;
        RECT 724.950 184.950 727.050 185.400 ;
        RECT 748.950 184.950 751.050 185.400 ;
        RECT 667.950 182.550 717.600 183.600 ;
        RECT 667.950 182.100 670.050 182.550 ;
        RECT 679.950 182.400 717.600 182.550 ;
        RECT 718.950 183.600 721.050 184.200 ;
        RECT 730.950 183.600 733.050 184.050 ;
        RECT 718.950 182.400 733.050 183.600 ;
        RECT 761.400 183.600 762.600 185.400 ;
        RECT 811.950 185.400 820.050 186.600 ;
        RECT 811.950 184.950 814.050 185.400 ;
        RECT 817.950 184.950 820.050 185.400 ;
        RECT 826.950 186.600 829.050 187.050 ;
        RECT 841.950 186.600 844.050 187.050 ;
        RECT 826.950 185.400 834.600 186.600 ;
        RECT 826.950 184.950 829.050 185.400 ;
        RECT 763.950 183.600 766.050 184.200 ;
        RECT 761.400 182.400 766.050 183.600 ;
        RECT 679.950 182.100 682.050 182.400 ;
        RECT 718.950 182.100 721.050 182.400 ;
        RECT 730.950 181.950 733.050 182.400 ;
        RECT 763.950 182.100 766.050 182.400 ;
        RECT 778.950 182.100 781.050 184.200 ;
        RECT 796.950 183.750 799.050 184.200 ;
        RECT 802.950 183.750 805.050 184.200 ;
        RECT 796.950 182.550 805.050 183.750 ;
        RECT 796.950 182.100 799.050 182.550 ;
        RECT 802.950 182.100 805.050 182.550 ;
        RECT 823.950 183.600 828.000 184.050 ;
        RECT 638.400 177.900 639.600 181.950 ;
        RECT 779.400 180.600 780.600 182.100 ;
        RECT 823.950 181.950 828.600 183.600 ;
        RECT 793.950 180.600 796.050 181.050 ;
        RECT 779.400 179.400 796.050 180.600 ;
        RECT 793.950 178.950 796.050 179.400 ;
        RECT 508.950 176.400 513.600 177.600 ;
        RECT 526.950 177.600 529.050 177.900 ;
        RECT 541.950 177.600 544.050 177.900 ;
        RECT 526.950 176.400 544.050 177.600 ;
        RECT 508.950 175.800 511.050 176.400 ;
        RECT 526.950 175.800 529.050 176.400 ;
        RECT 541.950 175.800 544.050 176.400 ;
        RECT 565.950 175.800 568.050 177.900 ;
        RECT 571.950 177.450 574.050 177.900 ;
        RECT 580.950 177.450 583.050 177.900 ;
        RECT 571.950 176.250 583.050 177.450 ;
        RECT 571.950 175.800 574.050 176.250 ;
        RECT 580.950 175.800 583.050 176.250 ;
        RECT 589.950 175.800 592.050 177.900 ;
        RECT 595.950 177.450 598.050 177.900 ;
        RECT 601.950 177.450 604.050 177.900 ;
        RECT 595.950 176.250 604.050 177.450 ;
        RECT 595.950 175.800 598.050 176.250 ;
        RECT 601.950 175.800 604.050 176.250 ;
        RECT 607.950 175.800 610.050 177.900 ;
        RECT 631.950 175.800 634.050 177.900 ;
        RECT 637.950 175.800 640.050 177.900 ;
        RECT 655.950 177.600 658.050 177.900 ;
        RECT 667.950 177.600 670.050 178.050 ;
        RECT 655.950 176.400 670.050 177.600 ;
        RECT 655.950 175.800 658.050 176.400 ;
        RECT 667.950 175.950 670.050 176.400 ;
        RECT 682.950 177.600 685.050 177.900 ;
        RECT 691.950 177.600 694.050 178.050 ;
        RECT 682.950 176.400 694.050 177.600 ;
        RECT 682.950 175.800 685.050 176.400 ;
        RECT 691.950 175.950 694.050 176.400 ;
        RECT 730.950 177.450 733.050 177.900 ;
        RECT 736.950 177.450 739.050 177.900 ;
        RECT 730.950 176.250 739.050 177.450 ;
        RECT 730.950 175.800 733.050 176.250 ;
        RECT 736.950 175.800 739.050 176.250 ;
        RECT 742.950 177.450 745.050 177.900 ;
        RECT 748.800 177.450 750.900 177.900 ;
        RECT 742.950 176.250 750.900 177.450 ;
        RECT 742.950 175.800 745.050 176.250 ;
        RECT 748.800 175.800 750.900 176.250 ;
        RECT 751.950 177.600 754.050 178.050 ;
        RECT 766.950 177.600 769.050 177.900 ;
        RECT 781.950 177.600 784.050 177.900 ;
        RECT 751.950 177.000 765.600 177.600 ;
        RECT 751.950 176.400 766.050 177.000 ;
        RECT 751.950 175.950 754.050 176.400 ;
        RECT 581.400 174.600 582.600 175.800 ;
        RECT 613.950 174.600 616.050 175.050 ;
        RECT 581.400 173.400 616.050 174.600 ;
        RECT 613.950 172.950 616.050 173.400 ;
        RECT 763.950 172.950 766.050 176.400 ;
        RECT 766.950 176.400 784.050 177.600 ;
        RECT 766.950 175.800 769.050 176.400 ;
        RECT 781.950 175.800 784.050 176.400 ;
        RECT 799.950 177.600 802.050 178.050 ;
        RECT 814.950 177.600 817.050 178.050 ;
        RECT 827.400 177.900 828.600 181.950 ;
        RECT 833.400 177.900 834.600 185.400 ;
        RECT 841.950 185.400 879.600 186.600 ;
        RECT 841.950 184.950 844.050 185.400 ;
        RECT 835.950 183.600 838.050 184.050 ;
        RECT 835.950 182.400 855.600 183.600 ;
        RECT 835.950 181.950 838.050 182.400 ;
        RECT 854.400 180.600 855.600 182.400 ;
        RECT 854.400 179.400 873.600 180.600 ;
        RECT 872.400 177.900 873.600 179.400 ;
        RECT 878.400 177.900 879.600 185.400 ;
        RECT 886.950 181.950 889.050 184.050 ;
        RECT 887.400 178.050 888.600 181.950 ;
        RECT 799.950 176.400 817.050 177.600 ;
        RECT 799.950 175.950 802.050 176.400 ;
        RECT 814.950 175.950 817.050 176.400 ;
        RECT 826.950 175.800 829.050 177.900 ;
        RECT 832.950 175.800 835.050 177.900 ;
        RECT 871.950 175.800 874.050 177.900 ;
        RECT 877.950 175.800 880.050 177.900 ;
        RECT 886.950 175.950 889.050 178.050 ;
        RECT 893.400 175.050 894.600 187.950 ;
        RECT 898.950 183.600 901.050 184.200 ;
        RECT 910.950 183.600 913.050 184.200 ;
        RECT 921.000 183.600 925.050 184.050 ;
        RECT 898.950 182.400 913.050 183.600 ;
        RECT 898.950 182.100 901.050 182.400 ;
        RECT 910.950 182.100 913.050 182.400 ;
        RECT 920.400 181.950 925.050 183.600 ;
        RECT 934.950 182.100 937.050 184.200 ;
        RECT 946.950 183.600 951.000 184.050 ;
        RECT 920.400 178.050 921.600 181.950 ;
        RECT 920.400 176.400 925.050 178.050 ;
        RECT 921.000 175.950 925.050 176.400 ;
        RECT 935.400 175.050 936.600 182.100 ;
        RECT 946.950 181.950 951.600 183.600 ;
        RECT 950.400 175.050 951.600 181.950 ;
        RECT 853.950 174.600 856.050 175.050 ;
        RECT 859.950 174.600 862.050 175.050 ;
        RECT 853.950 173.400 862.050 174.600 ;
        RECT 853.950 172.950 856.050 173.400 ;
        RECT 859.950 172.950 862.050 173.400 ;
        RECT 889.950 173.400 894.600 175.050 ;
        RECT 904.950 174.600 907.050 175.050 ;
        RECT 910.950 174.600 913.050 175.050 ;
        RECT 904.950 173.400 913.050 174.600 ;
        RECT 889.950 172.950 894.000 173.400 ;
        RECT 904.950 172.950 907.050 173.400 ;
        RECT 910.950 172.950 913.050 173.400 ;
        RECT 934.950 172.950 937.050 175.050 ;
        RECT 946.950 173.400 951.600 175.050 ;
        RECT 946.950 172.950 951.000 173.400 ;
        RECT 388.950 170.400 405.600 171.600 ;
        RECT 415.950 171.600 418.050 172.050 ;
        RECT 445.950 171.600 448.050 172.050 ;
        RECT 415.950 170.400 448.050 171.600 ;
        RECT 388.950 169.950 391.050 170.400 ;
        RECT 415.950 169.950 418.050 170.400 ;
        RECT 445.950 169.950 448.050 170.400 ;
        RECT 451.950 171.600 454.050 172.050 ;
        RECT 484.950 171.600 487.050 172.050 ;
        RECT 451.950 170.400 487.050 171.600 ;
        RECT 451.950 169.950 454.050 170.400 ;
        RECT 484.950 169.950 487.050 170.400 ;
        RECT 517.950 171.600 520.050 172.050 ;
        RECT 529.950 171.600 532.050 172.050 ;
        RECT 517.950 170.400 532.050 171.600 ;
        RECT 517.950 169.950 520.050 170.400 ;
        RECT 529.950 169.950 532.050 170.400 ;
        RECT 535.950 171.600 538.050 172.050 ;
        RECT 688.950 171.600 691.050 172.050 ;
        RECT 694.950 171.600 697.050 172.050 ;
        RECT 535.950 170.400 697.050 171.600 ;
        RECT 535.950 169.950 538.050 170.400 ;
        RECT 688.950 169.950 691.050 170.400 ;
        RECT 694.950 169.950 697.050 170.400 ;
        RECT 730.950 171.600 733.050 172.050 ;
        RECT 751.950 171.600 754.050 172.050 ;
        RECT 730.950 170.400 754.050 171.600 ;
        RECT 730.950 169.950 733.050 170.400 ;
        RECT 751.950 169.950 754.050 170.400 ;
        RECT 757.950 171.600 760.050 171.900 ;
        RECT 793.950 171.600 796.050 172.050 ;
        RECT 805.950 171.600 808.050 172.050 ;
        RECT 757.950 170.400 808.050 171.600 ;
        RECT 757.950 169.800 760.050 170.400 ;
        RECT 793.950 169.950 796.050 170.400 ;
        RECT 805.950 169.950 808.050 170.400 ;
        RECT 817.950 171.600 820.050 172.050 ;
        RECT 835.950 171.600 838.050 172.050 ;
        RECT 817.950 170.400 838.050 171.600 ;
        RECT 817.950 169.950 820.050 170.400 ;
        RECT 835.950 169.950 838.050 170.400 ;
        RECT 925.950 171.600 928.050 172.050 ;
        RECT 937.950 171.600 940.050 172.050 ;
        RECT 925.950 170.400 940.050 171.600 ;
        RECT 925.950 169.950 928.050 170.400 ;
        RECT 937.950 169.950 940.050 170.400 ;
        RECT 13.950 168.600 16.050 169.050 ;
        RECT 52.950 168.600 55.050 169.050 ;
        RECT 73.950 168.600 76.050 169.050 ;
        RECT 13.950 167.400 76.050 168.600 ;
        RECT 13.950 166.950 16.050 167.400 ;
        RECT 52.950 166.950 55.050 167.400 ;
        RECT 73.950 166.950 76.050 167.400 ;
        RECT 85.950 168.600 88.050 169.050 ;
        RECT 106.950 168.600 109.050 169.050 ;
        RECT 85.950 167.400 109.050 168.600 ;
        RECT 85.950 166.950 88.050 167.400 ;
        RECT 106.950 166.950 109.050 167.400 ;
        RECT 187.950 168.600 190.050 169.050 ;
        RECT 217.950 168.600 220.050 169.050 ;
        RECT 187.950 167.400 220.050 168.600 ;
        RECT 187.950 166.950 190.050 167.400 ;
        RECT 217.950 166.950 220.050 167.400 ;
        RECT 223.950 168.600 226.050 169.050 ;
        RECT 301.950 168.600 304.050 169.050 ;
        RECT 223.950 167.400 304.050 168.600 ;
        RECT 223.950 166.950 226.050 167.400 ;
        RECT 301.950 166.950 304.050 167.400 ;
        RECT 316.950 168.600 319.050 169.050 ;
        RECT 346.950 168.600 349.050 169.050 ;
        RECT 316.950 167.400 349.050 168.600 ;
        RECT 316.950 166.950 319.050 167.400 ;
        RECT 346.950 166.950 349.050 167.400 ;
        RECT 424.950 168.600 427.050 169.050 ;
        RECT 430.950 168.600 433.050 169.050 ;
        RECT 424.950 167.400 433.050 168.600 ;
        RECT 424.950 166.950 427.050 167.400 ;
        RECT 430.950 166.950 433.050 167.400 ;
        RECT 454.950 168.600 457.050 169.050 ;
        RECT 466.950 168.600 469.050 169.050 ;
        RECT 454.950 167.400 469.050 168.600 ;
        RECT 454.950 166.950 457.050 167.400 ;
        RECT 466.950 166.950 469.050 167.400 ;
        RECT 646.950 168.600 649.050 169.050 ;
        RECT 682.950 168.600 685.050 169.050 ;
        RECT 646.950 167.400 685.050 168.600 ;
        RECT 646.950 166.950 649.050 167.400 ;
        RECT 682.950 166.950 685.050 167.400 ;
        RECT 832.950 168.600 835.050 169.050 ;
        RECT 856.950 168.600 859.050 169.050 ;
        RECT 832.950 167.400 859.050 168.600 ;
        RECT 832.950 166.950 835.050 167.400 ;
        RECT 856.950 166.950 859.050 167.400 ;
        RECT 865.950 168.600 868.050 169.050 ;
        RECT 895.950 168.600 898.050 169.050 ;
        RECT 913.950 168.600 916.050 169.050 ;
        RECT 865.950 167.400 916.050 168.600 ;
        RECT 865.950 166.950 868.050 167.400 ;
        RECT 895.950 166.950 898.050 167.400 ;
        RECT 913.950 166.950 916.050 167.400 ;
        RECT 220.950 165.600 223.050 166.050 ;
        RECT 274.950 165.600 277.050 166.050 ;
        RECT 220.950 164.400 277.050 165.600 ;
        RECT 220.950 163.950 223.050 164.400 ;
        RECT 274.950 163.950 277.050 164.400 ;
        RECT 319.950 165.600 322.050 166.050 ;
        RECT 418.950 165.600 421.050 166.050 ;
        RECT 319.950 164.400 421.050 165.600 ;
        RECT 319.950 163.950 322.050 164.400 ;
        RECT 418.950 163.950 421.050 164.400 ;
        RECT 427.950 165.600 430.050 166.050 ;
        RECT 448.950 165.600 451.050 166.050 ;
        RECT 427.950 164.400 451.050 165.600 ;
        RECT 427.950 163.950 430.050 164.400 ;
        RECT 448.950 163.950 451.050 164.400 ;
        RECT 532.950 165.600 535.050 166.050 ;
        RECT 775.950 165.600 778.050 166.050 ;
        RECT 787.950 165.600 790.050 166.050 ;
        RECT 796.950 165.600 799.050 166.050 ;
        RECT 532.950 164.400 799.050 165.600 ;
        RECT 532.950 163.950 535.050 164.400 ;
        RECT 775.950 163.950 778.050 164.400 ;
        RECT 787.950 163.950 790.050 164.400 ;
        RECT 796.950 163.950 799.050 164.400 ;
        RECT 19.950 162.600 22.050 163.050 ;
        RECT 55.950 162.600 58.050 163.050 ;
        RECT 79.950 162.600 82.050 163.050 ;
        RECT 19.950 161.400 82.050 162.600 ;
        RECT 19.950 160.950 22.050 161.400 ;
        RECT 55.950 160.950 58.050 161.400 ;
        RECT 79.950 160.950 82.050 161.400 ;
        RECT 121.950 162.600 124.050 163.050 ;
        RECT 142.950 162.600 145.050 163.050 ;
        RECT 121.950 161.400 145.050 162.600 ;
        RECT 121.950 160.950 124.050 161.400 ;
        RECT 142.950 160.950 145.050 161.400 ;
        RECT 199.950 162.600 202.050 163.050 ;
        RECT 217.950 162.600 220.050 163.050 ;
        RECT 199.950 161.400 220.050 162.600 ;
        RECT 199.950 160.950 202.050 161.400 ;
        RECT 217.950 160.950 220.050 161.400 ;
        RECT 232.950 162.600 235.050 163.050 ;
        RECT 253.950 162.600 256.050 163.050 ;
        RECT 232.950 161.400 256.050 162.600 ;
        RECT 232.950 160.950 235.050 161.400 ;
        RECT 253.950 160.950 256.050 161.400 ;
        RECT 283.950 162.600 286.050 163.050 ;
        RECT 304.950 162.600 307.050 163.050 ;
        RECT 322.950 162.600 325.050 163.050 ;
        RECT 283.950 161.400 325.050 162.600 ;
        RECT 283.950 160.950 286.050 161.400 ;
        RECT 304.950 160.950 307.050 161.400 ;
        RECT 322.950 160.950 325.050 161.400 ;
        RECT 337.950 162.600 340.050 163.050 ;
        RECT 361.950 162.600 364.050 163.050 ;
        RECT 337.950 161.400 364.050 162.600 ;
        RECT 337.950 160.950 340.050 161.400 ;
        RECT 361.950 160.950 364.050 161.400 ;
        RECT 421.950 162.600 424.050 163.050 ;
        RECT 481.950 162.600 484.050 163.050 ;
        RECT 553.950 162.600 556.050 163.050 ;
        RECT 421.950 161.400 556.050 162.600 ;
        RECT 421.950 160.950 424.050 161.400 ;
        RECT 481.950 160.950 484.050 161.400 ;
        RECT 553.950 160.950 556.050 161.400 ;
        RECT 673.950 162.600 676.050 163.050 ;
        RECT 751.950 162.600 754.050 163.050 ;
        RECT 673.950 161.400 754.050 162.600 ;
        RECT 673.950 160.950 676.050 161.400 ;
        RECT 751.950 160.950 754.050 161.400 ;
        RECT 805.950 162.600 808.050 163.050 ;
        RECT 862.950 162.600 865.050 163.050 ;
        RECT 943.950 162.600 946.050 163.050 ;
        RECT 805.950 161.400 861.600 162.600 ;
        RECT 805.950 160.950 808.050 161.400 ;
        RECT 40.950 159.600 43.050 160.050 ;
        RECT 58.950 159.600 61.050 160.050 ;
        RECT 40.950 158.400 61.050 159.600 ;
        RECT 40.950 157.950 43.050 158.400 ;
        RECT 58.950 157.950 61.050 158.400 ;
        RECT 151.950 159.600 154.050 160.050 ;
        RECT 175.950 159.600 178.050 160.050 ;
        RECT 259.950 159.600 262.050 160.050 ;
        RECT 151.950 158.400 262.050 159.600 ;
        RECT 151.950 157.950 154.050 158.400 ;
        RECT 175.950 157.950 178.050 158.400 ;
        RECT 259.950 157.950 262.050 158.400 ;
        RECT 277.950 159.600 280.050 160.050 ;
        RECT 328.950 159.600 331.050 160.050 ;
        RECT 460.800 159.600 462.900 160.050 ;
        RECT 277.950 158.400 462.900 159.600 ;
        RECT 277.950 157.950 280.050 158.400 ;
        RECT 328.950 157.950 331.050 158.400 ;
        RECT 460.800 157.950 462.900 158.400 ;
        RECT 463.950 159.600 466.050 160.050 ;
        RECT 700.950 159.600 703.050 160.050 ;
        RECT 742.950 159.600 745.050 160.050 ;
        RECT 463.950 158.400 672.600 159.600 ;
        RECT 463.950 157.950 466.050 158.400 ;
        RECT 37.950 156.600 40.050 157.050 ;
        RECT 64.950 156.600 67.050 157.050 ;
        RECT 37.950 155.400 67.050 156.600 ;
        RECT 37.950 154.950 40.050 155.400 ;
        RECT 64.950 154.950 67.050 155.400 ;
        RECT 193.950 156.600 196.050 157.050 ;
        RECT 199.950 156.600 202.050 157.050 ;
        RECT 193.950 155.400 202.050 156.600 ;
        RECT 193.950 154.950 196.050 155.400 ;
        RECT 199.950 154.950 202.050 155.400 ;
        RECT 253.950 156.600 256.050 157.050 ;
        RECT 322.950 156.600 325.050 157.050 ;
        RECT 253.950 155.400 325.050 156.600 ;
        RECT 253.950 154.950 256.050 155.400 ;
        RECT 322.950 154.950 325.050 155.400 ;
        RECT 334.950 156.600 337.050 157.050 ;
        RECT 340.950 156.600 343.050 157.050 ;
        RECT 334.950 155.400 343.050 156.600 ;
        RECT 334.950 154.950 337.050 155.400 ;
        RECT 340.950 154.950 343.050 155.400 ;
        RECT 346.950 156.600 349.050 157.050 ;
        RECT 433.950 156.600 436.050 157.050 ;
        RECT 346.950 155.400 436.050 156.600 ;
        RECT 346.950 154.950 349.050 155.400 ;
        RECT 433.950 154.950 436.050 155.400 ;
        RECT 445.950 156.600 448.050 157.050 ;
        RECT 508.950 156.600 511.050 157.050 ;
        RECT 445.950 155.400 511.050 156.600 ;
        RECT 671.400 156.600 672.600 158.400 ;
        RECT 700.950 158.400 745.050 159.600 ;
        RECT 700.950 157.950 703.050 158.400 ;
        RECT 742.950 157.950 745.050 158.400 ;
        RECT 763.950 159.600 766.050 160.050 ;
        RECT 811.950 159.600 814.050 160.050 ;
        RECT 763.950 158.400 814.050 159.600 ;
        RECT 860.400 159.600 861.600 161.400 ;
        RECT 862.950 161.400 946.050 162.600 ;
        RECT 862.950 160.950 865.050 161.400 ;
        RECT 943.950 160.950 946.050 161.400 ;
        RECT 874.950 159.600 877.050 160.050 ;
        RECT 860.400 158.400 877.050 159.600 ;
        RECT 763.950 157.950 766.050 158.400 ;
        RECT 811.950 157.950 814.050 158.400 ;
        RECT 874.950 157.950 877.050 158.400 ;
        RECT 685.950 156.600 688.050 157.050 ;
        RECT 671.400 155.400 688.050 156.600 ;
        RECT 445.950 154.950 448.050 155.400 ;
        RECT 508.950 154.950 511.050 155.400 ;
        RECT 685.950 154.950 688.050 155.400 ;
        RECT 745.950 156.600 748.050 157.050 ;
        RECT 802.950 156.600 805.050 157.050 ;
        RECT 847.950 156.600 850.050 157.050 ;
        RECT 883.950 156.600 886.050 157.050 ;
        RECT 745.950 155.400 886.050 156.600 ;
        RECT 745.950 154.950 748.050 155.400 ;
        RECT 802.950 154.950 805.050 155.400 ;
        RECT 847.950 154.950 850.050 155.400 ;
        RECT 883.950 154.950 886.050 155.400 ;
        RECT 118.950 153.600 121.050 154.050 ;
        RECT 184.950 153.600 187.050 154.050 ;
        RECT 118.950 152.400 187.050 153.600 ;
        RECT 118.950 151.950 121.050 152.400 ;
        RECT 184.950 151.950 187.050 152.400 ;
        RECT 274.950 153.600 277.050 154.050 ;
        RECT 409.950 153.600 412.050 154.050 ;
        RECT 493.950 153.600 496.050 154.050 ;
        RECT 274.950 152.400 496.050 153.600 ;
        RECT 274.950 151.950 277.050 152.400 ;
        RECT 409.950 151.950 412.050 152.400 ;
        RECT 493.950 151.950 496.050 152.400 ;
        RECT 769.950 153.600 772.050 154.050 ;
        RECT 799.950 153.600 802.050 154.050 ;
        RECT 769.950 152.400 802.050 153.600 ;
        RECT 769.950 151.950 772.050 152.400 ;
        RECT 799.950 151.950 802.050 152.400 ;
        RECT 814.950 153.600 817.050 154.050 ;
        RECT 829.950 153.600 832.050 154.050 ;
        RECT 814.950 152.400 832.050 153.600 ;
        RECT 814.950 151.950 817.050 152.400 ;
        RECT 829.950 151.950 832.050 152.400 ;
        RECT 898.950 153.600 901.050 154.050 ;
        RECT 937.950 153.600 940.050 154.050 ;
        RECT 898.950 152.400 940.050 153.600 ;
        RECT 898.950 151.950 901.050 152.400 ;
        RECT 937.950 151.950 940.050 152.400 ;
        RECT 91.950 150.600 94.050 151.050 ;
        RECT 97.950 150.600 100.050 151.050 ;
        RECT 91.950 149.400 100.050 150.600 ;
        RECT 91.950 148.950 94.050 149.400 ;
        RECT 97.950 148.950 100.050 149.400 ;
        RECT 202.950 150.600 205.050 151.050 ;
        RECT 223.950 150.600 226.050 151.050 ;
        RECT 202.950 149.400 226.050 150.600 ;
        RECT 202.950 148.950 205.050 149.400 ;
        RECT 223.950 148.950 226.050 149.400 ;
        RECT 244.950 150.600 247.050 151.050 ;
        RECT 268.950 150.600 271.050 151.050 ;
        RECT 244.950 149.400 271.050 150.600 ;
        RECT 244.950 148.950 247.050 149.400 ;
        RECT 268.950 148.950 271.050 149.400 ;
        RECT 340.950 150.600 343.050 151.050 ;
        RECT 358.800 150.600 360.900 151.050 ;
        RECT 340.950 149.400 360.900 150.600 ;
        RECT 340.950 148.950 343.050 149.400 ;
        RECT 358.800 148.950 360.900 149.400 ;
        RECT 361.950 150.600 364.050 151.050 ;
        RECT 463.950 150.600 466.050 151.050 ;
        RECT 361.950 149.400 466.050 150.600 ;
        RECT 361.950 148.950 364.050 149.400 ;
        RECT 463.950 148.950 466.050 149.400 ;
        RECT 478.950 150.600 481.050 151.050 ;
        RECT 538.950 150.600 541.050 151.050 ;
        RECT 478.950 149.400 541.050 150.600 ;
        RECT 478.950 148.950 481.050 149.400 ;
        RECT 538.950 148.950 541.050 149.400 ;
        RECT 556.950 150.600 559.050 151.050 ;
        RECT 589.950 150.600 592.050 151.050 ;
        RECT 556.950 149.400 592.050 150.600 ;
        RECT 556.950 148.950 559.050 149.400 ;
        RECT 589.950 148.950 592.050 149.400 ;
        RECT 625.950 150.600 628.050 151.050 ;
        RECT 643.950 150.600 646.050 151.050 ;
        RECT 625.950 149.400 646.050 150.600 ;
        RECT 625.950 148.950 628.050 149.400 ;
        RECT 643.950 148.950 646.050 149.400 ;
        RECT 670.950 150.600 673.050 151.050 ;
        RECT 703.950 150.600 706.050 151.050 ;
        RECT 670.950 149.400 706.050 150.600 ;
        RECT 670.950 148.950 673.050 149.400 ;
        RECT 703.950 148.950 706.050 149.400 ;
        RECT 712.950 150.600 715.050 151.050 ;
        RECT 787.950 150.600 790.050 151.050 ;
        RECT 808.950 150.600 811.050 151.050 ;
        RECT 832.950 150.600 835.050 151.050 ;
        RECT 712.950 149.400 835.050 150.600 ;
        RECT 712.950 148.950 715.050 149.400 ;
        RECT 787.950 148.950 790.050 149.400 ;
        RECT 808.950 148.950 811.050 149.400 ;
        RECT 832.950 148.950 835.050 149.400 ;
        RECT 907.950 150.600 910.050 151.050 ;
        RECT 946.950 150.600 949.050 151.050 ;
        RECT 907.950 149.400 949.050 150.600 ;
        RECT 907.950 148.950 910.050 149.400 ;
        RECT 946.950 148.950 949.050 149.400 ;
        RECT 34.950 147.600 37.050 148.050 ;
        RECT 76.950 147.600 79.050 148.050 ;
        RECT 106.950 147.600 109.050 148.050 ;
        RECT 34.950 146.400 109.050 147.600 ;
        RECT 34.950 145.950 37.050 146.400 ;
        RECT 76.950 145.950 79.050 146.400 ;
        RECT 106.950 145.950 109.050 146.400 ;
        RECT 124.950 147.600 127.050 148.050 ;
        RECT 187.950 147.600 190.050 148.050 ;
        RECT 124.950 146.400 190.050 147.600 ;
        RECT 124.950 145.950 127.050 146.400 ;
        RECT 187.950 145.950 190.050 146.400 ;
        RECT 196.950 147.600 199.050 148.050 ;
        RECT 208.950 147.600 211.050 148.050 ;
        RECT 436.950 147.600 439.050 148.050 ;
        RECT 688.950 147.600 691.050 148.050 ;
        RECT 706.950 147.600 709.050 148.050 ;
        RECT 196.950 146.400 231.600 147.600 ;
        RECT 196.950 145.950 199.050 146.400 ;
        RECT 208.950 145.950 211.050 146.400 ;
        RECT 230.400 145.050 231.600 146.400 ;
        RECT 436.950 146.400 709.050 147.600 ;
        RECT 436.950 145.950 439.050 146.400 ;
        RECT 688.950 145.950 691.050 146.400 ;
        RECT 706.950 145.950 709.050 146.400 ;
        RECT 727.950 147.600 730.050 148.050 ;
        RECT 781.950 147.600 784.050 148.050 ;
        RECT 814.950 147.600 817.050 148.050 ;
        RECT 838.950 147.600 841.050 148.050 ;
        RECT 727.950 146.400 841.050 147.600 ;
        RECT 727.950 145.950 730.050 146.400 ;
        RECT 781.950 145.950 784.050 146.400 ;
        RECT 814.950 145.950 817.050 146.400 ;
        RECT 838.950 145.950 841.050 146.400 ;
        RECT 112.950 144.600 115.050 145.050 ;
        RECT 118.950 144.600 121.050 145.050 ;
        RECT 130.950 144.600 133.050 145.050 ;
        RECT 112.950 143.400 133.050 144.600 ;
        RECT 112.950 142.950 115.050 143.400 ;
        RECT 118.950 142.950 121.050 143.400 ;
        RECT 130.950 142.950 133.050 143.400 ;
        RECT 229.950 144.600 232.050 145.050 ;
        RECT 244.950 144.600 247.050 145.050 ;
        RECT 229.950 143.400 247.050 144.600 ;
        RECT 229.950 142.950 232.050 143.400 ;
        RECT 244.950 142.950 247.050 143.400 ;
        RECT 277.950 144.600 280.050 145.050 ;
        RECT 307.950 144.600 310.050 145.050 ;
        RECT 277.950 143.400 310.050 144.600 ;
        RECT 277.950 142.950 280.050 143.400 ;
        RECT 307.950 142.950 310.050 143.400 ;
        RECT 319.950 144.600 322.050 145.050 ;
        RECT 367.950 144.600 370.050 145.050 ;
        RECT 319.950 143.400 370.050 144.600 ;
        RECT 319.950 142.950 322.050 143.400 ;
        RECT 367.950 142.950 370.050 143.400 ;
        RECT 415.950 144.600 418.050 145.050 ;
        RECT 421.950 144.600 424.050 145.050 ;
        RECT 415.950 143.400 424.050 144.600 ;
        RECT 415.950 142.950 418.050 143.400 ;
        RECT 421.950 142.950 424.050 143.400 ;
        RECT 475.950 144.600 478.050 145.050 ;
        RECT 502.950 144.600 505.050 145.050 ;
        RECT 475.950 143.400 505.050 144.600 ;
        RECT 475.950 142.950 478.050 143.400 ;
        RECT 502.950 142.950 505.050 143.400 ;
        RECT 559.950 144.600 562.050 145.050 ;
        RECT 586.950 144.600 589.050 145.050 ;
        RECT 595.950 144.600 598.050 145.050 ;
        RECT 559.950 143.400 598.050 144.600 ;
        RECT 559.950 142.950 562.050 143.400 ;
        RECT 586.950 142.950 589.050 143.400 ;
        RECT 595.950 142.950 598.050 143.400 ;
        RECT 784.950 144.600 787.050 145.050 ;
        RECT 805.950 144.600 808.050 145.050 ;
        RECT 784.950 143.400 808.050 144.600 ;
        RECT 784.950 142.950 787.050 143.400 ;
        RECT 805.950 142.950 808.050 143.400 ;
        RECT 841.950 144.600 844.050 145.050 ;
        RECT 847.950 144.600 850.050 145.050 ;
        RECT 841.950 143.400 850.050 144.600 ;
        RECT 841.950 142.950 844.050 143.400 ;
        RECT 847.950 142.950 850.050 143.400 ;
        RECT 877.950 144.600 880.050 145.050 ;
        RECT 886.950 144.600 889.050 145.050 ;
        RECT 919.950 144.600 922.050 145.050 ;
        RECT 877.950 143.400 922.050 144.600 ;
        RECT 877.950 142.950 880.050 143.400 ;
        RECT 886.950 142.950 889.050 143.400 ;
        RECT 919.950 142.950 922.050 143.400 ;
        RECT 94.950 141.600 97.050 142.050 ;
        RECT 145.950 141.600 148.050 142.050 ;
        RECT 94.950 140.400 148.050 141.600 ;
        RECT 94.950 139.950 97.050 140.400 ;
        RECT 145.950 139.950 148.050 140.400 ;
        RECT 7.950 138.750 10.050 139.200 ;
        RECT 13.950 138.750 16.050 139.200 ;
        RECT 7.950 137.550 16.050 138.750 ;
        RECT 7.950 137.100 10.050 137.550 ;
        RECT 13.950 137.100 16.050 137.550 ;
        RECT 19.950 138.600 22.050 139.200 ;
        RECT 31.950 138.750 34.050 139.200 ;
        RECT 37.950 138.750 40.050 139.200 ;
        RECT 31.950 138.600 40.050 138.750 ;
        RECT 49.950 138.600 52.050 139.050 ;
        RECT 70.950 138.600 73.050 139.200 ;
        RECT 19.950 137.550 40.050 138.600 ;
        RECT 19.950 137.400 34.050 137.550 ;
        RECT 19.950 137.100 22.050 137.400 ;
        RECT 31.950 137.100 34.050 137.400 ;
        RECT 37.950 137.100 40.050 137.550 ;
        RECT 47.400 137.400 73.050 138.600 ;
        RECT 16.950 132.600 19.050 132.900 ;
        RECT 40.950 132.600 43.050 132.900 ;
        RECT 16.950 131.400 43.050 132.600 ;
        RECT 16.950 130.800 19.050 131.400 ;
        RECT 40.950 130.800 43.050 131.400 ;
        RECT 47.400 130.050 48.600 137.400 ;
        RECT 49.950 136.950 52.050 137.400 ;
        RECT 70.950 137.100 73.050 137.400 ;
        RECT 112.950 138.600 115.050 139.200 ;
        RECT 124.950 138.600 127.050 139.200 ;
        RECT 151.950 138.600 154.050 142.050 ;
        RECT 172.950 141.600 175.050 142.050 ;
        RECT 202.950 141.600 205.050 142.050 ;
        RECT 172.950 140.400 205.050 141.600 ;
        RECT 172.950 139.950 175.050 140.400 ;
        RECT 202.950 139.950 205.050 140.400 ;
        RECT 211.950 141.600 214.050 142.050 ;
        RECT 250.950 141.600 253.050 142.050 ;
        RECT 211.950 140.400 253.050 141.600 ;
        RECT 211.950 139.950 214.050 140.400 ;
        RECT 250.950 139.950 253.050 140.400 ;
        RECT 256.950 139.950 259.050 142.050 ;
        RECT 274.950 141.600 277.050 142.050 ;
        RECT 313.950 141.600 316.050 142.200 ;
        RECT 274.950 140.400 316.050 141.600 ;
        RECT 274.950 139.950 277.050 140.400 ;
        RECT 313.950 140.100 316.050 140.400 ;
        RECT 427.950 141.600 430.050 142.050 ;
        RECT 529.950 141.600 532.050 142.050 ;
        RECT 547.950 141.600 550.050 142.050 ;
        RECT 427.950 140.400 550.050 141.600 ;
        RECT 427.950 139.950 430.050 140.400 ;
        RECT 529.950 139.950 532.050 140.400 ;
        RECT 547.950 139.950 550.050 140.400 ;
        RECT 622.950 141.600 625.050 142.050 ;
        RECT 637.950 141.600 640.050 142.050 ;
        RECT 622.950 140.400 640.050 141.600 ;
        RECT 622.950 139.950 625.050 140.400 ;
        RECT 637.950 139.950 640.050 140.400 ;
        RECT 823.950 141.600 826.050 142.050 ;
        RECT 850.950 141.600 853.050 142.050 ;
        RECT 865.950 141.600 868.050 142.050 ;
        RECT 823.950 140.400 868.050 141.600 ;
        RECT 823.950 139.950 826.050 140.400 ;
        RECT 850.950 139.950 853.050 140.400 ;
        RECT 865.950 139.950 868.050 140.400 ;
        RECT 112.950 137.400 127.050 138.600 ;
        RECT 112.950 137.100 115.050 137.400 ;
        RECT 124.950 137.100 127.050 137.400 ;
        RECT 149.400 138.000 154.050 138.600 ;
        RECT 154.950 138.750 157.050 139.200 ;
        RECT 166.950 138.750 169.050 139.200 ;
        RECT 149.400 137.400 153.600 138.000 ;
        RECT 154.950 137.550 169.050 138.750 ;
        RECT 52.950 132.600 55.050 133.050 ;
        RECT 67.950 132.600 70.050 132.900 ;
        RECT 52.950 131.400 70.050 132.600 ;
        RECT 52.950 130.950 55.050 131.400 ;
        RECT 67.950 130.800 70.050 131.400 ;
        RECT 109.950 132.600 112.050 132.900 ;
        RECT 127.950 132.600 130.050 132.900 ;
        RECT 109.950 131.400 130.050 132.600 ;
        RECT 109.950 130.800 112.050 131.400 ;
        RECT 127.950 130.800 130.050 131.400 ;
        RECT 133.950 132.600 136.050 132.900 ;
        RECT 139.950 132.600 142.050 133.050 ;
        RECT 149.400 132.900 150.600 137.400 ;
        RECT 154.950 137.100 157.050 137.550 ;
        RECT 166.950 137.100 169.050 137.550 ;
        RECT 217.950 137.100 220.050 139.200 ;
        RECT 202.950 135.600 205.050 136.050 ;
        RECT 218.400 135.600 219.600 137.100 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 238.950 137.100 241.050 139.200 ;
        RECT 226.950 135.600 229.050 136.050 ;
        RECT 202.950 134.400 229.050 135.600 ;
        RECT 202.950 133.950 205.050 134.400 ;
        RECT 226.950 133.950 229.050 134.400 ;
        RECT 133.950 131.400 142.050 132.600 ;
        RECT 133.950 130.800 136.050 131.400 ;
        RECT 139.950 130.950 142.050 131.400 ;
        RECT 148.950 130.800 151.050 132.900 ;
        RECT 157.950 132.600 160.050 133.050 ;
        RECT 181.950 132.600 184.050 133.050 ;
        RECT 190.950 132.600 193.050 132.900 ;
        RECT 157.950 131.400 193.050 132.600 ;
        RECT 157.950 130.950 160.050 131.400 ;
        RECT 181.950 130.950 184.050 131.400 ;
        RECT 190.950 130.800 193.050 131.400 ;
        RECT 220.950 132.600 223.050 132.900 ;
        RECT 233.400 132.600 234.600 136.950 ;
        RECT 220.950 131.400 234.600 132.600 ;
        RECT 220.950 130.800 223.050 131.400 ;
        RECT 239.400 130.050 240.600 137.100 ;
        RECT 247.950 136.950 250.050 139.050 ;
        RECT 241.950 132.600 244.050 132.900 ;
        RECT 248.400 132.600 249.600 136.950 ;
        RECT 257.400 135.600 258.600 139.950 ;
        RECT 298.950 138.600 301.050 139.050 ;
        RECT 313.950 138.600 316.050 139.050 ;
        RECT 331.950 138.600 334.050 139.200 ;
        RECT 336.000 138.600 340.050 139.050 ;
        RECT 298.950 137.400 334.050 138.600 ;
        RECT 298.950 136.950 301.050 137.400 ;
        RECT 313.950 136.950 316.050 137.400 ;
        RECT 331.950 137.100 334.050 137.400 ;
        RECT 335.400 136.950 340.050 138.600 ;
        RECT 352.950 138.750 355.050 139.200 ;
        RECT 364.950 138.750 367.050 139.200 ;
        RECT 352.950 137.550 367.050 138.750 ;
        RECT 352.950 137.100 355.050 137.550 ;
        RECT 364.950 137.100 367.050 137.550 ;
        RECT 373.950 138.600 376.050 139.200 ;
        RECT 382.950 138.750 385.050 139.200 ;
        RECT 391.950 138.750 394.050 139.200 ;
        RECT 373.950 137.400 381.600 138.600 ;
        RECT 373.950 137.100 376.050 137.400 ;
        RECT 335.400 135.600 336.600 136.950 ;
        RECT 257.400 134.400 264.600 135.600 ;
        RECT 326.400 135.000 336.600 135.600 ;
        RECT 241.950 131.400 249.600 132.600 ;
        RECT 250.950 132.450 253.050 132.900 ;
        RECT 259.950 132.450 262.050 132.900 ;
        RECT 241.950 130.800 244.050 131.400 ;
        RECT 250.950 131.250 262.050 132.450 ;
        RECT 263.400 132.600 264.600 134.400 ;
        RECT 325.950 134.400 336.600 135.000 ;
        RECT 380.400 135.600 381.600 137.400 ;
        RECT 382.950 137.550 394.050 138.750 ;
        RECT 382.950 137.100 385.050 137.550 ;
        RECT 391.950 137.100 394.050 137.550 ;
        RECT 433.950 138.600 436.050 139.050 ;
        RECT 469.950 138.600 472.050 139.050 ;
        RECT 475.950 138.600 478.050 139.050 ;
        RECT 496.950 138.600 499.050 139.200 ;
        RECT 433.950 137.400 499.050 138.600 ;
        RECT 433.950 136.950 436.050 137.400 ;
        RECT 469.950 136.950 472.050 137.400 ;
        RECT 475.950 136.950 478.050 137.400 ;
        RECT 496.950 137.100 499.050 137.400 ;
        RECT 502.950 138.600 505.050 139.200 ;
        RECT 523.950 138.600 526.050 139.200 ;
        RECT 502.950 137.400 526.050 138.600 ;
        RECT 502.950 137.100 505.050 137.400 ;
        RECT 523.950 137.100 526.050 137.400 ;
        RECT 553.950 138.600 556.050 139.200 ;
        RECT 568.950 138.600 571.050 139.200 ;
        RECT 553.950 137.400 571.050 138.600 ;
        RECT 553.950 137.100 556.050 137.400 ;
        RECT 568.950 137.100 571.050 137.400 ;
        RECT 574.950 138.600 577.050 139.200 ;
        RECT 583.950 138.600 586.050 139.050 ;
        RECT 613.950 138.750 616.050 139.200 ;
        RECT 619.950 138.750 622.050 139.200 ;
        RECT 613.950 138.600 622.050 138.750 ;
        RECT 649.950 138.600 652.050 139.200 ;
        RECT 574.950 137.400 582.600 138.600 ;
        RECT 574.950 137.100 577.050 137.400 ;
        RECT 581.400 135.600 582.600 137.400 ;
        RECT 583.950 137.400 600.600 138.600 ;
        RECT 583.950 136.950 586.050 137.400 ;
        RECT 380.400 134.400 399.600 135.600 ;
        RECT 581.400 135.000 594.600 135.600 ;
        RECT 581.400 134.400 595.050 135.000 ;
        RECT 265.950 132.600 268.050 132.900 ;
        RECT 263.400 131.400 268.050 132.600 ;
        RECT 250.950 130.800 253.050 131.250 ;
        RECT 259.950 130.800 262.050 131.250 ;
        RECT 265.950 130.800 268.050 131.400 ;
        RECT 304.950 132.600 307.050 133.050 ;
        RECT 319.950 132.600 322.050 133.050 ;
        RECT 304.950 131.400 322.050 132.600 ;
        RECT 304.950 130.950 307.050 131.400 ;
        RECT 319.950 130.950 322.050 131.400 ;
        RECT 325.950 130.950 328.050 134.400 ;
        RECT 398.400 132.900 399.600 134.400 ;
        RECT 397.950 130.800 400.050 132.900 ;
        RECT 418.950 132.450 421.050 132.900 ;
        RECT 427.950 132.450 430.050 132.900 ;
        RECT 418.950 131.250 430.050 132.450 ;
        RECT 418.950 130.800 421.050 131.250 ;
        RECT 427.950 130.800 430.050 131.250 ;
        RECT 448.950 132.450 451.050 132.900 ;
        RECT 478.950 132.600 481.050 132.900 ;
        RECT 499.950 132.600 502.050 132.900 ;
        RECT 478.950 132.450 502.050 132.600 ;
        RECT 448.950 131.400 502.050 132.450 ;
        RECT 448.950 131.250 481.050 131.400 ;
        RECT 448.950 130.800 451.050 131.250 ;
        RECT 478.950 130.800 481.050 131.250 ;
        RECT 499.950 130.800 502.050 131.400 ;
        RECT 514.950 132.450 517.050 132.900 ;
        RECT 520.950 132.600 523.050 132.900 ;
        RECT 544.950 132.600 547.050 132.900 ;
        RECT 520.950 132.450 547.050 132.600 ;
        RECT 514.950 131.400 547.050 132.450 ;
        RECT 514.950 131.250 523.050 131.400 ;
        RECT 514.950 130.800 517.050 131.250 ;
        RECT 520.950 130.800 523.050 131.250 ;
        RECT 544.950 130.800 547.050 131.400 ;
        RECT 577.950 132.450 580.050 132.900 ;
        RECT 586.950 132.450 589.050 132.900 ;
        RECT 577.950 131.250 589.050 132.450 ;
        RECT 577.950 130.800 580.050 131.250 ;
        RECT 586.950 130.800 589.050 131.250 ;
        RECT 592.950 130.950 595.050 134.400 ;
        RECT 599.400 132.900 600.600 137.400 ;
        RECT 613.950 137.550 652.050 138.600 ;
        RECT 613.950 137.100 616.050 137.550 ;
        RECT 619.950 137.400 652.050 137.550 ;
        RECT 619.950 137.100 622.050 137.400 ;
        RECT 649.950 137.100 652.050 137.400 ;
        RECT 658.950 138.750 661.050 139.200 ;
        RECT 667.950 138.750 670.050 139.200 ;
        RECT 658.950 137.550 670.050 138.750 ;
        RECT 658.950 137.100 661.050 137.550 ;
        RECT 667.950 137.100 670.050 137.550 ;
        RECT 673.950 137.100 676.050 139.200 ;
        RECT 694.950 138.600 697.050 139.200 ;
        RECT 715.950 138.600 718.050 139.200 ;
        RECT 694.950 137.400 718.050 138.600 ;
        RECT 694.950 137.100 697.050 137.400 ;
        RECT 715.950 137.100 718.050 137.400 ;
        RECT 721.950 138.600 724.050 139.200 ;
        RECT 736.950 138.600 739.050 139.200 ;
        RECT 757.950 138.600 760.050 139.200 ;
        RECT 769.950 138.600 772.050 139.200 ;
        RECT 774.000 138.600 778.050 139.050 ;
        RECT 721.950 137.400 741.600 138.600 ;
        RECT 721.950 137.100 724.050 137.400 ;
        RECT 736.950 137.100 739.050 137.400 ;
        RECT 661.950 135.600 664.050 136.050 ;
        RECT 674.400 135.600 675.600 137.100 ;
        RECT 661.950 134.400 675.600 135.600 ;
        RECT 661.950 133.950 664.050 134.400 ;
        RECT 740.400 133.050 741.600 137.400 ;
        RECT 757.950 137.400 772.050 138.600 ;
        RECT 757.950 137.100 760.050 137.400 ;
        RECT 769.950 137.100 772.050 137.400 ;
        RECT 773.400 136.950 778.050 138.600 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 793.950 137.100 796.050 139.200 ;
        RECT 799.950 138.600 802.050 139.050 ;
        RECT 829.950 138.600 832.050 139.050 ;
        RECT 799.950 137.400 810.600 138.600 ;
        RECT 598.950 130.800 601.050 132.900 ;
        RECT 622.950 132.600 625.050 132.900 ;
        RECT 637.950 132.600 640.050 132.900 ;
        RECT 622.950 132.450 640.050 132.600 ;
        RECT 646.950 132.450 649.050 132.900 ;
        RECT 622.950 131.400 649.050 132.450 ;
        RECT 622.950 130.800 625.050 131.400 ;
        RECT 637.950 131.250 649.050 131.400 ;
        RECT 637.950 130.800 640.050 131.250 ;
        RECT 646.950 130.800 649.050 131.250 ;
        RECT 46.950 127.950 49.050 130.050 ;
        RECT 199.950 129.600 202.050 130.050 ;
        RECT 211.950 129.600 214.050 130.050 ;
        RECT 199.950 128.400 214.050 129.600 ;
        RECT 199.950 127.950 202.050 128.400 ;
        RECT 211.950 127.950 214.050 128.400 ;
        RECT 238.950 127.950 241.050 130.050 ;
        RECT 343.950 129.600 346.050 130.050 ;
        RECT 349.950 129.600 352.050 130.050 ;
        RECT 343.950 128.400 352.050 129.600 ;
        RECT 343.950 127.950 346.050 128.400 ;
        RECT 349.950 127.950 352.050 128.400 ;
        RECT 370.950 129.600 373.050 130.050 ;
        RECT 391.950 129.600 394.050 130.050 ;
        RECT 370.950 128.400 394.050 129.600 ;
        RECT 370.950 127.950 373.050 128.400 ;
        RECT 391.950 127.950 394.050 128.400 ;
        RECT 430.950 129.600 433.050 130.050 ;
        RECT 436.950 129.600 439.050 130.050 ;
        RECT 568.950 129.600 571.050 130.050 ;
        RECT 430.950 128.400 439.050 129.600 ;
        RECT 430.950 127.950 433.050 128.400 ;
        RECT 436.950 127.950 439.050 128.400 ;
        RECT 467.400 128.400 571.050 129.600 ;
        RECT 223.950 126.600 226.050 127.050 ;
        RECT 164.400 125.400 226.050 126.600 ;
        RECT 164.400 124.050 165.600 125.400 ;
        RECT 223.950 124.950 226.050 125.400 ;
        RECT 271.950 126.600 274.050 127.050 ;
        RECT 325.950 126.600 328.050 127.050 ;
        RECT 271.950 125.400 328.050 126.600 ;
        RECT 271.950 124.950 274.050 125.400 ;
        RECT 325.950 124.950 328.050 125.400 ;
        RECT 367.950 126.600 370.050 127.050 ;
        RECT 467.400 126.600 468.600 128.400 ;
        RECT 568.950 127.950 571.050 128.400 ;
        RECT 631.950 129.600 634.050 130.050 ;
        RECT 655.950 129.600 658.050 133.050 ;
        RECT 682.950 132.450 685.050 132.900 ;
        RECT 697.950 132.600 700.050 132.900 ;
        RECT 712.950 132.600 715.050 132.900 ;
        RECT 697.950 132.450 715.050 132.600 ;
        RECT 682.950 131.400 715.050 132.450 ;
        RECT 682.950 131.250 700.050 131.400 ;
        RECT 682.950 130.800 685.050 131.250 ;
        RECT 697.950 130.800 700.050 131.250 ;
        RECT 712.950 130.800 715.050 131.400 ;
        RECT 739.950 130.950 742.050 133.050 ;
        RECT 773.400 132.900 774.600 136.950 ;
        RECT 785.400 133.050 786.600 136.950 ;
        RECT 754.950 132.450 757.050 132.900 ;
        RECT 763.950 132.450 766.050 132.900 ;
        RECT 754.950 131.250 766.050 132.450 ;
        RECT 754.950 130.800 757.050 131.250 ;
        RECT 763.950 130.800 766.050 131.250 ;
        RECT 772.950 130.800 775.050 132.900 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 794.400 132.600 795.600 137.100 ;
        RECT 799.950 136.950 802.050 137.400 ;
        RECT 799.950 132.600 802.050 133.050 ;
        RECT 794.400 131.400 802.050 132.600 ;
        RECT 809.400 132.600 810.600 137.400 ;
        RECT 829.950 137.400 843.600 138.600 ;
        RECT 829.950 136.950 832.050 137.400 ;
        RECT 811.950 132.600 814.050 132.900 ;
        RECT 809.400 131.400 814.050 132.600 ;
        RECT 799.950 130.950 802.050 131.400 ;
        RECT 811.950 130.800 814.050 131.400 ;
        RECT 817.950 132.600 820.050 132.900 ;
        RECT 823.950 132.600 826.050 133.050 ;
        RECT 817.950 131.400 826.050 132.600 ;
        RECT 817.950 130.800 820.050 131.400 ;
        RECT 823.950 130.950 826.050 131.400 ;
        RECT 842.400 130.050 843.600 137.400 ;
        RECT 853.950 136.950 856.050 139.050 ;
        RECT 877.950 136.950 880.050 139.050 ;
        RECT 889.950 137.100 892.050 139.200 ;
        RECT 895.950 138.750 898.050 139.200 ;
        RECT 904.950 138.750 907.050 139.200 ;
        RECT 895.950 137.550 907.050 138.750 ;
        RECT 931.950 138.600 934.050 139.200 ;
        RECT 895.950 137.100 898.050 137.550 ;
        RECT 904.950 137.100 907.050 137.550 ;
        RECT 914.400 137.400 934.050 138.600 ;
        RECT 854.400 133.050 855.600 136.950 ;
        RECT 853.950 130.950 856.050 133.050 ;
        RECT 631.950 129.000 658.050 129.600 ;
        RECT 631.950 128.400 657.600 129.000 ;
        RECT 631.950 127.950 634.050 128.400 ;
        RECT 841.950 127.950 844.050 130.050 ;
        RECT 862.950 129.600 865.050 130.050 ;
        RECT 878.400 129.600 879.600 136.950 ;
        RECT 890.400 133.050 891.600 137.100 ;
        RECT 890.400 131.400 895.050 133.050 ;
        RECT 914.400 132.900 915.600 137.400 ;
        RECT 931.950 137.100 934.050 137.400 ;
        RECT 943.950 138.600 946.050 139.050 ;
        RECT 943.950 137.400 951.600 138.600 ;
        RECT 943.950 136.950 946.050 137.400 ;
        RECT 891.000 130.950 895.050 131.400 ;
        RECT 901.950 132.450 904.050 132.900 ;
        RECT 907.950 132.450 910.050 132.900 ;
        RECT 901.950 131.250 910.050 132.450 ;
        RECT 901.950 130.800 904.050 131.250 ;
        RECT 907.950 130.800 910.050 131.250 ;
        RECT 913.950 130.800 916.050 132.900 ;
        RECT 940.950 132.600 943.050 132.900 ;
        RECT 946.950 132.600 949.050 133.050 ;
        RECT 940.950 131.400 949.050 132.600 ;
        RECT 940.950 130.800 943.050 131.400 ;
        RECT 946.950 130.950 949.050 131.400 ;
        RECT 862.950 128.400 879.600 129.600 ;
        RECT 922.950 129.600 925.050 130.050 ;
        RECT 931.950 129.600 934.050 130.050 ;
        RECT 922.950 128.400 934.050 129.600 ;
        RECT 862.950 127.950 865.050 128.400 ;
        RECT 922.950 127.950 925.050 128.400 ;
        RECT 931.950 127.950 934.050 128.400 ;
        RECT 943.950 129.600 946.050 130.050 ;
        RECT 950.400 129.600 951.600 137.400 ;
        RECT 943.950 128.400 951.600 129.600 ;
        RECT 943.950 127.950 946.050 128.400 ;
        RECT 367.950 125.400 468.600 126.600 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 475.950 126.600 478.050 127.050 ;
        RECT 469.950 125.400 478.050 126.600 ;
        RECT 367.950 124.950 370.050 125.400 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 505.950 126.600 508.050 127.050 ;
        RECT 550.950 126.600 553.050 127.050 ;
        RECT 613.950 126.600 616.050 127.050 ;
        RECT 505.950 125.400 549.600 126.600 ;
        RECT 505.950 124.950 508.050 125.400 ;
        RECT 7.950 123.600 10.050 124.050 ;
        RECT 28.950 123.600 31.050 124.050 ;
        RECT 61.950 123.600 64.050 124.050 ;
        RECT 7.950 122.400 64.050 123.600 ;
        RECT 7.950 121.950 10.050 122.400 ;
        RECT 28.950 121.950 31.050 122.400 ;
        RECT 61.950 121.950 64.050 122.400 ;
        RECT 88.950 123.600 91.050 124.050 ;
        RECT 106.950 123.600 109.050 124.050 ;
        RECT 163.950 123.600 166.050 124.050 ;
        RECT 88.950 122.400 166.050 123.600 ;
        RECT 88.950 121.950 91.050 122.400 ;
        RECT 106.950 121.950 109.050 122.400 ;
        RECT 163.950 121.950 166.050 122.400 ;
        RECT 229.950 123.600 232.050 124.050 ;
        RECT 265.950 123.600 268.050 124.050 ;
        RECT 229.950 122.400 268.050 123.600 ;
        RECT 229.950 121.950 232.050 122.400 ;
        RECT 265.950 121.950 268.050 122.400 ;
        RECT 283.950 123.600 286.050 124.050 ;
        RECT 343.950 123.600 346.050 124.050 ;
        RECT 283.950 122.400 346.050 123.600 ;
        RECT 283.950 121.950 286.050 122.400 ;
        RECT 343.950 121.950 346.050 122.400 ;
        RECT 385.950 123.600 388.050 124.050 ;
        RECT 460.800 123.600 462.900 124.050 ;
        RECT 385.950 122.400 462.900 123.600 ;
        RECT 385.950 121.950 388.050 122.400 ;
        RECT 460.800 121.950 462.900 122.400 ;
        RECT 463.950 123.600 466.050 124.050 ;
        RECT 511.950 123.600 514.050 124.050 ;
        RECT 463.950 122.400 514.050 123.600 ;
        RECT 548.400 123.600 549.600 125.400 ;
        RECT 550.950 125.400 616.050 126.600 ;
        RECT 550.950 124.950 553.050 125.400 ;
        RECT 613.950 124.950 616.050 125.400 ;
        RECT 628.950 126.600 631.050 127.050 ;
        RECT 658.950 126.600 661.050 127.050 ;
        RECT 628.950 125.400 661.050 126.600 ;
        RECT 628.950 124.950 631.050 125.400 ;
        RECT 658.950 124.950 661.050 125.400 ;
        RECT 667.950 126.600 670.050 127.050 ;
        RECT 688.950 126.600 691.050 127.050 ;
        RECT 667.950 125.400 691.050 126.600 ;
        RECT 667.950 124.950 670.050 125.400 ;
        RECT 688.950 124.950 691.050 125.400 ;
        RECT 712.950 126.600 715.050 127.050 ;
        RECT 727.950 126.600 730.050 127.050 ;
        RECT 712.950 125.400 730.050 126.600 ;
        RECT 712.950 124.950 715.050 125.400 ;
        RECT 727.950 124.950 730.050 125.400 ;
        RECT 733.950 126.600 736.050 127.050 ;
        RECT 748.950 126.600 751.050 127.050 ;
        RECT 733.950 125.400 751.050 126.600 ;
        RECT 733.950 124.950 736.050 125.400 ;
        RECT 748.950 124.950 751.050 125.400 ;
        RECT 820.950 126.600 823.050 127.050 ;
        RECT 856.950 126.600 859.050 127.050 ;
        RECT 820.950 125.400 859.050 126.600 ;
        RECT 820.950 124.950 823.050 125.400 ;
        RECT 856.950 124.950 859.050 125.400 ;
        RECT 925.950 126.600 928.050 127.050 ;
        RECT 934.950 126.600 937.050 127.050 ;
        RECT 925.950 125.400 937.050 126.600 ;
        RECT 925.950 124.950 928.050 125.400 ;
        RECT 934.950 124.950 937.050 125.400 ;
        RECT 583.950 123.600 586.050 124.050 ;
        RECT 548.400 122.400 586.050 123.600 ;
        RECT 463.950 121.950 466.050 122.400 ;
        RECT 511.950 121.950 514.050 122.400 ;
        RECT 583.950 121.950 586.050 122.400 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 799.950 123.600 802.050 124.050 ;
        RECT 676.950 122.400 802.050 123.600 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 799.950 121.950 802.050 122.400 ;
        RECT 805.950 123.600 808.050 124.050 ;
        RECT 811.950 123.600 814.050 124.050 ;
        RECT 835.950 123.600 838.050 124.050 ;
        RECT 805.950 122.400 838.050 123.600 ;
        RECT 805.950 121.950 808.050 122.400 ;
        RECT 811.950 121.950 814.050 122.400 ;
        RECT 835.950 121.950 838.050 122.400 ;
        RECT 844.950 123.600 847.050 124.050 ;
        RECT 880.950 123.600 883.050 124.050 ;
        RECT 886.950 123.600 889.050 124.050 ;
        RECT 844.950 122.400 889.050 123.600 ;
        RECT 844.950 121.950 847.050 122.400 ;
        RECT 880.950 121.950 883.050 122.400 ;
        RECT 886.950 121.950 889.050 122.400 ;
        RECT 898.950 123.600 901.050 124.050 ;
        RECT 937.950 123.600 940.050 124.050 ;
        RECT 898.950 122.400 940.050 123.600 ;
        RECT 898.950 121.950 901.050 122.400 ;
        RECT 937.950 121.950 940.050 122.400 ;
        RECT 154.950 120.600 157.050 121.050 ;
        RECT 202.950 120.600 205.050 121.050 ;
        RECT 154.950 119.400 205.050 120.600 ;
        RECT 154.950 118.950 157.050 119.400 ;
        RECT 202.950 118.950 205.050 119.400 ;
        RECT 208.950 120.600 211.050 121.050 ;
        RECT 235.950 120.600 238.050 121.050 ;
        RECT 208.950 119.400 238.050 120.600 ;
        RECT 208.950 118.950 211.050 119.400 ;
        RECT 235.950 118.950 238.050 119.400 ;
        RECT 244.950 120.600 247.050 121.050 ;
        RECT 259.950 120.600 262.050 121.050 ;
        RECT 244.950 119.400 262.050 120.600 ;
        RECT 244.950 118.950 247.050 119.400 ;
        RECT 259.950 118.950 262.050 119.400 ;
        RECT 328.950 120.600 331.050 121.050 ;
        RECT 340.950 120.600 343.050 121.050 ;
        RECT 328.950 119.400 343.050 120.600 ;
        RECT 328.950 118.950 331.050 119.400 ;
        RECT 340.950 118.950 343.050 119.400 ;
        RECT 346.950 120.600 349.050 121.050 ;
        RECT 355.950 120.600 358.050 121.050 ;
        RECT 346.950 119.400 358.050 120.600 ;
        RECT 346.950 118.950 349.050 119.400 ;
        RECT 355.950 118.950 358.050 119.400 ;
        RECT 364.950 120.600 367.050 121.050 ;
        RECT 412.950 120.600 415.050 121.050 ;
        RECT 478.950 120.600 481.050 121.050 ;
        RECT 364.950 119.400 415.050 120.600 ;
        RECT 364.950 118.950 367.050 119.400 ;
        RECT 412.950 118.950 415.050 119.400 ;
        RECT 428.400 119.400 481.050 120.600 ;
        RECT 103.950 117.600 106.050 118.050 ;
        RECT 160.950 117.600 163.050 118.050 ;
        RECT 103.950 116.400 163.050 117.600 ;
        RECT 103.950 115.950 106.050 116.400 ;
        RECT 160.950 115.950 163.050 116.400 ;
        RECT 202.950 117.600 205.050 117.900 ;
        RECT 238.950 117.600 241.050 118.050 ;
        RECT 262.950 117.600 265.050 118.050 ;
        RECT 283.950 117.600 286.050 118.050 ;
        RECT 202.950 116.400 286.050 117.600 ;
        RECT 202.950 115.800 205.050 116.400 ;
        RECT 238.950 115.950 241.050 116.400 ;
        RECT 262.950 115.950 265.050 116.400 ;
        RECT 283.950 115.950 286.050 116.400 ;
        RECT 289.950 117.600 292.050 118.050 ;
        RECT 301.950 117.600 304.050 118.050 ;
        RECT 289.950 116.400 304.050 117.600 ;
        RECT 289.950 115.950 292.050 116.400 ;
        RECT 301.950 115.950 304.050 116.400 ;
        RECT 310.950 117.600 313.050 118.050 ;
        RECT 316.950 117.600 319.050 118.050 ;
        RECT 310.950 116.400 319.050 117.600 ;
        RECT 310.950 115.950 313.050 116.400 ;
        RECT 316.950 115.950 319.050 116.400 ;
        RECT 361.950 117.600 364.050 118.050 ;
        RECT 428.400 117.600 429.600 119.400 ;
        RECT 478.950 118.950 481.050 119.400 ;
        RECT 499.950 120.600 502.050 121.050 ;
        RECT 637.950 120.600 640.050 121.050 ;
        RECT 499.950 119.400 640.050 120.600 ;
        RECT 499.950 118.950 502.050 119.400 ;
        RECT 637.950 118.950 640.050 119.400 ;
        RECT 706.950 120.600 709.050 121.050 ;
        RECT 733.950 120.600 736.050 121.050 ;
        RECT 706.950 119.400 736.050 120.600 ;
        RECT 706.950 118.950 709.050 119.400 ;
        RECT 733.950 118.950 736.050 119.400 ;
        RECT 739.950 120.600 742.050 121.050 ;
        RECT 760.950 120.600 763.050 121.050 ;
        RECT 739.950 119.400 763.050 120.600 ;
        RECT 800.400 120.600 801.600 121.950 ;
        RECT 892.950 120.600 895.050 121.050 ;
        RECT 800.400 119.400 895.050 120.600 ;
        RECT 739.950 118.950 742.050 119.400 ;
        RECT 760.950 118.950 763.050 119.400 ;
        RECT 892.950 118.950 895.050 119.400 ;
        RECT 361.950 116.400 429.600 117.600 ;
        RECT 742.950 117.600 745.050 118.050 ;
        RECT 763.950 117.600 766.050 118.050 ;
        RECT 742.950 116.400 766.050 117.600 ;
        RECT 361.950 115.950 364.050 116.400 ;
        RECT 742.950 115.950 745.050 116.400 ;
        RECT 763.950 115.950 766.050 116.400 ;
        RECT 796.950 117.600 799.050 118.050 ;
        RECT 808.950 117.600 811.050 118.050 ;
        RECT 796.950 116.400 811.050 117.600 ;
        RECT 796.950 115.950 799.050 116.400 ;
        RECT 808.950 115.950 811.050 116.400 ;
        RECT 832.950 117.600 835.050 118.050 ;
        RECT 847.950 117.600 850.050 118.050 ;
        RECT 832.950 116.400 850.050 117.600 ;
        RECT 893.400 117.600 894.600 118.950 ;
        RECT 919.950 117.600 922.050 118.050 ;
        RECT 893.400 116.400 922.050 117.600 ;
        RECT 832.950 115.950 835.050 116.400 ;
        RECT 847.950 115.950 850.050 116.400 ;
        RECT 919.950 115.950 922.050 116.400 ;
        RECT 49.950 114.600 52.050 115.050 ;
        RECT 109.950 114.600 112.050 115.050 ;
        RECT 49.950 113.400 112.050 114.600 ;
        RECT 49.950 112.950 52.050 113.400 ;
        RECT 109.950 112.950 112.050 113.400 ;
        RECT 139.950 114.600 142.050 115.050 ;
        RECT 199.950 114.600 202.050 115.050 ;
        RECT 139.950 113.400 202.050 114.600 ;
        RECT 139.950 112.950 142.050 113.400 ;
        RECT 199.950 112.950 202.050 113.400 ;
        RECT 241.950 114.600 244.050 115.050 ;
        RECT 253.950 114.600 256.050 115.050 ;
        RECT 241.950 113.400 256.050 114.600 ;
        RECT 241.950 112.950 244.050 113.400 ;
        RECT 253.950 112.950 256.050 113.400 ;
        RECT 265.950 114.600 268.050 115.050 ;
        RECT 286.950 114.600 289.050 115.050 ;
        RECT 265.950 113.400 289.050 114.600 ;
        RECT 265.950 112.950 268.050 113.400 ;
        RECT 286.950 112.950 289.050 113.400 ;
        RECT 295.950 114.600 298.050 115.050 ;
        RECT 319.950 114.600 322.050 115.050 ;
        RECT 334.950 114.600 337.050 115.050 ;
        RECT 295.950 113.400 337.050 114.600 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 319.950 112.950 322.050 113.400 ;
        RECT 334.950 112.950 337.050 113.400 ;
        RECT 355.950 114.600 358.050 115.050 ;
        RECT 430.950 114.600 433.050 115.050 ;
        RECT 355.950 113.400 433.050 114.600 ;
        RECT 355.950 112.950 358.050 113.400 ;
        RECT 430.950 112.950 433.050 113.400 ;
        RECT 436.950 114.600 439.050 115.050 ;
        RECT 481.950 114.600 484.050 115.050 ;
        RECT 436.950 113.400 484.050 114.600 ;
        RECT 436.950 112.950 439.050 113.400 ;
        RECT 481.950 112.950 484.050 113.400 ;
        RECT 538.950 114.600 541.050 115.050 ;
        RECT 595.950 114.600 598.050 115.050 ;
        RECT 610.950 114.600 613.050 115.050 ;
        RECT 661.950 114.600 664.050 115.050 ;
        RECT 667.950 114.600 670.050 115.050 ;
        RECT 538.950 113.400 613.050 114.600 ;
        RECT 538.950 112.950 541.050 113.400 ;
        RECT 595.950 112.950 598.050 113.400 ;
        RECT 610.950 112.950 613.050 113.400 ;
        RECT 644.400 113.400 670.050 114.600 ;
        RECT 644.400 112.050 645.600 113.400 ;
        RECT 661.950 112.950 664.050 113.400 ;
        RECT 667.950 112.950 670.050 113.400 ;
        RECT 676.950 114.600 679.050 115.050 ;
        RECT 730.950 114.600 733.050 115.050 ;
        RECT 676.950 113.400 733.050 114.600 ;
        RECT 676.950 112.950 679.050 113.400 ;
        RECT 730.950 112.950 733.050 113.400 ;
        RECT 751.950 114.600 754.050 115.050 ;
        RECT 829.950 114.600 832.050 115.050 ;
        RECT 751.950 113.400 832.050 114.600 ;
        RECT 751.950 112.950 754.050 113.400 ;
        RECT 829.950 112.950 832.050 113.400 ;
        RECT 877.950 114.600 880.050 115.050 ;
        RECT 910.950 114.600 913.050 115.050 ;
        RECT 877.950 113.400 913.050 114.600 ;
        RECT 877.950 112.950 880.050 113.400 ;
        RECT 910.950 112.950 913.050 113.400 ;
        RECT 37.950 111.600 40.050 112.050 ;
        RECT 67.950 111.600 70.050 112.050 ;
        RECT 37.950 110.400 70.050 111.600 ;
        RECT 37.950 109.950 40.050 110.400 ;
        RECT 67.950 109.950 70.050 110.400 ;
        RECT 79.950 111.600 82.050 112.050 ;
        RECT 88.950 111.600 91.050 112.050 ;
        RECT 79.950 110.400 91.050 111.600 ;
        RECT 79.950 109.950 82.050 110.400 ;
        RECT 88.950 109.950 91.050 110.400 ;
        RECT 163.950 111.600 166.050 112.050 ;
        RECT 172.950 111.600 175.050 112.050 ;
        RECT 163.950 110.400 175.050 111.600 ;
        RECT 163.950 109.950 166.050 110.400 ;
        RECT 172.950 109.950 175.050 110.400 ;
        RECT 178.950 111.600 181.050 112.050 ;
        RECT 214.950 111.600 217.050 112.050 ;
        RECT 289.800 111.600 291.900 112.050 ;
        RECT 178.950 110.400 291.900 111.600 ;
        RECT 178.950 109.950 181.050 110.400 ;
        RECT 214.950 109.950 217.050 110.400 ;
        RECT 289.800 109.950 291.900 110.400 ;
        RECT 292.950 111.600 295.050 112.050 ;
        RECT 337.950 111.600 340.050 112.050 ;
        RECT 292.950 110.400 340.050 111.600 ;
        RECT 292.950 109.950 295.050 110.400 ;
        RECT 337.950 109.950 340.050 110.400 ;
        RECT 388.950 111.600 391.050 112.050 ;
        RECT 436.950 111.600 439.050 111.900 ;
        RECT 388.950 110.400 439.050 111.600 ;
        RECT 388.950 109.950 391.050 110.400 ;
        RECT 436.950 109.800 439.050 110.400 ;
        RECT 490.950 111.600 493.050 112.050 ;
        RECT 523.800 111.600 525.900 112.050 ;
        RECT 490.950 110.400 525.900 111.600 ;
        RECT 490.950 109.950 493.050 110.400 ;
        RECT 523.800 109.950 525.900 110.400 ;
        RECT 526.950 111.600 529.050 112.050 ;
        RECT 565.950 111.600 568.050 112.050 ;
        RECT 526.950 110.400 568.050 111.600 ;
        RECT 526.950 109.950 529.050 110.400 ;
        RECT 565.950 109.950 568.050 110.400 ;
        RECT 592.950 111.600 595.050 112.050 ;
        RECT 643.950 111.600 646.050 112.050 ;
        RECT 592.950 110.400 646.050 111.600 ;
        RECT 592.950 109.950 595.050 110.400 ;
        RECT 643.950 109.950 646.050 110.400 ;
        RECT 655.950 111.600 658.050 112.050 ;
        RECT 697.950 111.600 700.050 112.050 ;
        RECT 706.950 111.600 709.050 112.050 ;
        RECT 655.950 110.400 709.050 111.600 ;
        RECT 655.950 109.950 658.050 110.400 ;
        RECT 697.950 109.950 700.050 110.400 ;
        RECT 706.950 109.950 709.050 110.400 ;
        RECT 790.950 111.600 793.050 112.050 ;
        RECT 805.950 111.600 808.050 112.050 ;
        RECT 790.950 110.400 808.050 111.600 ;
        RECT 790.950 109.950 793.050 110.400 ;
        RECT 805.950 109.950 808.050 110.400 ;
        RECT 841.950 111.600 844.050 112.050 ;
        RECT 883.950 111.600 886.050 112.050 ;
        RECT 841.950 110.400 886.050 111.600 ;
        RECT 841.950 109.950 844.050 110.400 ;
        RECT 883.950 109.950 886.050 110.400 ;
        RECT 49.950 108.600 52.050 109.050 ;
        RECT 55.950 108.600 58.050 109.050 ;
        RECT 49.950 107.400 58.050 108.600 ;
        RECT 49.950 106.950 52.050 107.400 ;
        RECT 55.950 106.950 58.050 107.400 ;
        RECT 217.950 108.600 220.050 109.050 ;
        RECT 229.950 108.600 232.050 109.050 ;
        RECT 217.950 107.400 232.050 108.600 ;
        RECT 217.950 106.950 220.050 107.400 ;
        RECT 229.950 106.950 232.050 107.400 ;
        RECT 262.950 108.600 267.000 109.050 ;
        RECT 262.950 106.950 267.600 108.600 ;
        RECT 271.950 106.950 274.050 109.050 ;
        RECT 19.950 105.600 22.050 106.200 ;
        RECT 25.950 105.600 28.050 106.050 ;
        RECT 19.950 104.400 28.050 105.600 ;
        RECT 19.950 104.100 22.050 104.400 ;
        RECT 25.950 103.950 28.050 104.400 ;
        RECT 40.950 105.600 43.050 106.200 ;
        RECT 64.950 105.750 67.050 106.200 ;
        RECT 70.950 105.750 73.050 106.200 ;
        RECT 40.950 104.400 60.600 105.600 ;
        RECT 40.950 104.100 43.050 104.400 ;
        RECT 4.950 99.600 7.050 100.050 ;
        RECT 10.950 99.600 13.050 99.900 ;
        RECT 31.950 99.600 34.050 99.900 ;
        RECT 4.950 98.400 34.050 99.600 ;
        RECT 4.950 97.950 7.050 98.400 ;
        RECT 10.950 97.800 13.050 98.400 ;
        RECT 31.950 97.800 34.050 98.400 ;
        RECT 46.950 99.450 49.050 99.900 ;
        RECT 55.950 99.450 58.050 99.900 ;
        RECT 46.950 98.250 58.050 99.450 ;
        RECT 59.400 99.600 60.600 104.400 ;
        RECT 64.950 104.550 73.050 105.750 ;
        RECT 64.950 104.100 67.050 104.550 ;
        RECT 70.950 104.100 73.050 104.550 ;
        RECT 88.950 105.600 91.050 106.050 ;
        RECT 97.950 105.600 100.050 106.050 ;
        RECT 88.950 104.400 100.050 105.600 ;
        RECT 88.950 103.950 91.050 104.400 ;
        RECT 97.950 103.950 100.050 104.400 ;
        RECT 115.950 105.750 118.050 106.200 ;
        RECT 124.950 105.750 127.050 106.200 ;
        RECT 115.950 104.550 127.050 105.750 ;
        RECT 148.950 105.600 151.050 106.200 ;
        RECT 115.950 104.100 118.050 104.550 ;
        RECT 124.950 104.100 127.050 104.550 ;
        RECT 140.400 104.400 151.050 105.600 ;
        RECT 91.950 99.600 94.050 100.050 ;
        RECT 59.400 98.400 94.050 99.600 ;
        RECT 46.950 97.800 49.050 98.250 ;
        RECT 55.950 97.800 58.050 98.250 ;
        RECT 91.950 97.950 94.050 98.400 ;
        RECT 121.950 99.600 124.050 99.900 ;
        RECT 140.400 99.600 141.600 104.400 ;
        RECT 148.950 104.100 151.050 104.400 ;
        RECT 172.950 105.750 175.050 106.200 ;
        RECT 184.950 105.750 187.050 106.200 ;
        RECT 172.950 104.550 187.050 105.750 ;
        RECT 172.950 104.100 175.050 104.550 ;
        RECT 184.950 104.100 187.050 104.550 ;
        RECT 196.950 104.100 199.050 106.200 ;
        RECT 238.950 105.600 241.050 106.200 ;
        RECT 212.400 104.400 241.050 105.600 ;
        RECT 121.950 98.400 141.600 99.600 ;
        RECT 151.950 99.450 154.050 99.900 ;
        RECT 160.950 99.450 163.050 99.900 ;
        RECT 121.950 97.800 124.050 98.400 ;
        RECT 151.950 98.250 163.050 99.450 ;
        RECT 151.950 97.800 154.050 98.250 ;
        RECT 160.950 97.800 163.050 98.250 ;
        RECT 175.950 99.600 178.050 99.900 ;
        RECT 190.950 99.600 193.050 100.050 ;
        RECT 175.950 98.400 193.050 99.600 ;
        RECT 175.950 97.800 178.050 98.400 ;
        RECT 190.950 97.950 193.050 98.400 ;
        RECT 197.400 97.050 198.600 104.100 ;
        RECT 212.400 103.050 213.600 104.400 ;
        RECT 238.950 104.100 241.050 104.400 ;
        RECT 244.950 105.600 247.050 106.200 ;
        RECT 256.950 105.600 259.050 106.050 ;
        RECT 244.950 104.400 259.050 105.600 ;
        RECT 244.950 104.100 247.050 104.400 ;
        RECT 256.950 103.950 259.050 104.400 ;
        RECT 208.950 101.400 213.600 103.050 ;
        RECT 208.950 100.950 213.000 101.400 ;
        RECT 211.950 99.600 214.050 100.050 ;
        RECT 266.400 99.900 267.600 106.950 ;
        RECT 272.400 99.900 273.600 106.950 ;
        RECT 289.950 105.600 292.050 106.200 ;
        RECT 298.950 105.600 301.050 109.050 ;
        RECT 316.950 108.600 319.050 109.050 ;
        RECT 361.950 108.600 364.050 109.050 ;
        RECT 316.950 107.400 364.050 108.600 ;
        RECT 316.950 106.950 319.050 107.400 ;
        RECT 361.950 106.950 364.050 107.400 ;
        RECT 442.950 108.600 445.050 109.050 ;
        RECT 466.950 108.600 469.050 109.050 ;
        RECT 442.950 107.400 469.050 108.600 ;
        RECT 442.950 106.950 445.050 107.400 ;
        RECT 466.950 106.950 469.050 107.400 ;
        RECT 484.950 108.600 487.050 109.050 ;
        RECT 556.950 108.600 559.050 109.050 ;
        RECT 571.950 108.600 574.050 109.050 ;
        RECT 577.950 108.600 580.050 109.050 ;
        RECT 649.950 108.600 652.050 109.050 ;
        RECT 736.950 108.600 739.050 109.050 ;
        RECT 745.950 108.600 748.050 109.050 ;
        RECT 802.950 108.600 805.050 109.050 ;
        RECT 484.950 107.400 580.050 108.600 ;
        RECT 484.950 106.950 487.050 107.400 ;
        RECT 556.950 106.950 559.050 107.400 ;
        RECT 571.950 106.950 574.050 107.400 ;
        RECT 577.950 106.950 580.050 107.400 ;
        RECT 641.400 107.400 711.600 108.600 ;
        RECT 289.950 105.000 301.050 105.600 ;
        RECT 289.950 104.400 300.600 105.000 ;
        RECT 289.950 104.100 292.050 104.400 ;
        RECT 313.950 104.100 316.050 106.200 ;
        RECT 277.950 102.600 280.050 103.050 ;
        RECT 314.400 102.600 315.600 104.100 ;
        RECT 325.950 103.950 328.050 106.050 ;
        RECT 337.950 105.600 340.050 106.200 ;
        RECT 349.950 105.600 352.050 106.200 ;
        RECT 337.950 104.400 352.050 105.600 ;
        RECT 337.950 104.100 340.050 104.400 ;
        RECT 349.950 104.100 352.050 104.400 ;
        RECT 385.950 105.750 388.050 106.200 ;
        RECT 397.950 105.750 400.050 106.200 ;
        RECT 385.950 104.550 400.050 105.750 ;
        RECT 385.950 104.100 388.050 104.550 ;
        RECT 397.950 104.100 400.050 104.550 ;
        RECT 409.950 105.750 412.050 106.200 ;
        RECT 418.950 105.750 421.050 106.200 ;
        RECT 409.950 104.550 421.050 105.750 ;
        RECT 424.950 105.600 427.050 106.200 ;
        RECT 451.950 105.600 454.050 106.050 ;
        RECT 409.950 104.100 412.050 104.550 ;
        RECT 418.950 104.100 421.050 104.550 ;
        RECT 422.400 104.400 454.050 105.600 ;
        RECT 277.950 101.400 315.600 102.600 ;
        RECT 277.950 100.950 280.050 101.400 ;
        RECT 247.950 99.600 250.050 99.900 ;
        RECT 211.950 98.400 250.050 99.600 ;
        RECT 211.950 97.950 214.050 98.400 ;
        RECT 247.950 97.800 250.050 98.400 ;
        RECT 265.950 97.800 268.050 99.900 ;
        RECT 271.950 99.600 274.050 99.900 ;
        RECT 286.950 99.600 289.050 99.900 ;
        RECT 271.950 98.400 289.050 99.600 ;
        RECT 271.950 97.800 274.050 98.400 ;
        RECT 286.950 97.800 289.050 98.400 ;
        RECT 298.950 99.450 301.050 99.900 ;
        RECT 322.950 99.450 325.050 99.900 ;
        RECT 298.950 98.250 325.050 99.450 ;
        RECT 326.400 99.600 327.600 103.950 ;
        RECT 406.950 102.600 409.050 103.050 ;
        RECT 422.400 102.600 423.600 104.400 ;
        RECT 424.950 104.100 427.050 104.400 ;
        RECT 451.950 103.950 454.050 104.400 ;
        RECT 466.950 105.600 469.050 106.200 ;
        RECT 505.950 105.600 508.050 106.200 ;
        RECT 466.950 104.400 508.050 105.600 ;
        RECT 466.950 104.100 469.050 104.400 ;
        RECT 505.950 104.100 508.050 104.400 ;
        RECT 511.950 105.750 514.050 106.200 ;
        RECT 520.950 105.750 523.050 106.200 ;
        RECT 511.950 105.600 523.050 105.750 ;
        RECT 532.950 105.600 535.050 106.200 ;
        RECT 511.950 104.550 535.050 105.600 ;
        RECT 511.950 104.100 514.050 104.550 ;
        RECT 520.950 104.400 535.050 104.550 ;
        RECT 520.950 104.100 523.050 104.400 ;
        RECT 532.950 104.100 535.050 104.400 ;
        RECT 544.950 105.600 547.050 106.050 ;
        RECT 550.950 105.600 553.050 106.200 ;
        RECT 544.950 104.400 553.050 105.600 ;
        RECT 544.950 103.950 547.050 104.400 ;
        RECT 550.950 104.100 553.050 104.400 ;
        RECT 583.950 105.600 586.050 106.200 ;
        RECT 589.950 105.750 592.050 106.200 ;
        RECT 601.950 105.750 604.050 106.200 ;
        RECT 589.950 105.600 604.050 105.750 ;
        RECT 619.950 105.600 622.050 106.200 ;
        RECT 583.950 104.400 588.600 105.600 ;
        RECT 583.950 104.100 586.050 104.400 ;
        RECT 406.950 101.400 423.600 102.600 ;
        RECT 554.400 101.400 570.600 102.600 ;
        RECT 406.950 100.950 409.050 101.400 ;
        RECT 331.950 99.600 334.050 100.050 ;
        RECT 326.400 98.400 334.050 99.600 ;
        RECT 298.950 97.800 301.050 98.250 ;
        RECT 322.950 97.800 325.050 98.250 ;
        RECT 331.950 97.950 334.050 98.400 ;
        RECT 343.950 99.450 346.050 99.900 ;
        RECT 352.950 99.450 355.050 99.900 ;
        RECT 343.950 98.250 355.050 99.450 ;
        RECT 343.950 97.800 346.050 98.250 ;
        RECT 352.950 97.800 355.050 98.250 ;
        RECT 370.950 99.600 373.050 99.900 ;
        RECT 400.950 99.600 403.050 99.900 ;
        RECT 409.800 99.600 411.900 100.050 ;
        RECT 370.950 98.400 411.900 99.600 ;
        RECT 370.950 97.800 373.050 98.400 ;
        RECT 400.950 97.800 403.050 98.400 ;
        RECT 409.800 97.950 411.900 98.400 ;
        RECT 412.950 99.600 415.050 100.050 ;
        RECT 554.400 99.900 555.600 101.400 ;
        RECT 569.400 99.900 570.600 101.400 ;
        RECT 587.400 100.050 588.600 104.400 ;
        RECT 589.950 104.550 618.600 105.600 ;
        RECT 589.950 104.100 592.050 104.550 ;
        RECT 601.950 104.400 618.600 104.550 ;
        RECT 601.950 104.100 604.050 104.400 ;
        RECT 421.950 99.600 424.050 99.900 ;
        RECT 412.950 99.450 424.050 99.600 ;
        RECT 430.950 99.450 433.050 99.900 ;
        RECT 412.950 98.400 433.050 99.450 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 421.950 98.250 433.050 98.400 ;
        RECT 421.950 97.800 424.050 98.250 ;
        RECT 430.950 97.800 433.050 98.250 ;
        RECT 445.950 99.450 448.050 99.900 ;
        RECT 451.950 99.600 454.050 99.900 ;
        RECT 463.950 99.600 466.050 99.900 ;
        RECT 451.950 99.450 466.050 99.600 ;
        RECT 445.950 98.400 466.050 99.450 ;
        RECT 445.950 98.250 454.050 98.400 ;
        RECT 445.950 97.800 448.050 98.250 ;
        RECT 451.950 97.800 454.050 98.250 ;
        RECT 463.950 97.800 466.050 98.400 ;
        RECT 508.950 99.600 511.050 99.900 ;
        RECT 529.950 99.600 532.050 99.900 ;
        RECT 508.950 98.400 532.050 99.600 ;
        RECT 508.950 97.800 511.050 98.400 ;
        RECT 529.950 97.800 532.050 98.400 ;
        RECT 553.950 97.800 556.050 99.900 ;
        RECT 559.950 99.450 562.050 99.900 ;
        RECT 565.800 99.450 567.900 99.900 ;
        RECT 559.950 98.250 567.900 99.450 ;
        RECT 559.950 97.800 562.050 98.250 ;
        RECT 565.800 97.800 567.900 98.250 ;
        RECT 568.950 99.450 571.050 99.900 ;
        RECT 574.950 99.450 577.050 99.900 ;
        RECT 568.950 98.250 577.050 99.450 ;
        RECT 568.950 97.800 571.050 98.250 ;
        RECT 574.950 97.800 577.050 98.250 ;
        RECT 586.950 97.950 589.050 100.050 ;
        RECT 617.400 99.900 618.600 104.400 ;
        RECT 619.950 104.400 630.600 105.600 ;
        RECT 619.950 104.100 622.050 104.400 ;
        RECT 629.400 100.050 630.600 104.400 ;
        RECT 616.950 97.800 619.050 99.900 ;
        RECT 629.400 98.400 634.050 100.050 ;
        RECT 641.400 99.900 642.600 107.400 ;
        RECT 649.950 106.950 652.050 107.400 ;
        RECT 661.950 105.600 664.050 106.200 ;
        RECT 682.950 105.600 685.050 106.200 ;
        RECT 647.400 104.400 664.050 105.600 ;
        RECT 647.400 100.050 648.600 104.400 ;
        RECT 661.950 104.100 664.050 104.400 ;
        RECT 671.400 104.400 685.050 105.600 ;
        RECT 649.950 102.600 652.050 103.050 ;
        RECT 649.950 101.400 663.600 102.600 ;
        RECT 649.950 100.950 652.050 101.400 ;
        RECT 630.000 97.950 634.050 98.400 ;
        RECT 640.950 97.800 643.050 99.900 ;
        RECT 646.950 97.950 649.050 100.050 ;
        RECT 662.400 99.600 663.600 101.400 ;
        RECT 671.400 100.050 672.600 104.400 ;
        RECT 682.950 104.100 685.050 104.400 ;
        RECT 688.950 105.600 691.050 106.200 ;
        RECT 688.950 104.400 705.600 105.600 ;
        RECT 688.950 104.100 691.050 104.400 ;
        RECT 704.400 100.050 705.600 104.400 ;
        RECT 664.950 99.600 667.050 99.900 ;
        RECT 662.400 98.400 667.050 99.600 ;
        RECT 664.950 97.800 667.050 98.400 ;
        RECT 670.950 97.950 673.050 100.050 ;
        RECT 691.950 99.450 694.050 99.900 ;
        RECT 697.950 99.450 700.050 99.900 ;
        RECT 691.950 98.250 700.050 99.450 ;
        RECT 691.950 97.800 694.050 98.250 ;
        RECT 697.950 97.800 700.050 98.250 ;
        RECT 703.950 97.950 706.050 100.050 ;
        RECT 710.400 99.900 711.600 107.400 ;
        RECT 736.950 107.400 748.050 108.600 ;
        RECT 736.950 106.950 739.050 107.400 ;
        RECT 745.950 106.950 748.050 107.400 ;
        RECT 797.400 107.400 805.050 108.600 ;
        RECT 748.950 105.600 753.000 106.050 ;
        RECT 754.950 105.600 757.050 106.200 ;
        RECT 766.950 105.600 769.050 106.050 ;
        RECT 775.950 105.600 778.050 106.200 ;
        RECT 748.950 103.950 753.600 105.600 ;
        RECT 754.950 104.400 769.050 105.600 ;
        RECT 754.950 104.100 757.050 104.400 ;
        RECT 766.950 103.950 769.050 104.400 ;
        RECT 770.400 104.400 778.050 105.600 ;
        RECT 752.400 99.900 753.600 103.950 ;
        RECT 709.950 97.800 712.050 99.900 ;
        RECT 721.950 99.450 724.050 99.900 ;
        RECT 733.950 99.450 736.050 99.900 ;
        RECT 721.950 98.250 736.050 99.450 ;
        RECT 721.950 97.800 724.050 98.250 ;
        RECT 733.950 97.800 736.050 98.250 ;
        RECT 751.950 97.800 754.050 99.900 ;
        RECT 757.950 99.450 760.050 99.900 ;
        RECT 763.950 99.450 766.050 99.900 ;
        RECT 757.950 98.250 766.050 99.450 ;
        RECT 757.950 97.800 760.050 98.250 ;
        RECT 763.950 97.800 766.050 98.250 ;
        RECT 112.950 96.600 115.050 97.050 ;
        RECT 133.950 96.600 136.050 97.050 ;
        RECT 112.950 95.400 136.050 96.600 ;
        RECT 112.950 94.950 115.050 95.400 ;
        RECT 133.950 94.950 136.050 95.400 ;
        RECT 196.950 94.950 199.050 97.050 ;
        RECT 604.950 96.600 607.050 97.050 ;
        RECT 627.000 96.600 631.050 97.050 ;
        RECT 770.400 96.900 771.600 104.400 ;
        RECT 775.950 104.100 778.050 104.400 ;
        RECT 784.950 105.750 787.050 106.200 ;
        RECT 793.950 105.750 796.050 106.200 ;
        RECT 784.950 104.550 796.050 105.750 ;
        RECT 784.950 104.100 787.050 104.550 ;
        RECT 793.950 104.100 796.050 104.550 ;
        RECT 797.400 99.900 798.600 107.400 ;
        RECT 802.950 106.950 805.050 107.400 ;
        RECT 811.950 108.600 814.050 109.050 ;
        RECT 820.950 108.600 823.050 109.050 ;
        RECT 811.950 107.400 823.050 108.600 ;
        RECT 811.950 106.950 814.050 107.400 ;
        RECT 820.950 106.950 823.050 107.400 ;
        RECT 889.950 108.600 892.050 109.050 ;
        RECT 940.950 108.600 943.050 109.050 ;
        RECT 889.950 107.400 943.050 108.600 ;
        RECT 889.950 106.950 892.050 107.400 ;
        RECT 940.950 106.950 943.050 107.400 ;
        RECT 799.950 105.600 802.050 106.200 ;
        RECT 826.950 105.750 829.050 106.200 ;
        RECT 838.950 105.750 841.050 106.200 ;
        RECT 826.950 105.600 841.050 105.750 ;
        RECT 868.950 105.600 871.050 106.200 ;
        RECT 799.950 104.400 804.600 105.600 ;
        RECT 799.950 104.100 802.050 104.400 ;
        RECT 796.950 97.800 799.050 99.900 ;
        RECT 803.400 97.050 804.600 104.400 ;
        RECT 818.400 104.550 871.050 105.600 ;
        RECT 818.400 104.400 829.050 104.550 ;
        RECT 818.400 99.900 819.600 104.400 ;
        RECT 826.950 104.100 829.050 104.400 ;
        RECT 838.950 104.400 871.050 104.550 ;
        RECT 838.950 104.100 841.050 104.400 ;
        RECT 868.950 104.100 871.050 104.400 ;
        RECT 880.950 105.600 883.050 106.050 ;
        RECT 886.950 105.600 889.050 106.050 ;
        RECT 880.950 104.400 889.050 105.600 ;
        RECT 880.950 103.950 883.050 104.400 ;
        RECT 886.950 103.950 889.050 104.400 ;
        RECT 859.950 102.600 862.050 103.050 ;
        RECT 851.400 101.400 862.050 102.600 ;
        RECT 817.950 97.800 820.050 99.900 ;
        RECT 829.950 99.450 832.050 99.900 ;
        RECT 835.950 99.600 838.050 99.900 ;
        RECT 851.400 99.600 852.600 101.400 ;
        RECT 859.950 100.950 862.050 101.400 ;
        RECT 835.950 99.450 852.600 99.600 ;
        RECT 829.950 98.400 852.600 99.450 ;
        RECT 871.950 99.600 874.050 99.900 ;
        RECT 883.950 99.600 886.050 99.900 ;
        RECT 871.950 98.400 886.050 99.600 ;
        RECT 829.950 98.250 838.050 98.400 ;
        RECT 829.950 97.800 832.050 98.250 ;
        RECT 835.950 97.800 838.050 98.250 ;
        RECT 871.950 97.800 874.050 98.400 ;
        RECT 883.950 97.800 886.050 98.400 ;
        RECT 604.950 95.400 631.050 96.600 ;
        RECT 604.950 94.950 607.050 95.400 ;
        RECT 626.400 94.950 631.050 95.400 ;
        RECT 37.950 93.600 40.050 94.050 ;
        RECT 70.950 93.600 73.050 94.050 ;
        RECT 103.950 93.600 106.050 94.050 ;
        RECT 37.950 92.400 106.050 93.600 ;
        RECT 37.950 91.950 40.050 92.400 ;
        RECT 70.950 91.950 73.050 92.400 ;
        RECT 103.950 91.950 106.050 92.400 ;
        RECT 175.950 93.600 178.050 94.050 ;
        RECT 184.950 93.600 187.050 94.050 ;
        RECT 193.950 93.600 196.050 94.050 ;
        RECT 175.950 92.400 196.050 93.600 ;
        RECT 175.950 91.950 178.050 92.400 ;
        RECT 184.950 91.950 187.050 92.400 ;
        RECT 193.950 91.950 196.050 92.400 ;
        RECT 256.950 93.600 259.050 94.050 ;
        RECT 304.950 93.600 307.050 94.050 ;
        RECT 256.950 92.400 307.050 93.600 ;
        RECT 256.950 91.950 259.050 92.400 ;
        RECT 304.950 91.950 307.050 92.400 ;
        RECT 322.950 93.600 325.050 94.050 ;
        RECT 328.950 93.600 331.050 94.050 ;
        RECT 334.800 93.600 336.900 94.050 ;
        RECT 322.950 92.400 336.900 93.600 ;
        RECT 322.950 91.950 325.050 92.400 ;
        RECT 328.950 91.950 331.050 92.400 ;
        RECT 334.800 91.950 336.900 92.400 ;
        RECT 337.950 93.600 340.050 94.050 ;
        RECT 370.950 93.600 373.050 94.050 ;
        RECT 337.950 92.400 373.050 93.600 ;
        RECT 337.950 91.950 340.050 92.400 ;
        RECT 370.950 91.950 373.050 92.400 ;
        RECT 478.950 93.600 481.050 94.050 ;
        RECT 493.950 93.600 496.050 94.050 ;
        RECT 514.950 93.600 517.050 94.050 ;
        RECT 550.950 93.600 553.050 94.050 ;
        RECT 478.950 92.400 553.050 93.600 ;
        RECT 478.950 91.950 481.050 92.400 ;
        RECT 493.950 91.950 496.050 92.400 ;
        RECT 514.950 91.950 517.050 92.400 ;
        RECT 550.950 91.950 553.050 92.400 ;
        RECT 610.950 93.600 613.050 94.050 ;
        RECT 622.950 93.600 625.050 94.050 ;
        RECT 610.950 92.400 625.050 93.600 ;
        RECT 626.400 93.600 627.600 94.950 ;
        RECT 769.950 94.800 772.050 96.900 ;
        RECT 799.950 95.400 804.600 97.050 ;
        RECT 820.950 96.600 823.050 97.050 ;
        RECT 832.950 96.600 835.050 97.050 ;
        RECT 820.950 95.400 835.050 96.600 ;
        RECT 799.950 94.950 804.000 95.400 ;
        RECT 820.950 94.950 823.050 95.400 ;
        RECT 832.950 94.950 835.050 95.400 ;
        RECT 853.950 96.600 856.050 97.050 ;
        RECT 865.950 96.600 868.050 97.050 ;
        RECT 853.950 95.400 868.050 96.600 ;
        RECT 853.950 94.950 856.050 95.400 ;
        RECT 865.950 94.950 868.050 95.400 ;
        RECT 658.950 93.600 661.050 94.050 ;
        RECT 626.400 92.400 661.050 93.600 ;
        RECT 610.950 91.950 613.050 92.400 ;
        RECT 622.950 91.950 625.050 92.400 ;
        RECT 658.950 91.950 661.050 92.400 ;
        RECT 703.950 93.600 706.050 94.050 ;
        RECT 715.950 93.600 718.050 94.050 ;
        RECT 703.950 92.400 718.050 93.600 ;
        RECT 703.950 91.950 706.050 92.400 ;
        RECT 715.950 91.950 718.050 92.400 ;
        RECT 721.950 93.600 724.050 94.050 ;
        RECT 745.950 93.600 748.050 94.050 ;
        RECT 766.950 93.600 769.050 94.050 ;
        RECT 721.950 92.400 769.050 93.600 ;
        RECT 721.950 91.950 724.050 92.400 ;
        RECT 745.950 91.950 748.050 92.400 ;
        RECT 766.950 91.950 769.050 92.400 ;
        RECT 889.950 93.600 892.050 94.050 ;
        RECT 925.950 93.600 928.050 94.050 ;
        RECT 889.950 92.400 928.050 93.600 ;
        RECT 889.950 91.950 892.050 92.400 ;
        RECT 925.950 91.950 928.050 92.400 ;
        RECT 88.950 90.600 91.050 91.050 ;
        RECT 115.950 90.600 118.050 91.050 ;
        RECT 145.950 90.600 148.050 91.050 ;
        RECT 88.950 89.400 148.050 90.600 ;
        RECT 88.950 88.950 91.050 89.400 ;
        RECT 115.950 88.950 118.050 89.400 ;
        RECT 145.950 88.950 148.050 89.400 ;
        RECT 202.950 90.600 205.050 91.050 ;
        RECT 220.950 90.600 223.050 91.050 ;
        RECT 202.950 89.400 223.050 90.600 ;
        RECT 202.950 88.950 205.050 89.400 ;
        RECT 220.950 88.950 223.050 89.400 ;
        RECT 244.950 90.600 247.050 91.050 ;
        RECT 277.950 90.600 280.050 91.050 ;
        RECT 244.950 89.400 280.050 90.600 ;
        RECT 244.950 88.950 247.050 89.400 ;
        RECT 277.950 88.950 280.050 89.400 ;
        RECT 313.950 90.600 316.050 91.050 ;
        RECT 376.950 90.600 379.050 91.050 ;
        RECT 385.950 90.600 388.050 91.050 ;
        RECT 415.950 90.600 418.050 91.050 ;
        RECT 313.950 89.400 418.050 90.600 ;
        RECT 313.950 88.950 316.050 89.400 ;
        RECT 376.950 88.950 379.050 89.400 ;
        RECT 385.950 88.950 388.050 89.400 ;
        RECT 415.950 88.950 418.050 89.400 ;
        RECT 421.950 90.600 424.050 91.050 ;
        RECT 529.950 90.600 532.050 91.050 ;
        RECT 535.950 90.600 538.050 91.050 ;
        RECT 421.950 89.400 474.600 90.600 ;
        RECT 421.950 88.950 424.050 89.400 ;
        RECT 67.950 87.600 70.050 88.050 ;
        RECT 169.950 87.600 172.050 88.050 ;
        RECT 196.950 87.600 199.050 88.050 ;
        RECT 67.950 86.400 199.050 87.600 ;
        RECT 67.950 85.950 70.050 86.400 ;
        RECT 169.950 85.950 172.050 86.400 ;
        RECT 196.950 85.950 199.050 86.400 ;
        RECT 334.950 87.600 337.050 88.050 ;
        RECT 358.950 87.600 361.050 88.050 ;
        RECT 334.950 86.400 361.050 87.600 ;
        RECT 473.400 87.600 474.600 89.400 ;
        RECT 529.950 89.400 538.050 90.600 ;
        RECT 529.950 88.950 532.050 89.400 ;
        RECT 535.950 88.950 538.050 89.400 ;
        RECT 475.950 87.600 478.050 88.050 ;
        RECT 487.950 87.600 490.050 88.050 ;
        RECT 473.400 86.400 490.050 87.600 ;
        RECT 334.950 85.950 337.050 86.400 ;
        RECT 358.950 85.950 361.050 86.400 ;
        RECT 475.950 85.950 478.050 86.400 ;
        RECT 487.950 85.950 490.050 86.400 ;
        RECT 556.950 87.600 559.050 88.050 ;
        RECT 586.950 87.600 589.050 88.050 ;
        RECT 556.950 86.400 589.050 87.600 ;
        RECT 556.950 85.950 559.050 86.400 ;
        RECT 586.950 85.950 589.050 86.400 ;
        RECT 607.950 87.600 610.050 88.050 ;
        RECT 673.950 87.600 676.050 88.050 ;
        RECT 685.950 87.600 688.050 88.050 ;
        RECT 607.950 86.400 688.050 87.600 ;
        RECT 607.950 85.950 610.050 86.400 ;
        RECT 673.950 85.950 676.050 86.400 ;
        RECT 685.950 85.950 688.050 86.400 ;
        RECT 700.950 87.600 703.050 88.050 ;
        RECT 739.950 87.600 742.050 88.050 ;
        RECT 700.950 86.400 742.050 87.600 ;
        RECT 700.950 85.950 703.050 86.400 ;
        RECT 739.950 85.950 742.050 86.400 ;
        RECT 763.950 87.600 766.050 88.050 ;
        RECT 778.950 87.600 781.050 88.050 ;
        RECT 763.950 86.400 781.050 87.600 ;
        RECT 763.950 85.950 766.050 86.400 ;
        RECT 778.950 85.950 781.050 86.400 ;
        RECT 787.950 87.600 790.050 88.050 ;
        RECT 802.950 87.600 805.050 88.050 ;
        RECT 916.950 87.600 919.050 88.050 ;
        RECT 787.950 86.400 805.050 87.600 ;
        RECT 787.950 85.950 790.050 86.400 ;
        RECT 802.950 85.950 805.050 86.400 ;
        RECT 863.400 86.400 919.050 87.600 ;
        RECT 16.950 84.600 19.050 85.050 ;
        RECT 61.950 84.600 64.050 85.050 ;
        RECT 76.950 84.600 79.050 85.050 ;
        RECT 16.950 83.400 79.050 84.600 ;
        RECT 16.950 82.950 19.050 83.400 ;
        RECT 61.950 82.950 64.050 83.400 ;
        RECT 76.950 82.950 79.050 83.400 ;
        RECT 115.950 84.600 118.050 85.050 ;
        RECT 121.950 84.600 124.050 85.050 ;
        RECT 115.950 83.400 124.050 84.600 ;
        RECT 115.950 82.950 118.050 83.400 ;
        RECT 121.950 82.950 124.050 83.400 ;
        RECT 130.950 84.600 133.050 85.050 ;
        RECT 163.950 84.600 166.050 85.050 ;
        RECT 130.950 83.400 166.050 84.600 ;
        RECT 130.950 82.950 133.050 83.400 ;
        RECT 163.950 82.950 166.050 83.400 ;
        RECT 229.950 84.600 232.050 85.050 ;
        RECT 280.950 84.600 283.050 85.050 ;
        RECT 229.950 83.400 283.050 84.600 ;
        RECT 229.950 82.950 232.050 83.400 ;
        RECT 280.950 82.950 283.050 83.400 ;
        RECT 316.950 84.600 319.050 85.050 ;
        RECT 421.950 84.600 424.050 85.050 ;
        RECT 316.950 83.400 424.050 84.600 ;
        RECT 316.950 82.950 319.050 83.400 ;
        RECT 421.950 82.950 424.050 83.400 ;
        RECT 439.950 84.600 442.050 85.050 ;
        RECT 469.950 84.600 472.050 85.050 ;
        RECT 520.950 84.600 523.050 85.050 ;
        RECT 439.950 83.400 523.050 84.600 ;
        RECT 439.950 82.950 442.050 83.400 ;
        RECT 469.950 82.950 472.050 83.400 ;
        RECT 520.950 82.950 523.050 83.400 ;
        RECT 796.950 84.600 799.050 85.050 ;
        RECT 863.400 84.600 864.600 86.400 ;
        RECT 916.950 85.950 919.050 86.400 ;
        RECT 796.950 83.400 864.600 84.600 ;
        RECT 796.950 82.950 799.050 83.400 ;
        RECT 91.950 81.600 94.050 82.050 ;
        RECT 427.950 81.600 430.050 82.050 ;
        RECT 454.950 81.600 457.050 82.050 ;
        RECT 91.950 80.400 147.600 81.600 ;
        RECT 91.950 79.950 94.050 80.400 ;
        RECT 146.400 79.050 147.600 80.400 ;
        RECT 427.950 80.400 457.050 81.600 ;
        RECT 427.950 79.950 430.050 80.400 ;
        RECT 454.950 79.950 457.050 80.400 ;
        RECT 544.950 81.600 547.050 82.050 ;
        RECT 592.950 81.600 595.050 82.050 ;
        RECT 544.950 80.400 595.050 81.600 ;
        RECT 544.950 79.950 547.050 80.400 ;
        RECT 592.950 79.950 595.050 80.400 ;
        RECT 145.950 78.600 148.050 79.050 ;
        RECT 169.950 78.600 172.050 79.050 ;
        RECT 145.950 77.400 172.050 78.600 ;
        RECT 145.950 76.950 148.050 77.400 ;
        RECT 169.950 76.950 172.050 77.400 ;
        RECT 319.950 78.600 322.050 79.050 ;
        RECT 424.950 78.600 427.050 79.050 ;
        RECT 319.950 77.400 427.050 78.600 ;
        RECT 319.950 76.950 322.050 77.400 ;
        RECT 424.950 76.950 427.050 77.400 ;
        RECT 433.950 78.600 436.050 79.050 ;
        RECT 508.950 78.600 511.050 79.050 ;
        RECT 433.950 77.400 511.050 78.600 ;
        RECT 433.950 76.950 436.050 77.400 ;
        RECT 508.950 76.950 511.050 77.400 ;
        RECT 550.950 78.600 553.050 79.050 ;
        RECT 565.950 78.600 568.050 79.050 ;
        RECT 550.950 77.400 568.050 78.600 ;
        RECT 550.950 76.950 553.050 77.400 ;
        RECT 565.950 76.950 568.050 77.400 ;
        RECT 610.950 78.600 613.050 79.050 ;
        RECT 703.950 78.600 706.050 79.050 ;
        RECT 610.950 77.400 706.050 78.600 ;
        RECT 610.950 76.950 613.050 77.400 ;
        RECT 703.950 76.950 706.050 77.400 ;
        RECT 718.950 78.600 721.050 79.050 ;
        RECT 841.950 78.600 844.050 79.050 ;
        RECT 718.950 77.400 844.050 78.600 ;
        RECT 718.950 76.950 721.050 77.400 ;
        RECT 841.950 76.950 844.050 77.400 ;
        RECT 76.950 75.600 79.050 76.050 ;
        RECT 130.950 75.600 133.050 76.050 ;
        RECT 76.950 74.400 133.050 75.600 ;
        RECT 76.950 73.950 79.050 74.400 ;
        RECT 130.950 73.950 133.050 74.400 ;
        RECT 178.950 75.600 181.050 76.050 ;
        RECT 211.950 75.600 214.050 76.050 ;
        RECT 178.950 74.400 214.050 75.600 ;
        RECT 178.950 73.950 181.050 74.400 ;
        RECT 211.950 73.950 214.050 74.400 ;
        RECT 382.950 75.600 385.050 76.050 ;
        RECT 412.950 75.600 415.050 76.050 ;
        RECT 382.950 74.400 415.050 75.600 ;
        RECT 382.950 73.950 385.050 74.400 ;
        RECT 412.950 73.950 415.050 74.400 ;
        RECT 427.950 75.600 430.050 76.050 ;
        RECT 523.950 75.600 526.050 76.050 ;
        RECT 427.950 74.400 526.050 75.600 ;
        RECT 427.950 73.950 430.050 74.400 ;
        RECT 523.950 73.950 526.050 74.400 ;
        RECT 532.950 75.600 535.050 76.050 ;
        RECT 580.950 75.600 583.050 76.050 ;
        RECT 532.950 74.400 583.050 75.600 ;
        RECT 532.950 73.950 535.050 74.400 ;
        RECT 580.950 73.950 583.050 74.400 ;
        RECT 598.950 75.600 601.050 76.050 ;
        RECT 604.950 75.600 607.050 76.050 ;
        RECT 826.950 75.600 829.050 76.050 ;
        RECT 598.950 74.400 607.050 75.600 ;
        RECT 598.950 73.950 601.050 74.400 ;
        RECT 604.950 73.950 607.050 74.400 ;
        RECT 617.400 74.400 829.050 75.600 ;
        RECT 40.950 72.600 43.050 73.050 ;
        RECT 49.950 72.600 52.050 73.050 ;
        RECT 40.950 71.400 52.050 72.600 ;
        RECT 40.950 70.950 43.050 71.400 ;
        RECT 49.950 70.950 52.050 71.400 ;
        RECT 70.950 72.600 73.050 73.050 ;
        RECT 127.950 72.600 130.050 73.050 ;
        RECT 70.950 71.400 130.050 72.600 ;
        RECT 70.950 70.950 73.050 71.400 ;
        RECT 127.950 70.950 130.050 71.400 ;
        RECT 139.950 72.600 142.050 73.050 ;
        RECT 175.950 72.600 178.050 73.050 ;
        RECT 268.950 72.600 271.050 73.050 ;
        RECT 550.950 72.600 553.050 73.050 ;
        RECT 617.400 72.600 618.600 74.400 ;
        RECT 826.950 73.950 829.050 74.400 ;
        RECT 889.950 75.600 892.050 76.050 ;
        RECT 928.950 75.600 931.050 76.050 ;
        RECT 889.950 74.400 931.050 75.600 ;
        RECT 889.950 73.950 892.050 74.400 ;
        RECT 928.950 73.950 931.050 74.400 ;
        RECT 139.950 71.400 178.050 72.600 ;
        RECT 139.950 70.950 142.050 71.400 ;
        RECT 175.950 70.950 178.050 71.400 ;
        RECT 185.400 71.400 267.600 72.600 ;
        RECT 163.950 69.600 166.050 70.050 ;
        RECT 185.400 69.600 186.600 71.400 ;
        RECT 163.950 68.400 186.600 69.600 ;
        RECT 266.400 69.600 267.600 71.400 ;
        RECT 268.950 71.400 408.600 72.600 ;
        RECT 268.950 70.950 271.050 71.400 ;
        RECT 407.400 70.050 408.600 71.400 ;
        RECT 550.950 71.400 618.600 72.600 ;
        RECT 619.950 72.600 622.050 73.050 ;
        RECT 640.950 72.600 643.050 73.050 ;
        RECT 853.950 72.600 856.050 73.050 ;
        RECT 619.950 71.400 643.050 72.600 ;
        RECT 550.950 70.950 553.050 71.400 ;
        RECT 619.950 70.950 622.050 71.400 ;
        RECT 640.950 70.950 643.050 71.400 ;
        RECT 704.400 71.400 856.050 72.600 ;
        RECT 331.950 69.600 334.050 70.050 ;
        RECT 266.400 68.400 334.050 69.600 ;
        RECT 163.950 67.950 166.050 68.400 ;
        RECT 331.950 67.950 334.050 68.400 ;
        RECT 340.950 69.600 343.050 70.050 ;
        RECT 346.950 69.600 349.050 70.050 ;
        RECT 355.950 69.600 358.050 70.050 ;
        RECT 340.950 68.400 358.050 69.600 ;
        RECT 340.950 67.950 343.050 68.400 ;
        RECT 346.950 67.950 349.050 68.400 ;
        RECT 355.950 67.950 358.050 68.400 ;
        RECT 406.950 69.600 409.050 70.050 ;
        RECT 442.950 69.600 445.050 70.050 ;
        RECT 454.950 69.600 457.050 70.050 ;
        RECT 406.950 68.400 457.050 69.600 ;
        RECT 406.950 67.950 409.050 68.400 ;
        RECT 442.950 67.950 445.050 68.400 ;
        RECT 454.950 67.950 457.050 68.400 ;
        RECT 589.950 69.600 592.050 70.050 ;
        RECT 704.400 69.600 705.600 71.400 ;
        RECT 853.950 70.950 856.050 71.400 ;
        RECT 589.950 68.400 705.600 69.600 ;
        RECT 862.950 69.600 865.050 70.050 ;
        RECT 901.950 69.600 904.050 70.050 ;
        RECT 862.950 68.400 904.050 69.600 ;
        RECT 589.950 67.950 592.050 68.400 ;
        RECT 862.950 67.950 865.050 68.400 ;
        RECT 901.950 67.950 904.050 68.400 ;
        RECT 58.950 66.600 61.050 67.050 ;
        RECT 103.950 66.600 106.050 67.050 ;
        RECT 124.800 66.600 126.900 67.050 ;
        RECT 58.950 65.400 126.900 66.600 ;
        RECT 58.950 64.950 61.050 65.400 ;
        RECT 103.950 64.950 106.050 65.400 ;
        RECT 124.800 64.950 126.900 65.400 ;
        RECT 127.950 66.600 130.050 67.050 ;
        RECT 154.950 66.600 157.050 67.050 ;
        RECT 127.950 65.400 157.050 66.600 ;
        RECT 127.950 64.950 130.050 65.400 ;
        RECT 154.950 64.950 157.050 65.400 ;
        RECT 160.950 66.600 163.050 66.900 ;
        RECT 178.950 66.600 181.050 67.050 ;
        RECT 160.950 65.400 181.050 66.600 ;
        RECT 160.950 64.800 163.050 65.400 ;
        RECT 178.950 64.950 181.050 65.400 ;
        RECT 208.950 66.600 211.050 67.050 ;
        RECT 217.950 66.600 220.050 67.050 ;
        RECT 247.950 66.600 250.050 67.050 ;
        RECT 208.950 65.400 250.050 66.600 ;
        RECT 208.950 64.950 211.050 65.400 ;
        RECT 217.950 64.950 220.050 65.400 ;
        RECT 247.950 64.950 250.050 65.400 ;
        RECT 334.950 66.600 337.050 67.050 ;
        RECT 367.950 66.600 370.050 67.050 ;
        RECT 391.950 66.600 394.050 67.050 ;
        RECT 334.950 65.400 394.050 66.600 ;
        RECT 334.950 64.950 337.050 65.400 ;
        RECT 367.950 64.950 370.050 65.400 ;
        RECT 391.950 64.950 394.050 65.400 ;
        RECT 475.950 66.600 478.050 67.050 ;
        RECT 535.950 66.600 538.050 67.050 ;
        RECT 475.950 65.400 538.050 66.600 ;
        RECT 475.950 64.950 478.050 65.400 ;
        RECT 535.950 64.950 538.050 65.400 ;
        RECT 649.950 66.600 652.050 67.050 ;
        RECT 670.950 66.600 673.050 67.050 ;
        RECT 649.950 65.400 673.050 66.600 ;
        RECT 649.950 64.950 652.050 65.400 ;
        RECT 670.950 64.950 673.050 65.400 ;
        RECT 682.950 66.600 685.050 67.050 ;
        RECT 706.950 66.600 709.050 67.050 ;
        RECT 769.950 66.600 772.050 67.050 ;
        RECT 682.950 65.400 772.050 66.600 ;
        RECT 682.950 64.950 685.050 65.400 ;
        RECT 706.950 64.950 709.050 65.400 ;
        RECT 769.950 64.950 772.050 65.400 ;
        RECT 253.950 63.600 256.050 64.050 ;
        RECT 292.950 63.600 295.050 64.050 ;
        RECT 301.950 63.600 304.050 64.050 ;
        RECT 316.950 63.600 319.050 64.050 ;
        RECT 331.950 63.600 334.050 64.050 ;
        RECT 469.950 63.600 472.050 64.200 ;
        RECT 556.950 63.600 559.050 64.050 ;
        RECT 253.950 62.400 334.050 63.600 ;
        RECT 253.950 61.950 256.050 62.400 ;
        RECT 292.950 61.950 295.050 62.400 ;
        RECT 301.950 61.950 304.050 62.400 ;
        RECT 316.950 61.950 319.050 62.400 ;
        RECT 331.950 61.950 334.050 62.400 ;
        RECT 347.400 62.400 357.600 63.600 ;
        RECT 22.950 60.750 25.050 61.200 ;
        RECT 52.950 60.750 55.050 61.200 ;
        RECT 22.950 59.550 55.050 60.750 ;
        RECT 22.950 59.100 25.050 59.550 ;
        RECT 52.950 59.100 55.050 59.550 ;
        RECT 58.950 59.100 61.050 61.200 ;
        RECT 76.950 60.600 79.050 61.200 ;
        RECT 62.400 59.400 79.050 60.600 ;
        RECT 59.400 57.600 60.600 59.100 ;
        RECT 44.400 57.000 60.600 57.600 ;
        RECT 43.950 56.400 60.600 57.000 ;
        RECT 43.950 52.950 46.050 56.400 ;
        RECT 62.400 54.900 63.600 59.400 ;
        RECT 76.950 59.100 79.050 59.400 ;
        RECT 82.950 59.100 85.050 61.200 ;
        RECT 94.950 60.750 97.050 61.200 ;
        RECT 109.950 60.750 112.050 61.200 ;
        RECT 94.950 59.550 112.050 60.750 ;
        RECT 94.950 59.100 97.050 59.550 ;
        RECT 109.950 59.100 112.050 59.550 ;
        RECT 61.950 52.800 64.050 54.900 ;
        RECT 73.950 54.600 76.050 55.050 ;
        RECT 83.400 54.600 84.600 59.100 ;
        RECT 139.950 58.950 142.050 61.050 ;
        RECT 160.950 60.600 163.050 60.900 ;
        RECT 175.950 60.600 178.050 61.200 ;
        RECT 181.950 60.600 184.050 61.050 ;
        RECT 160.950 59.400 184.050 60.600 ;
        RECT 73.950 53.400 84.600 54.600 ;
        RECT 85.950 54.600 88.050 54.900 ;
        RECT 91.950 54.600 94.050 55.050 ;
        RECT 85.950 53.400 94.050 54.600 ;
        RECT 73.950 52.950 76.050 53.400 ;
        RECT 85.950 52.800 88.050 53.400 ;
        RECT 91.950 52.950 94.050 53.400 ;
        RECT 106.950 54.600 109.050 54.900 ;
        RECT 115.950 54.600 118.050 55.050 ;
        RECT 106.950 53.400 118.050 54.600 ;
        RECT 106.950 52.800 109.050 53.400 ;
        RECT 115.950 52.950 118.050 53.400 ;
        RECT 127.950 54.600 130.050 54.900 ;
        RECT 140.400 54.600 141.600 58.950 ;
        RECT 160.950 58.800 163.050 59.400 ;
        RECT 175.950 59.100 178.050 59.400 ;
        RECT 181.950 58.950 184.050 59.400 ;
        RECT 190.950 59.100 193.050 61.200 ;
        RECT 196.950 60.600 199.050 61.200 ;
        RECT 202.950 60.600 205.050 61.050 ;
        RECT 196.950 59.400 205.050 60.600 ;
        RECT 196.950 59.100 199.050 59.400 ;
        RECT 191.400 55.050 192.600 59.100 ;
        RECT 127.950 53.400 141.600 54.600 ;
        RECT 148.950 54.450 151.050 54.900 ;
        RECT 160.950 54.450 163.050 54.900 ;
        RECT 127.950 52.800 130.050 53.400 ;
        RECT 148.950 53.250 163.050 54.450 ;
        RECT 148.950 52.800 151.050 53.250 ;
        RECT 160.950 52.800 163.050 53.250 ;
        RECT 172.950 54.600 175.050 54.900 ;
        RECT 178.950 54.600 181.050 55.050 ;
        RECT 172.950 53.400 181.050 54.600 ;
        RECT 172.950 52.800 175.050 53.400 ;
        RECT 178.950 52.950 181.050 53.400 ;
        RECT 187.950 53.400 192.600 55.050 ;
        RECT 187.950 52.950 192.000 53.400 ;
        RECT 16.950 51.600 19.050 52.050 ;
        RECT 31.950 51.600 34.050 52.050 ;
        RECT 46.950 51.600 49.050 52.050 ;
        RECT 16.950 50.400 49.050 51.600 ;
        RECT 16.950 49.950 19.050 50.400 ;
        RECT 31.950 49.950 34.050 50.400 ;
        RECT 46.950 49.950 49.050 50.400 ;
        RECT 118.950 51.600 121.050 52.050 ;
        RECT 184.950 51.600 187.050 52.050 ;
        RECT 193.950 51.600 196.050 52.050 ;
        RECT 118.950 50.400 147.600 51.600 ;
        RECT 118.950 49.950 121.050 50.400 ;
        RECT 37.950 48.600 40.050 49.050 ;
        RECT 49.950 48.600 52.050 49.050 ;
        RECT 37.950 47.400 52.050 48.600 ;
        RECT 37.950 46.950 40.050 47.400 ;
        RECT 49.950 46.950 52.050 47.400 ;
        RECT 64.950 48.600 67.050 49.050 ;
        RECT 73.950 48.600 76.050 49.050 ;
        RECT 142.950 48.600 145.050 49.050 ;
        RECT 64.950 47.400 145.050 48.600 ;
        RECT 146.400 48.600 147.600 50.400 ;
        RECT 184.950 50.400 196.050 51.600 ;
        RECT 184.950 49.950 187.050 50.400 ;
        RECT 193.950 49.950 196.050 50.400 ;
        RECT 178.950 48.600 181.050 49.050 ;
        RECT 197.400 48.600 198.600 59.100 ;
        RECT 202.950 58.950 205.050 59.400 ;
        RECT 211.950 57.600 214.050 61.050 ;
        RECT 223.950 60.600 226.050 61.200 ;
        RECT 229.950 60.750 232.050 61.200 ;
        RECT 235.950 60.750 238.050 61.200 ;
        RECT 229.950 60.600 238.050 60.750 ;
        RECT 223.950 59.550 238.050 60.600 ;
        RECT 223.950 59.400 232.050 59.550 ;
        RECT 223.950 59.100 226.050 59.400 ;
        RECT 229.950 59.100 232.050 59.400 ;
        RECT 235.950 59.100 238.050 59.550 ;
        RECT 241.950 60.600 244.050 61.050 ;
        RECT 247.950 60.600 250.050 61.050 ;
        RECT 241.950 59.400 250.050 60.600 ;
        RECT 241.950 58.950 244.050 59.400 ;
        RECT 247.950 58.950 250.050 59.400 ;
        RECT 259.950 60.750 262.050 61.200 ;
        RECT 271.950 60.750 274.050 61.200 ;
        RECT 259.950 59.550 274.050 60.750 ;
        RECT 277.950 60.600 280.050 61.200 ;
        RECT 259.950 59.100 262.050 59.550 ;
        RECT 271.950 59.100 274.050 59.550 ;
        RECT 275.400 59.400 280.050 60.600 ;
        RECT 211.950 57.000 216.600 57.600 ;
        RECT 212.400 56.400 216.600 57.000 ;
        RECT 215.400 54.900 216.600 56.400 ;
        RECT 275.400 55.050 276.600 59.400 ;
        RECT 277.950 59.100 280.050 59.400 ;
        RECT 283.950 60.600 286.050 61.200 ;
        RECT 289.950 60.600 292.050 61.050 ;
        RECT 283.950 59.400 292.050 60.600 ;
        RECT 283.950 59.100 286.050 59.400 ;
        RECT 289.950 58.950 292.050 59.400 ;
        RECT 310.950 58.950 313.050 61.050 ;
        RECT 319.950 58.950 322.050 61.050 ;
        RECT 325.950 60.750 328.050 61.200 ;
        RECT 340.950 60.750 343.050 61.200 ;
        RECT 325.950 59.550 343.050 60.750 ;
        RECT 347.400 60.600 348.600 62.400 ;
        RECT 325.950 59.100 328.050 59.550 ;
        RECT 340.950 59.100 343.050 59.550 ;
        RECT 344.400 59.400 348.600 60.600 ;
        RECT 199.950 54.450 202.050 54.900 ;
        RECT 205.950 54.450 208.050 54.900 ;
        RECT 199.950 53.250 208.050 54.450 ;
        RECT 199.950 52.800 202.050 53.250 ;
        RECT 205.950 52.800 208.050 53.250 ;
        RECT 214.950 52.800 217.050 54.900 ;
        RECT 244.950 54.600 247.050 55.050 ;
        RECT 262.950 54.600 265.050 54.900 ;
        RECT 244.950 53.400 265.050 54.600 ;
        RECT 244.950 52.950 247.050 53.400 ;
        RECT 262.950 52.800 265.050 53.400 ;
        RECT 274.950 52.950 277.050 55.050 ;
        RECT 301.950 54.600 304.050 54.900 ;
        RECT 311.400 54.600 312.600 58.950 ;
        RECT 320.400 55.050 321.600 58.950 ;
        RECT 344.400 57.600 345.600 59.400 ;
        RECT 352.950 59.100 355.050 61.200 ;
        RECT 356.400 60.600 357.600 62.400 ;
        RECT 469.950 62.400 559.050 63.600 ;
        RECT 469.950 62.100 472.050 62.400 ;
        RECT 556.950 61.950 559.050 62.400 ;
        RECT 625.950 63.600 628.050 64.050 ;
        RECT 631.950 63.600 634.050 64.050 ;
        RECT 646.950 63.600 649.050 64.050 ;
        RECT 625.950 62.400 649.050 63.600 ;
        RECT 625.950 61.950 628.050 62.400 ;
        RECT 631.950 61.950 634.050 62.400 ;
        RECT 646.950 61.950 649.050 62.400 ;
        RECT 790.950 63.600 793.050 64.050 ;
        RECT 811.950 63.600 814.050 64.050 ;
        RECT 790.950 62.400 814.050 63.600 ;
        RECT 790.950 61.950 793.050 62.400 ;
        RECT 811.950 61.950 814.050 62.400 ;
        RECT 856.950 63.600 859.050 64.050 ;
        RECT 868.950 63.600 871.050 64.050 ;
        RECT 856.950 62.400 871.050 63.600 ;
        RECT 856.950 61.950 859.050 62.400 ;
        RECT 868.950 61.950 871.050 62.400 ;
        RECT 907.950 63.600 910.050 64.050 ;
        RECT 919.950 63.600 922.050 64.050 ;
        RECT 934.950 63.600 937.050 64.050 ;
        RECT 907.950 62.400 937.050 63.600 ;
        RECT 907.950 61.950 910.050 62.400 ;
        RECT 919.950 61.950 922.050 62.400 ;
        RECT 934.950 61.950 937.050 62.400 ;
        RECT 373.950 60.750 376.050 61.200 ;
        RECT 382.950 60.750 385.050 61.200 ;
        RECT 356.400 59.400 369.600 60.600 ;
        RECT 341.400 57.000 345.600 57.600 ;
        RECT 340.950 56.400 345.600 57.000 ;
        RECT 301.950 53.400 312.600 54.600 ;
        RECT 301.950 52.800 304.050 53.400 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 328.950 54.600 331.050 54.900 ;
        RECT 337.800 54.600 339.900 55.050 ;
        RECT 328.950 53.400 339.900 54.600 ;
        RECT 328.950 52.800 331.050 53.400 ;
        RECT 337.800 52.950 339.900 53.400 ;
        RECT 340.950 52.950 343.050 56.400 ;
        RECT 353.400 54.600 354.600 59.100 ;
        RECT 368.400 57.600 369.600 59.400 ;
        RECT 373.950 59.550 385.050 60.750 ;
        RECT 373.950 59.100 376.050 59.550 ;
        RECT 382.950 59.100 385.050 59.550 ;
        RECT 397.950 60.750 400.050 61.200 ;
        RECT 403.950 60.750 406.050 61.200 ;
        RECT 397.950 59.550 406.050 60.750 ;
        RECT 397.950 59.100 400.050 59.550 ;
        RECT 403.950 59.100 406.050 59.550 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 436.950 60.750 439.050 61.200 ;
        RECT 448.800 60.750 450.900 61.200 ;
        RECT 436.950 60.600 450.900 60.750 ;
        RECT 425.400 59.550 450.900 60.600 ;
        RECT 425.400 59.400 439.050 59.550 ;
        RECT 406.950 57.600 409.050 58.050 ;
        RECT 419.400 57.600 420.600 59.100 ;
        RECT 425.400 57.600 426.600 59.400 ;
        RECT 436.950 59.100 439.050 59.400 ;
        RECT 448.800 59.100 450.900 59.550 ;
        RECT 451.950 60.750 454.050 61.200 ;
        RECT 460.950 60.750 463.050 61.200 ;
        RECT 451.950 59.550 463.050 60.750 ;
        RECT 451.950 59.100 454.050 59.550 ;
        RECT 460.950 59.100 463.050 59.550 ;
        RECT 466.950 58.950 469.050 61.050 ;
        RECT 478.950 60.750 481.050 61.200 ;
        RECT 487.950 60.750 490.050 61.200 ;
        RECT 478.950 60.600 490.050 60.750 ;
        RECT 508.950 60.600 511.050 61.200 ;
        RECT 478.950 59.550 511.050 60.600 ;
        RECT 478.950 59.100 481.050 59.550 ;
        RECT 487.950 59.400 511.050 59.550 ;
        RECT 487.950 59.100 490.050 59.400 ;
        RECT 508.950 59.100 511.050 59.400 ;
        RECT 514.950 60.600 517.050 61.200 ;
        RECT 529.950 60.600 532.050 61.200 ;
        RECT 553.950 60.600 556.050 61.200 ;
        RECT 514.950 59.400 556.050 60.600 ;
        RECT 514.950 59.100 517.050 59.400 ;
        RECT 529.950 59.100 532.050 59.400 ;
        RECT 553.950 59.100 556.050 59.400 ;
        RECT 562.950 60.750 565.050 61.200 ;
        RECT 574.950 60.750 577.050 61.200 ;
        RECT 562.950 59.550 577.050 60.750 ;
        RECT 562.950 59.100 565.050 59.550 ;
        RECT 574.950 59.100 577.050 59.550 ;
        RECT 592.950 60.750 595.050 61.200 ;
        RECT 619.950 60.750 622.050 61.200 ;
        RECT 592.950 59.550 622.050 60.750 ;
        RECT 592.950 59.100 595.050 59.550 ;
        RECT 619.950 59.100 622.050 59.550 ;
        RECT 658.950 59.100 661.050 61.200 ;
        RECT 664.950 60.750 667.050 61.200 ;
        RECT 673.950 60.750 676.050 61.200 ;
        RECT 664.950 59.550 676.050 60.750 ;
        RECT 664.950 59.100 667.050 59.550 ;
        RECT 673.950 59.100 676.050 59.550 ;
        RECT 688.950 60.750 691.050 61.200 ;
        RECT 700.950 60.750 703.050 61.200 ;
        RECT 688.950 59.550 703.050 60.750 ;
        RECT 688.950 59.100 691.050 59.550 ;
        RECT 700.950 59.100 703.050 59.550 ;
        RECT 712.950 60.600 715.050 61.200 ;
        RECT 736.950 60.600 739.050 61.200 ;
        RECT 748.950 60.600 751.050 61.200 ;
        RECT 712.950 59.400 751.050 60.600 ;
        RECT 712.950 59.100 715.050 59.400 ;
        RECT 736.950 59.100 739.050 59.400 ;
        RECT 748.950 59.100 751.050 59.400 ;
        RECT 757.950 60.750 760.050 61.200 ;
        RECT 763.950 60.750 766.050 61.200 ;
        RECT 757.950 59.550 766.050 60.750 ;
        RECT 757.950 59.100 760.050 59.550 ;
        RECT 763.950 59.100 766.050 59.550 ;
        RECT 784.950 60.600 787.050 61.200 ;
        RECT 805.950 60.600 808.050 61.200 ;
        RECT 784.950 59.400 808.050 60.600 ;
        RECT 784.950 59.100 787.050 59.400 ;
        RECT 805.950 59.100 808.050 59.400 ;
        RECT 832.950 59.100 835.050 61.200 ;
        RECT 844.950 60.750 847.050 61.200 ;
        RECT 859.950 60.750 862.050 61.200 ;
        RECT 844.950 59.550 862.050 60.750 ;
        RECT 844.950 59.100 847.050 59.550 ;
        RECT 859.950 59.100 862.050 59.550 ;
        RECT 368.400 56.400 372.600 57.600 ;
        RECT 364.950 54.600 367.050 54.900 ;
        RECT 353.400 53.400 367.050 54.600 ;
        RECT 371.400 54.600 372.600 56.400 ;
        RECT 406.950 56.400 420.600 57.600 ;
        RECT 422.400 56.400 426.600 57.600 ;
        RECT 406.950 55.950 409.050 56.400 ;
        RECT 376.950 54.600 379.050 55.050 ;
        RECT 371.400 53.400 379.050 54.600 ;
        RECT 364.950 52.800 367.050 53.400 ;
        RECT 376.950 52.950 379.050 53.400 ;
        RECT 382.950 54.600 385.050 55.050 ;
        RECT 394.950 54.600 397.050 54.900 ;
        RECT 382.950 53.400 397.050 54.600 ;
        RECT 382.950 52.950 385.050 53.400 ;
        RECT 394.950 52.800 397.050 53.400 ;
        RECT 403.950 54.600 406.050 55.050 ;
        RECT 415.950 54.600 418.050 54.900 ;
        RECT 422.400 54.600 423.600 56.400 ;
        RECT 403.950 53.400 418.050 54.600 ;
        RECT 419.400 54.000 423.600 54.600 ;
        RECT 403.950 52.950 406.050 53.400 ;
        RECT 415.950 52.800 418.050 53.400 ;
        RECT 418.950 53.400 423.600 54.000 ;
        RECT 427.950 54.450 430.050 54.900 ;
        RECT 439.950 54.600 442.050 54.900 ;
        RECT 451.800 54.600 453.900 55.050 ;
        RECT 439.950 54.450 453.900 54.600 ;
        RECT 427.950 53.400 453.900 54.450 ;
        RECT 206.400 51.600 207.600 52.800 ;
        RECT 238.950 51.600 241.050 52.050 ;
        RECT 206.400 50.400 241.050 51.600 ;
        RECT 238.950 49.950 241.050 50.400 ;
        RECT 316.950 51.600 319.050 52.050 ;
        RECT 343.950 51.600 346.050 52.050 ;
        RECT 316.950 50.400 346.050 51.600 ;
        RECT 316.950 49.950 319.050 50.400 ;
        RECT 343.950 49.950 346.050 50.400 ;
        RECT 418.950 49.950 421.050 53.400 ;
        RECT 427.950 53.250 442.050 53.400 ;
        RECT 427.950 52.800 430.050 53.250 ;
        RECT 439.950 52.800 442.050 53.250 ;
        RECT 451.800 52.950 453.900 53.400 ;
        RECT 454.950 54.450 457.050 54.900 ;
        RECT 463.950 54.450 466.050 54.900 ;
        RECT 454.950 53.250 466.050 54.450 ;
        RECT 454.950 52.800 457.050 53.250 ;
        RECT 463.950 52.800 466.050 53.250 ;
        RECT 467.400 52.050 468.600 58.950 ;
        RECT 475.950 54.450 478.050 54.900 ;
        RECT 484.950 54.450 487.050 54.900 ;
        RECT 475.950 53.250 487.050 54.450 ;
        RECT 475.950 52.800 478.050 53.250 ;
        RECT 484.950 52.800 487.050 53.250 ;
        RECT 490.950 54.600 493.050 54.900 ;
        RECT 511.950 54.600 514.050 54.900 ;
        RECT 520.950 54.600 523.050 55.050 ;
        RECT 490.950 54.000 498.600 54.600 ;
        RECT 490.950 53.400 499.050 54.000 ;
        RECT 490.950 52.800 493.050 53.400 ;
        RECT 466.950 49.950 469.050 52.050 ;
        RECT 496.950 49.950 499.050 53.400 ;
        RECT 511.950 53.400 523.050 54.600 ;
        RECT 511.950 52.800 514.050 53.400 ;
        RECT 520.950 52.950 523.050 53.400 ;
        RECT 526.950 54.600 529.050 55.050 ;
        RECT 544.950 54.600 547.050 55.050 ;
        RECT 526.950 53.400 547.050 54.600 ;
        RECT 526.950 52.950 529.050 53.400 ;
        RECT 544.950 52.950 547.050 53.400 ;
        RECT 565.950 54.450 568.050 54.900 ;
        RECT 571.950 54.450 574.050 54.900 ;
        RECT 565.950 53.250 574.050 54.450 ;
        RECT 565.950 52.800 568.050 53.250 ;
        RECT 571.950 52.800 574.050 53.250 ;
        RECT 577.950 54.600 580.050 54.900 ;
        RECT 589.950 54.600 592.050 55.050 ;
        RECT 577.950 53.400 592.050 54.600 ;
        RECT 577.950 52.800 580.050 53.400 ;
        RECT 589.950 52.950 592.050 53.400 ;
        RECT 601.950 54.450 604.050 54.900 ;
        RECT 610.950 54.450 613.050 54.900 ;
        RECT 601.950 53.250 613.050 54.450 ;
        RECT 601.950 52.800 604.050 53.250 ;
        RECT 610.950 52.800 613.050 53.250 ;
        RECT 631.950 54.450 634.050 54.900 ;
        RECT 643.950 54.450 646.050 54.900 ;
        RECT 631.950 53.250 646.050 54.450 ;
        RECT 659.400 54.600 660.600 59.100 ;
        RECT 833.400 57.600 834.600 59.100 ;
        RECT 871.950 58.950 874.050 61.050 ;
        RECT 877.950 60.600 880.050 61.050 ;
        RECT 886.950 60.600 889.050 61.050 ;
        RECT 877.950 59.400 889.050 60.600 ;
        RECT 877.950 58.950 880.050 59.400 ;
        RECT 886.950 58.950 889.050 59.400 ;
        RECT 898.950 59.100 901.050 61.200 ;
        RECT 925.950 59.100 928.050 61.200 ;
        RECT 865.950 57.600 868.050 58.050 ;
        RECT 818.400 56.400 834.600 57.600 ;
        RECT 854.400 56.400 868.050 57.600 ;
        RECT 679.950 54.600 682.050 54.900 ;
        RECT 659.400 53.400 682.050 54.600 ;
        RECT 631.950 52.800 634.050 53.250 ;
        RECT 643.950 52.800 646.050 53.250 ;
        RECT 679.950 52.800 682.050 53.400 ;
        RECT 685.950 54.450 688.050 54.900 ;
        RECT 694.950 54.600 697.050 54.900 ;
        RECT 709.950 54.600 712.050 54.900 ;
        RECT 694.950 54.450 712.050 54.600 ;
        RECT 685.950 53.400 712.050 54.450 ;
        RECT 685.950 53.250 697.050 53.400 ;
        RECT 685.950 52.800 688.050 53.250 ;
        RECT 694.950 52.800 697.050 53.250 ;
        RECT 709.950 52.800 712.050 53.400 ;
        RECT 721.950 54.450 724.050 54.900 ;
        RECT 733.950 54.450 736.050 54.900 ;
        RECT 721.950 53.250 736.050 54.450 ;
        RECT 721.950 52.800 724.050 53.250 ;
        RECT 733.950 52.800 736.050 53.250 ;
        RECT 742.950 54.450 745.050 54.900 ;
        RECT 751.950 54.450 754.050 54.900 ;
        RECT 742.950 53.250 754.050 54.450 ;
        RECT 742.950 52.800 745.050 53.250 ;
        RECT 751.950 52.800 754.050 53.250 ;
        RECT 787.950 54.450 790.050 54.900 ;
        RECT 799.950 54.450 802.050 54.900 ;
        RECT 787.950 53.250 802.050 54.450 ;
        RECT 787.950 52.800 790.050 53.250 ;
        RECT 799.950 52.800 802.050 53.250 ;
        RECT 523.950 51.600 526.050 52.050 ;
        RECT 532.950 51.600 535.050 52.050 ;
        RECT 523.950 50.400 535.050 51.600 ;
        RECT 523.950 49.950 526.050 50.400 ;
        RECT 532.950 49.950 535.050 50.400 ;
        RECT 805.950 51.600 808.050 52.050 ;
        RECT 818.400 51.600 819.600 56.400 ;
        RECT 820.950 54.600 823.050 55.050 ;
        RECT 829.950 54.600 832.050 54.900 ;
        RECT 820.950 53.400 832.050 54.600 ;
        RECT 820.950 52.950 823.050 53.400 ;
        RECT 829.950 52.800 832.050 53.400 ;
        RECT 850.950 54.600 853.050 54.900 ;
        RECT 854.400 54.600 855.600 56.400 ;
        RECT 865.950 55.950 868.050 56.400 ;
        RECT 872.400 55.050 873.600 58.950 ;
        RECT 850.950 53.400 855.600 54.600 ;
        RECT 856.950 54.450 859.050 54.900 ;
        RECT 862.950 54.450 865.050 54.900 ;
        RECT 850.950 52.800 853.050 53.400 ;
        RECT 856.950 53.250 865.050 54.450 ;
        RECT 856.950 52.800 859.050 53.250 ;
        RECT 862.950 52.800 865.050 53.250 ;
        RECT 871.950 52.950 874.050 55.050 ;
        RECT 899.400 51.600 900.600 59.100 ;
        RECT 910.950 54.600 913.050 55.050 ;
        RECT 916.950 54.600 919.050 54.900 ;
        RECT 910.950 53.400 919.050 54.600 ;
        RECT 910.950 52.950 913.050 53.400 ;
        RECT 916.950 52.800 919.050 53.400 ;
        RECT 904.950 51.600 907.050 52.050 ;
        RECT 926.400 51.600 927.600 59.100 ;
        RECT 805.950 50.400 819.600 51.600 ;
        RECT 848.400 50.400 927.600 51.600 ;
        RECT 805.950 49.950 808.050 50.400 ;
        RECT 848.400 49.050 849.600 50.400 ;
        RECT 904.950 49.950 907.050 50.400 ;
        RECT 146.400 47.400 198.600 48.600 ;
        RECT 220.950 48.600 223.050 49.050 ;
        RECT 247.950 48.600 250.050 49.050 ;
        RECT 220.950 47.400 250.050 48.600 ;
        RECT 64.950 46.950 67.050 47.400 ;
        RECT 73.950 46.950 76.050 47.400 ;
        RECT 142.950 46.950 145.050 47.400 ;
        RECT 178.950 46.950 181.050 47.400 ;
        RECT 220.950 46.950 223.050 47.400 ;
        RECT 247.950 46.950 250.050 47.400 ;
        RECT 271.950 48.600 274.050 49.050 ;
        RECT 280.950 48.600 283.050 49.050 ;
        RECT 271.950 47.400 283.050 48.600 ;
        RECT 271.950 46.950 274.050 47.400 ;
        RECT 280.950 46.950 283.050 47.400 ;
        RECT 286.950 48.600 289.050 49.050 ;
        RECT 313.950 48.600 316.050 49.050 ;
        RECT 286.950 47.400 316.050 48.600 ;
        RECT 286.950 46.950 289.050 47.400 ;
        RECT 313.950 46.950 316.050 47.400 ;
        RECT 358.950 48.600 361.050 49.050 ;
        RECT 388.950 48.600 391.050 49.050 ;
        RECT 358.950 47.400 391.050 48.600 ;
        RECT 358.950 46.950 361.050 47.400 ;
        RECT 388.950 46.950 391.050 47.400 ;
        RECT 421.950 48.600 424.050 49.050 ;
        RECT 547.950 48.600 550.050 49.050 ;
        RECT 421.950 47.400 550.050 48.600 ;
        RECT 421.950 46.950 424.050 47.400 ;
        RECT 547.950 46.950 550.050 47.400 ;
        RECT 622.950 48.600 625.050 49.050 ;
        RECT 652.950 48.600 655.050 49.050 ;
        RECT 622.950 47.400 655.050 48.600 ;
        RECT 622.950 46.950 625.050 47.400 ;
        RECT 652.950 46.950 655.050 47.400 ;
        RECT 679.950 48.600 682.050 49.050 ;
        RECT 703.800 48.600 705.900 49.050 ;
        RECT 679.950 47.400 705.900 48.600 ;
        RECT 679.950 46.950 682.050 47.400 ;
        RECT 703.800 46.950 705.900 47.400 ;
        RECT 706.950 48.600 709.050 49.050 ;
        RECT 727.950 48.600 730.050 49.050 ;
        RECT 706.950 47.400 730.050 48.600 ;
        RECT 706.950 46.950 709.050 47.400 ;
        RECT 727.950 46.950 730.050 47.400 ;
        RECT 766.950 48.600 769.050 49.050 ;
        RECT 847.950 48.600 850.050 49.050 ;
        RECT 766.950 47.400 850.050 48.600 ;
        RECT 766.950 46.950 769.050 47.400 ;
        RECT 847.950 46.950 850.050 47.400 ;
        RECT 868.950 48.600 871.050 49.050 ;
        RECT 880.950 48.600 883.050 49.050 ;
        RECT 868.950 47.400 883.050 48.600 ;
        RECT 868.950 46.950 871.050 47.400 ;
        RECT 880.950 46.950 883.050 47.400 ;
        RECT 919.950 48.600 922.050 49.050 ;
        RECT 937.950 48.600 940.050 49.050 ;
        RECT 919.950 47.400 940.050 48.600 ;
        RECT 919.950 46.950 922.050 47.400 ;
        RECT 937.950 46.950 940.050 47.400 ;
        RECT 55.950 45.600 58.050 46.050 ;
        RECT 70.950 45.600 73.050 46.050 ;
        RECT 55.950 44.400 73.050 45.600 ;
        RECT 55.950 43.950 58.050 44.400 ;
        RECT 70.950 43.950 73.050 44.400 ;
        RECT 100.950 45.600 103.050 46.050 ;
        RECT 121.950 45.600 124.050 46.050 ;
        RECT 166.950 45.600 169.050 46.050 ;
        RECT 100.950 44.400 169.050 45.600 ;
        RECT 100.950 43.950 103.050 44.400 ;
        RECT 121.950 43.950 124.050 44.400 ;
        RECT 166.950 43.950 169.050 44.400 ;
        RECT 283.950 45.600 286.050 46.050 ;
        RECT 364.950 45.600 367.050 46.050 ;
        RECT 283.950 44.400 367.050 45.600 ;
        RECT 283.950 43.950 286.050 44.400 ;
        RECT 364.950 43.950 367.050 44.400 ;
        RECT 373.950 45.600 376.050 46.050 ;
        RECT 418.950 45.600 421.050 46.050 ;
        RECT 373.950 44.400 421.050 45.600 ;
        RECT 373.950 43.950 376.050 44.400 ;
        RECT 418.950 43.950 421.050 44.400 ;
        RECT 463.950 45.600 466.050 46.050 ;
        RECT 478.950 45.600 481.050 46.050 ;
        RECT 568.950 45.600 571.050 46.050 ;
        RECT 595.950 45.600 598.050 46.050 ;
        RECT 463.950 44.400 552.600 45.600 ;
        RECT 463.950 43.950 466.050 44.400 ;
        RECT 478.950 43.950 481.050 44.400 ;
        RECT 58.950 42.600 61.050 43.050 ;
        RECT 67.950 42.600 70.050 43.050 ;
        RECT 58.950 41.400 70.050 42.600 ;
        RECT 58.950 40.950 61.050 41.400 ;
        RECT 67.950 40.950 70.050 41.400 ;
        RECT 196.950 42.600 199.050 43.050 ;
        RECT 217.950 42.600 220.050 43.050 ;
        RECT 196.950 41.400 220.050 42.600 ;
        RECT 196.950 40.950 199.050 41.400 ;
        RECT 217.950 40.950 220.050 41.400 ;
        RECT 280.950 42.600 283.050 43.050 ;
        RECT 358.950 42.600 361.050 43.050 ;
        RECT 421.950 42.600 424.050 43.050 ;
        RECT 280.950 41.400 424.050 42.600 ;
        RECT 280.950 40.950 283.050 41.400 ;
        RECT 358.950 40.950 361.050 41.400 ;
        RECT 421.950 40.950 424.050 41.400 ;
        RECT 484.950 42.600 487.050 43.050 ;
        RECT 505.950 42.600 508.050 43.050 ;
        RECT 484.950 41.400 508.050 42.600 ;
        RECT 484.950 40.950 487.050 41.400 ;
        RECT 505.950 40.950 508.050 41.400 ;
        RECT 517.950 42.600 520.050 43.050 ;
        RECT 551.400 42.600 552.600 44.400 ;
        RECT 568.950 44.400 598.050 45.600 ;
        RECT 568.950 43.950 571.050 44.400 ;
        RECT 595.950 43.950 598.050 44.400 ;
        RECT 673.950 45.600 676.050 46.050 ;
        RECT 700.800 45.600 702.900 46.050 ;
        RECT 673.950 44.400 702.900 45.600 ;
        RECT 704.400 45.600 705.600 46.950 ;
        RECT 757.800 45.600 759.900 46.050 ;
        RECT 704.400 44.400 759.900 45.600 ;
        RECT 673.950 43.950 676.050 44.400 ;
        RECT 700.800 43.950 702.900 44.400 ;
        RECT 757.800 43.950 759.900 44.400 ;
        RECT 760.950 45.600 763.050 46.050 ;
        RECT 811.950 45.600 814.050 46.050 ;
        RECT 760.950 44.400 814.050 45.600 ;
        RECT 760.950 43.950 763.050 44.400 ;
        RECT 811.950 43.950 814.050 44.400 ;
        RECT 829.950 45.600 832.050 46.050 ;
        RECT 844.950 45.600 847.050 46.050 ;
        RECT 829.950 44.400 847.050 45.600 ;
        RECT 829.950 43.950 832.050 44.400 ;
        RECT 844.950 43.950 847.050 44.400 ;
        RECT 850.950 45.600 853.050 46.050 ;
        RECT 895.950 45.600 898.050 46.050 ;
        RECT 850.950 44.400 898.050 45.600 ;
        RECT 850.950 43.950 853.050 44.400 ;
        RECT 895.950 43.950 898.050 44.400 ;
        RECT 562.950 42.600 565.050 43.050 ;
        RECT 517.950 41.400 543.600 42.600 ;
        RECT 551.400 41.400 565.050 42.600 ;
        RECT 517.950 40.950 520.050 41.400 ;
        RECT 22.950 39.600 25.050 40.050 ;
        RECT 76.950 39.600 79.050 40.050 ;
        RECT 22.950 38.400 79.050 39.600 ;
        RECT 22.950 37.950 25.050 38.400 ;
        RECT 76.950 37.950 79.050 38.400 ;
        RECT 127.950 39.600 130.050 40.050 ;
        RECT 136.950 39.600 139.050 40.050 ;
        RECT 220.950 39.600 223.050 40.050 ;
        RECT 256.950 39.600 259.050 40.050 ;
        RECT 274.950 39.600 277.050 40.050 ;
        RECT 127.950 38.400 223.050 39.600 ;
        RECT 127.950 37.950 130.050 38.400 ;
        RECT 136.950 37.950 139.050 38.400 ;
        RECT 220.950 37.950 223.050 38.400 ;
        RECT 230.400 38.400 277.050 39.600 ;
        RECT 230.400 37.050 231.600 38.400 ;
        RECT 256.950 37.950 259.050 38.400 ;
        RECT 274.950 37.950 277.050 38.400 ;
        RECT 301.950 39.600 304.050 40.050 ;
        RECT 331.950 39.600 334.050 40.050 ;
        RECT 355.950 39.600 358.050 40.050 ;
        RECT 301.950 38.400 358.050 39.600 ;
        RECT 301.950 37.950 304.050 38.400 ;
        RECT 331.950 37.950 334.050 38.400 ;
        RECT 355.950 37.950 358.050 38.400 ;
        RECT 370.950 39.600 373.050 40.050 ;
        RECT 403.950 39.600 406.050 40.050 ;
        RECT 370.950 38.400 406.050 39.600 ;
        RECT 370.950 37.950 373.050 38.400 ;
        RECT 403.950 37.950 406.050 38.400 ;
        RECT 418.950 39.600 421.050 40.050 ;
        RECT 424.950 39.600 427.050 40.050 ;
        RECT 418.950 38.400 427.050 39.600 ;
        RECT 418.950 37.950 421.050 38.400 ;
        RECT 424.950 37.950 427.050 38.400 ;
        RECT 478.950 39.600 481.050 40.050 ;
        RECT 542.400 39.600 543.600 41.400 ;
        RECT 562.950 40.950 565.050 41.400 ;
        RECT 688.950 42.600 691.050 43.050 ;
        RECT 901.950 42.600 904.050 43.050 ;
        RECT 913.950 42.600 916.050 43.050 ;
        RECT 922.950 42.600 925.050 43.050 ;
        RECT 688.950 41.400 925.050 42.600 ;
        RECT 688.950 40.950 691.050 41.400 ;
        RECT 901.950 40.950 904.050 41.400 ;
        RECT 913.950 40.950 916.050 41.400 ;
        RECT 922.950 40.950 925.050 41.400 ;
        RECT 559.950 39.600 562.050 40.050 ;
        RECT 478.950 38.400 540.600 39.600 ;
        RECT 542.400 38.400 562.050 39.600 ;
        RECT 478.950 37.950 481.050 38.400 ;
        RECT 91.950 36.600 94.050 37.050 ;
        RECT 121.950 36.600 124.050 37.050 ;
        RECT 91.950 35.400 124.050 36.600 ;
        RECT 91.950 34.950 94.050 35.400 ;
        RECT 121.950 34.950 124.050 35.400 ;
        RECT 169.950 36.600 172.050 37.050 ;
        RECT 208.950 36.600 211.050 37.050 ;
        RECT 169.950 35.400 211.050 36.600 ;
        RECT 169.950 34.950 172.050 35.400 ;
        RECT 208.950 34.950 211.050 35.400 ;
        RECT 217.950 36.600 220.050 37.050 ;
        RECT 230.400 36.600 235.050 37.050 ;
        RECT 406.950 36.600 409.050 37.050 ;
        RECT 466.950 36.600 469.050 37.050 ;
        RECT 217.950 35.400 235.050 36.600 ;
        RECT 217.950 34.950 220.050 35.400 ;
        RECT 231.000 34.950 235.050 35.400 ;
        RECT 296.400 35.400 469.050 36.600 ;
        RECT 296.400 34.050 297.600 35.400 ;
        RECT 406.950 34.950 409.050 35.400 ;
        RECT 466.950 34.950 469.050 35.400 ;
        RECT 484.950 36.600 487.050 37.050 ;
        RECT 517.950 36.600 520.050 37.050 ;
        RECT 484.950 35.400 520.050 36.600 ;
        RECT 539.400 36.600 540.600 38.400 ;
        RECT 559.950 37.950 562.050 38.400 ;
        RECT 574.950 39.600 577.050 40.050 ;
        RECT 586.950 39.600 589.050 40.050 ;
        RECT 574.950 38.400 589.050 39.600 ;
        RECT 574.950 37.950 577.050 38.400 ;
        RECT 586.950 37.950 589.050 38.400 ;
        RECT 598.950 39.600 601.050 40.050 ;
        RECT 607.950 39.600 610.050 40.050 ;
        RECT 598.950 38.400 610.050 39.600 ;
        RECT 598.950 37.950 601.050 38.400 ;
        RECT 607.950 37.950 610.050 38.400 ;
        RECT 616.950 39.600 619.050 40.050 ;
        RECT 640.950 39.600 643.050 40.050 ;
        RECT 616.950 38.400 643.050 39.600 ;
        RECT 616.950 37.950 619.050 38.400 ;
        RECT 640.950 37.950 643.050 38.400 ;
        RECT 721.950 39.600 724.050 40.050 ;
        RECT 814.950 39.600 817.050 40.050 ;
        RECT 721.950 38.400 817.050 39.600 ;
        RECT 721.950 37.950 724.050 38.400 ;
        RECT 814.950 37.950 817.050 38.400 ;
        RECT 835.950 39.600 838.050 40.050 ;
        RECT 850.950 39.600 853.050 40.050 ;
        RECT 835.950 38.400 853.050 39.600 ;
        RECT 835.950 37.950 838.050 38.400 ;
        RECT 850.950 37.950 853.050 38.400 ;
        RECT 562.800 36.600 564.900 37.050 ;
        RECT 539.400 35.400 564.900 36.600 ;
        RECT 484.950 34.950 487.050 35.400 ;
        RECT 517.950 34.950 520.050 35.400 ;
        RECT 562.800 34.950 564.900 35.400 ;
        RECT 565.950 36.600 568.050 37.050 ;
        RECT 736.950 36.600 739.050 37.050 ;
        RECT 754.950 36.600 757.050 37.050 ;
        RECT 775.950 36.600 778.050 37.050 ;
        RECT 874.950 36.600 877.050 37.050 ;
        RECT 565.950 35.400 648.600 36.600 ;
        RECT 565.950 34.950 568.050 35.400 ;
        RECT 647.400 34.050 648.600 35.400 ;
        RECT 736.950 35.400 877.050 36.600 ;
        RECT 736.950 34.950 739.050 35.400 ;
        RECT 754.950 34.950 757.050 35.400 ;
        RECT 775.950 34.950 778.050 35.400 ;
        RECT 874.950 34.950 877.050 35.400 ;
        RECT 166.950 33.600 169.050 34.050 ;
        RECT 187.950 33.600 190.050 34.050 ;
        RECT 166.950 32.400 190.050 33.600 ;
        RECT 166.950 31.950 169.050 32.400 ;
        RECT 187.950 31.950 190.050 32.400 ;
        RECT 235.950 33.600 238.050 34.050 ;
        RECT 247.950 33.600 250.050 34.050 ;
        RECT 235.950 32.400 250.050 33.600 ;
        RECT 235.950 31.950 238.050 32.400 ;
        RECT 247.950 31.950 250.050 32.400 ;
        RECT 262.950 33.600 265.050 34.050 ;
        RECT 274.950 33.600 277.050 34.050 ;
        RECT 262.950 32.400 277.050 33.600 ;
        RECT 262.950 31.950 265.050 32.400 ;
        RECT 274.950 31.950 277.050 32.400 ;
        RECT 286.950 33.600 289.050 34.050 ;
        RECT 295.950 33.600 298.050 34.050 ;
        RECT 286.950 32.400 298.050 33.600 ;
        RECT 286.950 31.950 289.050 32.400 ;
        RECT 295.950 31.950 298.050 32.400 ;
        RECT 310.950 33.600 313.050 34.050 ;
        RECT 322.950 33.600 325.050 34.050 ;
        RECT 310.950 32.400 325.050 33.600 ;
        RECT 310.950 31.950 313.050 32.400 ;
        RECT 322.950 31.950 325.050 32.400 ;
        RECT 355.950 33.600 358.050 34.050 ;
        RECT 361.950 33.600 364.050 34.050 ;
        RECT 355.950 32.400 364.050 33.600 ;
        RECT 355.950 31.950 358.050 32.400 ;
        RECT 361.950 31.950 364.050 32.400 ;
        RECT 367.950 33.600 370.050 34.050 ;
        RECT 376.950 33.600 379.050 34.050 ;
        RECT 367.950 32.400 379.050 33.600 ;
        RECT 367.950 31.950 370.050 32.400 ;
        RECT 376.950 31.950 379.050 32.400 ;
        RECT 394.950 33.600 397.050 34.050 ;
        RECT 445.950 33.600 448.050 34.050 ;
        RECT 394.950 32.400 448.050 33.600 ;
        RECT 394.950 31.950 397.050 32.400 ;
        RECT 445.950 31.950 448.050 32.400 ;
        RECT 469.950 33.600 472.050 34.050 ;
        RECT 526.950 33.600 529.050 34.050 ;
        RECT 469.950 32.400 529.050 33.600 ;
        RECT 469.950 31.950 472.050 32.400 ;
        RECT 526.950 31.950 529.050 32.400 ;
        RECT 589.950 33.600 592.050 34.050 ;
        RECT 628.950 33.600 631.050 34.050 ;
        RECT 589.950 32.400 631.050 33.600 ;
        RECT 589.950 31.950 592.050 32.400 ;
        RECT 628.950 31.950 631.050 32.400 ;
        RECT 646.950 33.600 649.050 34.050 ;
        RECT 661.950 33.600 664.050 34.050 ;
        RECT 646.950 32.400 664.050 33.600 ;
        RECT 646.950 31.950 649.050 32.400 ;
        RECT 661.950 31.950 664.050 32.400 ;
        RECT 694.950 33.600 697.050 34.050 ;
        RECT 706.950 33.600 709.050 34.050 ;
        RECT 718.950 33.600 721.050 34.050 ;
        RECT 931.950 33.600 934.050 34.050 ;
        RECT 694.950 32.400 721.050 33.600 ;
        RECT 694.950 31.950 697.050 32.400 ;
        RECT 706.950 31.950 709.050 32.400 ;
        RECT 718.950 31.950 721.050 32.400 ;
        RECT 917.400 32.400 934.050 33.600 ;
        RECT 112.950 30.600 115.050 31.050 ;
        RECT 199.950 30.600 202.050 31.050 ;
        RECT 112.950 29.400 202.050 30.600 ;
        RECT 112.950 28.950 115.050 29.400 ;
        RECT 199.950 28.950 202.050 29.400 ;
        RECT 232.950 28.950 235.050 31.050 ;
        RECT 256.950 30.600 259.050 31.050 ;
        RECT 292.950 30.600 295.050 31.050 ;
        RECT 307.950 30.600 310.050 31.050 ;
        RECT 256.950 29.400 295.050 30.600 ;
        RECT 256.950 28.950 259.050 29.400 ;
        RECT 292.950 28.950 295.050 29.400 ;
        RECT 302.400 29.400 310.050 30.600 ;
        RECT 16.950 27.750 19.050 28.200 ;
        RECT 28.950 27.750 31.050 28.200 ;
        RECT 16.950 26.550 31.050 27.750 ;
        RECT 16.950 26.100 19.050 26.550 ;
        RECT 28.950 26.100 31.050 26.550 ;
        RECT 37.950 27.600 40.050 28.200 ;
        RECT 52.950 27.600 55.050 28.050 ;
        RECT 37.950 26.400 55.050 27.600 ;
        RECT 37.950 26.100 40.050 26.400 ;
        RECT 52.950 25.950 55.050 26.400 ;
        RECT 64.950 27.600 67.050 28.200 ;
        RECT 85.950 27.750 88.050 28.200 ;
        RECT 94.950 27.750 97.050 28.200 ;
        RECT 64.950 26.400 84.600 27.600 ;
        RECT 64.950 26.100 67.050 26.400 ;
        RECT 28.950 21.600 31.050 22.050 ;
        RECT 34.950 21.600 37.050 21.900 ;
        RECT 28.950 20.400 37.050 21.600 ;
        RECT 28.950 19.950 31.050 20.400 ;
        RECT 34.950 19.800 37.050 20.400 ;
        RECT 40.950 21.600 43.050 21.900 ;
        RECT 49.950 21.600 52.050 22.050 ;
        RECT 40.950 20.400 52.050 21.600 ;
        RECT 40.950 19.800 43.050 20.400 ;
        RECT 49.950 19.950 52.050 20.400 ;
        RECT 67.950 21.600 70.050 21.900 ;
        RECT 76.950 21.600 79.050 22.050 ;
        RECT 83.400 21.900 84.600 26.400 ;
        RECT 85.950 26.550 97.050 27.750 ;
        RECT 85.950 26.100 88.050 26.550 ;
        RECT 94.950 26.100 97.050 26.550 ;
        RECT 106.950 26.100 109.050 28.200 ;
        RECT 127.950 27.600 130.050 28.200 ;
        RECT 148.950 27.600 151.050 28.200 ;
        RECT 166.950 27.600 169.050 28.200 ;
        RECT 125.400 26.400 130.050 27.600 ;
        RECT 97.950 24.600 100.050 25.050 ;
        RECT 89.400 23.400 100.050 24.600 ;
        RECT 89.400 21.900 90.600 23.400 ;
        RECT 97.950 22.950 100.050 23.400 ;
        RECT 67.950 20.400 79.050 21.600 ;
        RECT 67.950 19.800 70.050 20.400 ;
        RECT 76.950 19.950 79.050 20.400 ;
        RECT 82.950 19.800 85.050 21.900 ;
        RECT 88.950 19.800 91.050 21.900 ;
        RECT 100.950 21.600 103.050 22.050 ;
        RECT 107.400 21.600 108.600 26.100 ;
        RECT 118.950 24.600 121.050 25.050 ;
        RECT 110.400 23.400 121.050 24.600 ;
        RECT 110.400 21.900 111.600 23.400 ;
        RECT 118.950 22.950 121.050 23.400 ;
        RECT 125.400 22.050 126.600 26.400 ;
        RECT 127.950 26.100 130.050 26.400 ;
        RECT 131.400 26.400 169.050 27.600 ;
        RECT 100.950 20.400 108.600 21.600 ;
        RECT 100.950 19.950 103.050 20.400 ;
        RECT 109.950 19.800 112.050 21.900 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 131.400 21.900 132.600 26.400 ;
        RECT 148.950 26.100 151.050 26.400 ;
        RECT 166.950 26.100 169.050 26.400 ;
        RECT 181.950 27.750 184.050 28.200 ;
        RECT 190.950 27.750 193.050 28.200 ;
        RECT 181.950 26.550 193.050 27.750 ;
        RECT 181.950 26.100 184.050 26.550 ;
        RECT 190.950 26.100 193.050 26.550 ;
        RECT 202.950 27.750 205.050 28.200 ;
        RECT 211.950 27.750 214.050 28.200 ;
        RECT 202.950 26.550 214.050 27.750 ;
        RECT 202.950 26.100 205.050 26.550 ;
        RECT 211.950 26.100 214.050 26.550 ;
        RECT 217.950 27.600 220.050 28.200 ;
        RECT 226.950 27.600 229.050 28.050 ;
        RECT 217.950 26.400 229.050 27.600 ;
        RECT 217.950 26.100 220.050 26.400 ;
        RECT 226.950 25.950 229.050 26.400 ;
        RECT 130.950 19.800 133.050 21.900 ;
        RECT 151.950 21.600 154.050 21.900 ;
        RECT 163.950 21.600 166.050 21.900 ;
        RECT 151.950 20.400 166.050 21.600 ;
        RECT 151.950 19.800 154.050 20.400 ;
        RECT 163.950 19.800 166.050 20.400 ;
        RECT 169.950 21.600 172.050 21.900 ;
        RECT 178.950 21.600 181.050 22.050 ;
        RECT 233.400 21.900 234.600 28.950 ;
        RECT 241.950 27.600 244.050 28.200 ;
        RECT 259.950 27.600 262.050 28.050 ;
        RECT 241.950 26.400 262.050 27.600 ;
        RECT 241.950 26.100 244.050 26.400 ;
        RECT 259.950 25.950 262.050 26.400 ;
        RECT 268.950 27.600 273.000 28.050 ;
        RECT 289.950 27.600 292.050 28.050 ;
        RECT 302.400 27.600 303.600 29.400 ;
        RECT 307.950 28.950 310.050 29.400 ;
        RECT 385.950 30.600 388.050 31.050 ;
        RECT 466.950 30.600 469.050 31.050 ;
        RECT 385.950 29.400 469.050 30.600 ;
        RECT 385.950 28.950 388.050 29.400 ;
        RECT 466.950 28.950 469.050 29.400 ;
        RECT 532.950 30.600 535.050 31.050 ;
        RECT 553.950 30.600 556.050 31.050 ;
        RECT 637.950 30.600 640.050 31.050 ;
        RECT 532.950 29.400 640.050 30.600 ;
        RECT 532.950 28.950 535.050 29.400 ;
        RECT 553.950 28.950 556.050 29.400 ;
        RECT 637.950 28.950 640.050 29.400 ;
        RECT 319.950 27.600 322.050 28.200 ;
        RECT 268.950 25.950 273.600 27.600 ;
        RECT 289.950 26.400 303.600 27.600 ;
        RECT 305.400 26.400 322.050 27.600 ;
        RECT 289.950 25.950 292.050 26.400 ;
        RECT 169.950 20.400 181.050 21.600 ;
        RECT 169.950 19.800 172.050 20.400 ;
        RECT 178.950 19.950 181.050 20.400 ;
        RECT 193.950 21.600 196.050 21.900 ;
        RECT 208.950 21.600 211.050 21.900 ;
        RECT 193.950 20.400 211.050 21.600 ;
        RECT 193.950 19.800 196.050 20.400 ;
        RECT 208.950 19.800 211.050 20.400 ;
        RECT 232.950 19.800 235.050 21.900 ;
        RECT 247.950 21.600 250.050 22.050 ;
        RECT 253.950 21.600 256.050 21.900 ;
        RECT 265.950 21.600 268.050 22.050 ;
        RECT 272.400 21.900 273.600 25.950 ;
        RECT 286.950 24.600 289.050 25.050 ;
        RECT 278.400 23.400 289.050 24.600 ;
        RECT 278.400 21.900 279.600 23.400 ;
        RECT 286.950 22.950 289.050 23.400 ;
        RECT 305.400 21.900 306.600 26.400 ;
        RECT 319.950 26.100 322.050 26.400 ;
        RECT 325.950 27.600 328.050 28.200 ;
        RECT 358.950 27.600 361.050 28.050 ;
        RECT 372.000 27.600 376.050 28.050 ;
        RECT 325.950 26.400 342.600 27.600 ;
        RECT 325.950 26.100 328.050 26.400 ;
        RECT 341.400 21.900 342.600 26.400 ;
        RECT 358.950 26.400 366.600 27.600 ;
        RECT 358.950 25.950 361.050 26.400 ;
        RECT 365.400 21.900 366.600 26.400 ;
        RECT 371.400 25.950 376.050 27.600 ;
        RECT 391.950 27.750 394.050 28.200 ;
        RECT 400.800 27.750 402.900 28.200 ;
        RECT 391.950 26.550 402.900 27.750 ;
        RECT 391.950 26.100 394.050 26.550 ;
        RECT 400.800 26.100 402.900 26.550 ;
        RECT 403.950 27.750 406.050 28.200 ;
        RECT 412.950 27.750 415.050 28.200 ;
        RECT 403.950 26.550 415.050 27.750 ;
        RECT 403.950 26.100 406.050 26.550 ;
        RECT 412.950 26.100 415.050 26.550 ;
        RECT 439.950 27.750 442.050 28.200 ;
        RECT 448.950 27.750 451.050 28.200 ;
        RECT 439.950 26.550 451.050 27.750 ;
        RECT 439.950 26.100 442.050 26.550 ;
        RECT 448.950 26.100 451.050 26.550 ;
        RECT 457.950 27.750 460.050 28.200 ;
        RECT 469.800 27.750 471.900 28.200 ;
        RECT 457.950 26.550 471.900 27.750 ;
        RECT 457.950 26.100 460.050 26.550 ;
        RECT 469.800 26.100 471.900 26.550 ;
        RECT 472.950 27.750 475.050 28.200 ;
        RECT 505.950 27.750 508.050 28.200 ;
        RECT 472.950 26.550 508.050 27.750 ;
        RECT 472.950 26.100 475.050 26.550 ;
        RECT 505.950 26.100 508.050 26.550 ;
        RECT 511.950 27.600 514.050 28.200 ;
        RECT 520.950 27.600 523.050 28.050 ;
        RECT 526.950 27.600 529.050 28.200 ;
        RECT 511.950 26.400 519.600 27.600 ;
        RECT 511.950 26.100 514.050 26.400 ;
        RECT 371.400 21.900 372.600 25.950 ;
        RECT 518.400 24.600 519.600 26.400 ;
        RECT 520.950 26.400 529.050 27.600 ;
        RECT 520.950 25.950 523.050 26.400 ;
        RECT 526.950 26.100 529.050 26.400 ;
        RECT 541.950 27.600 544.050 28.050 ;
        RECT 547.950 27.600 550.050 28.200 ;
        RECT 541.950 26.400 550.050 27.600 ;
        RECT 541.950 25.950 544.050 26.400 ;
        RECT 547.950 26.100 550.050 26.400 ;
        RECT 562.950 27.750 565.050 28.200 ;
        RECT 580.950 27.750 583.050 28.200 ;
        RECT 562.950 27.600 583.050 27.750 ;
        RECT 604.950 27.600 607.050 28.200 ;
        RECT 622.950 27.600 625.050 28.200 ;
        RECT 634.950 27.600 637.050 28.050 ;
        RECT 562.950 26.550 621.600 27.600 ;
        RECT 562.950 26.100 565.050 26.550 ;
        RECT 580.950 26.400 621.600 26.550 ;
        RECT 580.950 26.100 583.050 26.400 ;
        RECT 604.950 26.100 607.050 26.400 ;
        RECT 620.400 24.600 621.600 26.400 ;
        RECT 622.950 26.400 637.050 27.600 ;
        RECT 622.950 26.100 625.050 26.400 ;
        RECT 634.950 25.950 637.050 26.400 ;
        RECT 640.950 27.600 643.050 28.050 ;
        RECT 652.950 27.600 655.050 31.050 ;
        RECT 670.950 30.600 673.050 31.050 ;
        RECT 676.950 30.600 679.050 31.050 ;
        RECT 781.950 30.600 784.050 31.050 ;
        RECT 670.950 29.400 679.050 30.600 ;
        RECT 670.950 28.950 673.050 29.400 ;
        RECT 676.950 28.950 679.050 29.400 ;
        RECT 776.400 29.400 784.050 30.600 ;
        RECT 667.950 27.600 670.050 28.200 ;
        RECT 640.950 26.400 651.600 27.600 ;
        RECT 652.950 27.000 670.050 27.600 ;
        RECT 653.400 26.400 670.050 27.000 ;
        RECT 640.950 25.950 643.050 26.400 ;
        RECT 518.400 23.400 531.600 24.600 ;
        RECT 247.950 20.400 268.050 21.600 ;
        RECT 247.950 19.950 250.050 20.400 ;
        RECT 253.950 19.800 256.050 20.400 ;
        RECT 265.950 19.950 268.050 20.400 ;
        RECT 271.950 19.800 274.050 21.900 ;
        RECT 277.950 19.800 280.050 21.900 ;
        RECT 304.950 19.800 307.050 21.900 ;
        RECT 316.950 21.450 319.050 21.900 ;
        RECT 331.950 21.450 334.050 21.900 ;
        RECT 316.950 20.250 334.050 21.450 ;
        RECT 316.950 19.800 319.050 20.250 ;
        RECT 331.950 19.800 334.050 20.250 ;
        RECT 340.950 19.800 343.050 21.900 ;
        RECT 364.950 19.800 367.050 21.900 ;
        RECT 370.950 19.800 373.050 21.900 ;
        RECT 400.950 21.600 403.050 22.050 ;
        RECT 530.400 21.900 531.600 23.400 ;
        RECT 536.400 23.400 567.600 24.600 ;
        RECT 620.400 23.400 627.600 24.600 ;
        RECT 536.400 21.900 537.600 23.400 ;
        RECT 566.400 21.900 567.600 23.400 ;
        RECT 626.400 21.900 627.600 23.400 ;
        RECT 650.400 21.900 651.600 26.400 ;
        RECT 667.950 26.100 670.050 26.400 ;
        RECT 712.950 27.600 715.050 28.200 ;
        RECT 724.950 27.600 727.050 28.050 ;
        RECT 712.950 26.400 727.050 27.600 ;
        RECT 712.950 26.100 715.050 26.400 ;
        RECT 724.950 25.950 727.050 26.400 ;
        RECT 730.950 27.600 733.050 28.200 ;
        RECT 766.950 27.600 769.050 28.050 ;
        RECT 730.950 26.400 769.050 27.600 ;
        RECT 730.950 26.100 733.050 26.400 ;
        RECT 766.950 25.950 769.050 26.400 ;
        RECT 776.400 24.600 777.600 29.400 ;
        RECT 781.950 28.950 784.050 29.400 ;
        RECT 892.950 30.600 895.050 31.050 ;
        RECT 917.400 30.600 918.600 32.400 ;
        RECT 931.950 31.950 934.050 32.400 ;
        RECT 892.950 29.400 918.600 30.600 ;
        RECT 892.950 28.950 895.050 29.400 ;
        RECT 790.950 27.750 793.050 28.200 ;
        RECT 799.950 27.750 802.050 28.200 ;
        RECT 790.950 27.600 802.050 27.750 ;
        RECT 823.950 27.600 826.050 28.200 ;
        RECT 790.950 26.550 826.050 27.600 ;
        RECT 790.950 26.100 793.050 26.550 ;
        RECT 799.950 26.400 826.050 26.550 ;
        RECT 799.950 26.100 802.050 26.400 ;
        RECT 823.950 26.100 826.050 26.400 ;
        RECT 925.950 27.750 928.050 28.200 ;
        RECT 934.950 27.750 937.050 28.200 ;
        RECT 925.950 26.550 937.050 27.750 ;
        RECT 925.950 26.100 928.050 26.550 ;
        RECT 934.950 26.100 937.050 26.550 ;
        RECT 752.400 23.400 777.600 24.600 ;
        RECT 752.400 21.900 753.600 23.400 ;
        RECT 409.950 21.600 412.050 21.900 ;
        RECT 400.950 21.450 412.050 21.600 ;
        RECT 430.950 21.450 433.050 21.900 ;
        RECT 400.950 20.400 433.050 21.450 ;
        RECT 400.950 19.950 403.050 20.400 ;
        RECT 409.950 20.250 433.050 20.400 ;
        RECT 409.950 19.800 412.050 20.250 ;
        RECT 430.950 19.800 433.050 20.250 ;
        RECT 442.950 21.450 445.050 21.900 ;
        RECT 469.950 21.450 472.050 21.900 ;
        RECT 481.950 21.600 484.050 21.900 ;
        RECT 442.950 20.250 472.050 21.450 ;
        RECT 442.950 19.800 445.050 20.250 ;
        RECT 469.950 19.800 472.050 20.250 ;
        RECT 479.400 20.400 484.050 21.600 ;
        RECT 13.950 18.600 16.050 19.050 ;
        RECT 25.950 18.600 28.050 19.050 ;
        RECT 13.950 17.400 28.050 18.600 ;
        RECT 13.950 16.950 16.050 17.400 ;
        RECT 25.950 16.950 28.050 17.400 ;
        RECT 184.950 18.600 187.050 19.050 ;
        RECT 220.950 18.600 223.050 19.050 ;
        RECT 184.950 17.400 223.050 18.600 ;
        RECT 184.950 16.950 187.050 17.400 ;
        RECT 220.950 16.950 223.050 17.400 ;
        RECT 376.950 18.600 379.050 19.050 ;
        RECT 472.950 18.600 475.050 19.050 ;
        RECT 479.400 18.600 480.600 20.400 ;
        RECT 481.950 19.800 484.050 20.400 ;
        RECT 487.950 21.450 490.050 21.900 ;
        RECT 496.950 21.450 499.050 21.900 ;
        RECT 487.950 20.250 499.050 21.450 ;
        RECT 487.950 19.800 490.050 20.250 ;
        RECT 496.950 19.800 499.050 20.250 ;
        RECT 529.950 19.800 532.050 21.900 ;
        RECT 535.950 19.800 538.050 21.900 ;
        RECT 565.950 21.450 568.050 21.900 ;
        RECT 571.950 21.450 574.050 21.900 ;
        RECT 565.950 20.250 574.050 21.450 ;
        RECT 565.950 19.800 568.050 20.250 ;
        RECT 571.950 19.800 574.050 20.250 ;
        RECT 577.950 21.600 580.050 21.900 ;
        RECT 601.950 21.600 604.050 21.900 ;
        RECT 577.950 21.450 604.050 21.600 ;
        RECT 610.950 21.450 613.050 21.900 ;
        RECT 577.950 20.400 613.050 21.450 ;
        RECT 577.950 19.800 580.050 20.400 ;
        RECT 601.950 20.250 613.050 20.400 ;
        RECT 601.950 19.800 604.050 20.250 ;
        RECT 610.950 19.800 613.050 20.250 ;
        RECT 625.950 19.800 628.050 21.900 ;
        RECT 637.950 21.450 640.050 21.900 ;
        RECT 643.950 21.450 646.050 21.900 ;
        RECT 637.950 20.250 646.050 21.450 ;
        RECT 637.950 19.800 640.050 20.250 ;
        RECT 643.950 19.800 646.050 20.250 ;
        RECT 649.950 19.800 652.050 21.900 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 679.950 21.450 682.050 21.900 ;
        RECT 670.950 20.250 682.050 21.450 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 679.950 19.800 682.050 20.250 ;
        RECT 685.950 21.600 688.050 21.900 ;
        RECT 733.950 21.600 736.050 21.900 ;
        RECT 685.950 20.400 736.050 21.600 ;
        RECT 685.950 19.800 688.050 20.400 ;
        RECT 733.950 19.800 736.050 20.400 ;
        RECT 739.950 21.600 742.050 21.900 ;
        RECT 751.950 21.600 754.050 21.900 ;
        RECT 739.950 20.400 754.050 21.600 ;
        RECT 739.950 19.800 742.050 20.400 ;
        RECT 751.950 19.800 754.050 20.400 ;
        RECT 772.950 21.600 775.050 21.900 ;
        RECT 776.400 21.600 777.600 23.400 ;
        RECT 838.950 24.600 841.050 25.050 ;
        RECT 838.950 23.400 867.600 24.600 ;
        RECT 838.950 22.950 841.050 23.400 ;
        RECT 772.950 20.400 777.600 21.600 ;
        RECT 796.950 21.600 799.050 21.900 ;
        RECT 817.950 21.600 820.050 22.050 ;
        RECT 866.400 21.900 867.600 23.400 ;
        RECT 796.950 20.400 820.050 21.600 ;
        RECT 772.950 19.800 775.050 20.400 ;
        RECT 796.950 19.800 799.050 20.400 ;
        RECT 817.950 19.950 820.050 20.400 ;
        RECT 865.950 19.800 868.050 21.900 ;
        RECT 904.950 21.450 907.050 21.900 ;
        RECT 910.950 21.450 913.050 21.900 ;
        RECT 904.950 20.250 913.050 21.450 ;
        RECT 904.950 19.800 907.050 20.250 ;
        RECT 910.950 19.800 913.050 20.250 ;
        RECT 916.950 21.600 919.050 21.900 ;
        RECT 931.950 21.600 934.050 21.900 ;
        RECT 916.950 20.400 934.050 21.600 ;
        RECT 916.950 19.800 919.050 20.400 ;
        RECT 931.950 19.800 934.050 20.400 ;
        RECT 376.950 17.400 480.600 18.600 ;
        RECT 502.950 18.600 505.050 19.050 ;
        RECT 517.950 18.600 520.050 19.050 ;
        RECT 502.950 17.400 520.050 18.600 ;
        RECT 376.950 16.950 379.050 17.400 ;
        RECT 472.950 16.950 475.050 17.400 ;
        RECT 502.950 16.950 505.050 17.400 ;
        RECT 517.950 16.950 520.050 17.400 ;
        RECT 529.950 18.600 532.050 19.050 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 619.950 18.600 622.050 19.050 ;
        RECT 715.950 18.600 718.050 19.050 ;
        RECT 757.950 18.600 760.050 19.050 ;
        RECT 778.950 18.600 781.050 19.050 ;
        RECT 529.950 17.400 622.050 18.600 ;
        RECT 529.950 16.950 532.050 17.400 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 619.950 16.950 622.050 17.400 ;
        RECT 662.400 17.400 781.050 18.600 ;
        RECT 34.950 15.600 37.050 16.050 ;
        RECT 100.950 15.600 103.050 16.050 ;
        RECT 34.950 14.400 103.050 15.600 ;
        RECT 34.950 13.950 37.050 14.400 ;
        RECT 100.950 13.950 103.050 14.400 ;
        RECT 121.950 15.600 124.050 16.050 ;
        RECT 181.950 15.600 184.050 16.050 ;
        RECT 214.950 15.600 217.050 16.050 ;
        RECT 121.950 14.400 217.050 15.600 ;
        RECT 121.950 13.950 124.050 14.400 ;
        RECT 181.950 13.950 184.050 14.400 ;
        RECT 214.950 13.950 217.050 14.400 ;
        RECT 238.950 15.600 241.050 16.050 ;
        RECT 310.950 15.600 313.050 16.050 ;
        RECT 238.950 14.400 313.050 15.600 ;
        RECT 238.950 13.950 241.050 14.400 ;
        RECT 310.950 13.950 313.050 14.400 ;
        RECT 316.950 15.600 319.050 16.050 ;
        RECT 334.950 15.600 337.050 16.050 ;
        RECT 316.950 14.400 337.050 15.600 ;
        RECT 316.950 13.950 319.050 14.400 ;
        RECT 334.950 13.950 337.050 14.400 ;
        RECT 340.950 15.600 343.050 16.050 ;
        RECT 427.950 15.600 430.050 16.050 ;
        RECT 340.950 14.400 430.050 15.600 ;
        RECT 340.950 13.950 343.050 14.400 ;
        RECT 427.950 13.950 430.050 14.400 ;
        RECT 436.950 15.600 439.050 15.900 ;
        RECT 457.950 15.600 460.050 16.050 ;
        RECT 436.950 14.400 460.050 15.600 ;
        RECT 436.950 13.800 439.050 14.400 ;
        RECT 457.950 13.950 460.050 14.400 ;
        RECT 469.950 15.600 472.050 16.050 ;
        RECT 490.950 15.600 493.050 16.050 ;
        RECT 469.950 14.400 493.050 15.600 ;
        RECT 469.950 13.950 472.050 14.400 ;
        RECT 490.950 13.950 493.050 14.400 ;
        RECT 505.950 15.600 508.050 15.900 ;
        RECT 520.950 15.600 523.050 16.050 ;
        RECT 505.950 14.400 523.050 15.600 ;
        RECT 505.950 13.800 508.050 14.400 ;
        RECT 520.950 13.950 523.050 14.400 ;
        RECT 556.950 15.600 559.050 16.050 ;
        RECT 589.950 15.600 592.050 16.050 ;
        RECT 556.950 14.400 592.050 15.600 ;
        RECT 556.950 13.950 559.050 14.400 ;
        RECT 589.950 13.950 592.050 14.400 ;
        RECT 634.950 15.600 637.050 16.050 ;
        RECT 662.400 15.600 663.600 17.400 ;
        RECT 715.950 16.950 718.050 17.400 ;
        RECT 757.950 16.950 760.050 17.400 ;
        RECT 778.950 16.950 781.050 17.400 ;
        RECT 802.950 18.600 805.050 19.050 ;
        RECT 820.950 18.600 823.050 19.050 ;
        RECT 844.950 18.600 847.050 19.050 ;
        RECT 856.950 18.600 859.050 19.050 ;
        RECT 802.950 17.400 859.050 18.600 ;
        RECT 802.950 16.950 805.050 17.400 ;
        RECT 820.950 16.950 823.050 17.400 ;
        RECT 844.950 16.950 847.050 17.400 ;
        RECT 856.950 16.950 859.050 17.400 ;
        RECT 634.950 14.400 663.600 15.600 ;
        RECT 664.950 15.600 667.050 16.050 ;
        RECT 685.950 15.600 688.050 16.050 ;
        RECT 664.950 14.400 688.050 15.600 ;
        RECT 634.950 13.950 637.050 14.400 ;
        RECT 664.950 13.950 667.050 14.400 ;
        RECT 685.950 13.950 688.050 14.400 ;
        RECT 691.950 15.600 694.050 16.050 ;
        RECT 709.950 15.600 712.050 16.050 ;
        RECT 721.950 15.600 724.050 16.050 ;
        RECT 691.950 14.400 724.050 15.600 ;
        RECT 691.950 13.950 694.050 14.400 ;
        RECT 709.950 13.950 712.050 14.400 ;
        RECT 721.950 13.950 724.050 14.400 ;
        RECT 826.950 15.600 829.050 15.900 ;
        RECT 838.950 15.600 841.050 16.050 ;
        RECT 826.950 14.400 841.050 15.600 ;
        RECT 826.950 13.800 829.050 14.400 ;
        RECT 838.950 13.950 841.050 14.400 ;
        RECT 895.950 15.600 898.050 16.050 ;
        RECT 943.950 15.600 946.050 16.050 ;
        RECT 895.950 14.400 946.050 15.600 ;
        RECT 895.950 13.950 898.050 14.400 ;
        RECT 943.950 13.950 946.050 14.400 ;
        RECT 52.950 12.600 55.050 13.050 ;
        RECT 136.950 12.600 139.050 13.050 ;
        RECT 52.950 11.400 139.050 12.600 ;
        RECT 52.950 10.950 55.050 11.400 ;
        RECT 136.950 10.950 139.050 11.400 ;
        RECT 220.950 12.600 223.050 13.050 ;
        RECT 235.950 12.600 238.050 13.050 ;
        RECT 220.950 11.400 238.050 12.600 ;
        RECT 220.950 10.950 223.050 11.400 ;
        RECT 235.950 10.950 238.050 11.400 ;
        RECT 241.950 12.600 244.050 13.050 ;
        RECT 298.950 12.600 301.050 13.050 ;
        RECT 241.950 11.400 301.050 12.600 ;
        RECT 241.950 10.950 244.050 11.400 ;
        RECT 298.950 10.950 301.050 11.400 ;
        RECT 352.950 12.600 355.050 13.050 ;
        RECT 433.950 12.600 436.050 13.050 ;
        RECT 352.950 11.400 436.050 12.600 ;
        RECT 352.950 10.950 355.050 11.400 ;
        RECT 433.950 10.950 436.050 11.400 ;
        RECT 667.950 12.600 670.050 13.050 ;
        RECT 676.950 12.600 679.050 13.050 ;
        RECT 667.950 11.400 679.050 12.600 ;
        RECT 667.950 10.950 670.050 11.400 ;
        RECT 676.950 10.950 679.050 11.400 ;
        RECT 766.950 12.600 769.050 13.050 ;
        RECT 796.950 12.600 799.050 13.050 ;
        RECT 766.950 11.400 799.050 12.600 ;
        RECT 766.950 10.950 769.050 11.400 ;
        RECT 796.950 10.950 799.050 11.400 ;
        RECT 103.950 9.600 106.050 10.050 ;
        RECT 124.950 9.600 127.050 10.050 ;
        RECT 103.950 8.400 127.050 9.600 ;
        RECT 103.950 7.950 106.050 8.400 ;
        RECT 124.950 7.950 127.050 8.400 ;
        RECT 187.950 9.600 190.050 10.050 ;
        RECT 205.950 9.600 208.050 10.050 ;
        RECT 217.950 9.600 220.050 10.050 ;
        RECT 187.950 8.400 220.050 9.600 ;
        RECT 187.950 7.950 190.050 8.400 ;
        RECT 205.950 7.950 208.050 8.400 ;
        RECT 217.950 7.950 220.050 8.400 ;
        RECT 223.950 9.600 226.050 10.050 ;
        RECT 232.950 9.600 235.050 10.050 ;
        RECT 223.950 8.400 235.050 9.600 ;
        RECT 223.950 7.950 226.050 8.400 ;
        RECT 232.950 7.950 235.050 8.400 ;
        RECT 244.950 9.600 247.050 10.050 ;
        RECT 295.950 9.600 298.050 10.050 ;
        RECT 244.950 8.400 298.050 9.600 ;
        RECT 244.950 7.950 247.050 8.400 ;
        RECT 295.950 7.950 298.050 8.400 ;
        RECT 301.950 9.600 304.050 10.050 ;
        RECT 328.950 9.600 331.050 10.050 ;
        RECT 301.950 8.400 331.050 9.600 ;
        RECT 301.950 7.950 304.050 8.400 ;
        RECT 328.950 7.950 331.050 8.400 ;
        RECT 334.950 9.600 337.050 10.050 ;
        RECT 346.950 9.600 349.050 10.050 ;
        RECT 334.950 8.400 349.050 9.600 ;
        RECT 334.950 7.950 337.050 8.400 ;
        RECT 346.950 7.950 349.050 8.400 ;
        RECT 358.950 9.600 361.050 10.050 ;
        RECT 388.950 9.600 391.050 10.050 ;
        RECT 415.950 9.600 418.050 10.050 ;
        RECT 358.950 8.400 418.050 9.600 ;
        RECT 358.950 7.950 361.050 8.400 ;
        RECT 388.950 7.950 391.050 8.400 ;
        RECT 415.950 7.950 418.050 8.400 ;
        RECT 448.950 9.600 451.050 10.050 ;
        RECT 454.950 9.600 457.050 10.050 ;
        RECT 613.950 9.600 616.050 10.050 ;
        RECT 448.950 8.400 616.050 9.600 ;
        RECT 448.950 7.950 451.050 8.400 ;
        RECT 454.950 7.950 457.050 8.400 ;
        RECT 613.950 7.950 616.050 8.400 ;
        RECT 811.950 9.600 814.050 10.050 ;
        RECT 871.950 9.600 874.050 10.050 ;
        RECT 925.950 9.600 928.050 10.050 ;
        RECT 811.950 8.400 928.050 9.600 ;
        RECT 811.950 7.950 814.050 8.400 ;
        RECT 871.950 7.950 874.050 8.400 ;
        RECT 925.950 7.950 928.050 8.400 ;
        RECT 163.950 6.600 166.050 7.050 ;
        RECT 202.950 6.600 205.050 7.050 ;
        RECT 163.950 5.400 205.050 6.600 ;
        RECT 163.950 4.950 166.050 5.400 ;
        RECT 202.950 4.950 205.050 5.400 ;
        RECT 208.950 6.600 211.050 7.050 ;
        RECT 262.950 6.600 265.050 7.050 ;
        RECT 208.950 5.400 265.050 6.600 ;
        RECT 208.950 4.950 211.050 5.400 ;
        RECT 262.950 4.950 265.050 5.400 ;
        RECT 394.950 6.600 397.050 7.050 ;
        RECT 403.950 6.600 406.050 7.050 ;
        RECT 433.950 6.600 436.050 7.050 ;
        RECT 394.950 5.400 436.050 6.600 ;
        RECT 394.950 4.950 397.050 5.400 ;
        RECT 403.950 4.950 406.050 5.400 ;
        RECT 433.950 4.950 436.050 5.400 ;
        RECT 457.950 6.600 460.050 7.050 ;
        RECT 505.950 6.600 508.050 7.050 ;
        RECT 457.950 5.400 508.050 6.600 ;
        RECT 457.950 4.950 460.050 5.400 ;
        RECT 505.950 4.950 508.050 5.400 ;
        RECT 511.950 6.600 514.050 7.050 ;
        RECT 586.950 6.600 589.050 7.050 ;
        RECT 511.950 5.400 589.050 6.600 ;
        RECT 511.950 4.950 514.050 5.400 ;
        RECT 586.950 4.950 589.050 5.400 ;
        RECT 724.950 6.600 727.050 7.050 ;
        RECT 790.950 6.600 793.050 7.050 ;
        RECT 724.950 5.400 793.050 6.600 ;
        RECT 724.950 4.950 727.050 5.400 ;
        RECT 790.950 4.950 793.050 5.400 ;
        RECT 889.950 6.600 892.050 7.050 ;
        RECT 940.950 6.600 943.050 7.050 ;
        RECT 889.950 5.400 943.050 6.600 ;
        RECT 889.950 4.950 892.050 5.400 ;
        RECT 940.950 4.950 943.050 5.400 ;
        RECT 436.950 3.600 439.050 4.050 ;
        RECT 508.950 3.600 511.050 4.050 ;
        RECT 436.950 2.400 511.050 3.600 ;
        RECT 436.950 1.950 439.050 2.400 ;
        RECT 508.950 1.950 511.050 2.400 ;
        RECT 514.950 3.600 517.050 4.050 ;
        RECT 541.950 3.600 544.050 4.050 ;
        RECT 514.950 2.400 544.050 3.600 ;
        RECT 514.950 1.950 517.050 2.400 ;
        RECT 541.950 1.950 544.050 2.400 ;
  END
END ALU_wrapper
END LIBRARY

