magic
tech scmos
magscale 1 60
timestamp 1709416183
<< checkpaint >>
rect -1200 -1200 381200 381200
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 -1 342200 -1 0 175360
box -70 0 2070 50120
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1709081121
transform 1 0 120690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_1
timestamp 1709081121
transform 0 1 37800 -1 0 151309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_2
timestamp 1709081121
transform 1 0 174690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_3
timestamp 1709081121
transform 1 0 147690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_4
timestamp 1709081121
transform 1 0 228690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_5
timestamp 1709081121
transform 1 0 201690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_6
timestamp 1709081121
transform 0 1 37800 -1 0 124309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_8
timestamp 1709081121
transform 0 1 37800 -1 0 205309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_9
timestamp 1709081121
transform 0 1 37800 -1 0 178309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_10
timestamp 1709081121
transform 0 1 37800 -1 0 259309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_11
timestamp 1709081121
transform 0 1 37800 -1 0 232309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_14
timestamp 1709081121
transform 0 -1 342200 -1 0 205305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_15
timestamp 1709081121
transform 0 -1 342200 -1 0 178305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_16
timestamp 1709081121
transform 0 -1 342200 -1 0 259305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_17
timestamp 1709081121
transform 0 -1 342200 -1 0 232305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_18
timestamp 1709081121
transform 1 0 147690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_19
timestamp 1709081121
transform 1 0 120690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_20
timestamp 1709081121
transform 1 0 201690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_21
timestamp 1709081121
transform 1 0 174690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_22
timestamp 1709081121
transform 1 0 255690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_23
timestamp 1709081121
transform 1 0 228690 0 -1 342200
box 0 0 3620 50120
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 1 0 87287 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_1
timestamp 1692859860
transform 0 1 37800 -1 0 97233
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_2
timestamp 1692859860
transform 1 0 255648 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_3
timestamp 1692859860
transform 0 1 37800 -1 0 292759
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_4
timestamp 1692859860
transform 1 0 87417 0 -1 342200
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_5
timestamp 1692859860
transform 1 0 282662 0 -1 342199
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_6
timestamp 1692859860
transform 0 -1 342200 -1 0 97270
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_7
timestamp 1692859860
transform 0 -1 342200 -1 0 292717
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_8
timestamp 1692859860
transform 0 -1 342200 -1 0 164305
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_9
timestamp 1692859860
transform 0 -1 342200 -1 0 106780
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_10
timestamp 1692859860
transform 0 -1 342200 -1 0 116305
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_11
timestamp 1692859860
transform 0 -1 342200 -1 0 125905
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_12
timestamp 1692859860
transform 0 -1 342200 -1 0 135505
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_13
timestamp 1692859860
transform 0 -1 342200 -1 0 145105
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_14
timestamp 1692859860
transform 0 -1 342200 -1 0 154705
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_15
timestamp 1692859860
transform 0 -1 342200 -1 0 173905
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_16
timestamp 1692859860
transform 1 0 282762 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_17
timestamp 1692859860
transform 1 0 273362 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_18
timestamp 1692859860
transform 1 0 263968 0 1 37800
box -70 0 10070 50120
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 1 0 37800 0 1 37800
box 0 0 50600 50600
use PCORNER  PCORNER_1
timestamp 1692859860
transform -1 0 342200 0 1 37800
box 0 0 50600 50600
use PCORNER  PCORNER_2
timestamp 1692859860
transform 0 1 37800 -1 0 342200
box 0 0 50600 50600
use PCORNER  PCORNER_3
timestamp 1692859860
transform 0 -1 342200 -1 0 342200
box 0 0 50600 50600
use PAD80  PAD80_2 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1709379016
transform 1 0 262500 0 1 19500
box 0 0 17000 17000
use PAD80  PAD80_6
timestamp 1709379016
transform 1 0 343500 0 1 127500
box 0 0 17000 17000
use PAD80  PAD80_7
timestamp 1709379016
transform 1 0 343500 0 1 100500
box 0 0 17000 17000
use PAD80  PAD80_17
timestamp 1709379016
transform 1 0 343500 0 1 154500
box 0 0 17000 17000
use PIC  ABCMD_I_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1699925102
transform 1 0 259000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_1
timestamp 1699925102
transform 0 -1 342200 -1 0 229000
box -200 -18300 24200 50600
use PIC  ABCMD_I_2
timestamp 1699925102
transform 0 -1 342200 -1 0 256000
box -200 -18300 24200 50600
use PIC  ABCMD_I_3
timestamp 1699925102
transform 0 -1 342200 -1 0 283000
box -200 -18300 24200 50600
use PIC  ABCMD_I_4
timestamp 1699925102
transform 1 0 232000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_5
timestamp 1699925102
transform 1 0 205000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_6
timestamp 1699925102
transform 1 0 151000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_7
timestamp 1699925102
transform 1 0 178000 0 -1 342200
box -200 -18300 24200 50600
use PIC  CLK
timestamp 1699925102
transform 0 1 37800 -1 0 175000
box -200 -18300 24200 50600
use PIC  LOADA_I
timestamp 1699925102
transform 1 0 97000 0 -1 342200
box -200 -18300 24200 50600
use PIC  LOADB_I
timestamp 1699925102
transform 0 1 37800 -1 0 283000
box -200 -18300 24200 50600
use PIC  LOADCMD_I
timestamp 1699925102
transform 1 0 124000 0 -1 342200
box -200 -18300 24200 50600
use PIC  RESET
timestamp 1699925102
transform 0 1 37800 -1 0 256000
box -200 -18300 24200 50600
use POB8  ACC_O_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1699924048
transform 0 1 37800 -1 0 148000
box -200 -18300 24200 50600
use POB8  ACC_O_1
timestamp 1699924048
transform 0 1 37800 -1 0 121000
box -200 -18300 24200 50600
use POB8  ACC_O_2
timestamp 1699924048
transform 0 1 37800 -1 0 229000
box -200 -18300 24200 50600
use POB8  ACC_O_3
timestamp 1699924048
transform 1 0 205000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_4
timestamp 1699924048
transform 1 0 178000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_5
timestamp 1699924048
transform 1 0 151000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_6
timestamp 1699924048
transform 1 0 124000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_7
timestamp 1699924048
transform 1 0 97000 0 1 37800
box -200 -18300 24200 50600
use POB8  DONE_O
timestamp 1699924048
transform 1 0 232000 0 1 37800
box -200 -18300 24200 50600
use PVSS  PVSS_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 -1 342200 -1 0 202000
box 0 -18300 24000 50600
use PVDD  VDD_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 1 37800 -1 0 202000
box 0 -18300 24000 50600
use MY_LOGO  MY_LOGO_0
timestamp 1700409309
transform 1 0 299100 0 1 21600
box 0 0 40680 14580
<< end >>