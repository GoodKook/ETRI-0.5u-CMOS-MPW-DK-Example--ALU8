/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module ALU_wrapper(
    inout vdd,
    inout gnd,
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    output Done_o,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input clk,
    input reset
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire BI_0_bF$buf0 ;
wire BI_0_bF$buf1 ;
wire BI_0_bF$buf2 ;
wire BI_0_bF$buf3 ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire \u_ALU.AI7  ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire ABCmd_i_2_bF$buf0 ;
wire ABCmd_i_2_bF$buf1 ;
wire ABCmd_i_2_bF$buf2 ;
wire ABCmd_i_2_bF$buf3 ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _705__bF$buf0 ;
wire _705__bF$buf1 ;
wire _705__bF$buf2 ;
wire _705__bF$buf3 ;
wire _878_ ;
wire _458_ ;
wire _32__bF$buf0 ;
wire _32__bF$buf1 ;
wire _32__bF$buf2 ;
wire _32__bF$buf3 ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire Done_o ;
wire _740_ ;
wire _320_ ;
wire AI_5_bF$buf0 ;
wire AI_5_bF$buf1 ;
wire AI_5_bF$buf2 ;
wire AI_5_bF$buf3 ;
wire _56_ ;
wire _605_ ;
wire BI_4_bF$buf0 ;
wire BI_4_bF$buf1 ;
wire BI_4_bF$buf2 ;
wire BI_4_bF$buf3 ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire [7:0] _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _713_ ;
wire [6:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire BI_1_bF$buf0 ;
wire BI_1_bF$buf1 ;
wire BI_1_bF$buf2 ;
wire BI_1_bF$buf3 ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [2:0] state ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire [6:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire BI_3_bF$buf0 ;
wire BI_3_bF$buf1 ;
wire BI_3_bF$buf2 ;
wire BI_3_bF$buf3 ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire [2:0] _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _0__bF$buf0 ;
wire _0__bF$buf1 ;
wire _0__bF$buf2 ;
wire _0__bF$buf3 ;
wire _0__bF$buf4 ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_0__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf2),
    .B(_825_),
    .C(_863_),
    .Y(_864_)
);

AOI22X1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_324_),
    .C(_358_),
    .D(_359_),
    .Y(_363_)
);

FILL FILL_3__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(_712_),
    .C(_582_),
    .D(_588_),
    .Y(_12_)
);

NAND3X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_166_),
    .C(_171_),
    .Y(_172_)
);

FILL FILL_2__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_365_),
    .C(_399_),
    .Y(_400_)
);

FILL FILL_0__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(BI_3_bF$buf3),
    .Y(_493_)
);

FILL FILL_2__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_705__bF$buf3),
    .Y(_695_)
);

INVX1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .Y(_44_)
);

FILL FILL_1__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_123_),
    .C(_248_),
    .Y(_304_)
);

FILL FILL_2__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_513_),
    .C(_509_),
    .Y(_514_)
);

FILL FILL_1__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .Y(BI_4_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .Y(BI_4_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .Y(BI_4_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .Y(BI_4_bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(BI_1_bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(BI_1_bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(BI_1_bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(BI_1_bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf3)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf2)
);

FILL FILL_2__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_69_),
    .C(_72_),
    .Y(_76_)
);

FILL FILL_1__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_605_),
    .Y(_606_)
);

FILL FILL_3__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_744_),
    .C(_741_),
    .Y(_746_)
);

AND2X2 _1313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(BI_3_bF$buf3),
    .Y(_418_)
);

FILL FILL_1__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_167_),
    .C(_423_),
    .D(_597_),
    .Y(_643_)
);

NAND3X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

FILL FILL_1__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[1]),
    .Y(_42_)
);

OR2X2 _1771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_761_),
    .B(_844_),
    .Y(_782_)
);

OAI21X1 _1351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_455_),
    .C(_361_),
    .Y(_456_)
);

FILL FILL_1__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_498_),
    .Y(_511_)
);

FILL FILL92550x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_679_),
    .C(_712_),
    .Y(_680_)
);

NAND3X1 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_243_),
    .C(_244_),
    .Y(_266_)
);

FILL FILL_1__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf2),
    .Y(_824_)
);

AND2X2 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_317_),
    .Y(_322_)
);

FILL FILL_0__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf0),
    .Y(_73_)
);

FILL FILL_1__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_494_),
    .C(_492_),
    .D(_495_),
    .Y(_548_)
);

NAND2X1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf2),
    .B(AI[6]),
    .Y(_131_)
);

FILL FILL_1__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_860_),
    .B(_848_),
    .Y(_861_)
);

NAND3X1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(_358_),
    .C(_357_),
    .Y(_360_)
);

FILL FILL_0__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[3]),
    .B(_54_),
    .Y(_586_)
);

OAI21X1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_150_),
    .C(_111_),
    .Y(_169_)
);

FILL FILL_0__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_557_),
    .C(_596_),
    .Y(_640_)
);

NAND3X1 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_224_),
    .C(_222_),
    .Y(_225_)
);

FILL FILL_3__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_371_),
    .Y(_397_)
);

FILL FILL_0__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_875_),
    .C(_778_),
    .Y(_779_)
);

NAND3X1 _1348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_452_),
    .C(_451_),
    .Y(_453_)
);

FILL FILL_3__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_675_),
    .C(ABCmd_i[7]),
    .Y(_677_)
);

OAI21X1 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(_173_),
    .C(_171_),
    .Y(_263_)
);

FILL FILL_1__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_486_),
    .Y(_490_)
);

FILL FILL_2__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_289_),
    .C(_300_),
    .Y(_301_)
);

FILL FILL_1__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_176_),
    .C(_390_),
    .Y(_394_)
);

FILL FILL_2__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_600_),
    .Y(_603_)
);

FILL FILL_3__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_149_),
    .C(_198_),
    .Y(_204_)
);

FILL FILL_2__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_742_),
    .Y(_743_)
);

NAND2X1 _1310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(BI[5]),
    .Y(_415_)
);

FILL FILL_1__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .Y(_40_)
);

FILL FILL_1__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91350x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[6]),
    .Y(ACC_o[6])
);

NAND3X1 _1404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_507_),
    .C(_479_),
    .Y(_508_)
);

FILL FILL_1__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1633_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_888_[0]),
    .S(_0__bF$buf0),
    .R(vdd),
    .CLK(clk_bF$buf2),
    .Q(state[0])
);

NAND2X1 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

FILL FILL_0__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf1),
    .B(AI[3]),
    .Y(_70_)
);

FILL FILL_1__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(BI[7]),
    .Y(_545_)
);

NAND2X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_90_),
    .B(_127_),
    .Y(_128_)
);

FILL FILL_1__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .Y(_858_)
);

AND2X2 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_324_),
    .Y(_357_)
);

FILL FILL_0__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_734_),
    .C(_740_),
    .Y(HC)
);

NOR2X1 _1307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_339_),
    .Y(_412_)
);

FILL FILL_3__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .B(_300_),
    .Y(_583_)
);

NAND3X1 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_165_),
    .C(_163_),
    .Y(_166_)
);

FILL FILL_0__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_624_),
    .Y(_637_)
);

OAI21X1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_113_),
    .C(_221_),
    .Y(_222_)
);

FILL FILL_3__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_772_),
    .B(_774_),
    .C(_775_),
    .Y(_776_)
);

NAND3X1 _1345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_442_),
    .C(_449_),
    .Y(_450_)
);

FILL FILL_1__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_393_),
    .Y(_674_)
);

NAND3X1 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_100_),
    .C(_104_),
    .Y(_260_)
);

FILL FILL_1__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_482_),
    .Y(_487_)
);

FILL FILL_0__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_488_),
    .C(_484_),
    .Y(_542_)
);

AOI21X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_116_),
    .C(_118_),
    .Y(_125_)
);

FILL FILL_3__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_298_)
);

FILL FILL_1__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .B(_854_),
    .C(_849_),
    .Y(_855_)
);

AOI21X1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_342_),
    .B(_345_),
    .C(_338_),
    .Y(_354_)
);

FILL FILL_0__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(BI[5]),
    .Y(_105_)
);

FILL FILL_0__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .Y(_580_)
);

OAI21X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_119_),
    .C(_100_),
    .Y(_163_)
);

FILL FILL_0__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_175_),
    .Y(_391_)
);

FILL FILL_2__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .Y(_201_)
);

FILL FILL_0__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .B(_38_),
    .Y(_39_)
);

FILL FILL_1__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .Y(_295_)
);

FILL FILL_2__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[3]),
    .Y(ACC_o[3])
);

INVX1 _1401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_505_)
);

FILL FILL_1__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1630_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(AI[5])
);

INVX1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .Y(_316_)
);

OAI21X1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

FILL FILL_1__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .B(_737_),
    .Y(_738_)
);

OAI22X1 _1304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_408_),
    .C(_327_),
    .D(_335_),
    .Y(_409_)
);

FILL FILL_1__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(_712_),
    .C(_628_),
    .D(_634_),
    .Y(_13_)
);

INVX1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .Y(_219_)
);

FILL FILL_1__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[6]),
    .C(_825_),
    .Y(_773_)
);

OAI21X1 _1342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(_354_),
    .C(_432_),
    .Y(_447_)
);

FILL FILL_1__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[0]),
    .Y(ACC_o[0])
);

FILL FILL_3__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .Y(_671_)
);

NAND3X1 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_253_),
    .C(_254_),
    .Y(_257_)
);

FILL FILL_1__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1627_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf1),
    .Q(AI[2])
);

NAND2X1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_233_),
    .Y(_313_)
);

FILL FILL_0__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

FILL FILL_1__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_483_),
    .Y(_484_)
);

FILL FILL91650x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AV),
    .Y(_539_)
);

NAND3X1 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_121_),
    .C(_88_),
    .Y(_122_)
);

FILL FILL_1__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf1),
    .Y(_852_)
);

NAND3X1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_350_),
    .C(_326_),
    .Y(_351_)
);

FILL FILL_0__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_98_),
    .C(_95_),
    .Y(_102_)
);

FILL FILL_0__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(_573_),
    .Y(_577_)
);

NAND2X1 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_155_),
    .Y(_160_)
);

FILL FILL_0__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_715_),
    .C(_387_),
    .Y(_388_)
);

FILL FILL_0__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI[6]),
    .C(_769_),
    .D(_830_),
    .Y(_770_)
);

AOI21X1 _1339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_357_),
    .B(_359_),
    .C(_443_),
    .Y(_444_)
);

FILL FILL_3__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf2),
    .B(AI[4]),
    .Y(_198_)
);

FILL FILL_2__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(_667_),
    .Y(_668_)
);

NAND3X1 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_75_),
    .C(_72_),
    .Y(_254_)
);

FILL FILL_0__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_707_),
    .C(_887_),
    .Y(_708_)
);

FILL FILL_0__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_803_),
    .Y(AZ)
);

INVX1 _1377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .Y(_481_)
);

FILL FILL_0__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32__bF$buf1),
    .Y(_36_)
);

FILL FILL_1__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_273_),
    .Y(_292_)
);

FILL FILL_1__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(AI[2]),
    .Y(_195_)
);

FILL FILL_2__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_877_),
    .Y(_735_)
);

NOR2X1 _1301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_167_),
    .Y(_406_)
);

FILL FILL_1__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[4]),
    .B(_54_),
    .Y(_632_)
);

OAI21X1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_191_),
    .C(_211_),
    .Y(_216_)
);

FILL FILL_1__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_26_),
    .Y(_34_)
);

FILL FILL_1__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_815_),
    .C(_821_),
    .Y(_822_)
);

FILL FILL_1__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1624_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(_886_[7])
);

AOI21X1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_309_),
    .C(_287_),
    .Y(_310_)
);

FILL FILL_0__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_59_),
    .Y(_61_)
);

FILL FILL_1__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_536_),
    .C(_530_),
    .D(_532_),
    .Y(_537_)
);

AOI21X1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_96_),
    .C(_89_),
    .Y(_119_)
);

FILL FILL_1__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(AI[2]),
    .Y(_849_)
);

NAND2X1 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_341_),
    .Y(_348_)
);

FILL FILL_0__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_98_),
    .C(_94_),
    .Y(_99_)
);

FILL FILL_0__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_731_),
    .C(_732_),
    .Y(_733_)
);

AOI21X1 _1471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_507_),
    .C(_509_),
    .Y(_574_)
);

OAI21X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_143_),
    .C(_156_),
    .Y(_157_)
);

FILL FILL_2__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .Y(_629_)
);

NAND3X1 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_207_),
    .C(_180_),
    .Y(_213_)
);

FILL FILL_3__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[1]),
    .Y(_385_)
);

FILL FILL93150x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .Y(_767_)
);

NAND3X1 _1336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(_440_),
    .C(_439_),
    .Y(_441_)
);

FILL FILL_3__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_664_),
    .Y(_665_)
);

OAI21X1 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_149_),
    .C(_62_),
    .Y(_251_)
);

FILL FILL_0__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_704_),
    .Y(_705_)
);

FILL FILL_0__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(ACC[4]),
    .Y(_803_)
);

INVX1 _1374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .Y(_478_)
);

FILL FILL_0__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_277_),
    .C(_288_),
    .Y(_289_)
);

FILL FILL_1__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_828_),
    .Y(ACC[0])
);

NAND2X1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_344_),
    .Y(_345_)
);

FILL FILL_0__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

OAI21X1 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_109_),
    .C(_147_),
    .Y(_154_)
);

FILL FILL_3__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_882_),
    .C(_835_),
    .Y(_883_)
);

OAI21X1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_382_),
    .C(_380_),
    .Y(_383_)
);

FILL FILL_0__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_189_),
    .C(_186_),
    .Y(_192_)
);

FILL FILL_2__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_708_),
    .C(_25_),
    .Y(_31_)
);

FILL FILL_1__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .Y(_819_)
);

FILL FILL_1__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1621_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(_886_[4])
);

NAND3X1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_307_)
);

INVX2 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf3),
    .Y(_58_)
);

FILL FILL_1__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_298_),
    .C(ABCmd_i[7]),
    .Y(_534_)
);

AND2X2 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_111_),
    .Y(_116_)
);

FILL FILL_1__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

FILL FILL_2__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf0),
    .B(BI_3_bF$buf0),
    .C(_825_),
    .Y(_730_)
);

FILL FILL_1__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(_620_),
    .C(ABCmd_i[7]),
    .Y(_626_)
);

NAND3X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_187_),
    .C(_190_),
    .Y(_210_)
);

FILL FILL_3__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_764_),
    .Y(_765_)
);

XOR2X1 _1333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_405_),
    .Y(_438_)
);

FILL FILL_1__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_844_),
    .C(_794_),
    .Y(_816_)
);

FILL FILL92850x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_639_),
    .B(_646_),
    .C(_661_),
    .Y(_662_)
);

INVX1 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .Y(_248_)
);

FILL FILL_0__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .Y(_702_)
);

FILL FILL_0__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1618_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf2),
    .Q(_886_[1])
);

FILL FILL_0__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_32__bF$buf2),
    .C(_55_),
    .Y(_8_)
);

NAND2X1 _1791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(_797_),
    .Y(AN)
);

INVX1 _1371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .Y(_475_)
);

FILL FILL_2__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(AZ),
    .Y(_531_)
);

INVX1 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .Y(_113_)
);

FILL FILL_3__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_172_),
    .C(_124_),
    .Y(_286_)
);

FILL FILL_1__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .Y(_844_)
);

NAND2X1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_339_),
    .Y(_342_)
);

FILL FILL_0__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .Y(_93_)
);

FILL FILL_1__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_567_),
    .C(_564_),
    .Y(_568_)
);

OAI21X1 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_149_),
    .C(_150_),
    .Y(_151_)
);

FILL FILL93150x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI[2]),
    .C(_879_),
    .D(_830_),
    .Y(_880_)
);

OAI21X1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_377_),
    .C(_379_),
    .Y(_380_)
);

FILL FILL_0__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(_188_),
    .Y(_189_)
);

FILL FILL_0__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .Y(_659_)
);

NAND3X1 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_243_),
    .C(_244_),
    .Y(_245_)
);

FILL FILL_0__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_766_),
    .Y(_798_)
);

NOR2X1 _1368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(_470_),
    .Y(_472_)
);

FILL FILL_3__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_713_),
    .C(_28_),
    .D(_711_),
    .Y(_29_)
);

FILL FILL_1__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_705__bF$buf1),
    .Y(_693_)
);

AOI22X1 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_269_),
    .C(_259_),
    .D(_260_),
    .Y(_283_)
);

FILL FILL93150x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI_3_bF$buf0),
    .C(_726_),
    .D(_830_),
    .Y(_727_)
);

FILL FILL_1__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_573_),
    .B(_618_),
    .C(_474_),
    .Y(_623_)
);

OAI21X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_191_),
    .C(_206_),
    .Y(_207_)
);

FILL FILL_1__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .Y(_26_)
);

FILL FILL_1__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_761_),
    .C(_759_),
    .Y(_762_)
);

OAI21X1 _1330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_434_),
    .C(_348_),
    .Y(_435_)
);

FILL FILL_1__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_813_),
    .B(_810_),
    .Y(_814_)
);

FILL FILL_1__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .B(_699_),
    .Y(_700_)
);

FILL FILL_2__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1615_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf1),
    .Q(BI[6])
);

FILL FILL_0__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_52_),
    .B(_32__bF$buf1),
    .C(_53_),
    .Y(_7_)
);

FILL FILL_1__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .Y(_528_)
);

OAI21X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_109_),
    .C(_82_),
    .Y(_110_)
);

FILL FILL_3__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

AOI21X1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_186_),
    .C(_189_),
    .Y(_339_)
);

FILL FILL_0__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf2),
    .B(AI_5_bF$buf1),
    .Y(_90_)
);

FILL FILL_1__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(AI[4]),
    .Y(_724_)
);

FILL FILL_3__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_501_),
    .C(_506_),
    .Y(_565_)
);

NAND2X1 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_147_),
    .Y(_148_)
);

FILL FILL_0__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_617_),
    .C(_614_),
    .Y(_620_)
);

FILL FILL93150x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_871_),
    .C(_872_),
    .Y(_877_)
);

XOR2X1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_376_),
    .Y(_377_)
);

FILL FILL_0__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_),
    .B(_757_),
    .C(_754_),
    .Y(_759_)
);

NAND2X1 _1327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_427_),
    .Y(_432_)
);

FILL FILL_3__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .Y(_186_)
);

FILL FILL_0__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(_712_),
    .C(_651_),
    .D(_656_),
    .Y(_14_)
);

OAI21X1 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_237_),
    .C(_178_),
    .Y(_242_)
);

FILL FILL_1__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_794_),
    .C(_792_),
    .Y(_795_)
);

OAI21X1 _1365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .B(_699_),
    .C(_886_[2]),
    .Y(_469_)
);

FILL FILL_0__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_705__bF$buf2),
    .C(_691_),
    .Y(_17_)
);

OAI21X1 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_87_),
    .C(_86_),
    .Y(_280_)
);

FILL FILL_1__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_561_),
    .Y(_562_)
);

INVX1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .Y(_145_)
);

FILL FILL_1__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_861_),
    .Y(_875_)
);

NAND3X1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_365_),
    .C(_361_),
    .Y(_374_)
);

FILL FILL_0__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_596_),
    .Y(_599_)
);

AOI22X1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf2),
    .B(\u_ALU.AI7 ),
    .C(BI_1_bF$buf0),
    .D(AI[6]),
    .Y(_183_)
);

FILL FILL_2__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .Y(_714_)
);

FILL FILL_1__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_796_),
    .C(_795_),
    .Y(_811_)
);

FILL FILL_1__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1612_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(BI[3])
);

FILL FILL_0__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_32__bF$buf3),
    .C(_51_),
    .Y(_6_)
);

FILL FILL_1__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_475_),
    .C(_524_),
    .Y(_525_)
);

AND2X2 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf1),
    .B(AI[2]),
    .Y(_107_)
);

FILL FILL_1__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(_836_),
    .C(_837_),
    .Y(_838_)
);

INVX1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .Y(_336_)
);

AOI21X1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_79_),
    .C(_67_),
    .Y(_87_)
);

FILL FILL_1__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf0),
    .B(_825_),
    .C(_720_),
    .Y(_721_)
);

FILL FILL_3__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_616_),
    .C(_615_),
    .Y(_617_)
);

FILL FILL_1__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf0),
    .B(_755_),
    .Y(_756_)
);

NAND3X1 _1324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_421_),
    .C(_419_),
    .Y(_429_)
);

FILL FILL_1__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[5]),
    .Y(_654_)
);

OAI21X1 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_232_),
    .C(_229_),
    .Y(_239_)
);

FILL FILL_1__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1609_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(BI[0])
);

FILL FILL_0__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_790_),
    .C(_787_),
    .Y(_792_)
);

OAI21X1 _1362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_464_),
    .C(_465_),
    .Y(_467_)
);

FILL FILL_0__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_521_),
    .C(_442_),
    .Y(_522_)
);

FILL FILL_3__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_703_),
    .C(_712_),
    .Y(_690_)
);

NAND3X1 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_275_),
    .C(_270_),
    .Y(_277_)
);

FILL FILL_1__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .Y(_835_)
);

INVX1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .Y(_333_)
);

FILL FILL_0__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf1),
    .B(AI[1]),
    .Y(_84_)
);

FILL FILL_1__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_558_),
    .C(_494_),
    .Y(_559_)
);

NAND3X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_133_),
    .C(_128_),
    .Y(_142_)
);

FILL FILL_3__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_857_),
    .C(_855_),
    .Y(_872_)
);

OAI21X1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_366_),
    .B(_370_),
    .C(_312_),
    .Y(_371_)
);

FILL FILL_0__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .B(_593_),
    .Y(_596_)
);

AOI21X1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_156_),
    .C(_143_),
    .Y(_180_)
);

FILL FILL_0__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .Y(BI_3_bF$buf3)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .Y(BI_3_bF$buf2)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .Y(BI_3_bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .Y(BI_3_bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(BI_0_bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(BI_0_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(BI_0_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(BI_0_bF$buf0)
);

FILL FILL_0__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .Y(_789_)
);

AND2X2 _1359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_293_),
    .Y(_464_)
);

FILL FILL_3__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .Y(_711_)
);

FILL FILL_1__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_310_),
    .Y(_687_)
);

AOI22X1 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf1),
    .B(AI[2]),
    .C(BI_1_bF$buf1),
    .D(AI[1]),
    .Y(_274_)
);

FILL FILL_2__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_807_),
    .Y(_808_)
);

FILL FILL_1__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .Y(_501_)
);

FILL FILL_0__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(_32__bF$buf0),
    .C(_49_),
    .Y(_5_)
);

FILL FILL_1__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_718_),
    .Y(_719_)
);

FILL FILL_1__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_611_),
    .Y(_614_)
);

FILL FILL_3__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_751_),
    .C(_752_),
    .Y(_753_)
);

AOI21X1 _1321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_425_),
    .C(_415_),
    .Y(_426_)
);

FILL FILL_1__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

OAI21X1 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_232_),
    .C(_235_),
    .Y(_236_)
);

FILL FILL_1__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_52_),
    .B(_705__bF$buf1),
    .C(_697_),
    .Y(_23_)
);

FILL FILL_0__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(_32__bF$buf0),
    .C(_47_),
    .Y(_4_)
);

FILL FILL_1__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_515_),
    .Y(_519_)
);

FILL FILL_1__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf1),
    .B(_831_),
    .Y(_832_)
);

AND2X2 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf2),
    .B(BI_3_bF$buf2),
    .Y(_330_)
);

FILL FILL_0__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .Y(_81_)
);

FILL FILL_1__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(BI[5]),
    .Y(_556_)
);

AOI21X1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_135_),
    .C(_126_),
    .Y(_139_)
);

FILL FILL_1__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_571_),
    .C(_610_),
    .Y(_611_)
);

NAND2X1 _1682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_867_),
    .Y(_869_)
);

NAND3X1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_360_),
    .C(_362_),
    .Y(_368_)
);

FILL FILL_0__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .Y(_751_)
);

INVX2 _1318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .Y(_423_)
);

FILL FILL_3__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf3),
    .B(BI[7]),
    .Y(_593_)
);

NAND2X1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_169_),
    .Y(_177_)
);

FILL FILL_0__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_647_),
    .Y(_648_)
);

NAND3X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_227_),
    .C(_226_),
    .Y(_233_)
);

FILL FILL_1__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .B(_783_),
    .C(_775_),
    .Y(_786_)
);

AND2X2 _1356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_460_),
    .Y(_461_)
);

FILL FILL_1__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_683_),
    .Y(_684_)
);

NAND2X1 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf3),
    .B(AI[1]),
    .Y(_271_)
);

FILL FILL_1__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .B(_492_),
    .Y(_498_)
);

FILL FILL_0__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91350x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf1),
    .B(_833_),
    .Y(_866_)
);

OAI21X1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_364_),
    .C(_362_),
    .Y(_365_)
);

FILL FILL_3__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_550_),
    .C(_549_),
    .Y(_590_)
);

AOI21X1 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_161_),
    .C(_125_),
    .Y(_174_)
);

FILL FILL_2__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[2]),
    .C(_885_),
    .Y(_716_)
);

FILL FILL91950x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .Y(_402_)
);

FILL FILL_2__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf0),
    .B(_705__bF$buf2),
    .Y(_696_)
);

FILL FILL_0__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_32__bF$buf2),
    .C(_45_),
    .Y(_3_)
);

FILL FILL_1__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .B(_502_),
    .C(_509_),
    .Y(_516_)
);

FILL FILL_1__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[1]),
    .Y(_829_)
);

NAND2X1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(AI[3]),
    .Y(_327_)
);

AND2X2 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_71_),
    .Y(_78_)
);

FILL FILL_1__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_553_)
);

NOR2X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_131_),
    .Y(_136_)
);

FILL FILL_1__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_563_),
    .Y(_608_)
);

FILL FILL_3__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_4_bF$buf3),
    .C(_747_),
    .Y(_748_)
);

AOI22X1 _1315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(BI_3_bF$buf3),
    .C(AI_5_bF$buf3),
    .D(BI_4_bF$buf1),
    .Y(_420_)
);

FILL FILL_1__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_644_),
    .Y(_645_)
);

NAND3X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_213_),
    .C(_217_),
    .Y(_230_)
);

FILL FILL_1__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .Y(_784_)
);

NAND3X1 _1353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_452_),
    .C(_451_),
    .Y(_458_)
);

FILL FILL_1__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(_512_),
    .C(_490_),
    .Y(_513_)
);

INVX1 _1582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[7]),
    .Y(_681_)
);

AOI21X1 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_266_),
    .C(_265_),
    .Y(_268_)
);

FILL FILL_1__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(_825_),
    .C(ABCmd_i[4]),
    .Y(_826_)
);

OAI21X1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_322_),
    .C(_315_),
    .Y(_324_)
);

FILL FILL_0__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_74_),
    .C(_70_),
    .Y(_75_)
);

AOI22X1 _1391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(BI_3_bF$buf3),
    .C(AI[6]),
    .D(BI_4_bF$buf1),
    .Y(_495_)
);

FILL FILL_0__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_548_),
    .Y(_550_)
);

NAND2X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[4]),
    .Y(_133_)
);

FILL FILL_3__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_824_),
    .C(_862_),
    .Y(_863_)
);

AOI21X1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .B(_229_),
    .C(_232_),
    .Y(_362_)
);

FILL FILL_0__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_587_),
    .B(_703_),
    .C(_712_),
    .Y(_588_)
);

INVX1 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_171_)
);

FILL FILL_0__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .Y(_399_)
);

FILL FILL_0__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_25_),
    .Y(_679_)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_262_),
    .C(_263_),
    .D(_264_),
    .Y(_265_)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf3),
    .B(BI[5]),
    .Y(_492_)
);

FILL FILL_2__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(_705__bF$buf3),
    .C(_694_),
    .Y(_20_)
);

OAI21X1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_32__bF$buf3),
    .C(_43_),
    .Y(_2_)
);

FILL FILL_1__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_301_),
    .C(_282_),
    .Y(_303_)
);

FILL FILL_1__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_0__bF$buf1)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_0__bF$buf0)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .Y(AI_5_bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .Y(AI_5_bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .Y(AI_5_bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .Y(AI_5_bF$buf0)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .Y(_32__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .Y(_32__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .Y(_32__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .Y(_32__bF$buf0)
);

FILL FILL_2__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_603_),
    .Y(_605_)
);

FILL FILL_1__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_742_),
    .C(_835_),
    .Y(_745_)
);

AND2X2 _1312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf3),
    .B(BI_4_bF$buf1),
    .Y(_417_)
);

FILL FILL_1__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(BI[6]),
    .C(_641_),
    .Y(_642_)
);

OAI21X1 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_113_),
    .C(_220_),
    .Y(_227_)
);

FILL FILL_1__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_32__bF$buf3),
    .C(_41_),
    .Y(_1_)
);

FILL FILL_1__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_780_),
    .C(_749_),
    .Y(_781_)
);

AOI21X1 _1350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_455_)
);

FILL FILL_1__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(Done_o)
);

AOI22X1 _1406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .B(_489_),
    .C(_506_),
    .D(_500_),
    .Y(_510_)
);

FILL FILL_3__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1635_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_888_[2]),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf3),
    .Q(state[2])
);

NAND3X1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_319_),
    .C(_320_),
    .Y(_321_)
);

FILL FILL_0__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_71_),
    .Y(_72_)
);

FILL FILL_2_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_167_),
    .Y(_547_)
);

INVX2 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf3),
    .Y(_130_)
);

FILL FILL_1__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_858_),
    .S(_855_),
    .Y(_860_)
);

OAI21X1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_359_)
);

FILL FILL_0__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(BI_4_bF$buf3),
    .Y(_742_)
);

NAND2X1 _1309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(BI[2]),
    .Y(_414_)
);

FILL FILL_3__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_301_),
    .B(_584_),
    .Y(_585_)
);

NOR2X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_167_),
    .Y(_168_)
);

FILL FILL92550x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_605_),
    .C(_604_),
    .Y(_639_)
);

NAND2X1 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_220_),
    .Y(_224_)
);

FILL FILL_3__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_395_),
    .B(_389_),
    .C(_246_),
    .Y(_396_)
);

FILL FILL_2__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .Y(_778_)
);

OAI21X1 _1347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_448_),
    .C(_404_),
    .Y(_452_)
);

FILL FILL_3__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_309_),
    .C(_308_),
    .Y(_676_)
);

NAND3X1 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_122_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_488_),
    .B(_487_),
    .C(_480_),
    .Y(_489_)
);

FILL FILL_0__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_299_),
    .C(_81_),
    .Y(_300_)
);

FILL FILL_1__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_581_),
    .C(_540_),
    .Y(_582_)
);

OAI21X1 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_143_),
    .C(_160_),
    .Y(_165_)
);

FILL FILL_0__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_390_),
    .C(_392_),
    .Y(_393_)
);

FILL FILL_2__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_598_),
    .C(_596_),
    .Y(_602_)
);

FILL FILL_1__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_74_),
    .C(_197_),
    .Y(_203_)
);

FILL FILL_2__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .Y(_0_)
);

FILL FILL_1__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[5]),
    .Y(ACC_o[5])
);

NAND3X1 _1403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_500_),
    .C(_503_),
    .Y(_507_)
);

FILL FILL_1__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1632_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(\u_ALU.AI7 )
);

OAI21X1 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_200_),
    .C(_199_),
    .Y(_318_)
);

FILL FILL_0__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .Y(_69_)
);

FILL FILL_1__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_500_),
    .C(_499_),
    .Y(_544_)
);

AND2X2 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf0),
    .B(AI[6]),
    .Y(_127_)
);

FILL FILL_1__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_1_bF$buf3),
    .C(_856_),
    .Y(_857_)
);

NAND3X1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_355_),
    .C(_351_),
    .Y(_356_)
);

FILL FILL_0__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .Y(_740_)
);

XNOR2X1 _1306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_405_),
    .Y(_411_)
);

FILL FILL_3__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_387_),
    .Y(_636_)
);

INVX1 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .Y(_221_)
);

FILL FILL_1__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_774_),
    .C(_772_),
    .Y(_775_)
);

OAI21X1 _1344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_448_),
    .C(_444_),
    .Y(_449_)
);

FILL FILL_1__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_669_),
    .C(_672_),
    .Y(_673_)
);

OAI21X1 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_119_),
    .C(_116_),
    .Y(_259_)
);

FILL FILL_1__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1629_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(AI[4])
);

NAND2X1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .B(AI[1]),
    .Y(_315_)
);

FILL FILL_0__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(_484_),
    .C(_485_),
    .Y(_486_)
);

FILL FILL_0__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .Y(_541_)
);

OAI21X1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_123_),
    .C(_122_),
    .Y(_124_)
);

NAND3X1 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_296_),
    .C(_292_),
    .Y(_297_)
);

FILL FILL_1__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_853_),
    .C(_835_),
    .Y(_854_)
);

AOI22X1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_337_),
    .C(_349_),
    .D(_348_),
    .Y(_353_)
);

FILL FILL_0__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(_102_),
    .C(_101_),
    .Y(_104_)
);

FILL FILL_0__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_528_),
    .C(_541_),
    .Y(_579_)
);

NAND3X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_125_),
    .C(_157_),
    .Y(_162_)
);

FILL FILL_0__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .Y(_390_)
);

FILL FILL_0__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf2),
    .B(AI[4]),
    .C(BI_4_bF$buf2),
    .D(AI[3]),
    .Y(_200_)
);

FILL FILL_0__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_786_),
    .Y(_807_)
);

OAI21X1 _1379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_420_),
    .C(_419_),
    .Y(_483_)
);

FILL FILL_0__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_714_),
    .C(_715_),
    .Y(_38_)
);

FILL FILL_1__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_293_),
    .Y(_294_)
);

FILL FILL_2__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[2]),
    .Y(ACC_o[2])
);

NAND2X1 _1400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_431_),
    .Y(_504_)
);

FILL FILL_1__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_63_),
    .Y(_66_)
);

FILL FILL_1__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .B(_875_),
    .C(_736_),
    .Y(_737_)
);

NAND2X1 _1303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf2),
    .B(BI_4_bF$buf2),
    .Y(_408_)
);

FILL FILL93150x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_703_),
    .C(_712_),
    .Y(_634_)
);

NAND2X1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(BI[7]),
    .Y(_218_)
);

FILL FILL_1__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_35_),
    .Y(_888_[1])
);

OAI22X1 _1761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_767_),
    .C(_771_),
    .D(_770_),
    .Y(_772_)
);

NAND3X1 _1341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_431_),
    .C(_413_),
    .Y(_446_)
);

FILL FILL_1__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_822_),
    .B(_823_),
    .Y(AV)
);

FILL FILL_3__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_617_),
    .C(_658_),
    .Y(_670_)
);

AND2X2 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_85_),
    .Y(_256_)
);

FILL FILL_1__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1626_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(AI[1])
);

AOI21X1 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_243_),
    .C(_241_),
    .Y(_312_)
);

FILL FILL_0__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf0),
    .B(AI[3]),
    .Y(_63_)
);

FILL FILL_1__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[3]),
    .Y(_538_)
);

OAI21X1 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_119_),
    .C(_120_),
    .Y(_121_)
);

FILL FILL93150x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI_1_bF$buf3),
    .C(_850_),
    .D(_830_),
    .Y(_851_)
);

NAND3X1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_349_),
    .C(_347_),
    .Y(_350_)
);

FILL FILL_0__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_75_),
    .C(_77_),
    .Y(_101_)
);

FILL FILL_0__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .B(_571_),
    .C(_575_),
    .Y(_576_)
);

NAND3X1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_135_),
    .C(_138_),
    .Y(_159_)
);

FILL FILL_0__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_629_),
    .Y(_631_)
);

NAND3X1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_209_),
    .C(_206_),
    .Y(_215_)
);

FILL FILL_3__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_712_),
    .C(ABCmd_i[7]),
    .Y(_387_)
);

FILL FILL_0__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x50850 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_768_),
    .Y(_769_)
);

NOR3X1 _1338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_443_)
);

AND2X2 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf0),
    .B(AI[3]),
    .Y(_197_)
);

FILL FILL_2__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_167_),
    .C(_641_),
    .Y(_667_)
);

OAI21X1 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_78_),
    .C(_69_),
    .Y(_253_)
);

FILL FILL_0__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(_702_),
    .Y(_707_)
);

FILL FILL_0__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_804_),
    .B(AN),
    .Y(_805_)
);

NAND2X1 _1376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(BI[7]),
    .Y(_480_)
);

FILL FILL_0__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_271_),
    .C(_290_),
    .Y(_291_)
);

FILL FILL_1__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[2]),
    .C(_825_),
    .Y(_885_)
);

OAI21X1 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_700_),
    .C(_384_),
    .Y(_9_)
);

FILL FILL_0__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_135_),
    .C(_192_),
    .D(_193_),
    .Y(_194_)
);

FILL FILL_2__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _1720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_733_),
    .Y(_734_)
);

NAND2X1 _1300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(BI[7]),
    .Y(_405_)
);

FILL FILL_1__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_26_),
    .Y(_33_)
);

FILL FILL_1__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_820_),
    .Y(_821_)
);

FILL FILL_1__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1623_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(_886_[6])
);

OAI21X1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_286_),
    .C(_285_),
    .Y(_309_)
);

FILL FILL_0__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf0),
    .B(AI[1]),
    .Y(_60_)
);

FILL FILL_1__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .B(_25_),
    .Y(_536_)
);

AOI21X1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_103_),
    .C(_101_),
    .Y(_118_)
);

FILL FILL_1__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_847_),
    .C(_845_),
    .Y(_848_)
);

AND2X2 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_337_),
    .Y(_347_)
);

NOR2X1 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_97_),
    .Y(_98_)
);

FILL FILL_0__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_731_),
    .C(_729_),
    .Y(_732_)
);

FILL FILL_3__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_518_),
    .C(_572_),
    .Y(_573_)
);

AND2X2 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_152_),
    .Y(_156_)
);

FILL FILL_2__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_25_),
    .B(_627_),
    .C(_626_),
    .Y(_628_)
);

NAND3X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_210_),
    .C(_209_),
    .Y(_212_)
);

FILL FILL91950x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_753_),
    .C(_762_),
    .Y(_766_)
);

NAND2X1 _1335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(_413_),
    .Y(_440_)
);

FILL FILL_1__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .Y(_664_)
);

INVX1 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_65_),
    .Y(_250_)
);

FILL FILL_0__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(_703_),
    .Y(_704_)
);

FILL FILL_0__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_801_),
    .Y(_802_)
);

OAI21X1 _1373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_410_),
    .C(_476_),
    .Y(_477_)
);

FILL FILL_0__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_296_),
    .C(_294_),
    .Y(_533_)
);

NAND3X1 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_112_),
    .C(_114_),
    .Y(_115_)
);

FILL FILL_3__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .Y(_288_)
);

FILL FILL_1__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_843_),
    .C(_845_),
    .Y(_846_)
);

XNOR2X1 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_340_),
    .Y(_344_)
);

FILL FILL_0__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .Y(_95_)
);

FILL FILL_0__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_561_),
    .B(_566_),
    .C(_544_),
    .Y(_570_)
);

OAI21X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_149_),
    .C(_146_),
    .Y(_153_)
);

FILL FILL_0__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(_881_),
    .Y(_882_)
);

OAI21X1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[0]),
    .B(ABCmd_i[7]),
    .C(_715_),
    .Y(_382_)
);

FILL FILL_0__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_187_),
    .C(_181_),
    .Y(_191_)
);

FILL FILL_0__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(LoadB_i),
    .C(_26_),
    .Y(_30_)
);

FILL FILL_1__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_705__bF$buf3),
    .Y(_694_)
);

NAND3X1 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .B(_282_),
    .C(_284_),
    .Y(_285_)
);

FILL FILL_2__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(_817_),
    .C(_797_),
    .Y(_818_)
);

FILL FILL_1__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1620_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(_886_[3])
);

NAND3X1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .B(_305_),
    .C(_304_),
    .Y(_306_)
);

INVX1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .Y(_57_)
);

FILL FILL_1__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .B(_727_),
    .C(_724_),
    .Y(_729_)
);

FILL FILL_1__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_613_),
    .C(_624_),
    .D(_622_),
    .Y(_625_)
);

NAND3X1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .B(_192_),
    .C(_208_),
    .Y(_209_)
);

FILL FILL_1__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .Y(_764_)
);

OAI21X1 _1332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(_433_),
    .C(_411_),
    .Y(_437_)
);

FILL FILL_1__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .B(_804_),
    .C(AN),
    .Y(_815_)
);

NAND2X1 _1561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_647_),
    .Y(_661_)
);

INVX1 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .Y(_247_)
);

FILL FILL_1__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .Y(_887_)
);

FILL FILL_0__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1617_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(_886_[0])
);

FILL FILL_0__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .B(_32__bF$buf2),
    .Y(_55_)
);

FILL FILL_1__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_799_),
    .C(_798_),
    .Y(_800_)
);

AOI21X1 _1370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_459_),
    .C(_470_),
    .Y(_474_)
);

FILL FILL_2__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .B(_529_),
    .C(ABCmd_i[7]),
    .Y(_530_)
);

OAI21X1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_109_),
    .C(_60_),
    .Y(_112_)
);

FILL FILL_3__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf0),
    .B(ABCmd_i_2_bF$buf2),
    .C(_842_),
    .Y(_843_)
);

XOR2X1 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_340_),
    .Y(_341_)
);

FILL FILL_0__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf3),
    .B(AI_5_bF$buf1),
    .C(BI_1_bF$buf2),
    .D(AI[4]),
    .Y(_92_)
);

FILL FILL_1__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_561_),
    .B(_566_),
    .C(_565_),
    .Y(_567_)
);

NAND2X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf0),
    .B(AI[2]),
    .Y(_150_)
);

FILL FILL_0__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(BI[2]),
    .C(_831_),
    .Y(_879_)
);

NOR2X1 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_715_),
    .Y(_379_)
);

FILL FILL_0__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[5]),
    .C(_760_),
    .Y(_761_)
);

NOR2X1 _1329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_341_),
    .Y(_434_)
);

FILL FILL_3__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf0),
    .B(\u_ALU.AI7 ),
    .Y(_188_)
);

FILL FILL_0__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_647_),
    .C(_611_),
    .Y(_658_)
);

NAND3X1 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_236_),
    .C(_179_),
    .Y(_244_)
);

FILL FILL_3__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .Y(_699_)
);

FILL FILL_2__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_786_),
    .Y(_797_)
);

AOI22X1 _1367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_374_),
    .C(_453_),
    .D(_450_),
    .Y(_471_)
);

FILL FILL_0__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_25_),
    .C(_27_),
    .Y(_28_)
);

FILL FILL_1__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_705__bF$buf3),
    .C(_692_),
    .Y(_18_)
);

INVX1 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .Y(_282_)
);

FILL FILL_1__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .Y(_601_)
);

NAND2X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI_5_bF$buf2),
    .Y(_185_)
);

FILL FILL_2__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_725_),
    .Y(_726_)
);

FILL FILL_1__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_577_),
    .C(_621_),
    .Y(_622_)
);

AND2X2 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

FILL FILL_3__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .Y(_25_)
);

FILL FILL_1__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .B(_812_),
    .C(_811_),
    .Y(_813_)
);

FILL FILL_1__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1614_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(BI[5])
);

FILL FILL_0__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_32__bF$buf1),
    .Y(_53_)
);

FILL FILL_1__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_526_),
    .C(_475_),
    .Y(_527_)
);

INVX1 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .Y(_109_)
);

FILL FILL_1__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(ABCmd_i[5]),
    .Y(_840_)
);

NAND2X1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_337_),
    .B(_332_),
    .Y(_338_)
);

FILL FILL_0__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_78_),
    .C(_72_),
    .Y(_89_)
);

FILL FILL_1__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_721_),
    .C(_877_),
    .D(_722_),
    .Y(_723_)
);

FILL FILL_3__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_563_),
    .C(_544_),
    .Y(_564_)
);

AND2X2 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf1),
    .B(AI[3]),
    .Y(_147_)
);

FILL FILL_0__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_573_),
    .B(_618_),
    .C(_616_),
    .D(_474_),
    .Y(_619_)
);

FILL FILL_3__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_855_),
    .Y(_876_)
);

AND2X2 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_375_),
    .Y(_376_)
);

FILL FILL92250x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf0),
    .B(_755_),
    .C(_835_),
    .Y(_758_)
);

NAND3X1 _1326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_429_),
    .C(_428_),
    .Y(_431_)
);

FILL FILL_3__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_653_),
    .B(_655_),
    .C(_712_),
    .Y(_656_)
);

AOI21X1 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(_240_),
    .C(_238_),
    .Y(_241_)
);

FILL FILL_1__917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[7]),
    .C(_793_),
    .Y(_794_)
);

AOI22X1 _1364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_712_),
    .C(_463_),
    .D(_468_),
    .Y(_10_)
);

FILL FILL_0__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(_705__bF$buf2),
    .Y(_691_)
);

OAI21X1 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

FILL FILL_1__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .Y(_837_)
);

AOI22X1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI_5_bF$buf2),
    .B(BI_3_bF$buf2),
    .C(BI_4_bF$buf2),
    .D(AI[4]),
    .Y(_335_)
);

FILL FILL_0__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_554_),
    .C(_560_),
    .Y(_561_)
);

NAND2X1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(AI[1]),
    .Y(_144_)
);

FILL FILL_3__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_871_),
    .B(_873_),
    .Y(_874_)
);

NAND3X1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_369_),
    .C(_368_),
    .Y(_373_)
);

FILL FILL_3__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_597_),
    .C(_595_),
    .Y(_598_)
);

NAND3X1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf2),
    .B(\u_ALU.AI7 ),
    .C(_127_),
    .Y(_182_)
);

FILL FILL_2__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91350x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__901_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(state[0]),
    .C(_699_),
    .Y(_713_)
);

FILL FILL_1__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_837_),
    .B(_835_),
    .Y(_810_)
);

FILL FILL_1__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .B(_489_),
    .Y(_503_)
);

FILL FILL_0__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1611_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf1),
    .Q(BI[2])
);

NAND2X1 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(_32__bF$buf2),
    .Y(_51_)
);

FILL FILL_1__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

FILL FILL_1__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

NAND2X1 _1420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_520_),
    .Y(_524_)
);

INVX1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .Y(_106_)
);

FILL FILL_3__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_81_),
    .C(_85_),
    .Y(_86_)
);

FILL FILL_1__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .Y(_720_)
);

FILL FILL_1__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_524_),
    .Y(_616_)
);

FILL FILL_3__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(BI[5]),
    .Y(_755_)
);

NAND3X1 _1323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_424_),
    .C(_425_),
    .Y(_428_)
);

FILL FILL_1__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_308_),
    .C(ABCmd_i[7]),
    .Y(_653_)
);

AOI21X1 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_171_),
    .C(_174_),
    .Y(_238_)
);

FILL FILL_1__914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_705__bF$buf0),
    .C(_698_),
    .Y(_24_)
);

FILL FILL_0__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf3),
    .B(_32__bF$buf0),
    .Y(_49_)
);

OAI21X1 _1781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .C(_835_),
    .Y(_791_)
);

OAI21X1 _1361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_293_),
    .C(ABCmd_i[7]),
    .Y(_466_)
);

FILL FILL_0__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_441_),
    .C(_404_),
    .Y(_521_)
);

FILL FILL_1__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_687_),
    .C(_688_),
    .Y(_689_)
);

OAI21X1 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_66_),
    .C(_65_),
    .Y(_276_)
);

FILL FILL_1__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf1),
    .B(_833_),
    .C(_830_),
    .D(_832_),
    .Y(_834_)
);

NAND3X1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_329_),
    .C(_331_),
    .Y(_332_)
);

FILL FILL_0__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf2),
    .Y(_83_)
);

FILL FILL_1__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .Y(_558_)
);

OAI21X1 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_136_),
    .C(_134_),
    .Y(_141_)
);

FILL FILL92250x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_864_),
    .C(_870_),
    .D(_827_),
    .Y(_871_)
);

AOI21X1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_369_),
    .C(_367_),
    .Y(_370_)
);

FILL FILL_0__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_557_),
    .C(_594_),
    .Y(_595_)
);

OAI21X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_173_),
    .C(_166_),
    .Y(_179_)
);

FILL FILL_0__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_620_),
    .C(_647_),
    .Y(_650_)
);

NAND2X1 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

FILL FILL_0__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(BI[7]),
    .Y(_788_)
);

OAI21X1 _1358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_461_),
    .C(_388_),
    .Y(_463_)
);

FILL FILL_0__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .B(_709_),
    .C(LoadB_i),
    .Y(_710_)
);

FILL FILL_1__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_247_),
    .Y(_686_)
);

NAND2X1 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(BI[2]),
    .Y(_273_)
);

FILL FILL_1__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_500_)
);

FILL FILL_0__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_716_),
    .C(_717_),
    .Y(_718_)
);

FILL FILL_1__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_403_),
    .C(_358_),
    .Y(_404_)
);

FILL FILL_2__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_612_),
    .B(_609_),
    .C(_607_),
    .Y(_613_)
);

FILL FILL_1__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .Y(_752_)
);

OAI21X1 _1320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_83_),
    .C(_418_),
    .Y(_425_)
);

FILL FILL92550x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_705__bF$buf1),
    .Y(_697_)
);

FILL FILL_0__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf1),
    .B(_32__bF$buf0),
    .Y(_47_)
);

FILL FILL_1__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_516_),
    .C(_517_),
    .Y(_518_)
);

FILL FILL_1__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .Y(_831_)
);

OAI21X1 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_58_),
    .C(_328_),
    .Y(_329_)
);

FILL FILL_0__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_67_),
    .C(_76_),
    .Y(_80_)
);

FILL FILL_1__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(BI_4_bF$buf1),
    .Y(_555_)
);

OAI21X1 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_136_),
    .C(_133_),
    .Y(_138_)
);

FILL FILL_0_CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .B(_607_),
    .Y(_610_)
);

FILL FILL_3__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(_837_),
    .C(ABCmd_i[5]),
    .Y(_868_)
);

INVX1 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .Y(_367_)
);

FILL FILL_0__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .B(_748_),
    .C(_749_),
    .Y(_750_)
);

AOI21X1 _1317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_421_),
    .C(_416_),
    .Y(_422_)
);

FILL FILL_1__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .Y(_592_)
);

NAND3X1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_175_),
    .C(_124_),
    .Y(_176_)
);

FILL FILL_0__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_639_),
    .B(_646_),
    .Y(_647_)
);

AOI21X1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_212_),
    .C(_180_),
    .Y(_232_)
);

FILL FILL92250x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_785_),
    .Y(ACC[6])
);

NAND2X1 _1355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_454_),
    .Y(_460_)
);

FILL FILL_1__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_642_),
    .C(_666_),
    .Y(_683_)
);

NAND3X1 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_250_),
    .C(_64_),
    .Y(_270_)
);

FILL FILL_1__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_494_),
    .C(_496_),
    .Y(_497_)
);

FILL FILL_0__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__904_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_549_),
    .C(_551_),
    .Y(_552_)
);

NAND3X1 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

FILL FILL_3__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[1]),
    .B(_836_),
    .S(ABCmd_i[0]),
    .Y(_865_)
);

AOI21X1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_355_),
    .C(_325_),
    .Y(_364_)
);

FILL FILL_0__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[4]),
    .Y(_589_)
);

AOI21X1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_164_),
    .C(_163_),
    .Y(_173_)
);

FILL FILL_2__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_323_),
    .C(_319_),
    .Y(_401_)
);

FILL FILL_2__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(_705__bF$buf2),
    .C(_695_),
    .Y(_21_)
);

FILL FILL_0__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(_32__bF$buf2),
    .Y(_45_)
);

FILL FILL_1__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_122_),
    .C(_261_),
    .Y(_305_)
);

FILL FILL_2__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(_514_),
    .C(_508_),
    .Y(_515_)
);

FILL FILL_1__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf1)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf0)
);

FILL FILL_2__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_827_),
    .Y(_828_)
);

AOI21X1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_209_),
    .C(_194_),
    .Y(_326_)
);

NOR2X1 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_71_),
    .Y(_77_)
);

FILL FILL_1__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_606_),
    .C(_591_),
    .Y(_607_)
);

FILL FILL_1__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_4_bF$buf3),
    .C(_825_),
    .Y(_747_)
);

NAND2X1 _1314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_418_),
    .Y(_419_)
);

FILL FILL_1__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_642_),
    .Y(_644_)
);

NAND2X1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_225_),
    .Y(_229_)
);

FILL FILL_1__905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_782_),
    .C(_781_),
    .D(_764_),
    .Y(_783_)
);

NAND3X1 _1352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_442_),
    .C(_449_),
    .Y(_457_)
);

FILL FILL_1__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_504_),
    .Y(_512_)
);

FILL FILL_3__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_657_),
    .B(_712_),
    .C(_673_),
    .D(_680_),
    .Y(_15_)
);

OAI21X1 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_237_),
    .C(_177_),
    .Y(_267_)
);

FILL FILL_1__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _1637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[3]),
    .Y(_825_)
);

NOR2X1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_318_),
    .Y(_323_)
);

FILL FILL_0__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .Y(_74_)
);

FILL FILL_1__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(BI_4_bF$buf1),
    .Y(_494_)
);

FILL FILL_0__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_548_),
    .Y(_549_)
);

OAI21X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_130_),
    .C(_131_),
    .Y(_132_)
);

FILL FILL_3__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .Y(_862_)
);

NAND3X1 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_361_)
);

FILL FILL_0__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_585_),
    .C(_586_),
    .Y(_587_)
);

XNOR2X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_168_),
    .Y(_170_)
);

FILL FILL_0__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_396_),
    .C(_375_),
    .Y(_398_)
);

FILL FILL_0__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(ACC[3]),
    .C(_739_),
    .Y(_780_)
);

NAND3X1 _1349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(_453_),
    .C(_400_),
    .Y(_454_)
);

FILL FILL_3__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(ACC[6]),
    .Y(_678_)
);

NAND3X1 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_162_),
    .C(_166_),
    .Y(_264_)
);

FILL FILL_0__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_340_),
    .Y(_491_)
);

FILL FILL_2__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf2),
    .B(_32__bF$buf3),
    .Y(_43_)
);

FILL FILL_1__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_269_),
    .C(_279_),
    .Y(_302_)
);

FILL FILL_1__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .Y(_705__bF$buf3)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .Y(_705__bF$buf2)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .Y(_705__bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .Y(_705__bF$buf0)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_0__bF$buf4)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_0__bF$buf3)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(_0__bF$buf2)
);

FILL FILL_0__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_603_),
    .Y(_604_)
);

FILL FILL_1__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_203_),
    .C(_204_),
    .Y(_205_)
);

FILL FILL_2__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI_4_bF$buf3),
    .C(_743_),
    .D(_830_),
    .Y(_744_)
);

INVX1 _1311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .Y(_416_)
);

FILL FILL_1__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_597_),
    .Y(_641_)
);

NAND2X1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_221_),
    .Y(_226_)
);

FILL FILL_1__902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf3),
    .B(_32__bF$buf3),
    .Y(_41_)
);

FILL FILL_1__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[7]),
    .Y(ACC_o[7])
);

OAI21X1 _1405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_411_),
    .B(_436_),
    .C(_439_),
    .Y(_509_)
);

FILL FILL_1__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1634_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_888_[1]),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(state[1])
);

OR2X2 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_317_),
    .Y(_320_)
);

FILL FILL_0__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf3),
    .B(AI[4]),
    .Y(_71_)
);

FILL FILL_1__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .Y(_546_)
);

INVX1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf2),
    .Y(_129_)
);

FILL FILL_1__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf0),
    .B(_825_),
    .C(_858_),
    .Y(_859_)
);

NAND3X1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_358_)
);

FILL FILL_0__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(AI_5_bF$buf0),
    .Y(_741_)
);

AOI21X1 _1308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_349_),
    .C(_412_),
    .Y(_413_)
);

FILL FILL_3__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_583_),
    .Y(_584_)
);

INVX4 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .Y(_167_)
);

FILL FILL_2__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .Y(_638_)
);

NOR2X1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_113_),
    .Y(_223_)
);

FILL FILL_3__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_394_),
    .C(_393_),
    .Y(_395_)
);

FILL FILL_2__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .B(_766_),
    .Y(_777_)
);

NAND3X1 _1346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_441_),
    .C(_444_),
    .Y(_451_)
);

FILL FILL_1__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_674_),
    .Y(_675_)
);

NAND3X1 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_259_),
    .C(_258_),
    .Y(_261_)
);

FILL FILL_1__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_483_),
    .Y(_488_)
);

FILL FILL_0__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .Y(_299_)
);

FILL FILL_1__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_1_bF$buf3),
    .C(_825_),
    .Y(_856_)
);

OAI21X1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_354_),
    .C(_352_),
    .Y(_355_)
);

FILL FILL_0__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(_579_),
    .C(ABCmd_i[7]),
    .Y(_581_)
);

NAND3X1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_158_),
    .C(_156_),
    .Y(_164_)
);

FILL FILL_0__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_262_),
    .C(_391_),
    .Y(_392_)
);

FILL FILL_2__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_201_),
    .C(_199_),
    .Y(_202_)
);

FILL FILL92250x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_708_),
    .C(_39_),
    .Y(_888_[2])
);

FILL FILL_1__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[4]),
    .Y(ACC_o[4])
);

NAND2X1 _1402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_505_),
    .Y(_506_)
);

FILL FILL_1__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1631_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf1),
    .Q(AI[6])
);

NOR2X1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_167_),
    .Y(_317_)
);

NAND2X1 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[2]),
    .Y(_68_)
);

FILL FILL_1__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .Y(_543_)
);

OAI21X1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_94_),
    .C(_91_),
    .Y(_126_)
);

FILL FILL_1__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_723_),
    .C(_732_),
    .Y(_739_)
);

XNOR2X1 _1305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_406_),
    .Y(_410_)
);

FILL FILL_1__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[5]),
    .Y(_635_)
);

AOI22X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_197_),
    .C(_151_),
    .D(_145_),
    .Y(_220_)
);

FILL FILL_1__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[6]),
    .C(_773_),
    .Y(_774_)
);

AOI21X1 _1343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_447_),
    .C(_411_),
    .Y(_448_)
);

FILL FILL_1__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[1]),
    .Y(ACC_o[1])
);

FILL FILL_3__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_670_),
    .C(_671_),
    .Y(_672_)
);

AOI21X1 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

FILL FILL_1__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1628_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(AI[3])
);

OAI21X1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_231_),
    .C(_217_),
    .Y(_314_)
);

FILL FILL_0__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[1]),
    .Y(_65_)
);

OR2X2 _1381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_482_),
    .Y(_485_)
);

FILL FILL_2__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_715_),
    .C(_387_),
    .Y(_540_)
);

AOI21X1 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_117_),
    .C(_88_),
    .Y(_123_)
);

FILL FILL_3__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_295_),
    .C(_291_),
    .Y(_296_)
);

FILL FILL_1__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(_852_),
    .Y(_853_)
);

OAI21X1 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_191_),
    .C(_210_),
    .Y(_352_)
);

FILL FILL_0__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_94_),
    .C(_91_),
    .Y(_103_)
);

FILL FILL_0__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_577_),
    .C(_525_),
    .Y(_578_)
);

NAND3X1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_159_),
    .C(_158_),
    .Y(_161_)
);

FILL FILL_0__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_245_),
    .C(_242_),
    .Y(_389_)
);

FILL FILL_0__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_198_),
    .Y(_199_)
);

FILL FILL_2__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(_663_),
    .C(_660_),
    .Y(_669_)
);

AOI21X1 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_253_),
    .C(_252_),
    .Y(_255_)
);

FILL FILL_0__897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_796_),
    .C(_798_),
    .Y(_806_)
);

NOR2X1 _1378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(_167_),
    .Y(_482_)
);

FILL FILL_0__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_33_),
    .C(_706_),
    .D(_34_),
    .Y(_37_)
);

FILL FILL_1__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(BI_1_bF$buf3),
    .Y(_293_)
);

FILL FILL_1__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_722_),
    .C(_861_),
    .Y(_736_)
);

NAND2X1 _1302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_3_bF$buf2),
    .B(AI[4]),
    .Y(_407_)
);

FILL FILL_1__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_631_),
    .C(_632_),
    .Y(_633_)
);

NAND3X1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_214_),
    .C(_216_),
    .Y(_217_)
);

FILL FILL_1__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_33_),
    .B(_32__bF$buf1),
    .C(_705__bF$buf0),
    .D(_34_),
    .Y(_35_)
);

FILL FILL_1__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_768_),
    .C(_835_),
    .Y(_771_)
);

AOI21X1 _1340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_440_),
    .C(_438_),
    .Y(_445_)
);

FILL FILL_1__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_820_),
    .C(CO),
    .Y(_823_)
);

FILL FILL_1__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1625_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf1),
    .Q(AI[0])
);

OAI21X1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_310_),
    .C(_247_),
    .Y(_311_)
);

FILL FILL_0__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf1),
    .B(AI[2]),
    .Y(_62_)
);

FILL FILL_1__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_537_),
    .C(_469_),
    .Y(_11_)
);

NAND2X1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_115_),
    .Y(_120_)
);

FILL FILL_1__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(BI_1_bF$buf3),
    .C(_831_),
    .Y(_850_)
);

NAND2X1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_339_),
    .Y(_349_)
);

FILL FILL_0__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_99_),
    .C(_89_),
    .Y(_100_)
);

FILL FILL_0__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_733_),
    .Y(ACC[3])
);

FILL FILL_3__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(_574_),
    .C(_516_),
    .Y(_575_)
);

NAND3X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_141_),
    .C(_140_),
    .Y(_158_)
);

FILL FILL_0__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_282_),
    .C(_301_),
    .Y(_630_)
);

OAI21X1 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_139_),
    .C(_159_),
    .Y(_214_)
);

INVX1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .Y(_386_)
);

FILL FILL_2__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(BI[6]),
    .Y(_768_)
);

NAND3X1 _1337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_437_),
    .C(_404_),
    .Y(_442_)
);

FILL FILL_3__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .Y(_196_)
);

FILL FILL_2__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_644_),
    .C(_665_),
    .Y(_666_)
);

AOI21X1 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_251_),
    .C(_249_),
    .Y(_252_)
);

FILL FILL_0__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705__bF$buf0),
    .Y(_706_)
);

FILL FILL_0__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_777_),
    .C(_785_),
    .Y(_804_)
);

AOI21X1 _1375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(_440_),
    .C(_433_),
    .Y(_479_)
);

FILL FILL_0__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .Y(_290_)
);

FILL FILL_1__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91350x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_571_),
    .B(_568_),
    .Y(_572_)
);

NAND3X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_153_),
    .C(_154_),
    .Y(_155_)
);

FILL FILL_0__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_880_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

NAND2X1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_383_),
    .Y(_384_)
);

FILL FILL_0__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_193_)
);

FILL FILL_2__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__912_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_707_),
    .Y(_32_)
);

FILL FILL_1__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_819_),
    .C(_807_),
    .Y(_820_)
);

FILL FILL_1__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1622_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(_886_[5])
);

INVX1 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .Y(_308_)
);

FILL FILL_0__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_58_),
    .Y(_59_)
);

FILL FILL_1__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91650x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(ACC[2]),
    .Y(_535_)
);

NAND3X1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_104_),
    .C(_116_),
    .Y(_117_)
);

FILL FILL_1__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_841_),
    .Y(_847_)
);

NAND3X1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_338_),
    .C(_342_),
    .Y(_346_)
);

NAND2X1 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf2),
    .B(AI_5_bF$buf1),
    .Y(_97_)
);

FILL FILL92250x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf0),
    .B(BI_3_bF$buf0),
    .C(_730_),
    .Y(_731_)
);

FILL FILL_1__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(CO),
    .Y(_627_)
);

NAND2X1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_205_),
    .Y(_211_)
);

FILL FILL_1__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .Y(ACC[5])
);

NAND3X1 _1334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_439_)
);

FILL FILL_1__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .Y(_663_)
);

NOR2X1 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_63_),
    .Y(_249_)
);

FILL FILL_0__891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .Y(_703_)
);

FILL FILL_0__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1619_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(_886_[2])
);

FILL FILL_0__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[0]),
    .B(_737_),
    .Y(_801_)
);

NAND2X1 _1372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_409_),
    .Y(_476_)
);

FILL FILL_0__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_715_),
    .Y(_532_)
);

OAI21X1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_113_),
    .C(_107_),
    .Y(_114_)
);

NOR3X1 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_265_),
    .C(_286_),
    .Y(_287_)
);

FILL FILL_1__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_843_),
    .C(_841_),
    .Y(_845_)
);

OAI21X1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_185_),
    .C(_182_),
    .Y(_343_)
);

FILL FILL_0__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[3]),
    .Y(_94_)
);

FILL FILL_1__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_562_),
    .C(_565_),
    .Y(_569_)
);

NAND3X1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_145_),
    .C(_148_),
    .Y(_152_)
);

FILL FILL_3__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .Y(_881_)
);

AOI21X1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf3),
    .B(AI[0]),
    .C(_54_),
    .Y(_381_)
);

FILL FILL_0__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_189_),
    .C(_185_),
    .Y(_190_)
);

FILL FILL_0__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .Y(_799_)
);

NAND3X1 _1369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_472_),
    .C(_311_),
    .Y(_473_)
);

FILL FILL_0__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_710_),
    .Y(_888_[0])
);

FILL FILL_1__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_705__bF$buf1),
    .C(_693_),
    .Y(_19_)
);

OAI21X1 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_123_),
    .C(_61_),
    .Y(_284_)
);

FILL FILL_2__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_767_),
    .Y(_817_)
);

FILL FILL_1__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[0]),
    .Y(_56_)
);

FILL FILL_1__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_725_),
    .C(_835_),
    .Y(_728_)
);

FILL FILL_1__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_526_),
    .C(_623_),
    .Y(_624_)
);

AOI21X1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_134_),
    .C(_136_),
    .Y(_208_)
);

FILL FILL_3__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_887_),
    .C(_26_),
    .Y(_27_)
);

OAI21X1 _1751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_761_),
    .C(_762_),
    .Y(_763_)
);

AOI21X1 _1331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_436_)
);

FILL FILL_1__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_808_),
    .C(_814_),
    .Y(CO)
);

FILL FILL_3__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_659_),
    .C(_624_),
    .Y(_660_)
);

AOI21X1 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_242_),
    .B(_245_),
    .C(_176_),
    .Y(_246_)
);

FILL FILL_1__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_700_),
    .Y(_701_)
);

FILL FILL_0__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1616_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(BI[7])
);

FILL FILL_0__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .Y(_54_)
);

FILL FILL_1__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_527_),
    .Y(_529_)
);

NAND3X1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(_106_),
    .C(_108_),
    .Y(_111_)
);

FILL FILL_1__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf0),
    .B(ABCmd_i_2_bF$buf2),
    .C(_825_),
    .Y(_842_)
);

NAND2X1 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[6]),
    .Y(_340_)
);

FILL FILL_0__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_1_bF$buf2),
    .B(AI[4]),
    .C(_90_),
    .Y(_91_)
);

FILL FILL_1__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91950x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .Y(_566_)
);

INVX2 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .Y(_149_)
);

FILL FILL_0__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_573_),
    .B(_618_),
    .Y(_621_)
);

FILL FILL_3__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(AI[3]),
    .Y(_878_)
);

NOR2X1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(HC),
    .Y(_378_)
);

FILL FILL_0__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[5]),
    .C(_825_),
    .Y(_760_)
);

NOR2X1 _1328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(_413_),
    .Y(_433_)
);

FILL FILL_3__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_186_),
    .C(_182_),
    .Y(_187_)
);

FILL FILL_0__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_[6]),
    .Y(_657_)
);

NAND3X1 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_239_),
    .C(_238_),
    .Y(_243_)
);

FILL FILL_1__919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_794_),
    .C(_795_),
    .Y(_796_)
);

AOI21X1 _1366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_470_)
);

FILL FILL_3__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_705__bF$buf3),
    .Y(_692_)
);

NAND3X1 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_279_),
    .C(_280_),
    .Y(_281_)
);

FILL FILL_1__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .Y(ACC[1])
);

NAND3X1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_374_),
    .C(_372_),
    .Y(_375_)
);

FILL FILL_0__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_558_),
    .C(_599_),
    .Y(_600_)
);

INVX1 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .Y(_184_)
);

FILL FILL_2__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(BI_3_bF$buf0),
    .Y(_725_)
);

FILL FILL_1__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL93150x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__903_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_712_),
    .Y(_715_)
);

FILL FILL_1__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_776_),
    .Y(_812_)
);

FILL FILL_1__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92850x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1613_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf3),
    .Q(BI[4])
);

FILL FILL_0__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .Y(_52_)
);

FILL FILL_1__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_472_),
    .Y(_526_)
);

NAND2X1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_107_),
    .Y(_108_)
);

FILL FILL_3__894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_838_),
    .Y(_839_)
);

NAND3X1 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_336_),
    .C(_334_),
    .Y(_337_)
);

OAI21X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_87_),
    .C(_80_),
    .Y(_88_)
);

FILL FILL_1__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .Y(_722_)
);

FILL FILL_3__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_554_),
    .C(_552_),
    .Y(_563_)
);

AND2X2 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf0),
    .B(AI[2]),
    .Y(_146_)
);

FILL FILL_0__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(_523_),
    .Y(_618_)
);

FILL FILL_3__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI[5]),
    .C(_756_),
    .D(_830_),
    .Y(_757_)
);

NOR2X1 _1325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_127_),
    .Y(_430_)
);

FILL FILL_1__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_654_),
    .C(state[1]),
    .Y(_655_)
);

NAND3X1 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_213_),
    .C(_217_),
    .Y(_240_)
);

FILL FILL_1__916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[7]),
    .C(_825_),
    .Y(_793_)
);

AOI21X1 _1363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(_703_),
    .C(_712_),
    .Y(_468_)
);

FILL FILL_0__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_518_),
    .C(_522_),
    .Y(_523_)
);

FILL FILL92850x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_712_),
    .C(_685_),
    .D(_690_),
    .Y(_16_)
);

AOI21X1 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_276_),
    .C(_275_),
    .Y(_278_)
);

FILL FILL_1__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf1),
    .Y(_836_)
);

NAND2X1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_330_),
    .Y(_334_)
);

FILL FILL_0__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_83_),
    .C(_84_),
    .Y(_85_)
);

FILL FILL_0__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_559_),
    .Y(_560_)
);

AOI21X1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_142_),
    .C(_140_),
    .Y(_143_)
);

FILL FILL_1__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_857_),
    .C(_872_),
    .Y(_873_)
);

OAI21X1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_237_),
    .C(_244_),
    .Y(_372_)
);

FILL FILL_0__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .Y(_597_)
);

OAI21X1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_133_),
    .C(_128_),
    .Y(_181_)
);

FILL FILL93150x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__900_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .Y(_712_)
);

FILL FILL_1__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_54_),
    .Y(_688_)
);

OAI21X1 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(_275_)
);

FILL FILL_2__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .B(_804_),
    .Y(_809_)
);

FILL FILL_1__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_501_),
    .C(_490_),
    .Y(_502_)
);

FILL FILL_0__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1610_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(BI[1])
);

INVX1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .Y(_50_)
);

FILL FILL_1__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .Y(ACC[2])
);

FILL FILL_1__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_460_),
    .Y(_615_)
);

FILL FILL_1__1675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(AI[6]),
    .Y(_754_)
);

OAI22X1 _1322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_414_),
    .C(_422_),
    .D(_426_),
    .Y(_427_)
);

FILL FILL_1__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_652_)
);

AOI21X1 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_230_),
    .C(_179_),
    .Y(_237_)
);

FILL FILL_1__913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL92550x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU.AI7 ),
    .B(_705__bF$buf0),
    .Y(_698_)
);

FILL FILL_0__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[4]),
    .Y(_48_)
);

FILL FILL_1__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(BI[7]),
    .C(_789_),
    .D(_830_),
    .Y(_790_)
);

NAND2X1 _1360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[1]),
    .B(_54_),
    .Y(_465_)
);

FILL FILL_0__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_457_),
    .C(_519_),
    .Y(_520_)
);

FILL FILL_3__1660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(ABCmd_i[1]),
    .Y(_833_)
);

OAI21X1 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_74_),
    .C(_330_),
    .Y(_331_)
);

FILL FILL_0__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf0),
    .B(AI[1]),
    .Y(_82_)
);

FILL FILL_1__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_556_),
    .Y(_557_)
);

AOI21X1 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_95_),
    .C(_98_),
    .Y(_140_)
);

FILL FILL_1__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_863_),
    .C(_869_),
    .Y(_870_)
);

OAI21X1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_364_),
    .C(_314_),
    .Y(_369_)
);

FILL FILL_0__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_751_),
    .Y(ACC[4])
);

OAI21X1 _1319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_58_),
    .C(_417_),
    .Y(_424_)
);

OAI21X1 _1492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_167_),
    .C(_557_),
    .Y(_594_)
);

INVX1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .Y(_178_)
);

FILL FILL_0__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .B(_637_),
    .C(_648_),
    .Y(_649_)
);

NAND3X1 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_224_),
    .C(_222_),
    .Y(_234_)
);

FILL FILL_3__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(ABCmd_i[4]),
    .Y(_787_)
);

OAI21X1 _1357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_398_),
    .C(ABCmd_i[7]),
    .Y(_462_)
);

FILL FILL_3__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL91350x150 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_708_),
    .Y(_709_)
);

FILL FILL_1__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_682_),
    .C(_636_),
    .Y(_685_)
);

OR2X2 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_271_),
    .Y(_272_)
);

FILL FILL_1__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

AOI21X1 _1395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_499_)
);

FILL FILL_0__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .Y(_591_)
);

OAI21X1 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(_173_),
    .C(_170_),
    .Y(_175_)
);

FILL FILL_2__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_716_),
    .C(_884_),
    .Y(_717_)
);

FILL FILL_1__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_403_)
);

FILL FILL_2__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_571_),
    .Y(_612_)
);

FILL FILL_3__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_705__bF$buf2),
    .C(_696_),
    .Y(_22_)
);

FILL FILL_0__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[3]),
    .Y(_46_)
);

FILL FILL_1__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_513_),
    .C(_479_),
    .Y(_517_)
);

FILL FILL_1__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(_829_),
    .Y(_830_)
);

AND2X2 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_4_bF$buf2),
    .B(AI[4]),
    .Y(_328_)
);

FILL FILL_0__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_78_),
    .C(_68_),
    .Y(_79_)
);

FILL FILL_1__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_553_),
    .C(_545_),
    .Y(_554_)
);

AOI22X1 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI_0_bF$buf2),
    .B(AI[6]),
    .C(BI_1_bF$buf0),
    .D(AI_5_bF$buf1),
    .Y(_137_)
);

FILL FILL_1__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_605_),
    .C(_608_),
    .Y(_609_)
);

FILL FILL_1__1669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .B(_865_),
    .Y(_867_)
);

AOI21X1 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_365_),
    .C(_313_),
    .Y(_366_)
);

FILL FILL_0__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_748_),
    .C(_746_),
    .Y(_749_)
);

INVX1 _1316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .Y(_421_)
);

FILL FILL_3__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _1545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_640_),
    .Y(_646_)
);

AOI21X1 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_215_),
    .C(_214_),
    .Y(_231_)
);

FILL FILL_1__907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_783_),
    .Y(_785_)
);

NAND3X1 _1354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_459_)
);

FILL FILL_1__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_663_),
    .C(_668_),
    .Y(_682_)
);

NAND3X1 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .C(_80_),
    .Y(_269_)
);

FILL FILL_1__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(_826_),
    .Y(_827_)
);

NAND2X1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_321_),
    .Y(_325_)
);

FILL FILL_0__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_496_)
);

FILL FILL_0__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .Y(_551_)
);

INVX1 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .Y(_134_)
);

FILL FILL_3__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule
