* NGSPICE file created from ALU_wrapper.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR D S R CLK Q vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

.subckt ALU_wrapper gnd vdd ABCmd_i[7] ABCmd_i[6] ABCmd_i[5] ABCmd_i[4] ABCmd_i[3]
+ ABCmd_i[2] ABCmd_i[1] ABCmd_i[0] ACC_o[7] ACC_o[6] ACC_o[5] ACC_o[4] ACC_o[3] ACC_o[2]
+ ACC_o[1] ACC_o[0] Done_o LoadA_i LoadB_i LoadCmd_i clk reset
XFILL_1__1670_ vdd gnd FILL
XFILL_0__1759_ vdd gnd FILL
XFILL_3__1606_ vdd gnd FILL
XFILL_3__1468_ vdd gnd FILL
XFILL_3__1537_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL_3__1399_ vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_1__1799_ vdd gnd FILL
XFILL92250x150 vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL_2__1144_ vdd gnd FILL
XFILL_2__1075_ vdd gnd FILL
XFILL_3__957_ vdd gnd FILL
X_1270_ _1292_/B _1370_/A _1422_/A vdd gnd AND2X2
XFILL_0__1544_ vdd gnd FILL
XFILL_3__1322_ vdd gnd FILL
XFILL_3__1253_ vdd gnd FILL
XFILL_0__1475_ vdd gnd FILL
X_1606_ _946_/A _1606_/B _1606_/C _1631_/D vdd gnd OAI21X1
XFILL93150x89850 vdd gnd FILL
XFILL_1__1722_ vdd gnd FILL
XFILL_1__1653_ vdd gnd FILL
X_1468_ _1468_/A _1510_/A _1468_/C _1510_/B vdd gnd NAND3X1
X_1537_ _1558_/A _1561_/A vdd gnd INVX1
X_1399_ _1406_/A _1406_/B _1441_/A vdd gnd AND2X2
XFILL_1__1584_ vdd gnd FILL
XFILL_2__975_ vdd gnd FILL
X_981_ _981_/A _981_/B _981_/C _982_/B vdd gnd AOI21X1
XFILL_2__1762_ vdd gnd FILL
XFILL_1__1018_ vdd gnd FILL
XFILL_2__1693_ vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
XFILL_2__1058_ vdd gnd FILL
XFILL_2__1127_ vdd gnd FILL
XFILL_1__993_ vdd gnd FILL
X_1253_ _1338_/A _1342_/B _1338_/C _1339_/B vdd gnd OAI21X1
X_1322_ _1325_/B _1325_/A _1322_/C _1322_/D _1341_/A vdd gnd OAI22X1
X_1184_ _1184_/A _1185_/C vdd gnd INVX1
XFILL_0__1527_ vdd gnd FILL
XFILL_3__1305_ vdd gnd FILL
XFILL_3__1236_ vdd gnd FILL
XFILL_3__1167_ vdd gnd FILL
XFILL_3__1098_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_0__1458_ vdd gnd FILL
XFILL_1__1636_ vdd gnd FILL
XFILL_1__1705_ vdd gnd FILL
XFILL_1__1567_ vdd gnd FILL
XFILL_1__1498_ vdd gnd FILL
XFILL_2__958_ vdd gnd FILL
XFILL_2__889_ vdd gnd FILL
XFILL_2__1814_ vdd gnd FILL
XFILL_2__1745_ vdd gnd FILL
X_964_ _964_/A _988_/B _972_/A vdd gnd NAND2X1
X_895_ _898_/A _899_/A _896_/B vdd gnd NOR2X1
XFILL_2__1676_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
XFILL_0__1312_ vdd gnd FILL
XFILL_0__1243_ vdd gnd FILL
XFILL_1__976_ vdd gnd FILL
X_1305_ _1372_/B _1372_/A _1373_/B vdd gnd XNOR2X1
X_1236_ _1329_/B _1307_/B _1248_/A vdd gnd NAND2X1
X_1167_ _999_/A _988_/A _1186_/B vdd gnd NAND2X1
XBUFX2_insert0 _1612_/Q _952_/A vdd gnd BUFX2
X_1098_ _979_/B _1301_/A _1098_/C _1099_/C vdd gnd OAI21X1
XFILL_1__1283_ vdd gnd FILL
XFILL_3__1219_ vdd gnd FILL
XFILL_1__1352_ vdd gnd FILL
XFILL_1__1421_ vdd gnd FILL
XFILL_2__1530_ vdd gnd FILL
XFILL_2__1461_ vdd gnd FILL
XFILL_2__1392_ vdd gnd FILL
XFILL_3_CLKBUF1_insert12 vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
XFILL_2__1659_ vdd gnd FILL
XFILL_0__1792_ vdd gnd FILL
XFILL_2__1728_ vdd gnd FILL
X_947_ ABCmd_i[7] _949_/A vdd gnd INVX4
X_1021_ _1082_/A _1760_/A _1325_/B vdd gnd AND2X2
X_1785_ _1809_/B _1809_/C _1809_/A _1803_/C vdd gnd OAI21X1
XFILL_0__1157_ vdd gnd FILL
XFILL_3__1004_ vdd gnd FILL
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
XFILL_1__959_ vdd gnd FILL
X_1219_ _1257_/B _1257_/A _1299_/A vdd gnd NAND2X1
XFILL_1__1404_ vdd gnd FILL
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL92250x70350 vdd gnd FILL
XFILL_3__990_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
XFILL_2__1513_ vdd gnd FILL
XFILL_2__1375_ vdd gnd FILL
XFILL_2__1444_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
X_1570_ _1570_/A _1570_/B _1570_/C _1572_/B vdd gnd AOI21X1
XFILL_0__1775_ vdd gnd FILL
X_1004_ _953_/B _1211_/A _980_/A _1005_/A vdd gnd OAI21X1
XFILL_1__1120_ vdd gnd FILL
X_1768_ _1768_/A _1768_/B _1768_/C _1769_/A vdd gnd AOI21X1
XFILL_1__1051_ vdd gnd FILL
XFILL_0__1209_ vdd gnd FILL
X_1699_ _1716_/A _988_/A _1783_/C _1700_/C vdd gnd OAI21X1
XFILL_2__1160_ vdd gnd FILL
XFILL92250x82050 vdd gnd FILL
XFILL_0__900_ vdd gnd FILL
XFILL_2__1091_ vdd gnd FILL
XFILL_1__1318_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_3__973_ vdd gnd FILL
XFILL_0__1560_ vdd gnd FILL
XFILL_2__1427_ vdd gnd FILL
XFILL_2__1289_ vdd gnd FILL
XFILL_2__1358_ vdd gnd FILL
XFILL_0__1491_ vdd gnd FILL
X_1622_ _1622_/D vdd _1624_/R _1624_/CLK _1823_/A vdd gnd DFFSR
XFILL_2_BUFX2_insert36 vdd gnd FILL
X_1484_ _949_/A _1484_/B _1484_/C _1485_/A vdd gnd OAI21X1
X_1553_ _1754_/Y _1554_/B vdd gnd INVX1
XFILL_2_BUFX2_insert25 vdd gnd FILL
XFILL_2_BUFX2_insert14 vdd gnd FILL
XFILL_0__1758_ vdd gnd FILL
XFILL_0__1689_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_2__991_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_1__1798_ vdd gnd FILL
XFILL_1_BUFX2_insert0 vdd gnd FILL
XFILL_2__1143_ vdd gnd FILL
XFILL_2__1212_ vdd gnd FILL
XFILL_2__1074_ vdd gnd FILL
XFILL_0__1543_ vdd gnd FILL
XFILL_3__1183_ vdd gnd FILL
XFILL_0__1474_ vdd gnd FILL
X_1605_ _1760_/A _1606_/B _1606_/C vdd gnd NAND2X1
X_1536_ _1560_/A _1560_/C _1548_/B vdd gnd NAND2X1
XFILL_1__1721_ vdd gnd FILL
XFILL_1__1652_ vdd gnd FILL
X_1398_ _1441_/C _1462_/B _1462_/A _1471_/A vdd gnd OAI21X1
X_1467_ _1467_/A _1467_/B _1467_/C _1468_/C vdd gnd OAI21X1
XFILL_1__1583_ vdd gnd FILL
XFILL_2__974_ vdd gnd FILL
XFILL_1__1017_ vdd gnd FILL
XFILL_2__1692_ vdd gnd FILL
XFILL_2__1761_ vdd gnd FILL
X_980_ _980_/A _980_/B _980_/C _982_/A vdd gnd OAI21X1
XFILL_0__1190_ vdd gnd FILL
XFILL_2__1126_ vdd gnd FILL
XFILL_2__1057_ vdd gnd FILL
XFILL_1__992_ vdd gnd FILL
X_1321_ _1323_/B _1323_/C _1379_/A _1322_/D vdd gnd AOI21X1
X_1252_ _1298_/A _1298_/B _1298_/C _1299_/C vdd gnd NAND3X1
X_1183_ _975_/A _1193_/A _1183_/C _1480_/A vdd gnd NAND3X1
XFILL_0__1526_ vdd gnd FILL
XFILL_0__1457_ vdd gnd FILL
XFILL_0__1388_ vdd gnd FILL
X_1519_ _1521_/A _1521_/B _1520_/C vdd gnd NAND2X1
XFILL_1__1704_ vdd gnd FILL
XFILL_1__1566_ vdd gnd FILL
XFILL_2__957_ vdd gnd FILL
XFILL_1__1497_ vdd gnd FILL
X_963_ _983_/A _995_/A vdd gnd INVX1
XFILL_2__1813_ vdd gnd FILL
XFILL_2__1675_ vdd gnd FILL
XFILL_2__1744_ vdd gnd FILL
X_894_ _915_/A _899_/A vdd gnd INVX2
XFILL_3__1020_ vdd gnd FILL
XFILL_0__1311_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
XFILL_0__1242_ vdd gnd FILL
XFILL_2__1109_ vdd gnd FILL
XFILL_3__1784_ vdd gnd FILL
X_1166_ _960_/A _1361_/A _1169_/C vdd gnd OR2X2
XFILL_1__975_ vdd gnd FILL
XBUFX2_insert1 _1612_/Q _1302_/A vdd gnd BUFX2
XFILL_1__1420_ vdd gnd FILL
X_1235_ _1387_/A _1387_/B _1329_/B vdd gnd XOR2X1
X_1304_ _1304_/A _1304_/B _1304_/C _1304_/D _1372_/B vdd gnd OAI22X1
XFILL_1__1282_ vdd gnd FILL
X_1097_ _953_/B _969_/B _1114_/B _1099_/B vdd gnd OAI21X1
XFILL_1__1351_ vdd gnd FILL
XFILL_0__1509_ vdd gnd FILL
XFILL_2__1391_ vdd gnd FILL
XFILL_2__1460_ vdd gnd FILL
XFILL_1__1549_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
XFILL_2__1658_ vdd gnd FILL
XFILL_0__1791_ vdd gnd FILL
XFILL_2__1727_ vdd gnd FILL
X_1020_ _996_/A _997_/B _997_/C _1053_/A vdd gnd OAI21X1
X_946_ _946_/A _946_/B _946_/C _946_/Y vdd gnd OAI21X1
XFILL_2__1589_ vdd gnd FILL
X_1784_ _1784_/A _948_/A _1784_/C _1809_/C vdd gnd AOI21X1
XFILL_0__1156_ vdd gnd FILL
XFILL_0__1087_ vdd gnd FILL
XFILL_0__1225_ vdd gnd FILL
XFILL_3__1767_ vdd gnd FILL
XFILL_1__958_ vdd gnd FILL
X_1149_ _1151_/C _1151_/B _1151_/A _1174_/A vdd gnd AOI21X1
XFILL_3__1698_ vdd gnd FILL
XFILL_1__889_ vdd gnd FILL
X_1218_ _1296_/B _1218_/B _1296_/A _1257_/B vdd gnd OAI21X1
XFILL_1__1403_ vdd gnd FILL
XFILL_1__1196_ vdd gnd FILL
XFILL92550x54750 vdd gnd FILL
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
XFILL92250x89850 vdd gnd FILL
XFILL_2__1512_ vdd gnd FILL
XFILL_2__1374_ vdd gnd FILL
XFILL_2__1443_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_3__1552_ vdd gnd FILL
XFILL_0__1774_ vdd gnd FILL
X_929_ ABCmd_i[1] _931_/A vdd gnd INVX1
XFILL_3__1483_ vdd gnd FILL
X_1003_ _962_/B _1211_/A vdd gnd INVX1
XFILL_1__1050_ vdd gnd FILL
X_1698_ _1698_/A _1698_/B _1698_/C _1708_/A vdd gnd OAI21X1
X_1767_ ABCmd_i[6] _1768_/C vdd gnd INVX1
XFILL_0__1208_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
XFILL_3__1819_ vdd gnd FILL
XFILL92850x31350 vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_2__1090_ vdd gnd FILL
XFILL_0__1490_ vdd gnd FILL
XFILL_2__1426_ vdd gnd FILL
XFILL_2__1288_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_0__959_ vdd gnd FILL
XFILL_2_BUFX2_insert26 vdd gnd FILL
X_1552_ _1552_/A _1576_/C ABCmd_i[7] _1555_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert15 vdd gnd FILL
X_1621_ _1621_/D vdd _1624_/R _1624_/CLK _1822_/A vdd gnd DFFSR
X_1483_ _1769_/B _949_/A _1484_/C vdd gnd NAND2X1
XFILL_3__1604_ vdd gnd FILL
XFILL_2_BUFX2_insert37 vdd gnd FILL
XFILL_3__1535_ vdd gnd FILL
XFILL_0__1826_ vdd gnd FILL
XFILL_0__1688_ vdd gnd FILL
XFILL_0__1757_ vdd gnd FILL
XFILL_2__990_ vdd gnd FILL
XFILL_3__1397_ vdd gnd FILL
XFILL_3__1466_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
X_1819_ _1819_/A ACC_o[1] vdd gnd BUFX2
XFILL92550x78150 vdd gnd FILL
XFILL_1__1797_ vdd gnd FILL
XFILL_1_BUFX2_insert1 vdd gnd FILL
XFILL_2__1142_ vdd gnd FILL
XFILL_2__1073_ vdd gnd FILL
XFILL_2__1211_ vdd gnd FILL
XFILL_0_CLKBUF1_insert8 vdd gnd FILL
XFILL_3__955_ vdd gnd FILL
XFILL_0__1473_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
XFILL_0__1542_ vdd gnd FILL
XFILL_1__1720_ vdd gnd FILL
X_1604_ _943_/A _1604_/B _1604_/C _1630_/D vdd gnd OAI21X1
X_1535_ _1535_/A _1586_/C vdd gnd INVX1
XFILL_0__1809_ vdd gnd FILL
XFILL_1__1651_ vdd gnd FILL
X_1397_ _1441_/B _1462_/B vdd gnd INVX1
X_1466_ _1506_/B _1466_/B _1466_/C _1510_/A vdd gnd NAND3X1
XFILL_3__1518_ vdd gnd FILL
XFILL_1__1582_ vdd gnd FILL
XFILL_2__973_ vdd gnd FILL
XFILL_3__1449_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_2__1691_ vdd gnd FILL
XFILL_2__1760_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
XFILL_2__1125_ vdd gnd FILL
X_1320_ _1496_/A _979_/B _1320_/C _1323_/C vdd gnd OAI21X1
X_1182_ _1194_/A _1183_/C vdd gnd INVX1
XFILL_3__938_ vdd gnd FILL
XFILL_1__991_ vdd gnd FILL
X_1251_ _1257_/A _1257_/B _1339_/A vdd gnd AND2X2
XFILL_3__1165_ vdd gnd FILL
XFILL_0__1525_ vdd gnd FILL
XFILL_3__1234_ vdd gnd FILL
XFILL_0__1456_ vdd gnd FILL
XFILL_3__1303_ vdd gnd FILL
XFILL_3__1096_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
XFILL_1__1703_ vdd gnd FILL
X_1518_ _1570_/A _1570_/B _1548_/A _1549_/B vdd gnd AOI21X1
X_1449_ _1449_/A _1488_/C _1449_/C _1460_/C vdd gnd NAND3X1
XFILL_1__1565_ vdd gnd FILL
XFILL_1__1496_ vdd gnd FILL
XFILL_2__956_ vdd gnd FILL
XFILL_2__1812_ vdd gnd FILL
XFILL_2__1674_ vdd gnd FILL
X_962_ _988_/A _962_/B _983_/A vdd gnd NAND2X1
XFILL_2__1743_ vdd gnd FILL
X_893_ _904_/B _898_/B vdd gnd INVX1
XFILL_0__1241_ vdd gnd FILL
XFILL_0__1310_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
XFILL_2__1108_ vdd gnd FILL
XFILL_2__1039_ vdd gnd FILL
XFILL_1__974_ vdd gnd FILL
X_1303_ _1303_/A _977_/A _1304_/B vdd gnd NAND2X1
X_1165_ _986_/A _978_/B _1361_/A vdd gnd NAND2X1
XBUFX2_insert2 _1612_/Q _978_/A vdd gnd BUFX2
X_1234_ _988_/A _1760_/A _1387_/B vdd gnd NAND2X1
X_1096_ _1096_/A _1096_/B _1212_/C _1105_/A vdd gnd NAND3X1
XFILL_1__1350_ vdd gnd FILL
XFILL_3__1148_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_3__1217_ vdd gnd FILL
XFILL_0__1508_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_3__1079_ vdd gnd FILL
XFILL_2__1390_ vdd gnd FILL
XFILL_1__1548_ vdd gnd FILL
XFILL_1__1479_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
XFILL_2__939_ vdd gnd FILL
X_945_ _945_/A _946_/B _946_/C vdd gnd NAND2X1
XFILL_2__1657_ vdd gnd FILL
XFILL_0__1790_ vdd gnd FILL
XFILL_2__1726_ vdd gnd FILL
XFILL_2__1588_ vdd gnd FILL
XFILL_0__1224_ vdd gnd FILL
X_1783_ _1784_/A _948_/A _1783_/C _1784_/C vdd gnd OAI21X1
XFILL_0__1155_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
XFILL_1__957_ vdd gnd FILL
X_1148_ _983_/A _995_/B _983_/C _1151_/C vdd gnd NAND3X1
X_1079_ _988_/A _1303_/A _1237_/B vdd gnd NAND2X1
X_1217_ _1217_/A _1217_/B _1296_/B vdd gnd NOR2X1
XFILL_1__1402_ vdd gnd FILL
XFILL_1__1333_ vdd gnd FILL
XFILL_1__1195_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_2__1511_ vdd gnd FILL
XFILL_2__1442_ vdd gnd FILL
XFILL_2__1373_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
XFILL_0__1773_ vdd gnd FILL
X_928_ _928_/A _943_/B _928_/C _928_/Y vdd gnd OAI21X1
XFILL_2__1709_ vdd gnd FILL
X_1002_ _955_/A _1114_/A _1005_/C vdd gnd NAND2X1
XFILL_0__1207_ vdd gnd FILL
X_1697_ _962_/B _1697_/B _1802_/B _1698_/B vdd gnd OAI21X1
X_1766_ _1804_/B _1805_/A _1795_/B vdd gnd NAND2X1
XFILL_0__1069_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_1__1316_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_3__971_ vdd gnd FILL
XFILL_2__1425_ vdd gnd FILL
XFILL_2__1356_ vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
XFILL_2__1287_ vdd gnd FILL
XFILL_2_BUFX2_insert38 vdd gnd FILL
X_1551_ _1551_/A _1551_/B _1551_/C _1552_/A vdd gnd AOI21X1
X_1482_ _1528_/C _1482_/B _1484_/B vdd gnd NAND2X1
XFILL_2_BUFX2_insert27 vdd gnd FILL
XFILL_2_BUFX2_insert16 vdd gnd FILL
XFILL_0__889_ vdd gnd FILL
X_1620_ _1620_/D vdd _1624_/R _1624_/CLK _1821_/A vdd gnd DFFSR
XFILL_0__1756_ vdd gnd FILL
XFILL_0__1825_ vdd gnd FILL
XFILL_0__1687_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_1__1032_ vdd gnd FILL
X_1818_ _950_/A ACC_o[0] vdd gnd BUFX2
X_1749_ _932_/A _999_/B _1749_/C _1771_/A vdd gnd AOI21X1
XFILL_1__1796_ vdd gnd FILL
XFILL_1_BUFX2_insert2 vdd gnd FILL
XFILL_2__1210_ vdd gnd FILL
XFILL_2__1072_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_0_CLKBUF1_insert9 vdd gnd FILL
XFILL_3__1181_ vdd gnd FILL
XFILL_2__1339_ vdd gnd FILL
XFILL_0__1472_ vdd gnd FILL
XFILL_3__1250_ vdd gnd FILL
XFILL_2__1408_ vdd gnd FILL
XFILL_0__1541_ vdd gnd FILL
X_1603_ _1746_/A _1604_/B _1604_/C vdd gnd NAND2X1
X_1465_ _1465_/A _1465_/B _1465_/C _1473_/A vdd gnd NAND3X1
X_1534_ _1823_/A _1556_/A vdd gnd INVX1
XFILL_1__1650_ vdd gnd FILL
XFILL_0__1808_ vdd gnd FILL
XFILL_0__1739_ vdd gnd FILL
X_1396_ _1400_/A _1400_/B _1408_/A _1441_/B vdd gnd NAND3X1
XFILL_1__1581_ vdd gnd FILL
XFILL_2__972_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_2__1690_ vdd gnd FILL
XFILL_1__1779_ vdd gnd FILL
XFILL91650x54750 vdd gnd FILL
XFILL_2__1055_ vdd gnd FILL
XFILL_2__1124_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
X_1181_ _1551_/A _1203_/A _1203_/B _1204_/C vdd gnd NOR3X1
X_1250_ _1299_/A _1258_/B _1258_/A _1350_/A vdd gnd NAND3X1
XFILL_0__1524_ vdd gnd FILL
XFILL_0__1455_ vdd gnd FILL
XFILL_0__1386_ vdd gnd FILL
XFILL_1__1702_ vdd gnd FILL
X_1448_ _1488_/B _1449_/C vdd gnd INVX1
X_1517_ _1521_/A _1521_/B _1517_/C _1521_/C _1570_/A vdd gnd AOI22X1
XFILL_1__1564_ vdd gnd FILL
XFILL_1__1495_ vdd gnd FILL
X_1379_ _1379_/A _1379_/B _1379_/C _1384_/B vdd gnd OAI21X1
XFILL_2__955_ vdd gnd FILL
X_961_ _961_/A _961_/B _961_/C _981_/C vdd gnd OAI21X1
XFILL_2__1811_ vdd gnd FILL
XFILL_2__1742_ vdd gnd FILL
XFILL_2__1673_ vdd gnd FILL
X_892_ _892_/A _909_/B vdd gnd INVX1
XFILL_0__1240_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
XFILL_2__1038_ vdd gnd FILL
XFILL_2__1107_ vdd gnd FILL
XFILL_1__973_ vdd gnd FILL
XFILL_3__1782_ vdd gnd FILL
X_1233_ _1233_/A _1233_/B _1233_/C _1307_/B vdd gnd AOI21X1
X_1302_ _1302_/A _986_/D _1304_/A vdd gnd NAND2X1
X_1164_ _1164_/A _1164_/B _961_/C _1172_/A vdd gnd NAND3X1
XBUFX2_insert3 _1612_/Q _1716_/B vdd gnd BUFX2
XFILL_1__1280_ vdd gnd FILL
X_1095_ _1212_/B _1096_/B vdd gnd INVX1
XFILL_0__1507_ vdd gnd FILL
XFILL_0__1438_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_1_BUFX2_insert40 vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_1__1547_ vdd gnd FILL
XFILL_1__1478_ vdd gnd FILL
XFILL_2__938_ vdd gnd FILL
XFILL_2__1725_ vdd gnd FILL
X_944_ ABCmd_i[6] _946_/A vdd gnd INVX1
XFILL_2__1656_ vdd gnd FILL
XFILL_2__1587_ vdd gnd FILL
XFILL_0__1154_ vdd gnd FILL
XFILL_3__1001_ vdd gnd FILL
XFILL_0__1223_ vdd gnd FILL
X_1782_ _1782_/A _1782_/B _1782_/C _1809_/A vdd gnd OAI21X1
XFILL_0__1085_ vdd gnd FILL
XFILL_3__1696_ vdd gnd FILL
XFILL_1__956_ vdd gnd FILL
XFILL_3__1765_ vdd gnd FILL
X_1216_ _1217_/B _1217_/A _1218_/B vdd gnd AND2X2
X_1147_ _995_/C _983_/B _995_/A _1151_/B vdd gnd OAI21X1
XFILL93150x85950 vdd gnd FILL
X_1078_ _1237_/A _1233_/A vdd gnd INVX1
XFILL_1__1401_ vdd gnd FILL
XFILL_1__1332_ vdd gnd FILL
XFILL_1__1263_ vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL_2__1441_ vdd gnd FILL
XFILL_2__1510_ vdd gnd FILL
XFILL_2__1372_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
XFILL_2__1708_ vdd gnd FILL
XFILL_0__1772_ vdd gnd FILL
XFILL_3__1481_ vdd gnd FILL
X_927_ _986_/A _943_/B _928_/C vdd gnd NAND2X1
XFILL_3__1550_ vdd gnd FILL
XFILL_2__1639_ vdd gnd FILL
X_1001_ _978_/A _962_/B _1114_/A vdd gnd AND2X2
XCLKBUF1_insert10 clk _1634_/CLK vdd gnd CLKBUF1
X_1765_ _1765_/A _1765_/B _1803_/A _1804_/B vdd gnd OAI21X1
XFILL_0__1206_ vdd gnd FILL
XFILL_0__1137_ vdd gnd FILL
X_1696_ ABCmd_i[0] _1696_/B _1697_/B vdd gnd NOR2X1
XFILL_3__1817_ vdd gnd FILL
XFILL_3__1748_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
XFILL_3__1679_ vdd gnd FILL
XFILL_1__939_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_1__1315_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_2__1355_ vdd gnd FILL
XFILL_2__1424_ vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
XFILL_2__1286_ vdd gnd FILL
XFILL_2_BUFX2_insert39 vdd gnd FILL
X_1481_ _1481_/A _1481_/B _1482_/B vdd gnd NAND2X1
XFILL_2_BUFX2_insert28 vdd gnd FILL
XFILL_3__1602_ vdd gnd FILL
XFILL_2_BUFX2_insert17 vdd gnd FILL
X_1550_ _1586_/C _1550_/B _1550_/C _1556_/C vdd gnd NAND3X1
XFILL_0__1686_ vdd gnd FILL
XFILL_0__1755_ vdd gnd FILL
XFILL_3__1533_ vdd gnd FILL
XFILL_3__1464_ vdd gnd FILL
XFILL_0__1824_ vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_3__1395_ vdd gnd FILL
X_1817_ _1817_/A _1817_/B _1817_/Y vdd gnd NAND2X1
X_1748_ _932_/A _999_/B _1783_/C _1749_/C vdd gnd OAI21X1
XFILL_1__1031_ vdd gnd FILL
X_1679_ _1679_/A _1679_/B _1680_/A vdd gnd NAND2X1
XFILL_1__1795_ vdd gnd FILL
XFILL_1_BUFX2_insert3 vdd gnd FILL
XFILL_2__1140_ vdd gnd FILL
XFILL_2__1071_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_3__953_ vdd gnd FILL
XFILL_0__1540_ vdd gnd FILL
XFILL_2__1338_ vdd gnd FILL
XFILL_0__1471_ vdd gnd FILL
XFILL_2__1407_ vdd gnd FILL
XFILL_2__1269_ vdd gnd FILL
X_1602_ _940_/A _1604_/B _1602_/C _1629_/D vdd gnd OAI21X1
X_1533_ _1533_/A _911_/A _1533_/C _1533_/D _1621_/D vdd gnd AOI22X1
X_1464_ _1467_/A _1467_/B _1466_/C _1465_/B vdd gnd OAI21X1
X_1395_ _1400_/A _1400_/B _1408_/A _1441_/C vdd gnd AOI21X1
XFILL_0__1669_ vdd gnd FILL
XFILL_0__1807_ vdd gnd FILL
XFILL_0__1738_ vdd gnd FILL
XFILL_1__1580_ vdd gnd FILL
XFILL_3__1516_ vdd gnd FILL
XFILL_3__1447_ vdd gnd FILL
XFILL_3__1378_ vdd gnd FILL
XFILL_2__971_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL_1__1778_ vdd gnd FILL
XFILL_2__1123_ vdd gnd FILL
XFILL_2__1054_ vdd gnd FILL
XFILL_3__936_ vdd gnd FILL
X_1180_ _1286_/B _1286_/A _1180_/C _1203_/B vdd gnd AOI21X1
XFILL_0__1523_ vdd gnd FILL
XFILL_3__1232_ vdd gnd FILL
XFILL_3__1301_ vdd gnd FILL
XFILL_3__1163_ vdd gnd FILL
XFILL_3__1094_ vdd gnd FILL
XFILL_0__1454_ vdd gnd FILL
XFILL_0__1385_ vdd gnd FILL
X_1516_ _1516_/A _1516_/B _1521_/B vdd gnd NAND2X1
XFILL_1__1701_ vdd gnd FILL
X_1447_ _1447_/A _1447_/B _1488_/B vdd gnd NOR2X1
X_1378_ _969_/B _1567_/B _1384_/A vdd gnd NOR2X1
XFILL_1__1563_ vdd gnd FILL
XFILL_1__1494_ vdd gnd FILL
XFILL_2__954_ vdd gnd FILL
X_960_ _960_/A _960_/B _961_/B vdd gnd AND2X2
XFILL_2__1672_ vdd gnd FILL
XFILL_2__1810_ vdd gnd FILL
XFILL_2__1741_ vdd gnd FILL
X_891_ _915_/A _903_/A _892_/A vdd gnd NAND2X1
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1106_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
XFILL_3__919_ vdd gnd FILL
XFILL_1__972_ vdd gnd FILL
X_1232_ _1247_/B _1247_/A _1330_/A vdd gnd NAND2X1
X_1301_ _1301_/A _1567_/B _1372_/A vdd gnd NOR2X1
X_1163_ _1163_/A _1163_/B _982_/C _1196_/B vdd gnd NAND3X1
XBUFX2_insert4 _1609_/Q _986_/A vdd gnd BUFX2
XFILL_0__1437_ vdd gnd FILL
X_1094_ _1302_/A _986_/D _977_/A _988_/B _1212_/B vdd gnd AOI22X1
XFILL_3__1215_ vdd gnd FILL
XFILL_0__1506_ vdd gnd FILL
XFILL_3__1146_ vdd gnd FILL
XFILL_3__1077_ vdd gnd FILL
XFILL_0__1299_ vdd gnd FILL
XFILL_0__1368_ vdd gnd FILL
XFILL_1_BUFX2_insert41 vdd gnd FILL
XFILL_1_BUFX2_insert30 vdd gnd FILL
XFILL_1__1546_ vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_2__937_ vdd gnd FILL
XFILL_1__1477_ vdd gnd FILL
XFILL_2__1655_ vdd gnd FILL
XFILL_2__1724_ vdd gnd FILL
X_943_ _943_/A _943_/B _943_/C _943_/Y vdd gnd OAI21X1
XFILL_2__1586_ vdd gnd FILL
X_1781_ _1781_/A _1781_/B _1802_/B _1782_/A vdd gnd OAI21X1
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1222_ vdd gnd FILL
XFILL_0__1084_ vdd gnd FILL
X_1146_ _1164_/B _1164_/A _1170_/A _1151_/A vdd gnd AOI21X1
XFILL_1__955_ vdd gnd FILL
X_1215_ _1215_/A _1296_/C _1215_/C _1257_/A vdd gnd NAND3X1
XFILL_1__1400_ vdd gnd FILL
XFILL_1__1193_ vdd gnd FILL
X_1077_ _984_/A _1781_/A _1082_/A _1760_/A _1237_/A vdd gnd AOI22X1
XFILL_1__1331_ vdd gnd FILL
XFILL_1__1262_ vdd gnd FILL
XFILL_3__1129_ vdd gnd FILL
XFILL_1__1529_ vdd gnd FILL
XFILL_2__1440_ vdd gnd FILL
XFILL_2__1371_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
XFILL_2__1638_ vdd gnd FILL
XFILL_2__1707_ vdd gnd FILL
XFILL_0__1771_ vdd gnd FILL
X_926_ ABCmd_i[0] _928_/A vdd gnd INVX1
X_1000_ _999_/Y _1005_/B vdd gnd INVX1
XCLKBUF1_insert11 clk _1631_/CLK vdd gnd CLKBUF1
XFILL_2__1569_ vdd gnd FILL
X_1764_ _1809_/B _1765_/B _1765_/A _1803_/A vdd gnd OAI21X1
XFILL_0__1067_ vdd gnd FILL
XFILL_0__1205_ vdd gnd FILL
XFILL_0__1136_ vdd gnd FILL
X_1695_ _988_/A _1696_/B vdd gnd INVX1
XFILL_1__938_ vdd gnd FILL
X_1129_ _1207_/B _1129_/B _1208_/A vdd gnd NAND2X1
XFILL_1__1176_ vdd gnd FILL
XFILL_1__1314_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_2__1354_ vdd gnd FILL
XFILL_2__1423_ vdd gnd FILL
XFILL_0__956_ vdd gnd FILL
X_1480_ _1480_/A _1480_/B _1481_/B vdd gnd NAND2X1
XFILL_2_BUFX2_insert18 vdd gnd FILL
XFILL_2_BUFX2_insert29 vdd gnd FILL
XFILL_0__1823_ vdd gnd FILL
XFILL_0__1685_ vdd gnd FILL
XFILL_0__1754_ vdd gnd FILL
X_909_ _915_/B _909_/B _924_/A _910_/C vdd gnd OAI21X1
XFILL_1__1030_ vdd gnd FILL
X_1678_ ABCmd_i[1] _1678_/B ABCmd_i[0] _1680_/B vdd gnd MUX2X1
X_1816_ _1816_/A _1816_/B _1816_/C _1817_/B vdd gnd NAND3X1
X_1747_ _1747_/A _1747_/B _1747_/C _1772_/A vdd gnd OAI21X1
XFILL_0__1119_ vdd gnd FILL
XFILL_1__1794_ vdd gnd FILL
XFILL_1_BUFX2_insert4 vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_2__1070_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL_0__1470_ vdd gnd FILL
XFILL_2__1406_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
XFILL_2__1268_ vdd gnd FILL
XFILL_2__1199_ vdd gnd FILL
X_1601_ _986_/D _1601_/B _1602_/C vdd gnd NAND2X1
XFILL_0__939_ vdd gnd FILL
X_1532_ _1532_/A _899_/A _911_/A _1533_/D vdd gnd AOI21X1
XFILL_0__1806_ vdd gnd FILL
X_1463_ _1506_/B _1467_/B vdd gnd INVX1
X_1394_ _1394_/A _1445_/C _1408_/A vdd gnd XNOR2X1
XFILL_2__970_ vdd gnd FILL
XFILL_0__1668_ vdd gnd FILL
XFILL_0__1737_ vdd gnd FILL
XFILL_0__1599_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_1__1777_ vdd gnd FILL
XFILL_2__1053_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_0__1453_ vdd gnd FILL
XFILL_0__1522_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
XFILL_1__1700_ vdd gnd FILL
X_1515_ _1515_/A _1517_/C _1515_/C _1570_/B vdd gnd NAND3X1
XFILL_1__1562_ vdd gnd FILL
X_1446_ _1447_/A _1447_/B _1488_/C vdd gnd NAND2X1
X_1377_ _1439_/A _1382_/A vdd gnd INVX1
XFILL_2__953_ vdd gnd FILL
XFILL_1__1493_ vdd gnd FILL
XFILL92550x62550 vdd gnd FILL
XFILL_2__1671_ vdd gnd FILL
XFILL_2__1740_ vdd gnd FILL
X_890_ _904_/B _904_/C _903_/A vdd gnd NOR2X1
XFILL_2__1036_ vdd gnd FILL
XFILL_2__1105_ vdd gnd FILL
XFILL_3__1780_ vdd gnd FILL
XFILL_1__971_ vdd gnd FILL
X_1300_ _962_/B _948_/A _1373_/A vdd gnd NAND2X1
X_1231_ _1231_/A _1231_/B _1231_/C _1247_/B vdd gnd NAND3X1
X_1162_ _1162_/A _1162_/B _1203_/A _1205_/A vdd gnd AOI21X1
XFILL_0__1436_ vdd gnd FILL
XBUFX2_insert5 _1609_/Q _984_/A vdd gnd BUFX2
X_1093_ _1114_/B _1098_/C _1212_/C vdd gnd NAND2X1
XFILL_0__1505_ vdd gnd FILL
XFILL_0__1367_ vdd gnd FILL
XFILL_0__1298_ vdd gnd FILL
X_1429_ _1429_/A _1429_/B _1429_/C _1430_/A vdd gnd AOI21X1
XFILL_1_BUFX2_insert20 vdd gnd FILL
XFILL_1_BUFX2_insert31 vdd gnd FILL
XFILL_1__1545_ vdd gnd FILL
XFILL_1__1476_ vdd gnd FILL
XFILL92550x74250 vdd gnd FILL
XFILL_2__936_ vdd gnd FILL
XFILL_1_CLKBUF1_insert10 vdd gnd FILL
XFILL_2__1654_ vdd gnd FILL
XFILL_2__1723_ vdd gnd FILL
X_942_ _999_/B _949_/B _943_/C vdd gnd NAND2X1
XFILL_2__1585_ vdd gnd FILL
XFILL_0__1221_ vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
X_1780_ _1780_/A _948_/A _1780_/C _1780_/D _1782_/B vdd gnd AOI22X1
XFILL_2__1019_ vdd gnd FILL
XFILL_0__1083_ vdd gnd FILL
XFILL_3__1763_ vdd gnd FILL
XFILL_3__1694_ vdd gnd FILL
XFILL_1__954_ vdd gnd FILL
X_1145_ _969_/A _1301_/A _960_/A _1164_/A vdd gnd OAI21X1
X_1214_ _1217_/B _1217_/A _1215_/C vdd gnd OR2X2
XFILL_1__1330_ vdd gnd FILL
XFILL_1__1192_ vdd gnd FILL
X_1076_ _984_/A _1781_/A _1325_/B _1237_/C vdd gnd NAND3X1
XFILL_0__1419_ vdd gnd FILL
XFILL_1__1261_ vdd gnd FILL
XFILL_1__1528_ vdd gnd FILL
XFILL_1__1459_ vdd gnd FILL
XFILL_2__1370_ vdd gnd FILL
XFILL_2__919_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
X_925_ reset _925_/Y vdd gnd INVX8
XFILL_2__1637_ vdd gnd FILL
XFILL_2__1706_ vdd gnd FILL
XFILL_0__1770_ vdd gnd FILL
XFILL_2__1568_ vdd gnd FILL
XFILL_0__1204_ vdd gnd FILL
XFILL_2__1499_ vdd gnd FILL
XCLKBUF1_insert12 clk _1624_/CLK vdd gnd CLKBUF1
X_1763_ _1784_/A _945_/A _1763_/C _1765_/B vdd gnd AOI21X1
X_1694_ _1780_/A _988_/A _1694_/C _1780_/D _1698_/A vdd gnd AOI22X1
XFILL_0__1066_ vdd gnd FILL
XFILL_0__1135_ vdd gnd FILL
XFILL_3__1677_ vdd gnd FILL
XFILL_3__1815_ vdd gnd FILL
XFILL_3__1746_ vdd gnd FILL
XFILL_1__937_ vdd gnd FILL
X_1059_ _1108_/B _1074_/C _1108_/A _1067_/A vdd gnd OAI21X1
XFILL_1__1313_ vdd gnd FILL
X_1128_ _1128_/A _1128_/B _1128_/C _1129_/B vdd gnd NAND3X1
XFILL_1__1175_ vdd gnd FILL
XFILL_1__1244_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_2__1353_ vdd gnd FILL
XFILL_2__1284_ vdd gnd FILL
XFILL_0__955_ vdd gnd FILL
XFILL_0__1753_ vdd gnd FILL
XFILL_3__1531_ vdd gnd FILL
X_908_ LoadCmd_i _924_/A vdd gnd INVX1
XFILL_3__1600_ vdd gnd FILL
XFILL_2_BUFX2_insert19 vdd gnd FILL
XFILL_0__1822_ vdd gnd FILL
XFILL_0__1684_ vdd gnd FILL
XFILL_3__1462_ vdd gnd FILL
XFILL_3__1393_ vdd gnd FILL
X_1815_ _1815_/A _1815_/B _1815_/C _1817_/A vdd gnd NAND3X1
X_1677_ _1677_/A _1783_/C _1683_/B _1684_/B vdd gnd OAI21X1
X_1746_ _1746_/A _1746_/B _1802_/B _1747_/A vdd gnd OAI21X1
XFILL_0__1049_ vdd gnd FILL
XFILL_0__1118_ vdd gnd FILL
XFILL_1__1793_ vdd gnd FILL
XFILL_3__1729_ vdd gnd FILL
XFILL_1_BUFX2_insert5 vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_2__1405_ vdd gnd FILL
XFILL_2__1198_ vdd gnd FILL
XFILL_0__938_ vdd gnd FILL
XFILL_2__1336_ vdd gnd FILL
XFILL_2__1267_ vdd gnd FILL
X_1531_ _949_/A _1531_/B _1531_/C _1532_/A vdd gnd OAI21X1
X_1600_ _937_/A _1601_/B _1600_/C _1628_/D vdd gnd OAI21X1
X_1462_ _1462_/A _1462_/B _1462_/C _1466_/C vdd gnd OAI21X1
XFILL_0__1805_ vdd gnd FILL
XFILL_0__1736_ vdd gnd FILL
XFILL_3__1514_ vdd gnd FILL
XFILL_3__1445_ vdd gnd FILL
X_1393_ _1445_/A _1456_/C _1393_/C _1394_/A vdd gnd OAI21X1
XFILL_0__1667_ vdd gnd FILL
XFILL_0__1598_ vdd gnd FILL
XFILL_3__1376_ vdd gnd FILL
XFILL_1__1012_ vdd gnd FILL
X_1729_ _1778_/A _939_/A _1732_/B vdd gnd AND2X2
XFILL_1__1776_ vdd gnd FILL
XFILL_2__1052_ vdd gnd FILL
XFILL_2__1121_ vdd gnd FILL
XFILL_3__934_ vdd gnd FILL
XFILL_2__1319_ vdd gnd FILL
XFILL_0__1452_ vdd gnd FILL
XFILL_0__1521_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_3__1230_ vdd gnd FILL
X_1514_ _1520_/B _1520_/A _1517_/C vdd gnd NOR2X1
X_1445_ _1445_/A _1456_/C _1445_/C _1445_/D _1447_/B vdd gnd OAI22X1
XFILL_0__1719_ vdd gnd FILL
XFILL_3__1428_ vdd gnd FILL
XFILL_1__1561_ vdd gnd FILL
XFILL_1__1492_ vdd gnd FILL
X_1376_ _988_/B _948_/A _1439_/A vdd gnd NAND2X1
XFILL_3__1359_ vdd gnd FILL
XFILL_2__952_ vdd gnd FILL
XFILL_2__1670_ vdd gnd FILL
XFILL_1__1759_ vdd gnd FILL
XFILL_2__1035_ vdd gnd FILL
XFILL_2__1104_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
XFILL_2__1799_ vdd gnd FILL
XBUFX2_insert6 _1609_/Q _1679_/A vdd gnd BUFX2
XFILL_3__917_ vdd gnd FILL
X_1092_ _1302_/A _986_/D _1098_/C vdd gnd AND2X2
X_1230_ _1304_/D _1231_/B vdd gnd INVX1
X_1161_ _1206_/C _1266_/B _1266_/A _1162_/A vdd gnd OAI21X1
XFILL_3__1144_ vdd gnd FILL
XFILL_3__1075_ vdd gnd FILL
XFILL_3__1213_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_0__1504_ vdd gnd FILL
XFILL_0__1435_ vdd gnd FILL
XFILL92250x4050 vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
X_1428_ _1428_/A _922_/C _1433_/D vdd gnd NOR2X1
XFILL_1_BUFX2_insert21 vdd gnd FILL
XFILL_1_BUFX2_insert32 vdd gnd FILL
X_1359_ _1361_/A _1361_/B _1362_/B vdd gnd AND2X2
XFILL_1_CLKBUF1_insert11 vdd gnd FILL
XFILL_1__1475_ vdd gnd FILL
XFILL_1__1544_ vdd gnd FILL
XFILL_2__935_ vdd gnd FILL
XFILL_2__1722_ vdd gnd FILL
X_941_ ABCmd_i[5] _943_/A vdd gnd INVX1
XFILL_2__1653_ vdd gnd FILL
XFILL_2__1584_ vdd gnd FILL
XFILL_0__1220_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL_2__1018_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
XFILL_1__953_ vdd gnd FILL
X_1213_ _1217_/A _1217_/B _1296_/C vdd gnd NAND2X1
X_1144_ _961_/A _1164_/B vdd gnd INVX1
X_1075_ _1075_/A _1075_/B _1088_/A _1104_/A vdd gnd OAI21X1
XFILL_1__1260_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_3__1058_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_3__1127_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_1__1527_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_1__1458_ vdd gnd FILL
XFILL_2__918_ vdd gnd FILL
XFILL_2__1705_ vdd gnd FILL
X_924_ _924_/A _924_/B _924_/C _924_/Y vdd gnd OAI21X1
XFILL_2__1636_ vdd gnd FILL
XFILL_2__1567_ vdd gnd FILL
XFILL_2__1498_ vdd gnd FILL
XFILL_0__1203_ vdd gnd FILL
XFILL_0__1134_ vdd gnd FILL
X_1762_ _1784_/A _945_/A _1783_/C _1763_/C vdd gnd OAI21X1
X_1693_ _962_/B _988_/A _1778_/A _1694_/C vdd gnd NAND3X1
XFILL_0__1065_ vdd gnd FILL
XFILL_1__936_ vdd gnd FILL
X_1058_ _1108_/C _1074_/A _1074_/B _1067_/B vdd gnd NAND3X1
XFILL_1__1312_ vdd gnd FILL
XFILL_1__1243_ vdd gnd FILL
X_1127_ _1127_/A _1127_/B _1207_/A _1207_/B vdd gnd NAND3X1
XFILL_1__1174_ vdd gnd FILL
XFILL_2__1352_ vdd gnd FILL
XFILL_2__1421_ vdd gnd FILL
XFILL_0__954_ vdd gnd FILL
XFILL_2__1283_ vdd gnd FILL
XFILL_0__1752_ vdd gnd FILL
X_907_ _922_/C _914_/C vdd gnd INVX1
XFILL_0__1821_ vdd gnd FILL
XFILL_0__1683_ vdd gnd FILL
X_1814_ _1816_/A _1816_/B _1815_/C vdd gnd NAND2X1
X_1745_ _1780_/A _999_/B _1745_/C _1780_/D _1747_/B vdd gnd AOI22X1
XFILL_0__1117_ vdd gnd FILL
X_1676_ _1678_/B _1676_/B _1676_/C _1683_/B vdd gnd OAI21X1
XFILL_1__1792_ vdd gnd FILL
XFILL_0__1048_ vdd gnd FILL
XFILL_1_BUFX2_insert6 vdd gnd FILL
XFILL_1__919_ vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_3__950_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_2__1404_ vdd gnd FILL
XFILL_2__1335_ vdd gnd FILL
XFILL_2__1197_ vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
XFILL_2__1266_ vdd gnd FILL
X_1530_ _1794_/B _949_/A _1531_/C vdd gnd NAND2X1
X_1461_ _1466_/B _1506_/B _1467_/C _1465_/C vdd gnd NAND3X1
X_1392_ _1445_/D _1393_/C vdd gnd INVX1
XFILL_0__1804_ vdd gnd FILL
XFILL_0__1666_ vdd gnd FILL
XFILL_0__1735_ vdd gnd FILL
XFILL_0__1597_ vdd gnd FILL
XFILL_1__1011_ vdd gnd FILL
X_1728_ ABCmd_i[5] _1746_/A _1733_/C vdd gnd NAND2X1
X_1659_ _1659_/A _1661_/A _1792_/A vdd gnd XOR2X1
XFILL_1__1775_ vdd gnd FILL
XFILL_2__1051_ vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_2__1120_ vdd gnd FILL
XFILL_0__1520_ vdd gnd FILL
XFILL_3__1091_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
XFILL_2__1249_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_3__1160_ vdd gnd FILL
X_1375_ _1375_/A _1375_/B _1375_/C _1413_/C vdd gnd AOI21X1
X_1444_ _1496_/A _1567_/B _1447_/A vdd gnd NOR2X1
X_1513_ _1513_/A _1513_/B _1515_/C vdd gnd NOR2X1
XFILL_0__1649_ vdd gnd FILL
XFILL_0__1718_ vdd gnd FILL
XFILL_1__1560_ vdd gnd FILL
XFILL_1__1491_ vdd gnd FILL
XFILL_2__951_ vdd gnd FILL
XFILL_1__1758_ vdd gnd FILL
XFILL_1__1689_ vdd gnd FILL
XFILL_2__1103_ vdd gnd FILL
XFILL_2__1034_ vdd gnd FILL
XFILL_2__1798_ vdd gnd FILL
XBUFX2_insert7 _1609_/Q _967_/A vdd gnd BUFX2
X_1091_ _976_/A _988_/B _1114_/B vdd gnd AND2X2
XFILL_0__1503_ vdd gnd FILL
X_1160_ _1206_/A _1206_/B _1266_/C _1162_/B vdd gnd NAND3X1
XFILL_0__1434_ vdd gnd FILL
XFILL_0__1365_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
X_1427_ ABCmd_i[7] _1797_/Y _1428_/A vdd gnd NOR2X1
XFILL_1_BUFX2_insert33 vdd gnd FILL
XFILL_1_BUFX2_insert22 vdd gnd FILL
X_1358_ _1358_/A _1358_/B _1358_/C _1364_/C vdd gnd OAI21X1
X_1289_ _1289_/A _1289_/B _1289_/C _1290_/B vdd gnd AOI21X1
XFILL_1__1474_ vdd gnd FILL
XFILL_1__1543_ vdd gnd FILL
XFILL_1_CLKBUF1_insert12 vdd gnd FILL
XFILL_2__934_ vdd gnd FILL
XFILL_2__1721_ vdd gnd FILL
XFILL_2__1652_ vdd gnd FILL
X_940_ _940_/A _940_/B _940_/C _940_/Y vdd gnd OAI21X1
XFILL_2__1583_ vdd gnd FILL
XFILL_0__1150_ vdd gnd FILL
XFILL_3__1761_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
XFILL_3__1692_ vdd gnd FILL
XFILL_1__952_ vdd gnd FILL
X_1212_ _1212_/A _1212_/B _1212_/C _1217_/B vdd gnd OAI21X1
X_1143_ _960_/A _960_/B _1170_/A vdd gnd NOR2X1
X_1074_ _1074_/A _1074_/B _1074_/C _1126_/C vdd gnd AOI21X1
XFILL_0__1417_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_0__1348_ vdd gnd FILL
XFILL_1__1526_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
XFILL_2__917_ vdd gnd FILL
XFILL93150x150 vdd gnd FILL
XFILL_1__1457_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_2__1704_ vdd gnd FILL
X_923_ _923_/A _923_/B _924_/C vdd gnd AND2X2
XFILL_2__1566_ vdd gnd FILL
XFILL_2__1497_ vdd gnd FILL
X_1761_ _1802_/B _1810_/B _1761_/C _1761_/D _1765_/A vdd gnd OAI22X1
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
XFILL_3__1813_ vdd gnd FILL
X_1692_ ABCmd_i[5] _988_/B _1698_/C vdd gnd NAND2X1
XFILL_3__1744_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
XFILL_3__1675_ vdd gnd FILL
XFILL_1__935_ vdd gnd FILL
X_1126_ _1126_/A _1126_/B _1126_/C _1256_/C vdd gnd AOI21X1
XFILL_1__1173_ vdd gnd FILL
X_1057_ _1154_/A _1153_/B _994_/Y _1067_/C vdd gnd OAI21X1
XFILL_1__1242_ vdd gnd FILL
XFILL_1__1311_ vdd gnd FILL
XFILL_2__1282_ vdd gnd FILL
XFILL_2__1351_ vdd gnd FILL
XFILL_2__1420_ vdd gnd FILL
XFILL_1__1509_ vdd gnd FILL
XFILL_0__953_ vdd gnd FILL
XFILL_0__1820_ vdd gnd FILL
XFILL_0__1682_ vdd gnd FILL
XFILL_0__1751_ vdd gnd FILL
X_906_ _915_/A _911_/A _922_/C vdd gnd NOR2X1
XFILL_3__1391_ vdd gnd FILL
XFILL_3__1460_ vdd gnd FILL
XFILL_2__1549_ vdd gnd FILL
X_1813_ _1813_/A _1813_/B _1813_/C _1816_/B vdd gnd NAND3X1
X_1744_ _1746_/A _1746_/B _1745_/C vdd gnd NAND2X1
XFILL_0__1047_ vdd gnd FILL
XFILL_0__1116_ vdd gnd FILL
X_1675_ _1675_/A _1676_/C vdd gnd INVX1
XFILL_1__1791_ vdd gnd FILL
XFILL_3__1727_ vdd gnd FILL
XFILL_3__1658_ vdd gnd FILL
XFILL_1_BUFX2_insert7 vdd gnd FILL
XFILL_1__918_ vdd gnd FILL
XFILL_3__1589_ vdd gnd FILL
X_1109_ _1246_/C _1220_/B _1220_/A _1125_/B vdd gnd NAND3X1
XFILL_1__1156_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL_2__1403_ vdd gnd FILL
XFILL_2__1334_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL_2__1196_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
XFILL_0__1803_ vdd gnd FILL
X_1391_ _1781_/A _952_/A _1760_/A _1452_/B _1445_/D vdd gnd AOI22X1
X_1460_ _1460_/A _1460_/B _1460_/C _1506_/B vdd gnd NAND3X1
XFILL_0__1665_ vdd gnd FILL
XFILL_0__1734_ vdd gnd FILL
XFILL_0__1596_ vdd gnd FILL
XFILL_3__1374_ vdd gnd FILL
XFILL_3__1512_ vdd gnd FILL
XFILL_3__1443_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
X_1658_ _1684_/A _1660_/A _1661_/C _1659_/A vdd gnd OAI21X1
X_1727_ _1727_/A _1793_/A _1727_/C _1741_/A vdd gnd OAI21X1
XFILL_1__1774_ vdd gnd FILL
X_1589_ _1808_/C _949_/A _1590_/C vdd gnd NAND2X1
XFILL_2__1050_ vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_3__932_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_2__1248_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
XFILL_2__1317_ vdd gnd FILL
XFILL_2__1179_ vdd gnd FILL
XFILL_0__919_ vdd gnd FILL
X_1512_ _1558_/A _1558_/C _1548_/A vdd gnd NAND2X1
X_1374_ _1414_/A _1472_/A vdd gnd INVX1
X_1443_ _1488_/A _1449_/A vdd gnd INVX1
XFILL_0__1648_ vdd gnd FILL
XFILL_0__1717_ vdd gnd FILL
XFILL_0__1579_ vdd gnd FILL
XFILL_3__1288_ vdd gnd FILL
XFILL_2__950_ vdd gnd FILL
XFILL_1__1490_ vdd gnd FILL
XFILL_3__1426_ vdd gnd FILL
XFILL_3__1357_ vdd gnd FILL
XFILL_1__1688_ vdd gnd FILL
XFILL_1__1757_ vdd gnd FILL
XFILL_1__1826_ vdd gnd FILL
XFILL_2__1033_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_2__1797_ vdd gnd FILL
XFILL_3__915_ vdd gnd FILL
XFILL_3__1142_ vdd gnd FILL
XFILL_0__1433_ vdd gnd FILL
XFILL_0__1502_ vdd gnd FILL
XFILL_3__1211_ vdd gnd FILL
X_1090_ _1212_/A _1096_/A vdd gnd INVX1
XFILL_3__1073_ vdd gnd FILL
XFILL_0__1364_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
XFILL_1_BUFX2_insert34 vdd gnd FILL
X_1288_ _1289_/B _1289_/C _1289_/A _1576_/A vdd gnd NAND3X1
XFILL_1_BUFX2_insert23 vdd gnd FILL
X_1426_ _1475_/C _1426_/B ABCmd_i[7] _1433_/C vdd gnd OAI21X1
XFILL_1__1542_ vdd gnd FILL
X_1357_ _1513_/B _1357_/B ABCmd_i[7] _1358_/A vdd gnd OAI21X1
XFILL_2__933_ vdd gnd FILL
XFILL_1__1473_ vdd gnd FILL
XFILL_3__1409_ vdd gnd FILL
XFILL_1__1809_ vdd gnd FILL
XFILL_2__1651_ vdd gnd FILL
XFILL_2__1720_ vdd gnd FILL
XFILL_2__1582_ vdd gnd FILL
XFILL_2__1016_ vdd gnd FILL
XFILL_0__1080_ vdd gnd FILL
X_1142_ _955_/Y _1198_/C vdd gnd INVX1
XFILL_1__951_ vdd gnd FILL
X_999_ _999_/A _999_/B _999_/Y vdd gnd NAND2X1
X_1211_ _1211_/A _1567_/B _1217_/A vdd gnd NOR2X1
X_1073_ _1158_/A _1157_/B _1158_/C _1138_/C vdd gnd OAI21X1
XFILL_0__1416_ vdd gnd FILL
XFILL93150x19650 vdd gnd FILL
XFILL_3__1125_ vdd gnd FILL
XFILL_3__1056_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
XFILL_0__1347_ vdd gnd FILL
X_1409_ _1409_/A _1409_/B _1462_/A _1413_/B vdd gnd AOI21X1
XFILL_1__1525_ vdd gnd FILL
XFILL_2__916_ vdd gnd FILL
XFILL_1__1387_ vdd gnd FILL
XFILL_1__1456_ vdd gnd FILL
XFILL_2__1703_ vdd gnd FILL
X_922_ _922_/A _922_/B _922_/C _923_/B vdd gnd NAND3X1
XFILL_2__1565_ vdd gnd FILL
XFILL_0__1201_ vdd gnd FILL
XFILL_2__1496_ vdd gnd FILL
X_1691_ _1691_/A _1691_/B _1722_/A _1721_/B vdd gnd OAI21X1
X_1760_ _1760_/A _1760_/B _1802_/B _1761_/C vdd gnd OAI21X1
XFILL_0__1132_ vdd gnd FILL
XFILL_0__1063_ vdd gnd FILL
XFILL_1__934_ vdd gnd FILL
X_1125_ _1125_/A _1125_/B _1125_/C _1208_/B vdd gnd AOI21X1
XFILL_1__1310_ vdd gnd FILL
XFILL_1__1172_ vdd gnd FILL
X_1056_ _1068_/B _1068_/C _1068_/A _1158_/B vdd gnd NAND3X1
XFILL_3__1108_ vdd gnd FILL
XFILL_1__1241_ vdd gnd FILL
XFILL_3__1039_ vdd gnd FILL
XFILL_2__1281_ vdd gnd FILL
XFILL_1__1508_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_1_CLKBUF1_insert8 vdd gnd FILL
XFILL_0__952_ vdd gnd FILL
X_905_ LoadB_i _922_/B vdd gnd INVX1
XFILL_0__1681_ vdd gnd FILL
XFILL_0__1750_ vdd gnd FILL
XFILL_2__1548_ vdd gnd FILL
XFILL_2__1479_ vdd gnd FILL
X_1674_ _1674_/A _1674_/B _1722_/C vdd gnd NAND2X1
X_1812_ _1812_/A _1813_/B vdd gnd INVX1
X_1743_ _1778_/A _999_/B _1746_/B vdd gnd AND2X2
XFILL_0__1046_ vdd gnd FILL
XFILL_0__1115_ vdd gnd FILL
XFILL_1__1790_ vdd gnd FILL
XFILL_1__917_ vdd gnd FILL
X_1108_ _1108_/A _1108_/B _1108_/C _1125_/C vdd gnd OAI21X1
X_1039_ _1049_/A _1114_/D vdd gnd INVX1
XFILL92850x4050 vdd gnd FILL
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1086_ vdd gnd FILL
XFILL_1__1224_ vdd gnd FILL
XFILL92550x70350 vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_2__1195_ vdd gnd FILL
XFILL_2__1333_ vdd gnd FILL
XFILL_2__1264_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
XFILL_0__1802_ vdd gnd FILL
XFILL_0__1733_ vdd gnd FILL
X_1390_ _1781_/A _1452_/B _1456_/C vdd gnd NAND2X1
XFILL_0__1664_ vdd gnd FILL
XFILL_0__1595_ vdd gnd FILL
X_1657_ _1809_/B _1660_/A _1684_/A _1661_/C vdd gnd OAI21X1
X_1726_ _1769_/C _1727_/C vdd gnd INVX1
XFILL_0__1029_ vdd gnd FILL
X_1588_ _1588_/A _1588_/B _1590_/B vdd gnd XNOR2X1
XFILL_1__1773_ vdd gnd FILL
XFILL92550x82050 vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_2__1178_ vdd gnd FILL
XFILL_2__1316_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
XFILL_2__1247_ vdd gnd FILL
XFILL_0__918_ vdd gnd FILL
X_1511_ _1511_/A _1511_/B _1511_/C _1558_/A vdd gnd NAND3X1
X_1442_ _986_/D _948_/A _1488_/A vdd gnd NAND2X1
XFILL_0__1716_ vdd gnd FILL
X_1373_ _1373_/A _1373_/B _1373_/C _1414_/A vdd gnd OAI21X1
XFILL_0__1647_ vdd gnd FILL
XFILL_0__1578_ vdd gnd FILL
X_1709_ ABCmd_i[5] _986_/D _1714_/C vdd gnd NAND2X1
XFILL_1__1825_ vdd gnd FILL
XFILL_1__1687_ vdd gnd FILL
XFILL_1__1756_ vdd gnd FILL
XFILL_2__1032_ vdd gnd FILL
XFILL_2__1101_ vdd gnd FILL
XFILL_2__1796_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_0__1501_ vdd gnd FILL
XFILL_0__1294_ vdd gnd FILL
XFILL_1_BUFX2_insert24 vdd gnd FILL
XFILL_1_BUFX2_insert13 vdd gnd FILL
X_1425_ _1476_/B _1476_/A _1426_/B vdd gnd NOR2X1
X_1287_ _1287_/A _1287_/B _1287_/C _1289_/A vdd gnd NAND3X1
XFILL_1_BUFX2_insert35 vdd gnd FILL
XFILL_1__1472_ vdd gnd FILL
X_1356_ _1357_/B _1513_/B _1358_/B vdd gnd AND2X2
XFILL_1__1541_ vdd gnd FILL
XFILL_2__932_ vdd gnd FILL
XFILL_2__1650_ vdd gnd FILL
XFILL_1__1808_ vdd gnd FILL
XFILL_2__1581_ vdd gnd FILL
XFILL_1__1739_ vdd gnd FILL
XFILL_2__1015_ vdd gnd FILL
XFILL_3__1690_ vdd gnd FILL
XFILL_1__950_ vdd gnd FILL
XFILL_2__1779_ vdd gnd FILL
X_998_ _998_/A _998_/B _998_/C _998_/Y vdd gnd NAND3X1
X_1210_ _1296_/A _1215_/A vdd gnd INVX1
X_1072_ _1266_/A _1206_/A vdd gnd INVX1
X_1141_ _1291_/C _1587_/B vdd gnd INVX1
XFILL_0__1346_ vdd gnd FILL
XFILL_0__1415_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1408_/A _1408_/B _1409_/B vdd gnd NAND2X1
XFILL_1__1455_ vdd gnd FILL
X_1339_ _1339_/A _1339_/B _1339_/C _1346_/C vdd gnd AOI21X1
XFILL_1__1524_ vdd gnd FILL
XFILL_2__915_ vdd gnd FILL
XFILL_1__1386_ vdd gnd FILL
XFILL_2__1702_ vdd gnd FILL
X_921_ _921_/A _921_/B _921_/C _921_/D _923_/A vdd gnd AOI22X1
XFILL91650x7950 vdd gnd FILL
XFILL_2__1564_ vdd gnd FILL
XFILL_0__1200_ vdd gnd FILL
XFILL_2__1495_ vdd gnd FILL
X_1690_ _1690_/A _1690_/B _1691_/A vdd gnd NOR2X1
XFILL_3__1811_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
XFILL_0__1131_ vdd gnd FILL
XFILL_3__1673_ vdd gnd FILL
XFILL_3__1742_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
X_1055_ _1108_/A _1108_/C _1074_/A _1068_/B vdd gnd NAND3X1
X_1124_ _1256_/B _1256_/A _1208_/C _1138_/A vdd gnd NAND3X1
XFILL_1__1171_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
XFILL_0__1329_ vdd gnd FILL
XFILL_0__951_ vdd gnd FILL
XFILL_2__1280_ vdd gnd FILL
XFILL_1__1507_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
XFILL_1_CLKBUF1_insert9 vdd gnd FILL
X_904_ _915_/A _904_/B _904_/C _911_/B vdd gnd OAI21X1
XFILL_0__1680_ vdd gnd FILL
XFILL_2__1547_ vdd gnd FILL
XFILL_2__1478_ vdd gnd FILL
X_1811_ _1811_/A _1812_/A _1811_/C _1816_/A vdd gnd NAND3X1
XFILL_0__1114_ vdd gnd FILL
X_1673_ _1673_/A _1673_/B _1690_/B _1674_/A vdd gnd MUX2X1
X_1742_ ABCmd_i[5] _1760_/A _1747_/C vdd gnd NAND2X1
XFILL_0__1045_ vdd gnd FILL
XFILL_3__1656_ vdd gnd FILL
XFILL_3__1725_ vdd gnd FILL
XFILL_1__916_ vdd gnd FILL
XFILL_3__1587_ vdd gnd FILL
X_1038_ _999_/B _978_/B _1049_/A vdd gnd NAND2X1
XFILL_1__1223_ vdd gnd FILL
X_1107_ _1126_/B _1126_/A _1126_/C _1256_/A vdd gnd NAND3X1
XFILL_1__1154_ vdd gnd FILL
XFILL_1__1085_ vdd gnd FILL
XFILL92850x54750 vdd gnd FILL
XFILL92550x89850 vdd gnd FILL
XFILL_2__1401_ vdd gnd FILL
XFILL_2__1332_ vdd gnd FILL
XFILL_2__1194_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_2__1263_ vdd gnd FILL
XFILL_0__1801_ vdd gnd FILL
XFILL_0__1732_ vdd gnd FILL
XFILL_3__1441_ vdd gnd FILL
XFILL_3__1510_ vdd gnd FILL
XFILL_0__1663_ vdd gnd FILL
XFILL_0__1594_ vdd gnd FILL
XFILL_3__1372_ vdd gnd FILL
X_1725_ _1725_/A _1725_/B _1725_/C _1769_/C vdd gnd OAI21X1
X_1656_ _1784_/A _1783_/C _1809_/B vdd gnd NOR2X1
XFILL_1__1772_ vdd gnd FILL
XFILL_0__1028_ vdd gnd FILL
X_1587_ _1587_/A _1587_/B _1588_/A vdd gnd NAND2X1
XFILL_3__1639_ vdd gnd FILL
XFILL_3__1708_ vdd gnd FILL
XFILL92250x19650 vdd gnd FILL
XFILL_1__1206_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_3__930_ vdd gnd FILL
XFILL_2__1315_ vdd gnd FILL
XFILL_2__1177_ vdd gnd FILL
XFILL_0__917_ vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
X_1441_ _1441_/A _1441_/B _1441_/C _1467_/C vdd gnd AOI21X1
X_1510_ _1510_/A _1510_/B _1511_/A vdd gnd NAND2X1
XFILL_0__1715_ vdd gnd FILL
XFILL_0__1646_ vdd gnd FILL
XFILL_3__1424_ vdd gnd FILL
X_1372_ _1372_/A _1372_/B _1373_/C vdd gnd NAND2X1
XFILL_0__1577_ vdd gnd FILL
XFILL_3__1286_ vdd gnd FILL
XFILL_3__1355_ vdd gnd FILL
X_1708_ _1708_/A _1708_/B _1721_/B _1722_/B _1725_/B vdd gnd AOI22X1
X_1639_ ABCmd_i[5] _1639_/B _1684_/D vdd gnd NOR2X1
XFILL_1__1755_ vdd gnd FILL
XFILL_1__1824_ vdd gnd FILL
XFILL_1__1686_ vdd gnd FILL
XFILL92850x78150 vdd gnd FILL
XFILL_2__1031_ vdd gnd FILL
XFILL_2__1100_ vdd gnd FILL
XFILL_3__913_ vdd gnd FILL
XFILL_3_BUFX2_insert0 vdd gnd FILL
XFILL_2__1795_ vdd gnd FILL
XFILL_0__1500_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
XFILL_2__1229_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_3__1140_ vdd gnd FILL
XFILL_1_BUFX2_insert36 vdd gnd FILL
XFILL_1_BUFX2_insert25 vdd gnd FILL
XFILL_1_BUFX2_insert14 vdd gnd FILL
X_1355_ _1370_/B _1355_/B _1513_/B vdd gnd NAND2X1
X_1424_ _1520_/A _1476_/B vdd gnd INVX1
X_1286_ _1286_/A _1286_/B _1287_/C vdd gnd NAND2X1
XFILL_3__1338_ vdd gnd FILL
XFILL_1__1471_ vdd gnd FILL
XFILL_3__1407_ vdd gnd FILL
XFILL_1__1540_ vdd gnd FILL
XFILL_2__931_ vdd gnd FILL
XFILL_3__1269_ vdd gnd FILL
XFILL_1__1807_ vdd gnd FILL
XFILL_1__1738_ vdd gnd FILL
XFILL_2__1580_ vdd gnd FILL
XFILL_1__1669_ vdd gnd FILL
XFILL_2__1014_ vdd gnd FILL
XFILL91650x70350 vdd gnd FILL
X_997_ _997_/A _997_/B _997_/C _998_/A vdd gnd NAND3X1
XFILL_2__1778_ vdd gnd FILL
X_1071_ _1071_/A _1071_/B _1266_/A vdd gnd NAND2X1
X_1140_ _1284_/C _1284_/B _1289_/B _1291_/C vdd gnd AOI21X1
XFILL_0__1276_ vdd gnd FILL
XFILL_3__1054_ vdd gnd FILL
XFILL_0__1345_ vdd gnd FILL
XFILL_0__1414_ vdd gnd FILL
XFILL_3__1123_ vdd gnd FILL
X_1338_ _1338_/A _1342_/B _1338_/C _1339_/C vdd gnd NOR3X1
X_1407_ _1408_/B _1408_/A _1409_/A vdd gnd OR2X2
XFILL_1__1454_ vdd gnd FILL
XFILL_1__1523_ vdd gnd FILL
X_1269_ _1269_/A _1367_/B _1269_/C _1370_/A vdd gnd NAND3X1
XFILL_1__1385_ vdd gnd FILL
XFILL_2__914_ vdd gnd FILL
XFILL_2__1701_ vdd gnd FILL
X_920_ _946_/B _921_/A vdd gnd INVX1
XFILL_2__1563_ vdd gnd FILL
XFILL_2__1494_ vdd gnd FILL
XFILL_0__1130_ vdd gnd FILL
XFILL91650x82050 vdd gnd FILL
XFILL_0__1061_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
X_1054_ _1054_/A _1054_/B _1108_/A vdd gnd NAND2X1
X_1123_ _1123_/A _1123_/B _1256_/B vdd gnd NAND2X1
XFILL_1__1170_ vdd gnd FILL
XFILL_3__1037_ vdd gnd FILL
XFILL_3__1106_ vdd gnd FILL
XFILL_0__1328_ vdd gnd FILL
XFILL_0__1259_ vdd gnd FILL
XFILL92250x7950 vdd gnd FILL
XFILL_1__1506_ vdd gnd FILL
XFILL_0__950_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
X_903_ _903_/A _911_/A vdd gnd INVX4
XFILL_2__1546_ vdd gnd FILL
XFILL_2__1477_ vdd gnd FILL
X_1810_ _1810_/A _1810_/B _1812_/A vdd gnd XOR2X1
X_1741_ _1741_/A _1741_/B _1741_/C _1755_/B vdd gnd AOI21X1
XFILL_0__1113_ vdd gnd FILL
X_1672_ _1716_/A _1783_/C _1673_/B _1673_/A vdd gnd OAI21X1
XFILL_0__1044_ vdd gnd FILL
XFILL_1__915_ vdd gnd FILL
X_1106_ _1246_/A _1246_/C _1220_/B _1126_/B vdd gnd NAND3X1
XFILL_1__1153_ vdd gnd FILL
X_1037_ _1052_/B _1052_/A _1052_/C _1074_/C vdd gnd AOI21X1
XFILL_1__1222_ vdd gnd FILL
XFILL_1__1084_ vdd gnd FILL
XFILL_2__1400_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_2__1262_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_0__1800_ vdd gnd FILL
XFILL_0__1662_ vdd gnd FILL
XFILL_0__1731_ vdd gnd FILL
XFILL_2__1529_ vdd gnd FILL
XFILL_0__1593_ vdd gnd FILL
X_1724_ ABCmd_i[6] _1792_/B _1727_/A vdd gnd NAND2X1
XFILL_0__1027_ vdd gnd FILL
X_1655_ _967_/A _1677_/A _1675_/A _1660_/A vdd gnd AOI21X1
XFILL_1__1771_ vdd gnd FILL
X_1586_ _1586_/A _1586_/B _1586_/C _1592_/C vdd gnd OAI21X1
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
XFILL_2__1314_ vdd gnd FILL
XFILL_2__1245_ vdd gnd FILL
XFILL_2__1176_ vdd gnd FILL
XFILL_0__916_ vdd gnd FILL
X_1440_ _1468_/A _1465_/A vdd gnd INVX1
X_1371_ _1521_/C _1423_/C vdd gnd INVX1
XFILL_0__1645_ vdd gnd FILL
XFILL_0__1714_ vdd gnd FILL
XFILL_0__1576_ vdd gnd FILL
X_1638_ _1676_/B _1783_/C ABCmd_i[4] _1639_/B vdd gnd OAI21X1
X_1707_ _1721_/A _1722_/B vdd gnd INVX1
XFILL_1__1685_ vdd gnd FILL
XFILL_1__1754_ vdd gnd FILL
XFILL_1__1823_ vdd gnd FILL
X_1569_ _1583_/C _1583_/B _1583_/A _1573_/B vdd gnd NAND3X1
XFILL_2__1030_ vdd gnd FILL
XFILL_1__1119_ vdd gnd FILL
XFILL_2__1794_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
XFILL_3__1070_ vdd gnd FILL
XFILL_2__1228_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_2__1159_ vdd gnd FILL
X_1285_ _1551_/A _1289_/C vdd gnd INVX1
XFILL_1_BUFX2_insert26 vdd gnd FILL
XFILL_1_BUFX2_insert15 vdd gnd FILL
XFILL_1_BUFX2_insert37 vdd gnd FILL
X_1354_ _1416_/B _1366_/B _1366_/C _1370_/B vdd gnd NAND3X1
X_1423_ _1522_/A _1522_/B _1423_/C _1476_/A vdd gnd OAI21X1
XFILL_2__930_ vdd gnd FILL
XFILL_1__1470_ vdd gnd FILL
XFILL_0__1559_ vdd gnd FILL
XFILL_1__1806_ vdd gnd FILL
XFILL_1__1668_ vdd gnd FILL
XFILL_1__1737_ vdd gnd FILL
XFILL_1__1599_ vdd gnd FILL
XBUFX2_insert40 ABCmd_i[2] _1784_/A vdd gnd BUFX2
XFILL_2__1013_ vdd gnd FILL
XFILL91950x54750 vdd gnd FILL
XFILL_2__1777_ vdd gnd FILL
X_996_ _996_/A _996_/B _996_/C _998_/B vdd gnd OAI21X1
X_1070_ _1286_/A _1286_/B _1180_/C _1289_/B vdd gnd NAND3X1
XFILL_0__1413_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
XFILL_0__1344_ vdd gnd FILL
X_1337_ _1417_/B _1417_/A _1417_/C _1418_/C vdd gnd NAND3X1
X_1406_ _1406_/A _1406_/B _1462_/C _1441_/B _1413_/A vdd gnd AOI22X1
X_1268_ _1295_/A _1295_/B _1367_/A _1367_/B vdd gnd NAND3X1
XFILL_1__1522_ vdd gnd FILL
X_1199_ _955_/Y _1287_/A _1199_/C _1200_/B vdd gnd NAND3X1
XFILL_2__913_ vdd gnd FILL
XFILL_1__1453_ vdd gnd FILL
XFILL_1__1384_ vdd gnd FILL
XFILL_2__1700_ vdd gnd FILL
XFILL_2__1562_ vdd gnd FILL
XFILL_2__1493_ vdd gnd FILL
XFILL_0__1060_ vdd gnd FILL
XFILL_3__1740_ vdd gnd FILL
XFILL_3__1671_ vdd gnd FILL
XFILL_1__931_ vdd gnd FILL
X_979_ _979_/A _979_/B _979_/C _980_/C vdd gnd OAI21X1
X_1122_ _1128_/A _1127_/B _1207_/A _1123_/A vdd gnd NAND3X1
X_1053_ _1053_/A _1088_/B _1053_/C _1108_/C vdd gnd NAND3X1
XFILL_0__1189_ vdd gnd FILL
XFILL_0__1258_ vdd gnd FILL
XFILL_0__1327_ vdd gnd FILL
XFILL_1__1505_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
X_902_ LoadA_i _922_/A vdd gnd INVX1
XFILL_2__1545_ vdd gnd FILL
XFILL91950x78150 vdd gnd FILL
XFILL_2__1476_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
X_1671_ _1690_/A _1673_/B vdd gnd INVX1
X_1740_ _1770_/C _1741_/C vdd gnd INVX1
XFILL_0__1112_ vdd gnd FILL
XFILL_3__1654_ vdd gnd FILL
XFILL_3__1723_ vdd gnd FILL
XFILL_1__914_ vdd gnd FILL
X_1105_ _1105_/A _1105_/B _1246_/A vdd gnd NAND2X1
XFILL_3__1585_ vdd gnd FILL
XFILL_1__1152_ vdd gnd FILL
X_1036_ _1102_/A _1075_/B _1088_/A _1052_/A vdd gnd NAND3X1
XFILL_1__1221_ vdd gnd FILL
XFILL_1__1083_ vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_2__1330_ vdd gnd FILL
XFILL_2__1261_ vdd gnd FILL
XFILL_2__1192_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL_0__1661_ vdd gnd FILL
XFILL_2__1528_ vdd gnd FILL
XFILL_0__1730_ vdd gnd FILL
XFILL_3__1370_ vdd gnd FILL
XFILL_0__1592_ vdd gnd FILL
XFILL_2__1459_ vdd gnd FILL
X_1654_ _967_/A _1677_/A _1783_/C _1675_/A vdd gnd OAI21X1
X_1723_ _1723_/A _1768_/B _1723_/C _1792_/B vdd gnd NAND3X1
XFILL_0__1026_ vdd gnd FILL
XFILL93150x15750 vdd gnd FILL
XFILL_3__1637_ vdd gnd FILL
XFILL_3__1706_ vdd gnd FILL
XFILL_1__1770_ vdd gnd FILL
X_1585_ _1585_/A _1585_/B _1586_/A vdd gnd NAND2X1
X_1019_ _998_/Y _1153_/C _1153_/A _1068_/C vdd gnd AOI21X1
XFILL_3__1499_ vdd gnd FILL
XFILL_3__1568_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_1__1204_ vdd gnd FILL
XFILL_1__1135_ vdd gnd FILL
XFILL_2__1175_ vdd gnd FILL
XFILL_2__1313_ vdd gnd FILL
XFILL_2__1244_ vdd gnd FILL
XFILL_0__915_ vdd gnd FILL
XFILL_0__1713_ vdd gnd FILL
XFILL_3__988_ vdd gnd FILL
X_1370_ _1370_/A _1370_/B _1370_/C _1521_/C vdd gnd AOI21X1
XFILL_0__1644_ vdd gnd FILL
XFILL_0__1575_ vdd gnd FILL
XFILL_3__1353_ vdd gnd FILL
XFILL_3__1422_ vdd gnd FILL
XFILL_3__1284_ vdd gnd FILL
XFILL93150x27450 vdd gnd FILL
X_1637_ ABCmd_i[3] _1783_/C vdd gnd INVX4
X_1706_ _1716_/A _1783_/C _1706_/C _1708_/B vdd gnd OAI21X1
XFILL_0__1009_ vdd gnd FILL
XFILL_1__1822_ vdd gnd FILL
XFILL_1__1684_ vdd gnd FILL
XFILL_1__1753_ vdd gnd FILL
X_1499_ _1499_/A _1500_/A vdd gnd INVX1
X_1568_ _1584_/C _1568_/B _1583_/C vdd gnd XOR2X1
XFILL_1__1049_ vdd gnd FILL
XFILL_3_BUFX2_insert2 vdd gnd FILL
XFILL_1__1118_ vdd gnd FILL
XFILL_2__1793_ vdd gnd FILL
XFILL_3__911_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
XFILL_2__1158_ vdd gnd FILL
XFILL_2__1227_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
X_1422_ _1422_/A _1422_/B _1522_/B vdd gnd NAND2X1
XFILL_2__1089_ vdd gnd FILL
XFILL_1_BUFX2_insert38 vdd gnd FILL
XFILL_1_BUFX2_insert27 vdd gnd FILL
XFILL_1_BUFX2_insert16 vdd gnd FILL
XFILL93150x39150 vdd gnd FILL
X_1353_ _1418_/A _1353_/B _1353_/C _1366_/B vdd gnd NAND3X1
XFILL_3__1405_ vdd gnd FILL
X_1284_ _1289_/B _1284_/B _1284_/C _1587_/A vdd gnd NAND3X1
XFILL_3__1336_ vdd gnd FILL
XFILL_0__1489_ vdd gnd FILL
XFILL_0__1558_ vdd gnd FILL
XFILL_3__1267_ vdd gnd FILL
XFILL_3__1198_ vdd gnd FILL
XFILL_1__1805_ vdd gnd FILL
XFILL_1__1667_ vdd gnd FILL
XFILL_1__1736_ vdd gnd FILL
XFILL_1__1598_ vdd gnd FILL
XFILL_2__989_ vdd gnd FILL
XFILL_2__1012_ vdd gnd FILL
XBUFX2_insert41 ABCmd_i[2] _1716_/A vdd gnd BUFX2
XBUFX2_insert30 _1613_/Q _939_/A vdd gnd BUFX2
X_995_ _995_/A _995_/B _995_/C _998_/C vdd gnd AOI21X1
XFILL_2__1776_ vdd gnd FILL
XFILL_0__1412_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_3__1121_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
XFILL_3__1052_ vdd gnd FILL
X_1405_ _1405_/A _1405_/B _1405_/C _1471_/C vdd gnd OAI21X1
X_1198_ _1198_/A _1198_/B _1198_/C _1200_/C vdd gnd OAI21X1
XFILL_1__1452_ vdd gnd FILL
X_1336_ _1375_/A _1375_/B _1405_/C _1417_/B vdd gnd NAND3X1
XFILL_1__1521_ vdd gnd FILL
X_1267_ _1351_/A _1267_/B _1267_/C _1269_/A vdd gnd NAND3X1
XFILL_2__912_ vdd gnd FILL
XFILL_3__1319_ vdd gnd FILL
XFILL_1__1383_ vdd gnd FILL
XFILL_2__1561_ vdd gnd FILL
XFILL_1__1719_ vdd gnd FILL
XFILL_2__1492_ vdd gnd FILL
XFILL_1__930_ vdd gnd FILL
XFILL_2__1759_ vdd gnd FILL
X_978_ _978_/A _978_/B _979_/C vdd gnd NAND2X1
X_1052_ _1052_/A _1052_/B _1052_/C _1074_/A vdd gnd NAND3X1
X_1121_ _1567_/B _1121_/B _1121_/C _1127_/B vdd gnd OAI21X1
XFILL_3__1035_ vdd gnd FILL
XFILL_3__1104_ vdd gnd FILL
XFILL_0__1326_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
XFILL_0__1257_ vdd gnd FILL
X_1319_ _1567_/A _953_/B _1319_/C _1323_/B vdd gnd OAI21X1
XFILL_1__1504_ vdd gnd FILL
XFILL_1__1435_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
XFILL_1__1366_ vdd gnd FILL
X_901_ _921_/C _901_/B LoadB_i _912_/B vdd gnd OAI21X1
XFILL_2__1544_ vdd gnd FILL
XFILL_2__1475_ vdd gnd FILL
X_1670_ _1677_/A _1670_/B _1670_/C _1690_/A vdd gnd AOI21X1
XFILL_0__1042_ vdd gnd FILL
XFILL_0__1111_ vdd gnd FILL
XFILL_1__913_ vdd gnd FILL
X_1035_ _1075_/A _1102_/C _1102_/B _1052_/B vdd gnd OAI21X1
X_1104_ _1104_/A _1104_/B _1104_/C _1246_/C vdd gnd NAND3X1
XFILL_1__1151_ vdd gnd FILL
XFILL_3__1018_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
XFILL_0__1309_ vdd gnd FILL
XFILL_1__1220_ vdd gnd FILL
X_1799_ _1799_/A _1799_/B _1813_/C vdd gnd NAND2X1
XFILL_0_BUFX2_insert40 vdd gnd FILL
XFILL_2__1191_ vdd gnd FILL
XFILL_0__931_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_1__1349_ vdd gnd FILL
XFILL_2__1260_ vdd gnd FILL
XFILL_0__1660_ vdd gnd FILL
XFILL_2__1527_ vdd gnd FILL
XFILL_0__1591_ vdd gnd FILL
XFILL_2__1458_ vdd gnd FILL
XFILL_2__1389_ vdd gnd FILL
X_1722_ _1722_/A _1722_/B _1722_/C _1723_/C vdd gnd NAND3X1
X_1653_ _1653_/A _1653_/B _1683_/A _1684_/A vdd gnd OAI21X1
XFILL_0__1025_ vdd gnd FILL
X_1584_ _1584_/A _1585_/A _1584_/C _1585_/B vdd gnd NAND3X1
XFILL_0__1789_ vdd gnd FILL
X_1018_ _955_/Y _1198_/B _1287_/A _1180_/C vdd gnd OAI21X1
XFILL_1__1203_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_1__1134_ vdd gnd FILL
XFILL_2__1312_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_0__914_ vdd gnd FILL
XFILL_2__1243_ vdd gnd FILL
XFILL_0__1712_ vdd gnd FILL
XFILL_0__1643_ vdd gnd FILL
XFILL_0__1574_ vdd gnd FILL
X_1705_ _1705_/A _1706_/C vdd gnd INVX1
X_1636_ _1677_/A _1676_/B vdd gnd INVX1
XFILL_0__1008_ vdd gnd FILL
XFILL_1__1821_ vdd gnd FILL
X_1567_ _1567_/A _1567_/B _1584_/A _1568_/B vdd gnd OAI21X1
XFILL_1__1683_ vdd gnd FILL
XFILL_1__1752_ vdd gnd FILL
XFILL92850x7950 vdd gnd FILL
X_1498_ _1542_/A _1498_/B _1498_/C _1501_/B vdd gnd OAI21X1
XFILL_1__1048_ vdd gnd FILL
XFILL_1__1117_ vdd gnd FILL
XFILL_2__1792_ vdd gnd FILL
XFILL_2__1157_ vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_2__1088_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
X_1421_ _1421_/A _1423_/C _1520_/A _1475_/C vdd gnd AOI21X1
XFILL_1_BUFX2_insert39 vdd gnd FILL
XFILL_1_BUFX2_insert28 vdd gnd FILL
XFILL_1_BUFX2_insert17 vdd gnd FILL
X_1283_ _1283_/A _922_/C _1535_/A _1358_/C vdd gnd OAI21X1
X_1352_ _1352_/A _1418_/C _1352_/C _1416_/B vdd gnd NAND3X1
XFILL_0__1488_ vdd gnd FILL
XFILL_0__1557_ vdd gnd FILL
XFILL_1__1804_ vdd gnd FILL
XFILL_1__1735_ vdd gnd FILL
X_1619_ _1619_/D vdd _1635_/R _1634_/CLK _1820_/A vdd gnd DFFSR
XFILL_1__1666_ vdd gnd FILL
XFILL_1__1597_ vdd gnd FILL
XFILL92550x85950 vdd gnd FILL
XFILL_2__1011_ vdd gnd FILL
XFILL_2__988_ vdd gnd FILL
XBUFX2_insert20 _925_/Y _1631_/R vdd gnd BUFX2
XBUFX2_insert31 _1613_/Q _977_/A vdd gnd BUFX2
X_994_ _994_/A _994_/B _994_/C _994_/Y vdd gnd NAND3X1
XFILL_2__1775_ vdd gnd FILL
XFILL_0__1273_ vdd gnd FILL
XFILL_0__1411_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_2__1209_ vdd gnd FILL
X_1404_ _1471_/A _1471_/B _1413_/C _1411_/C vdd gnd NAND3X1
X_1335_ _1342_/C _1341_/C _1375_/B vdd gnd NAND2X1
X_1197_ _1528_/A _1528_/C _1528_/B _1551_/C vdd gnd NOR3X1
XFILL_1__1451_ vdd gnd FILL
XFILL_1__1520_ vdd gnd FILL
XFILL_1__1382_ vdd gnd FILL
X_1266_ _1266_/A _1266_/B _1266_/C _1269_/C vdd gnd OAI21X1
XFILL_2__911_ vdd gnd FILL
XFILL92250x15750 vdd gnd FILL
XFILL92850x62550 vdd gnd FILL
XFILL_1__1718_ vdd gnd FILL
XFILL_2__1560_ vdd gnd FILL
XFILL_2__1491_ vdd gnd FILL
XFILL_1__1649_ vdd gnd FILL
X_977_ _977_/A _979_/B vdd gnd INVX2
XFILL_2__1758_ vdd gnd FILL
XFILL_2__1689_ vdd gnd FILL
X_1051_ _1108_/B _1074_/C _1074_/B _1068_/A vdd gnd OAI21X1
X_1120_ _1120_/A _1120_/B _1207_/A vdd gnd NAND2X1
XFILL_0__1325_ vdd gnd FILL
XFILL_0__1256_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
XFILL_3__1798_ vdd gnd FILL
XFILL_1__989_ vdd gnd FILL
X_1318_ _1760_/A _1567_/A vdd gnd INVX2
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
XFILL_1__1503_ vdd gnd FILL
X_1249_ _1338_/A _1342_/B _1298_/C _1258_/B vdd gnd OAI21X1
XFILL92250x27450 vdd gnd FILL
XFILL92850x74250 vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
X_900_ LoadCmd_i _924_/B _901_/B vdd gnd NOR2X1
XFILL_2__1474_ vdd gnd FILL
XFILL_2__1543_ vdd gnd FILL
XFILL_0__1110_ vdd gnd FILL
XFILL_3__1721_ vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_3__1652_ vdd gnd FILL
XFILL_1__912_ vdd gnd FILL
XFILL_3__1583_ vdd gnd FILL
X_1034_ _997_/A _996_/C _996_/B _1052_/C vdd gnd AOI21X1
X_1103_ _1103_/A _1103_/B _1103_/C _1220_/B vdd gnd NAND3X1
XFILL_1__1150_ vdd gnd FILL
XFILL_1__1081_ vdd gnd FILL
XFILL_0__1308_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
X_1798_ _1803_/A _1804_/A _1798_/C _1813_/A vdd gnd NAND3X1
XFILL_0_BUFX2_insert41 vdd gnd FILL
XFILL_0_BUFX2_insert30 vdd gnd FILL
XFILL_2__1190_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_1__1417_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
XFILL_2__1526_ vdd gnd FILL
XFILL_0__1590_ vdd gnd FILL
XFILL_2__1457_ vdd gnd FILL
X_1721_ _1721_/A _1721_/B _1723_/A vdd gnd NAND2X1
XFILL_2__1388_ vdd gnd FILL
X_1652_ _978_/B ABCmd_i[5] _1683_/A vdd gnd NAND2X1
XFILL_3__1704_ vdd gnd FILL
XFILL_0__1024_ vdd gnd FILL
X_1583_ _1583_/A _1583_/B _1583_/C _1586_/B vdd gnd AOI21X1
XFILL_0__1788_ vdd gnd FILL
XFILL_3__1566_ vdd gnd FILL
XFILL_3__1497_ vdd gnd FILL
X_1017_ _1017_/A _1017_/B _982_/Y _1198_/B vdd gnd AOI21X1
XFILL_1__1202_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_1__1133_ vdd gnd FILL
XFILL_2__1242_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_2__1173_ vdd gnd FILL
XFILL_0__913_ vdd gnd FILL
XFILL_0__1711_ vdd gnd FILL
XFILL_0__1642_ vdd gnd FILL
XFILL_3__986_ vdd gnd FILL
XFILL_3__1351_ vdd gnd FILL
XFILL_3__1420_ vdd gnd FILL
XFILL_0_BUFX2_insert0 vdd gnd FILL
XFILL_3__1282_ vdd gnd FILL
XFILL_2__1509_ vdd gnd FILL
XFILL_0__1573_ vdd gnd FILL
X_1704_ _1768_/A _1704_/Y vdd gnd INVX1
XFILL_0__1007_ vdd gnd FILL
XFILL_1__1751_ vdd gnd FILL
XFILL_1__1820_ vdd gnd FILL
X_1635_ _924_/Y vdd _1635_/R _1635_/CLK _898_/A vdd gnd DFFSR
X_1566_ _1566_/A _1566_/B _1566_/C _1584_/C vdd gnd OAI21X1
X_1497_ _1500_/B _1539_/C _1498_/C vdd gnd NAND2X1
XFILL_1__1682_ vdd gnd FILL
XFILL_1__1116_ vdd gnd FILL
XFILL_3_BUFX2_insert4 vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
XFILL_2__1791_ vdd gnd FILL
XFILL_2__1225_ vdd gnd FILL
XFILL_2__1156_ vdd gnd FILL
XFILL_2__1087_ vdd gnd FILL
XFILL_1_BUFX2_insert18 vdd gnd FILL
XFILL_1_BUFX2_insert29 vdd gnd FILL
X_1351_ _1351_/A _1351_/B _1367_/A _1366_/C vdd gnd OAI21X1
X_1420_ _1516_/B _1420_/B _1520_/A vdd gnd NAND2X1
XFILL_3__969_ vdd gnd FILL
X_1282_ _915_/A _911_/A ABCmd_i[7] _1535_/A vdd gnd OAI21X1
XFILL_3__1403_ vdd gnd FILL
XFILL_3__1334_ vdd gnd FILL
XFILL_3__1196_ vdd gnd FILL
XFILL_3__1265_ vdd gnd FILL
XFILL_0__1556_ vdd gnd FILL
XFILL_0__1487_ vdd gnd FILL
X_1618_ _1618_/D vdd _1624_/R _1634_/CLK _1819_/A vdd gnd DFFSR
XFILL_1__1803_ vdd gnd FILL
XFILL_1__1665_ vdd gnd FILL
XFILL_1__1734_ vdd gnd FILL
X_1549_ _1561_/A _1549_/B _1561_/B _1550_/C vdd gnd OAI21X1
XFILL_1__1596_ vdd gnd FILL
XFILL_2__987_ vdd gnd FILL
XFILL_2__1010_ vdd gnd FILL
XBUFX2_insert21 _925_/Y _1635_/R vdd gnd BUFX2
XBUFX2_insert32 _1613_/Q _1452_/B vdd gnd BUFX2
XFILL_2__1774_ vdd gnd FILL
X_993_ _996_/A _996_/B _997_/B _994_/B vdd gnd OAI21X1
XFILL_0__1410_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_3__1050_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
XFILL_2__1208_ vdd gnd FILL
XFILL_2__1139_ vdd gnd FILL
X_1403_ _1462_/C _1441_/B _1441_/A _1471_/B vdd gnd NAND3X1
X_1334_ _1341_/A _1400_/B _1334_/C _1405_/C vdd gnd NAND3X1
X_1265_ _1265_/A _1265_/B _1265_/C _1292_/B vdd gnd OAI21X1
X_1196_ _1196_/A _1196_/B _1196_/C _1528_/A vdd gnd AOI21X1
XFILL_2__910_ vdd gnd FILL
XFILL_0__1608_ vdd gnd FILL
XFILL_1__1450_ vdd gnd FILL
XFILL_1__1381_ vdd gnd FILL
XFILL_0__1539_ vdd gnd FILL
XFILL_3__1317_ vdd gnd FILL
XFILL_3__1179_ vdd gnd FILL
XFILL_3__1248_ vdd gnd FILL
XFILL_1__1648_ vdd gnd FILL
XFILL_1__1717_ vdd gnd FILL
XFILL_2__1490_ vdd gnd FILL
XFILL_1__1579_ vdd gnd FILL
XFILL_2__1757_ vdd gnd FILL
X_976_ _976_/A _978_/B _980_/A vdd gnd NAND2X1
XFILL_2__1826_ vdd gnd FILL
XFILL_2__1688_ vdd gnd FILL
X_1050_ _1054_/B _1054_/A _1074_/B vdd gnd AND2X2
XFILL_3__1102_ vdd gnd FILL
XFILL_0__1186_ vdd gnd FILL
XFILL_3__1033_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
XFILL_0__1255_ vdd gnd FILL
XFILL_1__988_ vdd gnd FILL
XFILL_1__1502_ vdd gnd FILL
X_1248_ _1248_/A _1248_/B _1330_/A _1342_/B vdd gnd AOI21X1
X_1317_ _1379_/C _1324_/B _1324_/A _1322_/C vdd gnd AOI21X1
X_1179_ _1287_/B _1528_/B _1179_/C _1551_/A vdd gnd NAND3X1
XFILL_1__1433_ vdd gnd FILL
XFILL_1__1364_ vdd gnd FILL
XFILL_1__1295_ vdd gnd FILL
XFILL_2__1473_ vdd gnd FILL
XFILL_2__1542_ vdd gnd FILL
XFILL_0__1040_ vdd gnd FILL
X_959_ _988_/A _978_/B _961_/A vdd gnd NAND2X1
XFILL_2__1809_ vdd gnd FILL
XFILL_1__911_ vdd gnd FILL
X_1102_ _1102_/A _1102_/B _1102_/C _1103_/C vdd gnd AOI21X1
X_1033_ _1053_/C _1088_/B _1053_/A _1108_/B vdd gnd AOI21X1
XFILL_0__1169_ vdd gnd FILL
XFILL_3__1016_ vdd gnd FILL
X_1797_ _1797_/A _1797_/B _1797_/Y vdd gnd AND2X2
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_0_BUFX2_insert20 vdd gnd FILL
XFILL_0_BUFX2_insert31 vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_2__1525_ vdd gnd FILL
XFILL_2__1387_ vdd gnd FILL
XFILL_2__1456_ vdd gnd FILL
X_1651_ _1802_/B _1651_/B _1653_/B vdd gnd NAND2X1
X_1720_ _1725_/B _1725_/A _1793_/A vdd gnd XNOR2X1
XFILL_0__989_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
X_1582_ _1825_/A _1592_/A vdd gnd INVX1
XFILL_0__1787_ vdd gnd FILL
X_1016_ _1017_/B _1017_/A _982_/Y _1287_/A vdd gnd NAND3X1
XFILL_1__1201_ vdd gnd FILL
XFILL_1__1132_ vdd gnd FILL
XFILL_1__1063_ vdd gnd FILL
XFILL_2__1241_ vdd gnd FILL
XFILL_2__1310_ vdd gnd FILL
XFILL_2__1172_ vdd gnd FILL
XFILL_0__912_ vdd gnd FILL
XFILL91950x62550 vdd gnd FILL
XFILL_0__1710_ vdd gnd FILL
XFILL_0__1641_ vdd gnd FILL
XFILL_2__1508_ vdd gnd FILL
XFILL_0__1572_ vdd gnd FILL
XFILL_0_BUFX2_insert1 vdd gnd FILL
XFILL_2__1439_ vdd gnd FILL
X_1703_ _1721_/B _1721_/A _1768_/A vdd gnd XOR2X1
XFILL_0__1006_ vdd gnd FILL
X_1634_ _919_/Y vdd _1635_/R _1634_/CLK _915_/A vdd gnd DFFSR
XFILL_1__1681_ vdd gnd FILL
XFILL_1__1750_ vdd gnd FILL
X_1565_ _1565_/A _1565_/B _1566_/C vdd gnd NAND2X1
X_1496_ _1496_/A _1542_/D _1496_/C _1500_/B vdd gnd OAI21X1
XFILL_3__1548_ vdd gnd FILL
XFILL_3__1479_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_2__1790_ vdd gnd FILL
XFILL_2__1155_ vdd gnd FILL
XFILL_2__1224_ vdd gnd FILL
XFILL91350x27450 vdd gnd FILL
XFILL_2__1086_ vdd gnd FILL
XFILL_1_BUFX2_insert19 vdd gnd FILL
X_1281_ _1808_/C _1283_/A vdd gnd INVX1
X_1350_ _1350_/A _1350_/B _1350_/C _1351_/B vdd gnd AOI21X1
XFILL_0__1555_ vdd gnd FILL
XFILL_0__1486_ vdd gnd FILL
XFILL_1__1802_ vdd gnd FILL
X_1617_ _1617_/D vdd _1635_/R _1634_/CLK _950_/A vdd gnd DFFSR
XFILL_1__1733_ vdd gnd FILL
XFILL_1__1664_ vdd gnd FILL
X_1548_ _1548_/A _1548_/B _1548_/C _1550_/B vdd gnd OAI21X1
X_1479_ _1479_/A _1479_/B _1479_/C _1486_/C vdd gnd OAI21X1
XFILL_1__1595_ vdd gnd FILL
XFILL_2__986_ vdd gnd FILL
XBUFX2_insert33 _1613_/Q _976_/A vdd gnd BUFX2
XBUFX2_insert22 _1630_/Q _1491_/A vdd gnd BUFX2
XFILL_1__1029_ vdd gnd FILL
XFILL_2__1773_ vdd gnd FILL
X_992_ _992_/A _992_/B _996_/B vdd gnd NOR2X1
XFILL_0__1340_ vdd gnd FILL
XFILL_2__1207_ vdd gnd FILL
XFILL_2__1138_ vdd gnd FILL
XFILL_0__1271_ vdd gnd FILL
XFILL_2__1069_ vdd gnd FILL
X_1402_ _1408_/B _1402_/B _1462_/C vdd gnd NAND2X1
X_1333_ _1373_/B _1373_/A _1375_/A vdd gnd XOR2X1
X_1264_ _1267_/C _1267_/B _1351_/A _1265_/B vdd gnd AOI21X1
XFILL93150x11850 vdd gnd FILL
X_1195_ _1430_/B _1480_/A _1480_/B _1528_/C vdd gnd NAND3X1
XFILL_0__1607_ vdd gnd FILL
XFILL_0__1469_ vdd gnd FILL
XFILL_0__1538_ vdd gnd FILL
XFILL_1__1380_ vdd gnd FILL
XFILL_1__1716_ vdd gnd FILL
XFILL_1__1647_ vdd gnd FILL
XFILL_1__1578_ vdd gnd FILL
XFILL_2__969_ vdd gnd FILL
XFILL_2_CLKBUF1_insert8 vdd gnd FILL
XFILL_2__1687_ vdd gnd FILL
XFILL_2__1756_ vdd gnd FILL
X_975_ _975_/A _980_/B vdd gnd INVX1
XFILL_2__1825_ vdd gnd FILL
XFILL_0__1323_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
XFILL_0__1254_ vdd gnd FILL
XFILL93150x23550 vdd gnd FILL
XFILL_3__1796_ vdd gnd FILL
XFILL_1__987_ vdd gnd FILL
X_1178_ _1198_/A _1198_/B _955_/Y _1179_/C vdd gnd OAI21X1
XFILL_1__1432_ vdd gnd FILL
X_1316_ _1379_/B _1324_/B vdd gnd INVX1
X_1247_ _1247_/A _1247_/B _1308_/B _1330_/C _1338_/A vdd gnd AOI22X1
XFILL_1__1501_ vdd gnd FILL
XFILL_1__1363_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
XFILL_2__1541_ vdd gnd FILL
XFILL_2__1472_ vdd gnd FILL
XFILL_3__1650_ vdd gnd FILL
XFILL_1__910_ vdd gnd FILL
X_958_ _960_/A _960_/B _961_/C vdd gnd OR2X2
XFILL_2__1808_ vdd gnd FILL
XFILL_2__1739_ vdd gnd FILL
X_889_ _898_/A _904_/C vdd gnd INVX1
X_1032_ _1075_/A _1102_/C _1075_/B _1053_/C vdd gnd OAI21X1
X_1101_ _1220_/C _1246_/B _1220_/A _1126_/A vdd gnd OAI21X1
XFILL_3__1581_ vdd gnd FILL
XFILL93150x35250 vdd gnd FILL
XFILL_0__1306_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
X_1796_ _1808_/B _1808_/C _1797_/A vdd gnd NOR2X1
XFILL_0__1237_ vdd gnd FILL
XFILL_0__1099_ vdd gnd FILL
XFILL_0_BUFX2_insert21 vdd gnd FILL
XFILL_0_BUFX2_insert32 vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_2__1524_ vdd gnd FILL
XFILL_2__1455_ vdd gnd FILL
XFILL_2__1386_ vdd gnd FILL
X_1650_ ABCmd_i[0] _1678_/B _1802_/A _1651_/B vdd gnd OAI21X1
XFILL_0__988_ vdd gnd FILL
XFILL_0__1022_ vdd gnd FILL
X_1581_ _1581_/A _911_/A _1581_/C _1581_/D _1623_/D vdd gnd AOI22X1
XFILL_3__1702_ vdd gnd FILL
XFILL_0__1786_ vdd gnd FILL
X_1015_ _1153_/A _1153_/B _1154_/A _1017_/A vdd gnd OAI21X1
XFILL_3__1564_ vdd gnd FILL
XFILL_3__1495_ vdd gnd FILL
XFILL_1__1200_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
X_1779_ _1781_/A _1781_/B _1780_/C vdd gnd NAND2X1
XFILL_2__1171_ vdd gnd FILL
XFILL_2__1240_ vdd gnd FILL
XFILL_0__911_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_3__984_ vdd gnd FILL
XFILL_0__1640_ vdd gnd FILL
XFILL_0_BUFX2_insert2 vdd gnd FILL
XFILL_3__1280_ vdd gnd FILL
XFILL_2__1507_ vdd gnd FILL
XFILL_2__1438_ vdd gnd FILL
XFILL_0__1571_ vdd gnd FILL
XFILL_2__1369_ vdd gnd FILL
X_1702_ _1708_/A _1705_/A _1702_/C _1721_/A vdd gnd OAI21X1
XFILL_0__1005_ vdd gnd FILL
X_1633_ _912_/Y _1635_/R vdd _1634_/CLK _904_/B vdd gnd DFFSR
X_1564_ _1564_/A _1565_/B vdd gnd INVX1
XFILL_1__1680_ vdd gnd FILL
X_1495_ _948_/A _1542_/D vdd gnd INVX1
XFILL_0__1769_ vdd gnd FILL
XFILL_3_BUFX2_insert6 vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
XFILL_2__1223_ vdd gnd FILL
XFILL_2__1085_ vdd gnd FILL
XFILL_3__967_ vdd gnd FILL
XFILL_3__898_ vdd gnd FILL
X_1280_ _1819_/A _1364_/A vdd gnd INVX1
XFILL_3__1401_ vdd gnd FILL
XFILL_3__1194_ vdd gnd FILL
XFILL_0__1554_ vdd gnd FILL
XFILL_3__1332_ vdd gnd FILL
XFILL_3__1263_ vdd gnd FILL
XFILL_0__1485_ vdd gnd FILL
XFILL_1__1801_ vdd gnd FILL
X_1616_ _949_/Y vdd _1632_/R _1635_/CLK _948_/A vdd gnd DFFSR
X_1547_ _1561_/A _1561_/B _1548_/C vdd gnd NOR2X1
XFILL_1__1663_ vdd gnd FILL
XFILL_1__1732_ vdd gnd FILL
XFILL_1__1594_ vdd gnd FILL
X_1478_ _1478_/A _1478_/B ABCmd_i[7] _1479_/B vdd gnd OAI21X1
XFILL_2__985_ vdd gnd FILL
XBUFX2_insert34 _1610_/Q _1670_/B vdd gnd BUFX2
XFILL_1__1028_ vdd gnd FILL
XBUFX2_insert23 _1630_/Q _1303_/A vdd gnd BUFX2
XFILL_2__1772_ vdd gnd FILL
X_991_ _991_/A _991_/B _992_/B vdd gnd NAND2X1
XFILL_2__1068_ vdd gnd FILL
XFILL_0__1270_ vdd gnd FILL
XFILL_2__1206_ vdd gnd FILL
XFILL_2__1137_ vdd gnd FILL
X_1401_ _1408_/A _1402_/B vdd gnd INVX1
X_1194_ _1194_/A _1194_/B _980_/B _1480_/B vdd gnd OAI21X1
XFILL_0__1606_ vdd gnd FILL
X_1332_ _1405_/B _1375_/C _1405_/A _1417_/A vdd gnd OAI21X1
X_1263_ _1263_/A _1263_/B _1350_/C _1267_/B vdd gnd OAI21X1
XFILL_3__1177_ vdd gnd FILL
XFILL_3__1246_ vdd gnd FILL
XFILL_3__1315_ vdd gnd FILL
XFILL_0__1468_ vdd gnd FILL
XFILL_0__1537_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL_1__1715_ vdd gnd FILL
XFILL_1__1646_ vdd gnd FILL
XFILL_1__1577_ vdd gnd FILL
XFILL_2__968_ vdd gnd FILL
XFILL_2_CLKBUF1_insert9 vdd gnd FILL
XFILL_2__899_ vdd gnd FILL
XCLKBUF1_insert8 clk _1628_/CLK vdd gnd CLKBUF1
XFILL_2__1824_ vdd gnd FILL
X_974_ _981_/B _981_/C _981_/A _982_/C vdd gnd NAND3X1
XFILL_2__1686_ vdd gnd FILL
XFILL_2__1755_ vdd gnd FILL
XFILL_3__1031_ vdd gnd FILL
XFILL_3__1100_ vdd gnd FILL
XFILL_0__1322_ vdd gnd FILL
XFILL_0__1184_ vdd gnd FILL
XFILL_0__1253_ vdd gnd FILL
XFILL_1__986_ vdd gnd FILL
X_1315_ _1760_/A _952_/A _1491_/A _1452_/B _1379_/B vdd gnd AOI22X1
X_1177_ _982_/C _1196_/B _1177_/C _1177_/D _1198_/A vdd gnd AOI22X1
XFILL_1__1362_ vdd gnd FILL
XFILL_1__1431_ vdd gnd FILL
X_1246_ _1246_/A _1246_/B _1246_/C _1298_/C vdd gnd OAI21X1
XFILL_1__1500_ vdd gnd FILL
XFILL_1__1293_ vdd gnd FILL
XFILL_2__1471_ vdd gnd FILL
XFILL_2__1540_ vdd gnd FILL
X_957_ _967_/A _988_/B _960_/B vdd gnd NAND2X1
XFILL_2__1807_ vdd gnd FILL
XFILL_2__1669_ vdd gnd FILL
XFILL_2__1738_ vdd gnd FILL
X_1031_ _984_/A _1760_/A _1082_/A _991_/B _1075_/A vdd gnd AOI22X1
X_1100_ _1105_/B _1105_/A _1220_/A vdd gnd AND2X2
XFILL_3__1014_ vdd gnd FILL
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1236_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
X_1795_ _1795_/A _1795_/B _1795_/C _1808_/B vdd gnd NAND3X1
XFILL_0__1098_ vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_3__1778_ vdd gnd FILL
XFILL_0_BUFX2_insert33 vdd gnd FILL
XFILL_0_BUFX2_insert22 vdd gnd FILL
X_1229_ _1303_/A _1302_/A _977_/A _986_/D _1304_/D vdd gnd AOI22X1
XFILL_1__1345_ vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
XFILL_1__1276_ vdd gnd FILL
XFILL_2__1454_ vdd gnd FILL
XFILL_2__1523_ vdd gnd FILL
XFILL_2__1385_ vdd gnd FILL
XFILL_0__987_ vdd gnd FILL
X_1580_ _1580_/A _1580_/B _911_/A _1581_/D vdd gnd AOI21X1
XFILL_0__1021_ vdd gnd FILL
XFILL_0__1785_ vdd gnd FILL
X_1014_ _1063_/C _1014_/B _1154_/A vdd gnd NAND2X1
XFILL_1__1061_ vdd gnd FILL
XFILL_0__1219_ vdd gnd FILL
XFILL_1__1130_ vdd gnd FILL
X_1778_ _1778_/A _948_/A _1781_/B vdd gnd AND2X2
XFILL92250x11850 vdd gnd FILL
XFILL_2__1170_ vdd gnd FILL
XFILL_0__910_ vdd gnd FILL
XFILL_1__1328_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL_0_BUFX2_insert3 vdd gnd FILL
XFILL_2__1437_ vdd gnd FILL
XFILL_2__1506_ vdd gnd FILL
XFILL_0__1570_ vdd gnd FILL
X_1701_ _1809_/B _1705_/A _1708_/A _1702_/C vdd gnd OAI21X1
XFILL_2__1299_ vdd gnd FILL
XFILL_2__1368_ vdd gnd FILL
XFILL_0__1004_ vdd gnd FILL
X_1632_ _1632_/D vdd _1632_/R _1635_/CLK _1781_/A vdd gnd DFFSR
X_1563_ _1572_/A _1583_/B vdd gnd INVX1
X_1494_ _1496_/C _1494_/B _1539_/C vdd gnd OR2X2
XFILL_0__1768_ vdd gnd FILL
XFILL_0__1699_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL92850x70350 vdd gnd FILL
XFILL_2__1222_ vdd gnd FILL
XFILL_2__1153_ vdd gnd FILL
XFILL_2__1084_ vdd gnd FILL
XFILL_0__1484_ vdd gnd FILL
XFILL_0__1553_ vdd gnd FILL
XFILL_1__1800_ vdd gnd FILL
XFILL_1__1731_ vdd gnd FILL
X_1615_ _946_/Y vdd _1631_/R _1631_/CLK _945_/A vdd gnd DFFSR
X_1546_ _1562_/A _1562_/B _1561_/B vdd gnd XOR2X1
X_1477_ _1520_/B _1478_/A vdd gnd INVX1
XFILL_1__1662_ vdd gnd FILL
XFILL_3__1529_ vdd gnd FILL
XFILL_1__1593_ vdd gnd FILL
XBUFX2_insert24 _1630_/Q _991_/B vdd gnd BUFX2
XBUFX2_insert13 _896_/Y _1601_/B vdd gnd BUFX2
XFILL_2__984_ vdd gnd FILL
XFILL92250x35250 vdd gnd FILL
XFILL92850x82050 vdd gnd FILL
X_990_ _997_/A _996_/C _997_/C _994_/A vdd gnd NAND3X1
XBUFX2_insert35 _1610_/Q _991_/A vdd gnd BUFX2
XFILL_1__1027_ vdd gnd FILL
XFILL_2__1771_ vdd gnd FILL
XFILL_2__1205_ vdd gnd FILL
XFILL_2__1067_ vdd gnd FILL
XFILL_2__1136_ vdd gnd FILL
X_1400_ _1400_/A _1400_/B _1408_/B vdd gnd NAND2X1
X_1331_ _1341_/A _1400_/B _1334_/C _1405_/B vdd gnd AOI21X1
X_1193_ _1193_/A _1194_/B vdd gnd INVX1
XFILL_0__1605_ vdd gnd FILL
X_1262_ _1350_/A _1350_/B _1262_/C _1267_/C vdd gnd NAND3X1
XFILL_0__1398_ vdd gnd FILL
XFILL_0__1467_ vdd gnd FILL
XFILL_0__1536_ vdd gnd FILL
XFILL_1__1645_ vdd gnd FILL
XFILL_1__1714_ vdd gnd FILL
X_1529_ _1529_/A _1529_/B _1531_/B vdd gnd NAND2X1
XFILL_1__1576_ vdd gnd FILL
XFILL_2__967_ vdd gnd FILL
XFILL_2__898_ vdd gnd FILL
X_973_ _995_/C _983_/B _983_/A _981_/B vdd gnd OAI21X1
XFILL_2__1754_ vdd gnd FILL
XCLKBUF1_insert9 clk _1635_/CLK vdd gnd CLKBUF1
XFILL_2__1823_ vdd gnd FILL
XFILL_2__1685_ vdd gnd FILL
XFILL_0__1321_ vdd gnd FILL
XFILL_0__1252_ vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
XFILL_2__1119_ vdd gnd FILL
XFILL_3__1794_ vdd gnd FILL
XFILL_1__985_ vdd gnd FILL
X_1314_ _1319_/C _1320_/C _1379_/C vdd gnd NAND2X1
X_1176_ _1200_/A _1528_/B vdd gnd INVX1
XFILL_1__1430_ vdd gnd FILL
XFILL_1__1361_ vdd gnd FILL
XFILL_0__1519_ vdd gnd FILL
X_1245_ _1298_/A _1298_/B _1338_/C _1258_/A vdd gnd NAND3X1
XFILL_1__1292_ vdd gnd FILL
XFILL_2__1470_ vdd gnd FILL
XFILL_1__1559_ vdd gnd FILL
XFILL_2__1806_ vdd gnd FILL
X_956_ _964_/A _962_/B _960_/A vdd gnd NAND2X1
XFILL_2__1737_ vdd gnd FILL
XFILL_2__1668_ vdd gnd FILL
XFILL_2__1599_ vdd gnd FILL
X_1030_ _992_/B _1083_/A _1102_/C vdd gnd NOR2X1
XFILL_0__1166_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
XFILL_0__1304_ vdd gnd FILL
X_1794_ _1794_/A _1794_/B _1797_/B vdd gnd NOR2X1
XFILL_0__1097_ vdd gnd FILL
XFILL_0_BUFX2_insert34 vdd gnd FILL
XFILL_1__899_ vdd gnd FILL
XFILL_0_BUFX2_insert23 vdd gnd FILL
XFILL_1__968_ vdd gnd FILL
X_1228_ _1228_/A _1228_/B _1231_/C vdd gnd NAND2X1
X_1159_ _1287_/A _1287_/B _1159_/C _1159_/D _1203_/A vdd gnd AOI22X1
XFILL_1__1275_ vdd gnd FILL
XFILL_1__1344_ vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
XFILL_2__1453_ vdd gnd FILL
XFILL_2__1522_ vdd gnd FILL
XFILL_2__1384_ vdd gnd FILL
XFILL_0__1020_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
XFILL_3__1700_ vdd gnd FILL
XFILL_0__1784_ vdd gnd FILL
X_939_ _939_/A _940_/B _940_/C vdd gnd NAND2X1
XFILL_3__1562_ vdd gnd FILL
XFILL_3__1493_ vdd gnd FILL
X_1013_ _994_/B _994_/A _994_/C _1153_/B vdd gnd AOI21X1
XFILL_0__1149_ vdd gnd FILL
X_1777_ ABCmd_i[5] ABCmd_i[4] _1782_/C vdd gnd NAND2X1
XFILL_1__1060_ vdd gnd FILL
XFILL_0__1218_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
XFILL_3__982_ vdd gnd FILL
XFILL_2__1436_ vdd gnd FILL
XFILL_0_BUFX2_insert4 vdd gnd FILL
XFILL_2__1505_ vdd gnd FILL
XFILL_2__1367_ vdd gnd FILL
XFILL_0__969_ vdd gnd FILL
X_1700_ _932_/A _988_/A _1700_/C _1705_/A vdd gnd AOI21X1
X_1631_ _1631_/D vdd _1631_/R _1631_/CLK _1760_/A vdd gnd DFFSR
XFILL_0__1003_ vdd gnd FILL
XFILL_2__1298_ vdd gnd FILL
X_1562_ _1562_/A _1562_/B _1562_/C _1572_/A vdd gnd OAI21X1
X_1493_ _1567_/B _1539_/B _1493_/C _1496_/C vdd gnd OAI21X1
XFILL_0__1698_ vdd gnd FILL
XFILL_0__1767_ vdd gnd FILL
XFILL_3__1545_ vdd gnd FILL
XFILL_3__1476_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
XFILL_1__1043_ vdd gnd FILL
XFILL92850x89850 vdd gnd FILL
XFILL_2__1221_ vdd gnd FILL
XFILL_2__1152_ vdd gnd FILL
XFILL_2__1083_ vdd gnd FILL
XFILL_3__965_ vdd gnd FILL
XFILL_0__1552_ vdd gnd FILL
XFILL_3__896_ vdd gnd FILL
XFILL_3__1330_ vdd gnd FILL
XFILL_3__1192_ vdd gnd FILL
XFILL_0__1483_ vdd gnd FILL
XFILL_2__1419_ vdd gnd FILL
XFILL_3__1261_ vdd gnd FILL
X_1614_ _943_/Y vdd _1631_/R _1628_/CLK _999_/B vdd gnd DFFSR
XFILL_1__1661_ vdd gnd FILL
XFILL_1__1730_ vdd gnd FILL
X_1545_ _1564_/A _1565_/A _1562_/B vdd gnd XOR2X1
X_1476_ _1476_/A _1476_/B _1476_/C _1478_/B vdd gnd AOI21X1
XFILL_0__1819_ vdd gnd FILL
XFILL_1__1592_ vdd gnd FILL
XFILL_2__983_ vdd gnd FILL
XBUFX2_insert36 _1610_/Q _964_/A vdd gnd BUFX2
XBUFX2_insert25 _1630_/Q _1746_/A vdd gnd BUFX2
XBUFX2_insert14 _896_/Y _1604_/B vdd gnd BUFX2
XFILL92550x19650 vdd gnd FILL
XFILL_2__1770_ vdd gnd FILL
XFILL_1__1026_ vdd gnd FILL
XFILL_2__1204_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
XFILL_2__1066_ vdd gnd FILL
XFILL_3__948_ vdd gnd FILL
X_1330_ _1330_/A _1330_/B _1330_/C _1334_/C vdd gnd OAI21X1
X_1261_ _1295_/A _1351_/A vdd gnd INVX1
X_1192_ _1481_/A _1430_/B vdd gnd INVX1
XFILL_0__1604_ vdd gnd FILL
XFILL_3__1313_ vdd gnd FILL
XFILL_0__1535_ vdd gnd FILL
XFILL_3__1244_ vdd gnd FILL
XFILL_3__1175_ vdd gnd FILL
XFILL_0__1397_ vdd gnd FILL
XFILL_0__1466_ vdd gnd FILL
XFILL_1__1644_ vdd gnd FILL
XFILL_1__1713_ vdd gnd FILL
X_1528_ _1528_/A _1528_/B _1528_/C _1529_/A vdd gnd OAI21X1
X_1459_ _1467_/A _1466_/B vdd gnd INVX1
XFILL_1__1575_ vdd gnd FILL
XFILL_2__966_ vdd gnd FILL
XFILL_2__897_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
XFILL_2__1753_ vdd gnd FILL
X_972_ _972_/A _992_/A _983_/B vdd gnd AND2X2
XFILL_2__1822_ vdd gnd FILL
XFILL91350x11850 vdd gnd FILL
XFILL_2__1684_ vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_0__1320_ vdd gnd FILL
XFILL_0__1251_ vdd gnd FILL
XFILL_2__1118_ vdd gnd FILL
XFILL_2__1049_ vdd gnd FILL
XFILL_1__984_ vdd gnd FILL
X_1313_ _1760_/A _952_/A _1320_/C vdd gnd AND2X2
X_1244_ _1330_/C _1308_/B _1308_/A _1298_/B vdd gnd NAND3X1
X_1175_ _1196_/B _1196_/C _1196_/A _1200_/A vdd gnd NAND3X1
XFILL_1__1360_ vdd gnd FILL
XFILL_0__1518_ vdd gnd FILL
XFILL_3__1227_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
XFILL_3__1158_ vdd gnd FILL
XFILL_0__1449_ vdd gnd FILL
XFILL_3__1089_ vdd gnd FILL
XFILL_1__1558_ vdd gnd FILL
XFILL_2__949_ vdd gnd FILL
XFILL_1__1489_ vdd gnd FILL
XFILL_2__1805_ vdd gnd FILL
XFILL_2__1667_ vdd gnd FILL
XFILL_2__1736_ vdd gnd FILL
XFILL91950x70350 vdd gnd FILL
X_955_ _955_/A _975_/A _955_/Y vdd gnd NAND2X1
XFILL_2__1598_ vdd gnd FILL
XFILL_0__1303_ vdd gnd FILL
X_1793_ _1793_/A _1793_/B _1794_/A vdd gnd NAND2X1
XFILL_3__1012_ vdd gnd FILL
XFILL_0__1165_ vdd gnd FILL
XFILL_0__1234_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
XFILL_1__967_ vdd gnd FILL
X_1158_ _1158_/A _1158_/B _1158_/C _1159_/D vdd gnd NAND3X1
XFILL_0_BUFX2_insert35 vdd gnd FILL
XFILL_0_BUFX2_insert24 vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
XFILL_1__898_ vdd gnd FILL
XFILL_1__1412_ vdd gnd FILL
X_1227_ _1304_/C _1231_/A vdd gnd INVX1
XFILL_1__1274_ vdd gnd FILL
XFILL_1__1343_ vdd gnd FILL
X_1089_ _999_/B _962_/B _1212_/A vdd gnd NAND2X1
XFILL_2__1521_ vdd gnd FILL
XFILL_2__1452_ vdd gnd FILL
XFILL_2__1383_ vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
XFILL91950x82050 vdd gnd FILL
XFILL_0__1783_ vdd gnd FILL
XFILL_2__1719_ vdd gnd FILL
X_1012_ _998_/B _998_/A _998_/C _1153_/A vdd gnd AOI21X1
X_938_ ABCmd_i[4] _940_/A vdd gnd INVX1
XFILL_0__1148_ vdd gnd FILL
X_1776_ _1804_/B _1776_/B _1803_/A _1799_/B vdd gnd OAI21X1
XFILL_0__1079_ vdd gnd FILL
XFILL_0__1217_ vdd gnd FILL
XFILL_3__1759_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_2__1504_ vdd gnd FILL
XFILL_0_BUFX2_insert5 vdd gnd FILL
XFILL_2__1297_ vdd gnd FILL
XFILL_2__1366_ vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_0__1002_ vdd gnd FILL
XFILL_0__899_ vdd gnd FILL
XFILL_0__968_ vdd gnd FILL
X_1630_ _1630_/D vdd _1632_/R _1635_/CLK _1630_/Q vdd gnd DFFSR
X_1561_ _1561_/A _1561_/B _1562_/C vdd gnd NAND2X1
X_1492_ _1567_/A _1567_/B _1539_/B _1493_/C vdd gnd OAI21X1
XFILL_0__1697_ vdd gnd FILL
XFILL_0__1766_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
X_1759_ _1780_/A _945_/A _1759_/C _1780_/D _1761_/D vdd gnd AOI22X1
XFILL_2__1151_ vdd gnd FILL
XFILL_2__1220_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_0__1551_ vdd gnd FILL
XFILL_0__1482_ vdd gnd FILL
XFILL_2__1418_ vdd gnd FILL
XFILL_2__1349_ vdd gnd FILL
X_1613_ _940_/Y vdd _1628_/R _1635_/CLK _1613_/Q vdd gnd DFFSR
XFILL93150x31350 vdd gnd FILL
X_1544_ _1566_/A _1566_/B _1564_/A vdd gnd XNOR2X1
XFILL_1__1660_ vdd gnd FILL
XFILL_3__1527_ vdd gnd FILL
XFILL_0__1818_ vdd gnd FILL
XFILL_1__1591_ vdd gnd FILL
X_1475_ _1476_/C _1520_/B _1475_/C _1479_/A vdd gnd NOR3X1
XFILL_2__982_ vdd gnd FILL
XFILL_0__1749_ vdd gnd FILL
XFILL_3__1389_ vdd gnd FILL
XFILL_3__1458_ vdd gnd FILL
XBUFX2_insert26 _915_/Y _943_/B vdd gnd BUFX2
XBUFX2_insert15 _896_/Y _1606_/B vdd gnd BUFX2
XFILL_1__1025_ vdd gnd FILL
XBUFX2_insert37 _1610_/Q _1082_/A vdd gnd BUFX2
XFILL_1__1789_ vdd gnd FILL
XFILL_2__1203_ vdd gnd FILL
XFILL_2__1134_ vdd gnd FILL
XFILL_2__1065_ vdd gnd FILL
X_1191_ _1429_/C _1429_/B _1429_/A _1481_/A vdd gnd NAND3X1
X_1260_ _1367_/A _1295_/B _1295_/A _1265_/A vdd gnd AOI21X1
XFILL_0__1603_ vdd gnd FILL
XFILL_0__1465_ vdd gnd FILL
XFILL_0__1534_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ _1551_/C _1529_/B vdd gnd INVX1
XFILL_1__1643_ vdd gnd FILL
XFILL_1__1712_ vdd gnd FILL
XFILL_1__1574_ vdd gnd FILL
X_1389_ _1760_/A _952_/A _1445_/A vdd gnd NAND2X1
X_1458_ _1460_/C _1460_/B _1460_/A _1467_/A vdd gnd AOI21X1
XFILL_2__965_ vdd gnd FILL
XFILL_2__896_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
XFILL_2__1683_ vdd gnd FILL
X_971_ _972_/A _992_/A _995_/C vdd gnd NOR2X1
XFILL_2__1752_ vdd gnd FILL
XFILL_2__1821_ vdd gnd FILL
XFILL_0__1181_ vdd gnd FILL
XFILL_2__1048_ vdd gnd FILL
XFILL_0__1250_ vdd gnd FILL
XFILL_2__1117_ vdd gnd FILL
XFILL_3__1792_ vdd gnd FILL
XFILL_1__983_ vdd gnd FILL
X_1174_ _1174_/A _982_/B _982_/A _1196_/A vdd gnd OAI21X1
X_1312_ _1491_/A _1452_/B _1319_/C vdd gnd AND2X2
X_1243_ _1307_/A _1307_/B _1308_/B vdd gnd NAND2X1
XFILL_1__1290_ vdd gnd FILL
XFILL_0__1448_ vdd gnd FILL
XFILL_0__1517_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_1__1557_ vdd gnd FILL
XFILL_2__948_ vdd gnd FILL
XFILL_1__1488_ vdd gnd FILL
XFILL_2__1804_ vdd gnd FILL
XFILL_2__1666_ vdd gnd FILL
XFILL_2__1735_ vdd gnd FILL
XFILL_2__1597_ vdd gnd FILL
X_954_ _976_/A _978_/B _955_/A vdd gnd AND2X2
XFILL91950x89850 vdd gnd FILL
XFILL_0__1302_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
X_1792_ _1792_/A _1792_/B _1793_/B vdd gnd NOR2X1
XFILL_2_CLKBUF1_insert10 vdd gnd FILL
XFILL_0__1233_ vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_3__1775_ vdd gnd FILL
XFILL_0_BUFX2_insert36 vdd gnd FILL
XFILL_1__897_ vdd gnd FILL
X_1157_ _1157_/A _1157_/B _1157_/C _1159_/C vdd gnd OAI21X1
XFILL_0_BUFX2_insert25 vdd gnd FILL
XFILL_0_BUFX2_insert14 vdd gnd FILL
X_1226_ _1304_/C _1226_/B _1226_/C _1247_/A vdd gnd NAND3X1
XFILL_1__1411_ vdd gnd FILL
XFILL_1__1342_ vdd gnd FILL
XFILL_1__1273_ vdd gnd FILL
X_1088_ _1088_/A _1088_/B _1103_/B _1103_/A _1220_/C vdd gnd AOI22X1
XFILL_3__1209_ vdd gnd FILL
XFILL_2__1451_ vdd gnd FILL
XFILL_2__1520_ vdd gnd FILL
XFILL_2__1382_ vdd gnd FILL
XFILL91650x19650 vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_3__1560_ vdd gnd FILL
XFILL_2__1649_ vdd gnd FILL
XFILL_0__1782_ vdd gnd FILL
XFILL_2__1718_ vdd gnd FILL
X_1011_ _994_/Y _998_/Y _1153_/C _1017_/B vdd gnd NAND3X1
X_937_ _937_/A _940_/B _937_/C _937_/Y vdd gnd OAI21X1
XFILL_3__1491_ vdd gnd FILL
XFILL_0__1216_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
X_1775_ _1795_/B _1795_/C _1775_/Y vdd gnd NAND2X1
XFILL_0__1078_ vdd gnd FILL
XFILL_1__949_ vdd gnd FILL
XFILL_1__1325_ vdd gnd FILL
X_1209_ _948_/A _978_/B _1296_/A vdd gnd NAND2X1
XFILL_1__1187_ vdd gnd FILL
XFILL_1__1256_ vdd gnd FILL
XFILL_3__980_ vdd gnd FILL
XFILL_2__1434_ vdd gnd FILL
XFILL_2__1503_ vdd gnd FILL
XFILL_0_BUFX2_insert6 vdd gnd FILL
XFILL_2__1365_ vdd gnd FILL
XFILL_2__1296_ vdd gnd FILL
XFILL_0__967_ vdd gnd FILL
XFILL_0__898_ vdd gnd FILL
XFILL_0__1001_ vdd gnd FILL
X_1560_ _1560_/A _1560_/B _1560_/C _1583_/A vdd gnd NAND3X1
XFILL_0__1765_ vdd gnd FILL
XFILL_3__1543_ vdd gnd FILL
X_1491_ _1491_/A _948_/A _1494_/B vdd gnd NAND2X1
XFILL_0__1696_ vdd gnd FILL
XFILL_3__1474_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
XFILL_1__1110_ vdd gnd FILL
X_1758_ _1760_/A _1760_/B _1759_/C vdd gnd NAND2X1
X_1689_ _1768_/B _1689_/Y vdd gnd INVX1
XFILL_2__1150_ vdd gnd FILL
XFILL_2__1081_ vdd gnd FILL
XFILL_1__1308_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_3__963_ vdd gnd FILL
XFILL_3__894_ vdd gnd FILL
XFILL_0__1481_ vdd gnd FILL
XFILL_3__1190_ vdd gnd FILL
XFILL_2__1417_ vdd gnd FILL
XFILL_0__1550_ vdd gnd FILL
XFILL_2__1279_ vdd gnd FILL
XFILL_2__1348_ vdd gnd FILL
X_1612_ _937_/Y vdd _1628_/R _1628_/CLK _1612_/Q vdd gnd DFFSR
X_1474_ _1516_/A _1521_/A _1520_/B vdd gnd NAND2X1
X_1543_ _1543_/A _1585_/A _1566_/B vdd gnd NAND2X1
XFILL_0__1817_ vdd gnd FILL
XFILL_0__1748_ vdd gnd FILL
XFILL_1__1590_ vdd gnd FILL
XFILL_2__981_ vdd gnd FILL
XFILL_0__1679_ vdd gnd FILL
XBUFX2_insert38 ABCmd_i[2] _932_/A vdd gnd BUFX2
XBUFX2_insert27 _915_/Y _949_/B vdd gnd BUFX2
XBUFX2_insert16 _896_/Y _918_/C vdd gnd BUFX2
XFILL_1__1024_ vdd gnd FILL
XFILL_1__1788_ vdd gnd FILL
XFILL_2__1202_ vdd gnd FILL
XFILL_2__1064_ vdd gnd FILL
XFILL91950x150 vdd gnd FILL
XFILL_2__1133_ vdd gnd FILL
X_1190_ _979_/A _1190_/B _1190_/C _1429_/B vdd gnd OAI21X1
XFILL_3__946_ vdd gnd FILL
XFILL_0__1602_ vdd gnd FILL
XFILL_3__1311_ vdd gnd FILL
XFILL_3__1173_ vdd gnd FILL
XFILL_0__1533_ vdd gnd FILL
XFILL_0__1464_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
XFILL_3__1242_ vdd gnd FILL
XFILL_1__1711_ vdd gnd FILL
X_1526_ _914_/C _1526_/B _1526_/C _1533_/C vdd gnd NAND3X1
X_1457_ _1539_/B _1457_/B _1460_/A vdd gnd AND2X2
XFILL_1__1642_ vdd gnd FILL
XFILL_1__1573_ vdd gnd FILL
X_1388_ _1491_/A _999_/B _1445_/C vdd gnd NAND2X1
XFILL_2__964_ vdd gnd FILL
XFILL_2__895_ vdd gnd FILL
X_970_ _995_/B _995_/A _983_/C _981_/A vdd gnd NAND3X1
XFILL_2__1820_ vdd gnd FILL
XFILL_1__1007_ vdd gnd FILL
XFILL_2__1682_ vdd gnd FILL
XFILL_2__1751_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
XFILL_2__1047_ vdd gnd FILL
XFILL_2__1116_ vdd gnd FILL
XFILL_1__982_ vdd gnd FILL
X_1311_ _1379_/A _1324_/A vdd gnd INVX1
X_1173_ _980_/B _1194_/A _1193_/A _1196_/C vdd gnd OAI21X1
X_1242_ _1329_/A _1329_/B _1330_/C vdd gnd NAND2X1
XFILL_3__1156_ vdd gnd FILL
XFILL_3__1087_ vdd gnd FILL
XFILL_3__1225_ vdd gnd FILL
XFILL_0__1516_ vdd gnd FILL
XFILL_0__1447_ vdd gnd FILL
XFILL_0__1378_ vdd gnd FILL
X_1509_ _1510_/A _1510_/B _1509_/C _1558_/C vdd gnd NAND3X1
XFILL_1__1556_ vdd gnd FILL
XFILL_1__1487_ vdd gnd FILL
XFILL_2__947_ vdd gnd FILL
XFILL_2__1803_ vdd gnd FILL
XFILL_2__1734_ vdd gnd FILL
X_953_ _979_/A _953_/B _975_/A vdd gnd NOR2X1
XFILL_2__1665_ vdd gnd FILL
XFILL_2__1596_ vdd gnd FILL
XFILL_3__1010_ vdd gnd FILL
XFILL_0__1232_ vdd gnd FILL
XFILL_0__1301_ vdd gnd FILL
X_1791_ _1811_/A _1811_/C _1808_/C vdd gnd NAND2X1
XFILL_0__1163_ vdd gnd FILL
XFILL_2_CLKBUF1_insert11 vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
XFILL_1__965_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
X_1156_ _1198_/C _1287_/A _1199_/C _1287_/B vdd gnd NAND3X1
XFILL_0_BUFX2_insert26 vdd gnd FILL
XFILL_1__896_ vdd gnd FILL
XFILL_0_BUFX2_insert37 vdd gnd FILL
X_1087_ _1233_/A _1237_/B _1237_/C _1103_/A vdd gnd NAND3X1
X_1225_ _979_/B _969_/B _1228_/B _1226_/C vdd gnd OAI21X1
XFILL_1__1410_ vdd gnd FILL
XFILL_1__1341_ vdd gnd FILL
XFILL_1__1272_ vdd gnd FILL
XFILL_1__1608_ vdd gnd FILL
XFILL_2__1450_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
XFILL_2__1381_ vdd gnd FILL
XFILL_1__1539_ vdd gnd FILL
XFILL_0__1781_ vdd gnd FILL
XFILL_2__1717_ vdd gnd FILL
X_936_ _978_/A _940_/B _937_/C vdd gnd NAND2X1
XFILL_2__1648_ vdd gnd FILL
XFILL_2__1579_ vdd gnd FILL
X_1010_ _1014_/B _1063_/C _1153_/C vdd gnd AND2X2
XFILL_0__1215_ vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
X_1774_ _1788_/A _1776_/B _1795_/C vdd gnd NAND2X1
XFILL_0__1077_ vdd gnd FILL
XFILL_3__1826_ vdd gnd FILL
XFILL_3__1688_ vdd gnd FILL
XFILL_3__1757_ vdd gnd FILL
XFILL_1__948_ vdd gnd FILL
X_1208_ _1208_/A _1208_/B _1208_/C _1350_/C vdd gnd OAI21X1
XFILL_1__1324_ vdd gnd FILL
XFILL_1__1255_ vdd gnd FILL
X_1139_ _1266_/A _1206_/B _1266_/C _1284_/B vdd gnd NAND3X1
XFILL_1__1186_ vdd gnd FILL
XFILL_0_BUFX2_insert7 vdd gnd FILL
XFILL_2__1433_ vdd gnd FILL
XFILL_2__1364_ vdd gnd FILL
XFILL_2__1502_ vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
XFILL_2__1295_ vdd gnd FILL
XFILL_0__897_ vdd gnd FILL
X_1490_ _1781_/A _1542_/A vdd gnd INVX1
XFILL_0__1764_ vdd gnd FILL
X_919_ _919_/A _919_/B _919_/Y vdd gnd OR2X2
XFILL_0__1695_ vdd gnd FILL
XFILL_1__1040_ vdd gnd FILL
X_1826_ _909_/B Done_o vdd gnd BUFX2
XFILL_0__1129_ vdd gnd FILL
X_1688_ _1688_/A _1722_/C _1768_/B vdd gnd NAND2X1
XFILL_3_BUFX2_insert41 vdd gnd FILL
XFILL_3__1809_ vdd gnd FILL
X_1757_ _1778_/A _945_/A _1760_/B vdd gnd AND2X2
XFILL_2__1080_ vdd gnd FILL
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_0__1480_ vdd gnd FILL
XFILL_2__1347_ vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
X_1611_ _934_/Y vdd _1631_/R _1631_/CLK _988_/A vdd gnd DFFSR
XFILL_2__1278_ vdd gnd FILL
XFILL_0__949_ vdd gnd FILL
X_1473_ _1473_/A _1510_/B _1473_/C _1516_/A vdd gnd NAND3X1
X_1542_ _1542_/A _1567_/B _1567_/A _1542_/D _1543_/A vdd gnd OAI22X1
XFILL_0__1678_ vdd gnd FILL
XFILL_0__1816_ vdd gnd FILL
XFILL_0__1747_ vdd gnd FILL
XFILL_3__1525_ vdd gnd FILL
XFILL_2__980_ vdd gnd FILL
XBUFX2_insert39 ABCmd_i[2] _1677_/A vdd gnd BUFX2
X_1809_ _1809_/A _1809_/B _1809_/C _1810_/A vdd gnd AOI21X1
XBUFX2_insert28 _915_/Y _946_/B vdd gnd BUFX2
XFILL_1__1023_ vdd gnd FILL
XBUFX2_insert17 _925_/Y _1624_/R vdd gnd BUFX2
XFILL_1__1787_ vdd gnd FILL
XFILL_2__1201_ vdd gnd FILL
XFILL_2__1132_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_0__1601_ vdd gnd FILL
XFILL_0__1532_ vdd gnd FILL
XFILL_0__1463_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
XFILL_1__1710_ vdd gnd FILL
XFILL_1__1641_ vdd gnd FILL
X_1525_ ABCmd_i[7] _1816_/C _1526_/B vdd gnd OR2X2
X_1387_ _1387_/A _1387_/B _1400_/A vdd gnd OR2X2
X_1456_ _1567_/A _1498_/B _1456_/C _1457_/B vdd gnd OAI21X1
XFILL_3__1508_ vdd gnd FILL
XFILL_1__1572_ vdd gnd FILL
XFILL_3__1439_ vdd gnd FILL
XFILL_2__963_ vdd gnd FILL
XFILL_2__894_ vdd gnd FILL
XFILL_2__1750_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_2__1681_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
XFILL_2__1046_ vdd gnd FILL
XFILL_1__981_ vdd gnd FILL
XFILL_3__1790_ vdd gnd FILL
X_1241_ _1247_/A _1247_/B _1308_/A vdd gnd AND2X2
X_1310_ _986_/D _999_/B _1379_/A vdd gnd NAND2X1
X_1172_ _1172_/A _1172_/B _1172_/C _1194_/A vdd gnd AOI21X1
XFILL_0__1515_ vdd gnd FILL
XFILL_0__1446_ vdd gnd FILL
XFILL_0__1377_ vdd gnd FILL
X_1508_ _1511_/B _1511_/C _1509_/C vdd gnd NAND2X1
X_1439_ _1439_/A _1439_/B _1439_/C _1468_/A vdd gnd OAI21X1
XFILL_1__1555_ vdd gnd FILL
XFILL_1__1486_ vdd gnd FILL
XFILL92850x85950 vdd gnd FILL
XFILL_2__946_ vdd gnd FILL
XFILL_2__1802_ vdd gnd FILL
XFILL_2__1733_ vdd gnd FILL
X_952_ _952_/A _953_/B vdd gnd INVX2
XFILL_2__1664_ vdd gnd FILL
XFILL_2__1595_ vdd gnd FILL
X_1790_ _1803_/A _1799_/A _1798_/C _1811_/A vdd gnd NAND3X1
XFILL_0__1300_ vdd gnd FILL
XFILL_0__1231_ vdd gnd FILL
XFILL_0__1162_ vdd gnd FILL
XFILL_3__1773_ vdd gnd FILL
XFILL_2__1029_ vdd gnd FILL
XFILL_0__1093_ vdd gnd FILL
XFILL_2_CLKBUF1_insert12 vdd gnd FILL
XFILL_0_BUFX2_insert38 vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
XFILL_0_BUFX2_insert27 vdd gnd FILL
XFILL_0_BUFX2_insert16 vdd gnd FILL
XFILL_1__895_ vdd gnd FILL
X_1224_ _1303_/A _1302_/A _1228_/B vdd gnd AND2X2
X_1155_ _1177_/D _1177_/C _1155_/C _1199_/C vdd gnd NAND3X1
X_1086_ _1237_/A _1233_/C _1233_/B _1103_/B vdd gnd OAI21X1
XFILL_1__1340_ vdd gnd FILL
XFILL_1__1271_ vdd gnd FILL
XFILL_0__1429_ vdd gnd FILL
XFILL92550x15750 vdd gnd FILL
XFILL_1__1607_ vdd gnd FILL
XFILL_1__1538_ vdd gnd FILL
XFILL_2__1380_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
XFILL_1__1469_ vdd gnd FILL
XFILL_2__929_ vdd gnd FILL
XFILL_2__1716_ vdd gnd FILL
X_935_ ABCmd_i[3] _937_/A vdd gnd INVX1
XFILL_0__1780_ vdd gnd FILL
XFILL_2__1647_ vdd gnd FILL
XFILL_2__1578_ vdd gnd FILL
XFILL_0__1145_ vdd gnd FILL
X_1773_ _1804_/B _1788_/A vdd gnd INVX1
XFILL_0__1214_ vdd gnd FILL
XFILL_0__1076_ vdd gnd FILL
XFILL_1__947_ vdd gnd FILL
X_1207_ _1207_/A _1207_/B _1295_/A vdd gnd NAND2X1
X_1069_ _1157_/A _1157_/B _1158_/A _1286_/B vdd gnd OAI21X1
XFILL_1__1323_ vdd gnd FILL
XFILL_1__1254_ vdd gnd FILL
X_1138_ _1138_/A _1138_/B _1138_/C _1266_/C vdd gnd NAND3X1
XFILL92550x27450 vdd gnd FILL
XFILL_1__1185_ vdd gnd FILL
XFILL_2__1501_ vdd gnd FILL
XFILL_2__1432_ vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_2__1294_ vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
XFILL_0__896_ vdd gnd FILL
XFILL_0__1763_ vdd gnd FILL
XFILL_0__1694_ vdd gnd FILL
X_918_ _921_/B _946_/B _918_/C _921_/D _919_/B vdd gnd OAI22X1
XFILL_3__1472_ vdd gnd FILL
XFILL_3__1541_ vdd gnd FILL
X_1756_ _1781_/A _1810_/B vdd gnd INVX1
XFILL_0__1059_ vdd gnd FILL
XFILL_3_BUFX2_insert31 vdd gnd FILL
X_1825_ _1825_/A ACC_o[7] vdd gnd BUFX2
XFILL_0__1128_ vdd gnd FILL
X_1687_ _1691_/B _1687_/B _1688_/A vdd gnd NAND2X1
XFILL_1__1168_ vdd gnd FILL
XFILL_1__1237_ vdd gnd FILL
XFILL_1__1306_ vdd gnd FILL
XFILL_3__961_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_3__892_ vdd gnd FILL
XFILL_2__1277_ vdd gnd FILL
XFILL_2__1346_ vdd gnd FILL
XFILL_2__1415_ vdd gnd FILL
X_1610_ _931_/Y vdd _1628_/R _1628_/CLK _1610_/Q vdd gnd DFFSR
XFILL_0__948_ vdd gnd FILL
XFILL_0__1815_ vdd gnd FILL
X_1472_ _1472_/A _1472_/B _1472_/C _1473_/C vdd gnd OAI21X1
X_1541_ _1760_/A _945_/A _1584_/A _1585_/A vdd gnd NAND3X1
XFILL_0__1677_ vdd gnd FILL
XFILL_0__1746_ vdd gnd FILL
XFILL_3__1455_ vdd gnd FILL
XFILL_3__1386_ vdd gnd FILL
XBUFX2_insert18 _925_/Y _1628_/R vdd gnd BUFX2
XBUFX2_insert29 _915_/Y _940_/B vdd gnd BUFX2
XFILL_1__1022_ vdd gnd FILL
X_1808_ ABCmd_i[6] _1808_/B _1808_/C _1815_/B vdd gnd NAND3X1
X_1739_ _1741_/A _1741_/B _1794_/B vdd gnd XOR2X1
XFILL_1__1786_ vdd gnd FILL
XFILL_3_CLKBUF1_insert8 vdd gnd FILL
XFILL_2__1200_ vdd gnd FILL
XFILL_2__1131_ vdd gnd FILL
XFILL_2__1062_ vdd gnd FILL
XFILL_3__944_ vdd gnd FILL
XFILL_0__1531_ vdd gnd FILL
XFILL_0__1600_ vdd gnd FILL
XFILL_0__1462_ vdd gnd FILL
XFILL_3__1240_ vdd gnd FILL
XFILL_3__1171_ vdd gnd FILL
XFILL_2__1329_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
X_1524_ _1524_/A _1549_/B ABCmd_i[7] _1526_/C vdd gnd OAI21X1
XFILL_1__1640_ vdd gnd FILL
X_1455_ _999_/B _1498_/B vdd gnd INVX1
X_1386_ _1406_/B _1406_/A _1462_/A vdd gnd NAND2X1
XFILL_1__1571_ vdd gnd FILL
XFILL_2__962_ vdd gnd FILL
XFILL_0__1729_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_2__893_ vdd gnd FILL
XFILL_2__1680_ vdd gnd FILL
XFILL_1__1769_ vdd gnd FILL
XFILL_2__1114_ vdd gnd FILL
XFILL_2__1045_ vdd gnd FILL
X_1171_ _1172_/B _1172_/C _1172_/A _1193_/A vdd gnd NAND3X1
XFILL_1__980_ vdd gnd FILL
XFILL_3__927_ vdd gnd FILL
X_1240_ _1248_/B _1330_/A _1248_/A _1298_/A vdd gnd NAND3X1
XFILL_3__1154_ vdd gnd FILL
XFILL_3__1223_ vdd gnd FILL
XFILL_0__1514_ vdd gnd FILL
XFILL_0__1445_ vdd gnd FILL
XFILL_3__1085_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
X_1507_ _1538_/A _1538_/B _1507_/C _1511_/B vdd gnd NAND3X1
XFILL_1__1554_ vdd gnd FILL
X_1438_ _1516_/B _1476_/C vdd gnd INVX1
X_1369_ _1422_/A _1422_/B _1515_/A _1421_/A vdd gnd NAND3X1
XFILL_2__945_ vdd gnd FILL
XFILL_1__1485_ vdd gnd FILL
XFILL_2__1801_ vdd gnd FILL
XFILL_2__1663_ vdd gnd FILL
XFILL_2__1732_ vdd gnd FILL
X_951_ _999_/A _979_/A vdd gnd INVX1
XFILL_2__1594_ vdd gnd FILL
XFILL_2__1028_ vdd gnd FILL
XFILL_0__1092_ vdd gnd FILL
XFILL_0__1230_ vdd gnd FILL
XFILL_0__1161_ vdd gnd FILL
XFILL_1__963_ vdd gnd FILL
XFILL_0_BUFX2_insert39 vdd gnd FILL
X_1154_ _1154_/A _994_/Y _998_/Y _1177_/D vdd gnd NAND3X1
XFILL_0_BUFX2_insert28 vdd gnd FILL
XFILL_1__894_ vdd gnd FILL
XFILL_0_BUFX2_insert17 vdd gnd FILL
X_1223_ _1496_/A _953_/B _1228_/A _1226_/B vdd gnd OAI21X1
XFILL_0__1428_ vdd gnd FILL
X_1085_ _1104_/C _1104_/B _1104_/A _1246_/B vdd gnd AOI21X1
XFILL_1__1270_ vdd gnd FILL
XFILL_3__1206_ vdd gnd FILL
XFILL_3__1137_ vdd gnd FILL
XFILL_0__1359_ vdd gnd FILL
XFILL_3__1068_ vdd gnd FILL
XFILL_1__1606_ vdd gnd FILL
XFILL_1__1537_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
XFILL_2__928_ vdd gnd FILL
XFILL_1__1468_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_2__1715_ vdd gnd FILL
XFILL_2__1646_ vdd gnd FILL
X_934_ _934_/A _949_/B _934_/C _934_/Y vdd gnd OAI21X1
XFILL_2__1577_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
X_1772_ _1772_/A _1772_/B _1772_/C _1772_/D _1776_/B vdd gnd AOI22X1
XFILL_0__1075_ vdd gnd FILL
XFILL_0__1213_ vdd gnd FILL
XFILL_3__1755_ vdd gnd FILL
XFILL_3__1824_ vdd gnd FILL
XFILL_1__946_ vdd gnd FILL
X_1206_ _1206_/A _1206_/B _1206_/C _1265_/C vdd gnd AOI21X1
X_1137_ _1137_/A _1137_/B _1137_/C _1206_/B vdd gnd NAND3X1
XFILL_1__1184_ vdd gnd FILL
X_1068_ _1068_/A _1068_/B _1068_/C _1157_/A vdd gnd AOI21X1
XFILL_1__1253_ vdd gnd FILL
XFILL_1__1322_ vdd gnd FILL
XFILL_2__1431_ vdd gnd FILL
XFILL_2__1500_ vdd gnd FILL
XFILL_2__1362_ vdd gnd FILL
XFILL_2__1293_ vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_0__895_ vdd gnd FILL
XFILL_0__1762_ vdd gnd FILL
XFILL_0__1693_ vdd gnd FILL
X_917_ LoadB_i _924_/A _921_/D vdd gnd NOR2X1
X_1686_ _1690_/B _1690_/A _1722_/A _1687_/B vdd gnd OAI21X1
X_1755_ _1755_/A _1755_/B _1755_/C _1805_/A vdd gnd OAI21X1
XFILL_0__1058_ vdd gnd FILL
XFILL_3_BUFX2_insert21 vdd gnd FILL
X_1824_ _1824_/A ACC_o[6] vdd gnd BUFX2
XFILL_0__1127_ vdd gnd FILL
XFILL_3__1669_ vdd gnd FILL
XFILL_3__1807_ vdd gnd FILL
XFILL_3__1738_ vdd gnd FILL
XFILL_1__929_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_2__1414_ vdd gnd FILL
XFILL_2__1276_ vdd gnd FILL
XFILL_2__1345_ vdd gnd FILL
XFILL_0__947_ vdd gnd FILL
X_1540_ _1542_/A _1542_/D _1584_/A vdd gnd NOR2X1
XFILL_0__1814_ vdd gnd FILL
X_1471_ _1471_/A _1471_/B _1471_/C _1472_/B vdd gnd AOI21X1
XFILL_0__1676_ vdd gnd FILL
XFILL_0__1745_ vdd gnd FILL
X_1807_ _1807_/A _1807_/B _1815_/A _1816_/C vdd gnd OAI21X1
XBUFX2_insert19 _925_/Y _1632_/R vdd gnd BUFX2
XFILL_1__1021_ vdd gnd FILL
X_1669_ _1677_/A _1670_/B _1783_/C _1670_/C vdd gnd OAI21X1
X_1738_ _1770_/A _1741_/B vdd gnd INVX1
XFILL_1__1785_ vdd gnd FILL
XFILL_2__1061_ vdd gnd FILL
XFILL_2__1130_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL_0__1530_ vdd gnd FILL
XFILL_0__1461_ vdd gnd FILL
XFILL_2__1328_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2_BUFX2_insert0 vdd gnd FILL
X_1454_ _1454_/A _1499_/A _1539_/B vdd gnd OR2X2
X_1523_ _1558_/C _1558_/A _1560_/C _1560_/A _1524_/A vdd gnd AOI22X1
XFILL_0__1728_ vdd gnd FILL
XFILL_3__1506_ vdd gnd FILL
XFILL_1__1570_ vdd gnd FILL
X_1385_ _1439_/B _1385_/B _1439_/A _1406_/B vdd gnd OAI21X1
XFILL_2__961_ vdd gnd FILL
XFILL_0__1659_ vdd gnd FILL
XFILL_3__1437_ vdd gnd FILL
XFILL_3__1299_ vdd gnd FILL
XFILL_3__1368_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_2__892_ vdd gnd FILL
XFILL_1__1699_ vdd gnd FILL
XFILL_1__1768_ vdd gnd FILL
XFILL_2__1044_ vdd gnd FILL
XFILL_2__1113_ vdd gnd FILL
XFILL91650x27450 vdd gnd FILL
X_1170_ _1170_/A _961_/B _961_/A _1172_/B vdd gnd OAI21X1
XFILL_0__1375_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
XFILL_0__1513_ vdd gnd FILL
X_1437_ _1437_/A _922_/C _1535_/A _1479_/C vdd gnd OAI21X1
X_1506_ _1506_/A _1506_/B _1507_/C vdd gnd OR2X2
XFILL_1__1484_ vdd gnd FILL
XFILL_1__1553_ vdd gnd FILL
X_1299_ _1299_/A _1299_/B _1299_/C _1417_/C vdd gnd OAI21X1
X_1368_ _1368_/A _1370_/C _1422_/B vdd gnd NOR2X1
XFILL_2__944_ vdd gnd FILL
XFILL_2__1800_ vdd gnd FILL
X_950_ _950_/A _950_/Y vdd gnd INVX1
XFILL_2__1662_ vdd gnd FILL
XFILL_2__1731_ vdd gnd FILL
XFILL_2__1593_ vdd gnd FILL
XFILL_2__1027_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
XFILL_3__1771_ vdd gnd FILL
X_1153_ _1153_/A _1153_/B _1153_/C _1177_/C vdd gnd OAI21X1
XFILL_0_BUFX2_insert18 vdd gnd FILL
XFILL_1__893_ vdd gnd FILL
XFILL_3__909_ vdd gnd FILL
XFILL_0_BUFX2_insert29 vdd gnd FILL
X_1222_ _977_/A _986_/D _1228_/A vdd gnd AND2X2
X_1084_ _1237_/A _1233_/C _1237_/B _1104_/C vdd gnd OAI21X1
XFILL_0__1427_ vdd gnd FILL
XFILL93150x46950 vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL_1__1605_ vdd gnd FILL
XFILL_1__1467_ vdd gnd FILL
XFILL_1__1536_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
XFILL_2__1714_ vdd gnd FILL
X_933_ _988_/A _949_/B _934_/C vdd gnd NAND2X1
XFILL_2__1645_ vdd gnd FILL
XFILL_2__1576_ vdd gnd FILL
XFILL_0__1212_ vdd gnd FILL
XFILL_0__1143_ vdd gnd FILL
X_1771_ _1771_/A _1809_/B _1772_/B vdd gnd OR2X2
XFILL_0__1074_ vdd gnd FILL
XFILL_3__1685_ vdd gnd FILL
XFILL_1__945_ vdd gnd FILL
X_1067_ _1067_/A _1067_/B _1067_/C _1157_/B vdd gnd AOI21X1
XFILL_1__1321_ vdd gnd FILL
X_1205_ _1205_/A _1588_/B _1587_/B _1515_/A vdd gnd OAI21X1
X_1136_ _1206_/C _1266_/B _1206_/A _1284_/C vdd gnd OAI21X1
XFILL_1__1183_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_3__1119_ vdd gnd FILL
XFILL_2__1430_ vdd gnd FILL
XFILL_2__1361_ vdd gnd FILL
XFILL_1__1519_ vdd gnd FILL
XFILL_2__1292_ vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
XFILL_0__894_ vdd gnd FILL
XFILL_0__1761_ vdd gnd FILL
X_916_ LoadA_i _924_/A _921_/B vdd gnd NOR2X1
XFILL_3__1470_ vdd gnd FILL
XFILL_0__1692_ vdd gnd FILL
XFILL_2__1559_ vdd gnd FILL
X_1823_ _1823_/A ACC_o[5] vdd gnd BUFX2
X_1685_ _1809_/B _1690_/A _1690_/B _1722_/A vdd gnd OAI21X1
X_1754_ _1795_/A _1754_/Y vdd gnd INVX1
XFILL_0__1057_ vdd gnd FILL
XFILL_3_BUFX2_insert33 vdd gnd FILL
XFILL_0__1126_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__1235_ vdd gnd FILL
X_1119_ _1127_/A _1128_/B _1128_/C _1123_/B vdd gnd NAND3X1
XFILL_1__1304_ vdd gnd FILL
XFILL_1__1166_ vdd gnd FILL
XFILL_1__1097_ vdd gnd FILL
XFILL_3__890_ vdd gnd FILL
XFILL91650x150 vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL_2__1413_ vdd gnd FILL
XFILL_2__1275_ vdd gnd FILL
XFILL_0__946_ vdd gnd FILL
X_1470_ _1472_/C _1470_/B _1470_/C _1521_/A vdd gnd NAND3X1
XFILL_0__1813_ vdd gnd FILL
XFILL_0__1744_ vdd gnd FILL
XFILL_3__1453_ vdd gnd FILL
XFILL_3__1522_ vdd gnd FILL
XFILL_0__1675_ vdd gnd FILL
XFILL_3__1384_ vdd gnd FILL
X_1806_ _1806_/A _1806_/B _1815_/A vdd gnd XOR2X1
XFILL_1__1020_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
X_1668_ _1668_/A _1668_/B _1668_/C _1690_/B vdd gnd OAI21X1
X_1737_ _1737_/A _1737_/B _1770_/C _1770_/A vdd gnd OAI21X1
X_1599_ _988_/B _1601_/B _1600_/C vdd gnd NAND2X1
XFILL_1__1784_ vdd gnd FILL
XFILL_2__1060_ vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_3__942_ vdd gnd FILL
XFILL91950x4050 vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_0__1460_ vdd gnd FILL
XFILL_2__1327_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
XFILL_2__1189_ vdd gnd FILL
XFILL_2__1258_ vdd gnd FILL
XFILL_2_BUFX2_insert1 vdd gnd FILL
X_1453_ _1781_/A _999_/B _1499_/A vdd gnd NAND2X1
X_1522_ _1522_/A _1522_/B _1522_/C _1560_/C vdd gnd OAI21X1
XFILL_0__1658_ vdd gnd FILL
XFILL_0__1727_ vdd gnd FILL
X_1384_ _1384_/A _1384_/B _1439_/B vdd gnd NOR2X1
XFILL_2__960_ vdd gnd FILL
XFILL_2__891_ vdd gnd FILL
XFILL_0__1589_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_1__1767_ vdd gnd FILL
XFILL_1__1698_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL_2__1112_ vdd gnd FILL
XFILL_3__925_ vdd gnd FILL
XFILL_0__1512_ vdd gnd FILL
XFILL_3__1152_ vdd gnd FILL
XFILL_3__1083_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
XFILL_3__1221_ vdd gnd FILL
X_1436_ _1817_/Y _1437_/A vdd gnd INVX1
X_1505_ _1538_/C _1505_/B _1505_/C _1511_/C vdd gnd OAI21X1
X_1367_ _1367_/A _1367_/B _1367_/C _1367_/D _1368_/A vdd gnd AOI22X1
XFILL_1__1483_ vdd gnd FILL
XFILL_1__1552_ vdd gnd FILL
X_1298_ _1298_/A _1298_/B _1298_/C _1299_/B vdd gnd AOI21X1
XFILL_2__943_ vdd gnd FILL
XFILL_2__1730_ vdd gnd FILL
XFILL_2__1661_ vdd gnd FILL
XFILL_1__1819_ vdd gnd FILL
XFILL_2__1592_ vdd gnd FILL
XFILL_2__1026_ vdd gnd FILL
XFILL_0__1090_ vdd gnd FILL
XFILL_1__961_ vdd gnd FILL
XFILL_1__892_ vdd gnd FILL
X_1221_ _999_/B _988_/B _1304_/C vdd gnd NAND2X1
X_1152_ _1163_/A _1163_/B _1174_/A _1155_/C vdd gnd AOI21X1
XFILL_3__1204_ vdd gnd FILL
XFILL_0_BUFX2_insert19 vdd gnd FILL
X_1083_ _1083_/A _1387_/A _1233_/C vdd gnd NOR2X1
XFILL_0__1288_ vdd gnd FILL
XFILL_3__1066_ vdd gnd FILL
XFILL_0__1426_ vdd gnd FILL
XFILL_0__1357_ vdd gnd FILL
XFILL_3__1135_ vdd gnd FILL
XFILL_1__1604_ vdd gnd FILL
X_1419_ _1419_/A _1470_/B _1419_/C _1516_/B vdd gnd NAND3X1
XFILL_1__1535_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL_1__1466_ vdd gnd FILL
XFILL_2__926_ vdd gnd FILL
XFILL_2__1713_ vdd gnd FILL
X_932_ _932_/A _934_/A vdd gnd INVX1
XFILL_2__1644_ vdd gnd FILL
XFILL_2__1575_ vdd gnd FILL
X_1770_ _1770_/A _1770_/B _1770_/C _1772_/C vdd gnd OAI21X1
XFILL_0__1142_ vdd gnd FILL
XFILL_0__1211_ vdd gnd FILL
XFILL_2__1009_ vdd gnd FILL
XFILL_0__1073_ vdd gnd FILL
XFILL_1__944_ vdd gnd FILL
X_1204_ _1576_/C _1576_/B _1204_/C _1588_/B vdd gnd AOI21X1
X_1066_ _1158_/B _1158_/C _1157_/C _1286_/A vdd gnd NAND3X1
XFILL_1__1320_ vdd gnd FILL
XFILL_1__1251_ vdd gnd FILL
X_1135_ _1137_/B _1137_/A _1137_/C _1206_/C vdd gnd AOI21X1
XFILL_1__1182_ vdd gnd FILL
XFILL_0__1409_ vdd gnd FILL
XFILL_2__1360_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_1__1518_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_0__893_ vdd gnd FILL
XFILL_2__909_ vdd gnd FILL
XFILL_0__1691_ vdd gnd FILL
XFILL_0__1760_ vdd gnd FILL
X_915_ _915_/A _915_/B _915_/Y vdd gnd NAND2X1
XFILL_2__1489_ vdd gnd FILL
XFILL_2__1558_ vdd gnd FILL
X_1753_ _1755_/B _1772_/D _1795_/A vdd gnd XOR2X1
X_1822_ _1822_/A ACC_o[4] vdd gnd BUFX2
XFILL_0__1125_ vdd gnd FILL
X_1684_ _1684_/A _1684_/B _1684_/C _1684_/D _1691_/B vdd gnd AOI22X1
XFILL_3__1805_ vdd gnd FILL
XFILL_3__1736_ vdd gnd FILL
XFILL_0__1056_ vdd gnd FILL
XFILL_3_BUFX2_insert23 vdd gnd FILL
XFILL_3__1667_ vdd gnd FILL
XFILL_1__927_ vdd gnd FILL
XFILL_3__1598_ vdd gnd FILL
X_1049_ _1049_/A _1049_/B _1049_/C _1054_/B vdd gnd NAND3X1
XFILL_1__1234_ vdd gnd FILL
X_1118_ _1120_/A _1121_/C _1128_/B vdd gnd NAND2X1
XFILL_1__1303_ vdd gnd FILL
XFILL_1__1165_ vdd gnd FILL
XFILL_1__1096_ vdd gnd FILL
XFILL_2__1274_ vdd gnd FILL
XFILL_2__1412_ vdd gnd FILL
XFILL_2__1343_ vdd gnd FILL
XFILL_0__945_ vdd gnd FILL
XFILL_0__1674_ vdd gnd FILL
XFILL_0__1812_ vdd gnd FILL
XFILL_0__1743_ vdd gnd FILL
X_1805_ _1805_/A _1805_/B _1805_/C _1806_/A vdd gnd AOI21X1
X_1736_ _1809_/B _1737_/B _1737_/A _1770_/C vdd gnd OAI21X1
XFILL_0__1108_ vdd gnd FILL
XFILL_0__1039_ vdd gnd FILL
XFILL_1__1783_ vdd gnd FILL
XFILL_3__1719_ vdd gnd FILL
X_1667_ _978_/B _1667_/B _1802_/B _1668_/B vdd gnd OAI21X1
X_1598_ _934_/A _1606_/B _1598_/C _1627_/D vdd gnd OAI21X1
XFILL92550x11850 vdd gnd FILL
XFILL_1__1148_ vdd gnd FILL
XFILL_1__1217_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_2__1326_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_2__1257_ vdd gnd FILL
XFILL_2__1188_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
XFILL_2_BUFX2_insert2 vdd gnd FILL
X_1452_ _1760_/A _1452_/B _1454_/A vdd gnd NAND2X1
X_1521_ _1521_/A _1521_/B _1521_/C _1522_/C vdd gnd AOI21X1
X_1383_ _1384_/B _1384_/A _1385_/B vdd gnd AND2X2
XFILL_0__1657_ vdd gnd FILL
XFILL_0__1726_ vdd gnd FILL
XFILL_3__1366_ vdd gnd FILL
XFILL_3__1504_ vdd gnd FILL
XFILL_3__1435_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_2__890_ vdd gnd FILL
XFILL92550x4050 vdd gnd FILL
XFILL_0__1588_ vdd gnd FILL
X_1719_ _1725_/B _1725_/A _1769_/B vdd gnd XOR2X1
XFILL92550x23550 vdd gnd FILL
XFILL_1__1766_ vdd gnd FILL
XFILL_1__1697_ vdd gnd FILL
XFILL_2__1111_ vdd gnd FILL
XFILL_2__1042_ vdd gnd FILL
XFILL_0__1511_ vdd gnd FILL
XFILL_2__1309_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
X_1504_ _1538_/B _1505_/B vdd gnd INVX1
XFILL_1__1551_ vdd gnd FILL
X_1366_ _1416_/B _1366_/B _1366_/C _1370_/C vdd gnd AOI21X1
X_1435_ _1821_/A _1486_/A vdd gnd INVX1
XFILL_1__1482_ vdd gnd FILL
XFILL_0__1709_ vdd gnd FILL
XFILL_2__942_ vdd gnd FILL
X_1297_ _1352_/A _1418_/A vdd gnd INVX1
XFILL_3__1418_ vdd gnd FILL
XFILL_3__1349_ vdd gnd FILL
XFILL92550x35250 vdd gnd FILL
XFILL_2__1660_ vdd gnd FILL
XFILL_1__1749_ vdd gnd FILL
XFILL_1__1818_ vdd gnd FILL
XFILL_2__1591_ vdd gnd FILL
XFILL_2__1025_ vdd gnd FILL
XFILL_1__960_ vdd gnd FILL
X_1151_ _1151_/A _1151_/B _1151_/C _1163_/B vdd gnd NAND3X1
XFILL_2__1789_ vdd gnd FILL
XFILL_1__891_ vdd gnd FILL
X_1220_ _1220_/A _1220_/B _1220_/C _1338_/C vdd gnd AOI21X1
X_1082_ _1082_/A _1781_/A _1387_/A vdd gnd NAND2X1
XFILL_0__1425_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
XFILL_0__1356_ vdd gnd FILL
XFILL_1__1603_ vdd gnd FILL
X_1418_ _1418_/A _1418_/B _1418_/C _1419_/C vdd gnd OAI21X1
X_1349_ _1367_/D _1367_/C _1349_/C _1355_/B vdd gnd NAND3X1
XFILL_1__1534_ vdd gnd FILL
XFILL_2__925_ vdd gnd FILL
XFILL_1__1465_ vdd gnd FILL
XFILL_1__1396_ vdd gnd FILL
XFILL_2__1643_ vdd gnd FILL
XFILL_2__1712_ vdd gnd FILL
X_931_ _931_/A _943_/B _931_/C _931_/Y vdd gnd OAI21X1
XFILL_2__1574_ vdd gnd FILL
XFILL_2__1008_ vdd gnd FILL
XFILL_0__1210_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
XFILL_0__1141_ vdd gnd FILL
XFILL_3__1752_ vdd gnd FILL
XFILL_3__1821_ vdd gnd FILL
XFILL_3__1683_ vdd gnd FILL
XFILL_1__943_ vdd gnd FILL
X_1203_ _1203_/A _1203_/B _1551_/A _1576_/B vdd gnd OAI21X1
X_1134_ _1208_/A _1256_/A _1208_/C _1137_/A vdd gnd NAND3X1
X_1065_ _1158_/A _1157_/C vdd gnd INVX1
XFILL_1__1181_ vdd gnd FILL
XFILL_1__1250_ vdd gnd FILL
XFILL_0__1408_ vdd gnd FILL
XFILL_3__1117_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
XFILL_2__1290_ vdd gnd FILL
XFILL_1__1517_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_2__908_ vdd gnd FILL
XFILL_0__892_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_0__1690_ vdd gnd FILL
X_914_ _914_/A _924_/B _914_/C _919_/A vdd gnd OAI21X1
XFILL_2__1488_ vdd gnd FILL
XFILL_2__1557_ vdd gnd FILL
X_1683_ _1683_/A _1683_/B _1683_/C _1684_/C vdd gnd NAND3X1
X_1752_ _1755_/A _1772_/D vdd gnd INVX1
XFILL_3_BUFX2_insert35 vdd gnd FILL
XFILL_0__1055_ vdd gnd FILL
X_1821_ _1821_/A ACC_o[3] vdd gnd BUFX2
XFILL_0__1124_ vdd gnd FILL
XFILL_1__926_ vdd gnd FILL
X_1117_ _1567_/B _1121_/B _1120_/A vdd gnd NOR2X1
XFILL_1__1164_ vdd gnd FILL
X_1048_ _979_/B _1211_/A _1048_/C _1049_/C vdd gnd OAI21X1
XFILL_1__1233_ vdd gnd FILL
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1095_ vdd gnd FILL
XFILL_2__1411_ vdd gnd FILL
XFILL91350x7950 vdd gnd FILL
XFILL_2__1273_ vdd gnd FILL
XFILL_2__1342_ vdd gnd FILL
XFILL_0__944_ vdd gnd FILL
XFILL_0__1811_ vdd gnd FILL
XFILL_3__1520_ vdd gnd FILL
XFILL_0__1673_ vdd gnd FILL
XFILL_0__1742_ vdd gnd FILL
XFILL_3__1451_ vdd gnd FILL
XFILL_3__1382_ vdd gnd FILL
X_1804_ _1804_/A _1804_/B _1805_/B vdd gnd NOR2X1
X_1666_ ABCmd_i[0] _1666_/B _1667_/B vdd gnd NOR2X1
X_1735_ _932_/A _939_/A _1735_/C _1737_/B vdd gnd AOI21X1
XFILL_0__1038_ vdd gnd FILL
XFILL_0__1107_ vdd gnd FILL
XFILL_1__1782_ vdd gnd FILL
X_1597_ _962_/B _1606_/B _1598_/C vdd gnd NAND2X1
XFILL_1__909_ vdd gnd FILL
XFILL_1__1147_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_3__940_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
XFILL_2__1325_ vdd gnd FILL
XFILL_2__1256_ vdd gnd FILL
XFILL_0__927_ vdd gnd FILL
X_1520_ _1520_/A _1520_/B _1520_/C _1560_/A vdd gnd OAI21X1
XFILL_2_BUFX2_insert3 vdd gnd FILL
X_1451_ _1488_/B _1451_/B _1488_/A _1460_/B vdd gnd OAI21X1
X_1382_ _1382_/A _1439_/C _1382_/C _1406_/A vdd gnd NAND3X1
XFILL_0__1656_ vdd gnd FILL
XFILL_0__1725_ vdd gnd FILL
XFILL_3__1296_ vdd gnd FILL
XFILL_0__1587_ vdd gnd FILL
XFILL_1__1001_ vdd gnd FILL
X_1649_ _999_/A _1802_/A vdd gnd INVX1
X_1718_ _1718_/A _1718_/B _1725_/C _1725_/A vdd gnd OAI21X1
XFILL_1__1696_ vdd gnd FILL
XFILL_1__1765_ vdd gnd FILL
XFILL_2__1041_ vdd gnd FILL
XFILL_2__1110_ vdd gnd FILL
XFILL_3__923_ vdd gnd FILL
XFILL_3__1150_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_0__1510_ vdd gnd FILL
XFILL93150x4050 vdd gnd FILL
XFILL_3__1081_ vdd gnd FILL
XFILL_2__1308_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
X_1503_ _1506_/B _1506_/A _1538_/B vdd gnd NAND2X1
XFILL_0__1708_ vdd gnd FILL
X_1434_ _911_/A _1434_/B _1434_/C _1619_/D vdd gnd OAI21X1
X_1365_ _904_/B _904_/C _1820_/A _1434_/C vdd gnd OAI21X1
X_1296_ _1296_/A _1296_/B _1296_/C _1352_/A vdd gnd OAI21X1
XFILL_1__1550_ vdd gnd FILL
XFILL_0__1639_ vdd gnd FILL
XFILL_1__1481_ vdd gnd FILL
XFILL_2__941_ vdd gnd FILL
XFILL92850x19650 vdd gnd FILL
XFILL_1__1817_ vdd gnd FILL
XFILL_2__1590_ vdd gnd FILL
XFILL_1__1679_ vdd gnd FILL
XFILL_1__1748_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
XFILL_2__1788_ vdd gnd FILL
X_1150_ _955_/Y _980_/C _1163_/A vdd gnd AND2X2
XFILL_1__890_ vdd gnd FILL
XFILL_3__906_ vdd gnd FILL
XFILL_0_CLKBUF1_insert10 vdd gnd FILL
XFILL_3__1202_ vdd gnd FILL
X_1081_ _1233_/A _1233_/B _1237_/C _1104_/B vdd gnd NAND3X1
XFILL_0__1355_ vdd gnd FILL
XFILL_0__1424_ vdd gnd FILL
XFILL_3__1133_ vdd gnd FILL
XFILL_0__1286_ vdd gnd FILL
XFILL_3__1064_ vdd gnd FILL
X_1417_ _1417_/A _1417_/B _1417_/C _1418_/B vdd gnd AOI21X1
XFILL_1__1602_ vdd gnd FILL
X_1279_ _950_/Y _903_/A _1279_/C _1617_/D vdd gnd OAI21X1
XFILL_1__1533_ vdd gnd FILL
X_1348_ _1352_/A _1353_/B _1353_/C _1367_/C vdd gnd NAND3X1
XFILL_1__1464_ vdd gnd FILL
XFILL_2__924_ vdd gnd FILL
XFILL_1__1395_ vdd gnd FILL
X_930_ _991_/A _943_/B _931_/C vdd gnd NAND2X1
XFILL_2__1711_ vdd gnd FILL
XFILL_2__1642_ vdd gnd FILL
XFILL91650x11850 vdd gnd FILL
XFILL_2__1573_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
XFILL_2__1007_ vdd gnd FILL
XFILL_0__1140_ vdd gnd FILL
XFILL_1__942_ vdd gnd FILL
X_1202_ _1575_/A _1576_/C vdd gnd INVX1
X_1064_ _1071_/B _1071_/A _1158_/A vdd gnd XNOR2X1
X_1133_ _1208_/B _1256_/C _1256_/B _1137_/B vdd gnd OAI21X1
XFILL_1__1180_ vdd gnd FILL
XFILL_3__1047_ vdd gnd FILL
XFILL_0__1338_ vdd gnd FILL
XFILL_0__1407_ vdd gnd FILL
XFILL_0__1269_ vdd gnd FILL
XFILL_1__1516_ vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL_2__907_ vdd gnd FILL
XFILL_0__891_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
X_913_ LoadA_i LoadB_i _924_/A _914_/A vdd gnd OAI21X1
XFILL_2__1556_ vdd gnd FILL
X_1820_ _1820_/A ACC_o[2] vdd gnd BUFX2
XFILL_2__1487_ vdd gnd FILL
XFILL_3__1803_ vdd gnd FILL
X_1682_ _1682_/A _1682_/B _1683_/C vdd gnd NAND2X1
X_1751_ _1772_/A _1771_/A _1755_/C _1755_/A vdd gnd OAI21X1
XFILL_3_BUFX2_insert25 vdd gnd FILL
XFILL_3_BUFX2_insert14 vdd gnd FILL
XFILL_0__1054_ vdd gnd FILL
XFILL_0__1123_ vdd gnd FILL
XFILL_3__1665_ vdd gnd FILL
XFILL_3__1734_ vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_3__1596_ vdd gnd FILL
X_1047_ _953_/B _1301_/A _1047_/C _1049_/B vdd gnd OAI21X1
XFILL_1__1301_ vdd gnd FILL
X_1116_ _1567_/B _1121_/B _1120_/B _1128_/C vdd gnd OAI21X1
XFILL_1__1163_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL_1__1232_ vdd gnd FILL
XFILL_2__1410_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_2__1341_ vdd gnd FILL
XFILL_0__943_ vdd gnd FILL
XFILL91650x35250 vdd gnd FILL
XFILL_0__1810_ vdd gnd FILL
XFILL_0__1741_ vdd gnd FILL
XFILL_0__1672_ vdd gnd FILL
XFILL_2__1608_ vdd gnd FILL
XFILL_2__1539_ vdd gnd FILL
X_1803_ _1803_/A _1804_/A _1803_/C _1805_/C vdd gnd OAI21X1
X_1665_ _964_/A _1666_/B vdd gnd INVX1
X_1734_ _932_/A _939_/A _1783_/C _1735_/C vdd gnd OAI21X1
X_1596_ _931_/A _1601_/B _1596_/C _1626_/D vdd gnd OAI21X1
XFILL_0__1037_ vdd gnd FILL
XFILL_0__1106_ vdd gnd FILL
XFILL_3__1648_ vdd gnd FILL
XFILL_1__1781_ vdd gnd FILL
XFILL_3__1717_ vdd gnd FILL
XFILL_1__908_ vdd gnd FILL
XFILL_3__1579_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_2__1186_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
XFILL_2__1255_ vdd gnd FILL
XFILL_2_BUFX2_insert4 vdd gnd FILL
X_1450_ _1488_/C _1451_/B vdd gnd INVX1
XFILL_0__1724_ vdd gnd FILL
XFILL_3__999_ vdd gnd FILL
XFILL_3__1502_ vdd gnd FILL
X_1381_ _1384_/B _1384_/A _1382_/C vdd gnd OR2X2
XFILL_0__1655_ vdd gnd FILL
XFILL_0__1586_ vdd gnd FILL
XFILL93150x54750 vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
X_1648_ _1679_/A _1678_/B vdd gnd INVX1
X_1717_ _1809_/B _1718_/B _1718_/A _1725_/C vdd gnd OAI21X1
X_1579_ _1579_/A _914_/C _1580_/B vdd gnd NOR2X1
XFILL_1__1695_ vdd gnd FILL
XFILL_1__1764_ vdd gnd FILL
XFILL_2__1040_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
XFILL_2__1307_ vdd gnd FILL
XFILL_2__1169_ vdd gnd FILL
XFILL_0__909_ vdd gnd FILL
XFILL_2__1238_ vdd gnd FILL
X_1433_ _1433_/A _1433_/B _1433_/C _1433_/D _1434_/B vdd gnd AOI22X1
X_1502_ _1506_/B _1506_/A _1538_/C vdd gnd NOR2X1
XFILL_0__1707_ vdd gnd FILL
XFILL_1__1480_ vdd gnd FILL
X_1364_ _1364_/A _911_/A _1364_/C _1364_/D _1618_/D vdd gnd AOI22X1
XFILL_3__1416_ vdd gnd FILL
X_1295_ _1295_/A _1295_/B _1295_/C _1349_/C vdd gnd AOI21X1
XFILL_0__1638_ vdd gnd FILL
XFILL_2__940_ vdd gnd FILL
XFILL_3__1278_ vdd gnd FILL
XFILL_3__1347_ vdd gnd FILL
XFILL_0__1569_ vdd gnd FILL
XFILL_1__1816_ vdd gnd FILL
XFILL_1__1747_ vdd gnd FILL
XFILL_1__1678_ vdd gnd FILL
XFILL_2__1023_ vdd gnd FILL
XFILL_2__1787_ vdd gnd FILL
XFILL_0_CLKBUF1_insert11 vdd gnd FILL
X_1080_ _1237_/B _1233_/B vdd gnd INVX1
XFILL_0__1354_ vdd gnd FILL
XFILL_0__1423_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
XFILL93150x78150 vdd gnd FILL
XFILL_1__1601_ vdd gnd FILL
X_1347_ _1347_/A _1347_/B _1417_/C _1353_/B vdd gnd OAI21X1
X_1416_ _1418_/C _1416_/B _1416_/C _1420_/B vdd gnd NAND3X1
X_1278_ _903_/A _1278_/B _1279_/C vdd gnd NAND2X1
XFILL_1__1532_ vdd gnd FILL
XFILL_1__1463_ vdd gnd FILL
XFILL_1__1394_ vdd gnd FILL
XFILL_2__923_ vdd gnd FILL
XFILL_2__1710_ vdd gnd FILL
XFILL_2__1641_ vdd gnd FILL
XFILL_2__1572_ vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
XFILL_2__1006_ vdd gnd FILL
XFILL_3__1681_ vdd gnd FILL
XFILL_3__1750_ vdd gnd FILL
X_1201_ _1551_/A _1551_/B _1551_/C _1575_/A vdd gnd NAND3X1
XFILL_1__941_ vdd gnd FILL
X_989_ _997_/B _996_/C vdd gnd INVX1
X_1132_ _1158_/B _1157_/C _1157_/A _1137_/C vdd gnd AOI21X1
X_1063_ _979_/C _1063_/B _1063_/C _1071_/B vdd gnd OAI21X1
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1406_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
XFILL_0__1199_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_1__1515_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL_0__890_ vdd gnd FILL
XFILL_2__906_ vdd gnd FILL
XFILL91350x150 vdd gnd FILL
X_912_ _912_/A _912_/B _912_/Y vdd gnd NAND2X1
XFILL92850x150 vdd gnd FILL
XFILL_2__1555_ vdd gnd FILL
XFILL_2__1486_ vdd gnd FILL
X_1750_ _1809_/B _1771_/A _1772_/A _1755_/C vdd gnd OAI21X1
XFILL_0__1122_ vdd gnd FILL
X_1681_ _1681_/A _1802_/A ABCmd_i[5] _1682_/A vdd gnd AOI21X1
XFILL_0__1053_ vdd gnd FILL
XFILL_3_BUFX2_insert37 vdd gnd FILL
XFILL_1__924_ vdd gnd FILL
X_1046_ _1114_/C _1114_/D _1046_/C _1054_/A vdd gnd NAND3X1
XFILL_1__1300_ vdd gnd FILL
XFILL_1__1231_ vdd gnd FILL
X_1115_ _1121_/C _1120_/B vdd gnd INVX1
XFILL_3__1029_ vdd gnd FILL
XFILL_1__1093_ vdd gnd FILL
XFILL_1__1162_ vdd gnd FILL
XFILL_2__1340_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_0__942_ vdd gnd FILL
XFILL91950x19650 vdd gnd FILL
XFILL_2__1271_ vdd gnd FILL
XFILL_0__1671_ vdd gnd FILL
XFILL_0__1740_ vdd gnd FILL
XFILL_2__1607_ vdd gnd FILL
XFILL_2__1469_ vdd gnd FILL
XFILL_2__1538_ vdd gnd FILL
XFILL_3__1380_ vdd gnd FILL
X_1802_ _1802_/A _1802_/B _1806_/B vdd gnd NOR2X1
X_1733_ _1733_/A _1733_/B _1733_/C _1737_/A vdd gnd OAI21X1
XFILL_0__1105_ vdd gnd FILL
XFILL_1__1780_ vdd gnd FILL
X_1664_ _1780_/A _1670_/B _1664_/C _1780_/D _1668_/A vdd gnd AOI22X1
X_1595_ _978_/B _1601_/B _1596_/C vdd gnd NAND2X1
XFILL_0__1036_ vdd gnd FILL
XFILL_1__907_ vdd gnd FILL
X_1029_ _1102_/A _1102_/B _1088_/A _1088_/B vdd gnd NAND3X1
XFILL_1__1214_ vdd gnd FILL
XFILL_1__1145_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_2__1323_ vdd gnd FILL
XFILL_2__1185_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
XFILL_2__1254_ vdd gnd FILL
XFILL_2_BUFX2_insert5 vdd gnd FILL
X_1380_ _1384_/A _1384_/B _1439_/C vdd gnd NAND2X1
XFILL_0__1654_ vdd gnd FILL
XFILL_0__1723_ vdd gnd FILL
XFILL_3__1432_ vdd gnd FILL
XFILL_3__1363_ vdd gnd FILL
XFILL_3__1294_ vdd gnd FILL
XFILL_0__1585_ vdd gnd FILL
X_1716_ _1716_/A _1716_/B _1716_/C _1718_/B vdd gnd AOI21X1
XFILL_1__1763_ vdd gnd FILL
X_1647_ ABCmd_i[5] _1802_/B vdd gnd INVX2
X_1578_ ABCmd_i[7] _1775_/Y _1579_/A vdd gnd NOR2X1
XFILL_0__1019_ vdd gnd FILL
XFILL_1__1694_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_3__921_ vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_2__1237_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
XFILL_2__1306_ vdd gnd FILL
XFILL_2__1168_ vdd gnd FILL
XFILL_0__908_ vdd gnd FILL
XFILL_2__1099_ vdd gnd FILL
X_1432_ _1432_/A _914_/C _1433_/B vdd gnd NOR2X1
X_1363_ _1363_/A _899_/A _911_/A _1364_/D vdd gnd AOI21X1
X_1501_ _1566_/A _1501_/B _1506_/A vdd gnd NAND2X1
XFILL_0__1637_ vdd gnd FILL
XFILL_0__1706_ vdd gnd FILL
X_1294_ _1367_/A _1295_/C vdd gnd INVX1
XFILL_0__1499_ vdd gnd FILL
XFILL_0__1568_ vdd gnd FILL
XFILL_1__1815_ vdd gnd FILL
XFILL_1__1746_ vdd gnd FILL
XFILL_1__1677_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL_2__1022_ vdd gnd FILL
XFILL91950x7950 vdd gnd FILL
XFILL_2__1786_ vdd gnd FILL
XFILL_3__904_ vdd gnd FILL
XFILL_0_CLKBUF1_insert12 vdd gnd FILL
XFILL_3__1200_ vdd gnd FILL
XFILL_3__1062_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_3__1131_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
XFILL_1__1531_ vdd gnd FILL
XFILL_1__1600_ vdd gnd FILL
X_1346_ _1417_/A _1417_/B _1346_/C _1353_/C vdd gnd NAND3X1
X_1415_ _1470_/B _1419_/A _1416_/C vdd gnd NAND2X1
X_1277_ _1277_/A _1277_/B _1277_/C _1278_/B vdd gnd OAI21X1
XFILL_2__922_ vdd gnd FILL
XFILL_1__1462_ vdd gnd FILL
XFILL_1__1393_ vdd gnd FILL
XFILL_2__1640_ vdd gnd FILL
XFILL_1__1729_ vdd gnd FILL
XFILL_2__1571_ vdd gnd FILL
XFILL_2__1005_ vdd gnd FILL
XFILL_2__1769_ vdd gnd FILL
X_1200_ _1200_/A _1200_/B _1200_/C _1551_/B vdd gnd NAND3X1
X_988_ _988_/A _988_/B _997_/B vdd gnd NAND2X1
XFILL_1__940_ vdd gnd FILL
X_1062_ _979_/A _1567_/B _1071_/A vdd gnd NOR2X1
XFILL_0__1405_ vdd gnd FILL
X_1131_ _1138_/B _1138_/A _1138_/C _1266_/B vdd gnd AOI21X1
XFILL_3__1045_ vdd gnd FILL
XFILL_3__1114_ vdd gnd FILL
XFILL_0__1336_ vdd gnd FILL
XFILL_0__1267_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
XFILL_1__1514_ vdd gnd FILL
X_1329_ _1329_/A _1329_/B _1330_/B vdd gnd NOR2X1
XFILL92250x54750 vdd gnd FILL
XFILL_2__905_ vdd gnd FILL
XFILL_1__1445_ vdd gnd FILL
XFILL_1__1376_ vdd gnd FILL
X_911_ _911_/A _911_/B _911_/C _922_/A _912_/A vdd gnd AOI22X1
XFILL_2__1554_ vdd gnd FILL
XFILL_2__1485_ vdd gnd FILL
XFILL_0__1052_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
X_1680_ _1680_/A _1680_/B _1682_/B vdd gnd NAND2X1
XFILL_3__1801_ vdd gnd FILL
XFILL_3_BUFX2_insert27 vdd gnd FILL
XFILL_3_BUFX2_insert16 vdd gnd FILL
XFILL_3__1594_ vdd gnd FILL
XFILL_1__923_ vdd gnd FILL
X_1114_ _1114_/A _1114_/B _1114_/C _1114_/D _1121_/C vdd gnd AOI22X1
X_1045_ _953_/B _1301_/A _1063_/B _1114_/C vdd gnd OAI21X1
XFILL_1__1230_ vdd gnd FILL
XFILL_1__1161_ vdd gnd FILL
XFILL_1__1092_ vdd gnd FILL
XFILL_0__1319_ vdd gnd FILL
XFILL_2__1270_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_0__941_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_0__1670_ vdd gnd FILL
XFILL_2__1606_ vdd gnd FILL
XFILL_2__1468_ vdd gnd FILL
XFILL_2__1537_ vdd gnd FILL
XFILL_2__1399_ vdd gnd FILL
X_1801_ ABCmd_i[6] _1808_/B _1807_/A vdd gnd NAND2X1
X_1663_ _978_/B _1670_/B _1778_/A _1664_/C vdd gnd NAND3X1
X_1732_ _986_/D _1732_/B _1802_/B _1733_/A vdd gnd OAI21X1
XFILL_0__1035_ vdd gnd FILL
XFILL_0__1104_ vdd gnd FILL
XFILL_3__1715_ vdd gnd FILL
X_1594_ _928_/A _1604_/B _1594_/C _1625_/D vdd gnd OAI21X1
XFILL_0__1799_ vdd gnd FILL
XFILL_3__1646_ vdd gnd FILL
XFILL_3__1577_ vdd gnd FILL
XFILL_1__906_ vdd gnd FILL
XFILL_1__1144_ vdd gnd FILL
X_1028_ _1075_/B _1102_/B vdd gnd INVX1
XFILL_1__1213_ vdd gnd FILL
XFILL_1__1075_ vdd gnd FILL
XFILL92250x78150 vdd gnd FILL
XFILL_2__1253_ vdd gnd FILL
XFILL_2__1322_ vdd gnd FILL
XFILL_2__1184_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_2_BUFX2_insert6 vdd gnd FILL
XFILL_0__1722_ vdd gnd FILL
XFILL_0__1653_ vdd gnd FILL
XFILL_0__1584_ vdd gnd FILL
X_1715_ _1716_/A _1716_/B _1783_/C _1716_/C vdd gnd OAI21X1
X_1646_ _1679_/A _1679_/B _1780_/D _1681_/A _1653_/A vdd gnd AOI22X1
XFILL_0__1018_ vdd gnd FILL
XFILL_1__1762_ vdd gnd FILL
XFILL_1__1693_ vdd gnd FILL
X_1577_ _1577_/A _1577_/B ABCmd_i[7] _1580_/A vdd gnd OAI21X1
XFILL_1__1127_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL_2__1236_ vdd gnd FILL
XFILL_0__907_ vdd gnd FILL
XFILL_2__1098_ vdd gnd FILL
X_1500_ _1500_/A _1500_/B _1539_/C _1566_/A vdd gnd NAND3X1
X_1362_ _1362_/A _1362_/B _1362_/C _1363_/A vdd gnd OAI21X1
X_1431_ ABCmd_i[7] _1704_/Y _1432_/A vdd gnd NOR2X1
X_1293_ _1513_/A _1522_/A _1370_/A _1357_/B vdd gnd OAI21X1
XFILL_0__1636_ vdd gnd FILL
XFILL_0__1705_ vdd gnd FILL
XFILL_3__1276_ vdd gnd FILL
XFILL_3__1345_ vdd gnd FILL
XFILL_3__1414_ vdd gnd FILL
XFILL_0__1567_ vdd gnd FILL
XFILL_0__1498_ vdd gnd FILL
XFILL_2_BUFX2_insert40 vdd gnd FILL
X_1629_ _1629_/D vdd _1632_/R _1635_/CLK _986_/D vdd gnd DFFSR
XFILL_1__1676_ vdd gnd FILL
XFILL_1__1814_ vdd gnd FILL
XFILL_1__1745_ vdd gnd FILL
XFILL_2__1021_ vdd gnd FILL
XFILL_2__998_ vdd gnd FILL
XFILL_2__1785_ vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
XFILL_2__1219_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
X_1276_ _1792_/A ABCmd_i[7] _922_/C _1277_/B vdd gnd OAI21X1
XFILL_1__1530_ vdd gnd FILL
X_1345_ _1418_/A _1418_/C _1352_/C _1367_/D vdd gnd NAND3X1
X_1414_ _1414_/A _1472_/C _1414_/C _1470_/B vdd gnd NAND3X1
XFILL_2__921_ vdd gnd FILL
XFILL_1__1461_ vdd gnd FILL
XFILL_3__1328_ vdd gnd FILL
XFILL_3__1259_ vdd gnd FILL
XFILL92550x7950 vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_1__1659_ vdd gnd FILL
XFILL_1__1728_ vdd gnd FILL
XFILL_2__1570_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
XFILL_2__1699_ vdd gnd FILL
XFILL_2__1768_ vdd gnd FILL
X_987_ _996_/A _997_/A vdd gnd INVX1
X_1130_ _1208_/B _1256_/C _1208_/A _1138_/B vdd gnd OAI21X1
X_1061_ _945_/A _1567_/B vdd gnd INVX4
XFILL_0__1404_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
XFILL_0__1197_ vdd gnd FILL
XFILL_0__1266_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
X_1328_ _1342_/C _1341_/C _1375_/C vdd gnd NOR2X1
X_1259_ _1263_/A _1263_/B _1262_/C _1295_/B vdd gnd OAI21X1
XFILL_1__1444_ vdd gnd FILL
XFILL_1__1513_ vdd gnd FILL
XFILL_2__904_ vdd gnd FILL
XFILL_1__1375_ vdd gnd FILL
XFILL_2__1553_ vdd gnd FILL
X_910_ _922_/B _914_/C _910_/C _911_/C vdd gnd OAI21X1
XFILL_2__1484_ vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_0__1120_ vdd gnd FILL
XFILL_3_BUFX2_insert39 vdd gnd FILL
XFILL_3__1662_ vdd gnd FILL
XFILL_3__1731_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
X_1044_ _976_/A _962_/B _1063_/B vdd gnd NAND2X1
X_1113_ _1128_/A _1127_/A vdd gnd INVX1
XFILL_1__1091_ vdd gnd FILL
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1160_ vdd gnd FILL
XFILL_3__1027_ vdd gnd FILL
XFILL_0__1249_ vdd gnd FILL
XFILL92850x15750 vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_0__940_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
XFILL_2__1605_ vdd gnd FILL
XFILL_2__1536_ vdd gnd FILL
X_1800_ _1813_/A _1813_/C _1807_/B vdd gnd NAND2X1
XFILL_2__1398_ vdd gnd FILL
XFILL_2__1467_ vdd gnd FILL
X_1662_ ABCmd_i[5] _962_/B _1668_/C vdd gnd NAND2X1
X_1731_ _1780_/A _939_/A _1731_/C _1780_/D _1733_/B vdd gnd AOI22X1
XFILL_0__1034_ vdd gnd FILL
XFILL_0__1103_ vdd gnd FILL
X_1593_ _999_/A _1604_/B _1594_/C vdd gnd NAND2X1
XFILL_1__905_ vdd gnd FILL
XFILL_0__1798_ vdd gnd FILL
X_1027_ _988_/A _986_/D _1075_/B vdd gnd NAND2X1
XFILL_1__1143_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_1__1212_ vdd gnd FILL
XFILL92850x27450 vdd gnd FILL
XFILL_2__1183_ vdd gnd FILL
XFILL_2__1321_ vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
XFILL_0__1721_ vdd gnd FILL
XFILL_2_BUFX2_insert7 vdd gnd FILL
XFILL_3__996_ vdd gnd FILL
XFILL_0__1652_ vdd gnd FILL
XFILL_3__1430_ vdd gnd FILL
XFILL_3__1361_ vdd gnd FILL
XFILL_2__1519_ vdd gnd FILL
XFILL_0__1583_ vdd gnd FILL
XFILL_3__1292_ vdd gnd FILL
X_1645_ _999_/A ABCmd_i[1] _1679_/B vdd gnd NAND2X1
X_1714_ _1714_/A _1714_/B _1714_/C _1718_/A vdd gnd OAI21X1
XFILL_0__1017_ vdd gnd FILL
X_1576_ _1576_/A _1576_/B _1576_/C _1577_/A vdd gnd AOI21X1
XFILL_1__1692_ vdd gnd FILL
XFILL_1__1761_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
XFILL_2__1304_ vdd gnd FILL
XFILL_2__1166_ vdd gnd FILL
XFILL91350x54750 vdd gnd FILL
XFILL_0__906_ vdd gnd FILL
XFILL_2__1235_ vdd gnd FILL
X_1430_ _1430_/A _1430_/B ABCmd_i[7] _1433_/A vdd gnd OAI21X1
XFILL_2__1097_ vdd gnd FILL
XFILL_0__1704_ vdd gnd FILL
X_1361_ _1361_/A _1361_/B ABCmd_i[7] _1362_/A vdd gnd OAI21X1
X_1292_ _1370_/A _1292_/B _1513_/A vdd gnd NAND2X1
XFILL_0__1566_ vdd gnd FILL
XFILL_0__1497_ vdd gnd FILL
XFILL_1__1813_ vdd gnd FILL
XFILL_2_BUFX2_insert41 vdd gnd FILL
X_1628_ _1628_/D vdd _1628_/R _1628_/CLK _988_/B vdd gnd DFFSR
XFILL_2_BUFX2_insert30 vdd gnd FILL
X_1559_ _1570_/C _1560_/B vdd gnd INVX1
XFILL_1__1675_ vdd gnd FILL
XFILL_1__1744_ vdd gnd FILL
XFILL_2__1020_ vdd gnd FILL
XFILL_2__997_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_2__1784_ vdd gnd FILL
XFILL_3__902_ vdd gnd FILL
XFILL_3__1060_ vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_2__1149_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
XFILL_2__1218_ vdd gnd FILL
X_1413_ _1413_/A _1413_/B _1413_/C _1414_/C vdd gnd OAI21X1
X_1275_ _986_/A _999_/A _949_/A _1277_/A vdd gnd AOI21X1
X_1344_ _1347_/A _1347_/B _1346_/C _1352_/C vdd gnd OAI21X1
XFILL_1__1460_ vdd gnd FILL
XFILL_2__920_ vdd gnd FILL
XFILL_1__1391_ vdd gnd FILL
XFILL_0__1549_ vdd gnd FILL
XFILL_1__1727_ vdd gnd FILL
XFILL_1__1658_ vdd gnd FILL
XFILL_1__1589_ vdd gnd FILL
XFILL_2__1003_ vdd gnd FILL
XFILL93150x7950 vdd gnd FILL
XFILL_2__1698_ vdd gnd FILL
XFILL_2__1767_ vdd gnd FILL
X_986_ _986_/A _991_/B _991_/A _986_/D _996_/A vdd gnd AOI22X1
X_1060_ _1067_/B _1067_/A _1067_/C _1158_/C vdd gnd NAND3X1
XFILL_3__1043_ vdd gnd FILL
XFILL_3__1112_ vdd gnd FILL
XFILL_0__1403_ vdd gnd FILL
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1196_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
XFILL93150x50850 vdd gnd FILL
XFILL_1__998_ vdd gnd FILL
X_1189_ _988_/A _1190_/B vdd gnd INVX1
XFILL_1__1512_ vdd gnd FILL
X_1258_ _1258_/A _1258_/B _1299_/A _1263_/B vdd gnd AOI21X1
XFILL_1__1443_ vdd gnd FILL
X_1327_ _1400_/B _1341_/A _1342_/C vdd gnd NAND2X1
XFILL_2__903_ vdd gnd FILL
XFILL_1__1374_ vdd gnd FILL
XFILL_2__1483_ vdd gnd FILL
XFILL_2__1552_ vdd gnd FILL
XFILL_3_BUFX2_insert18 vdd gnd FILL
XFILL_3_BUFX2_insert29 vdd gnd FILL
XFILL_0__1050_ vdd gnd FILL
XFILL_1__921_ vdd gnd FILL
XFILL_2__1819_ vdd gnd FILL
XFILL_3__1592_ vdd gnd FILL
X_1043_ _988_/B _1301_/A vdd gnd INVX2
X_969_ _969_/A _969_/B _972_/A _995_/B vdd gnd OAI21X1
X_1112_ _999_/A _948_/A _1128_/A vdd gnd NAND2X1
XFILL93150x62550 vdd gnd FILL
XFILL_0__1248_ vdd gnd FILL
XFILL_0__1317_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
XFILL_2__1604_ vdd gnd FILL
XFILL_2__1535_ vdd gnd FILL
XFILL_2__1466_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_2__1397_ vdd gnd FILL
X_1661_ _1661_/A _1661_/B _1661_/C _1674_/B vdd gnd OAI21X1
X_1730_ _986_/D _1732_/B _1731_/C vdd gnd NAND2X1
XFILL_0__999_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
X_1592_ _1592_/A _911_/A _1592_/C _1592_/D _1624_/D vdd gnd AOI22X1
XFILL_3__1644_ vdd gnd FILL
XFILL_3__1713_ vdd gnd FILL
XFILL_3__1575_ vdd gnd FILL
XFILL_1__904_ vdd gnd FILL
XFILL93150x74250 vdd gnd FILL
XFILL_0__1797_ vdd gnd FILL
X_1026_ _1026_/A _1496_/A _1083_/A _1102_/A vdd gnd OAI21X1
XFILL_1__1211_ vdd gnd FILL
XFILL_1__1142_ vdd gnd FILL
XFILL_1__1073_ vdd gnd FILL
XFILL_2__1320_ vdd gnd FILL
XFILL_2__1182_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_2__1251_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_0__1651_ vdd gnd FILL
XFILL_0__1720_ vdd gnd FILL
XFILL_2__1518_ vdd gnd FILL
XFILL_2__1449_ vdd gnd FILL
XFILL_0__1582_ vdd gnd FILL
X_1713_ _988_/B _1713_/B _1802_/B _1714_/A vdd gnd OAI21X1
X_1644_ _1679_/A _1778_/A _1681_/A vdd gnd NAND2X1
XFILL_1__1760_ vdd gnd FILL
XFILL_0__1016_ vdd gnd FILL
X_1575_ _1575_/A _1575_/B _1577_/B vdd gnd NOR2X1
XFILL_1__1691_ vdd gnd FILL
XFILL_3__1558_ vdd gnd FILL
X_1009_ _999_/Y _1009_/B _1009_/C _1014_/B vdd gnd NAND3X1
XFILL_3__1489_ vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_2__1303_ vdd gnd FILL
XFILL_2__1165_ vdd gnd FILL
XFILL_0__905_ vdd gnd FILL
XFILL_2__1234_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
X_1360_ _1689_/Y _949_/A _1362_/C vdd gnd NAND2X1
XFILL_0__1703_ vdd gnd FILL
XFILL_3__978_ vdd gnd FILL
XFILL_3__1412_ vdd gnd FILL
XFILL_3__1343_ vdd gnd FILL
X_1291_ _1291_/A _1587_/A _1291_/C _1522_/A vdd gnd AOI21X1
XFILL_0__1565_ vdd gnd FILL
XFILL_0__1496_ vdd gnd FILL
XFILL_1__1812_ vdd gnd FILL
XFILL_1__1743_ vdd gnd FILL
XFILL_2_BUFX2_insert20 vdd gnd FILL
X_1627_ _1627_/D vdd _1632_/R _1631_/CLK _962_/B vdd gnd DFFSR
XFILL_2_BUFX2_insert31 vdd gnd FILL
X_1489_ _1538_/A _1505_/C vdd gnd INVX1
X_1558_ _1558_/A _1561_/B _1558_/C _1570_/C vdd gnd NAND3X1
XFILL_1__1674_ vdd gnd FILL
XFILL_2__996_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_2__1783_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_2__1217_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
XFILL_2__1079_ vdd gnd FILL
X_1412_ _1471_/B _1471_/A _1471_/C _1472_/C vdd gnd NAND3X1
X_1343_ _1343_/A _1343_/B _1405_/A _1347_/B vdd gnd AOI21X1
X_1274_ _949_/A _1274_/B _1274_/C _1277_/C vdd gnd OAI21X1
XFILL_3__1326_ vdd gnd FILL
XFILL_1__1390_ vdd gnd FILL
XFILL_3__1188_ vdd gnd FILL
XFILL_3__1257_ vdd gnd FILL
XFILL_0__1548_ vdd gnd FILL
XFILL_0__1479_ vdd gnd FILL
XFILL_1__1726_ vdd gnd FILL
XFILL_1__1657_ vdd gnd FILL
XFILL_1__1588_ vdd gnd FILL
XFILL_2__1002_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
XFILL92550x150 vdd gnd FILL
XFILL91950x27450 vdd gnd FILL
X_985_ _991_/A _986_/D _985_/C _997_/C vdd gnd NAND3X1
XFILL_2__1697_ vdd gnd FILL
XFILL_2__1766_ vdd gnd FILL
XFILL_0__1402_ vdd gnd FILL
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
XFILL_1__997_ vdd gnd FILL
X_1326_ _1326_/A _1326_/B _1326_/C _1400_/B vdd gnd NAND3X1
XFILL_1__1511_ vdd gnd FILL
X_1188_ _1361_/A _1361_/B _1429_/C vdd gnd NOR2X1
XFILL_3__1309_ vdd gnd FILL
X_1257_ _1257_/A _1257_/B _1299_/C _1339_/B _1263_/A vdd gnd AOI22X1
XFILL_1__1373_ vdd gnd FILL
XFILL_1__1442_ vdd gnd FILL
XFILL_2__902_ vdd gnd FILL
XFILL_2__1551_ vdd gnd FILL
XFILL_2__1482_ vdd gnd FILL
XFILL_1__1709_ vdd gnd FILL
XFILL_3__1660_ vdd gnd FILL
XFILL_2__1749_ vdd gnd FILL
XFILL_1__920_ vdd gnd FILL
X_968_ _986_/D _969_/B vdd gnd INVX1
XFILL_2__1818_ vdd gnd FILL
X_899_ _899_/A _915_/B _909_/B _924_/B vdd gnd AOI21X1
X_1042_ _1047_/C _1048_/C _1046_/C vdd gnd NAND2X1
X_1111_ _1125_/B _1125_/C _1125_/A _1208_/C vdd gnd NAND3X1
XFILL_0__1316_ vdd gnd FILL
XFILL_0__1247_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
X_1309_ _1781_/A _988_/A _1325_/A vdd gnd NAND2X1
XFILL_1__1287_ vdd gnd FILL
XFILL_1__1425_ vdd gnd FILL
XFILL_1__1356_ vdd gnd FILL
XFILL_2__1603_ vdd gnd FILL
XFILL_2__1465_ vdd gnd FILL
XFILL_2__1396_ vdd gnd FILL
XFILL_2__1534_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_0__1032_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
X_1660_ _1660_/A _1684_/A _1661_/B vdd gnd NOR2X1
X_1591_ _1591_/A _899_/A _911_/A _1592_/D vdd gnd AOI21X1
XFILL_0__1796_ vdd gnd FILL
XFILL_1__903_ vdd gnd FILL
X_1025_ _984_/A _1760_/A _1083_/A vdd gnd NAND2X1
XFILL_1__1210_ vdd gnd FILL
XFILL_1__1141_ vdd gnd FILL
XFILL_3__1008_ vdd gnd FILL
XFILL_1__1072_ vdd gnd FILL
X_1789_ _1804_/A _1799_/A vdd gnd INVX1
XFILL_2__1250_ vdd gnd FILL
XFILL_0__921_ vdd gnd FILL
XFILL_2__1181_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_1__1408_ vdd gnd FILL
XFILL_0__1650_ vdd gnd FILL
XFILL_3__994_ vdd gnd FILL
XFILL_3__1290_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
XFILL_2__1517_ vdd gnd FILL
XFILL_0__1581_ vdd gnd FILL
XFILL_2__1379_ vdd gnd FILL
X_1643_ ABCmd_i[0] _1778_/A vdd gnd INVX2
X_1712_ _1780_/A _1716_/B _1712_/C _1780_/D _1714_/B vdd gnd AOI22X1
XFILL_0__1015_ vdd gnd FILL
X_1574_ _1576_/B _1576_/A _1575_/B vdd gnd NAND2X1
XFILL_1__1690_ vdd gnd FILL
XFILL_0__1779_ vdd gnd FILL
X_1008_ _979_/B _1121_/B _1114_/A _1009_/C vdd gnd OAI21X1
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_2__1302_ vdd gnd FILL
XFILL_2__1164_ vdd gnd FILL
XFILL_0__904_ vdd gnd FILL
XFILL_2__1095_ vdd gnd FILL
XFILL_0__1702_ vdd gnd FILL
X_1290_ _1575_/A _1290_/B _1576_/A _1291_/A vdd gnd OAI21X1
XFILL_0__1564_ vdd gnd FILL
XFILL_3__1273_ vdd gnd FILL
XFILL_0__1495_ vdd gnd FILL
X_1626_ _1626_/D vdd _1628_/R _1628_/CLK _978_/B vdd gnd DFFSR
XFILL_1__1673_ vdd gnd FILL
XFILL_1__1811_ vdd gnd FILL
XFILL_1__1742_ vdd gnd FILL
XFILL_2_BUFX2_insert21 vdd gnd FILL
XFILL_2_BUFX2_insert32 vdd gnd FILL
X_1488_ _1488_/A _1488_/B _1488_/C _1538_/A vdd gnd OAI21X1
X_1557_ _1824_/A _1581_/A vdd gnd INVX1
XFILL_2__995_ vdd gnd FILL
XFILL92250x62550 vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_2__1782_ vdd gnd FILL
XFILL_3__900_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_2__1216_ vdd gnd FILL
XFILL_2__1147_ vdd gnd FILL
XFILL_2__1078_ vdd gnd FILL
X_1273_ _1273_/A _922_/C _1274_/C vdd gnd NOR2X1
X_1411_ _1472_/A _1411_/B _1411_/C _1419_/A vdd gnd NAND3X1
X_1342_ _1342_/A _1342_/B _1342_/C _1343_/B vdd gnd OAI21X1
XFILL_0__1547_ vdd gnd FILL
XFILL_0__1478_ vdd gnd FILL
X_1609_ _928_/Y vdd _1628_/R _1628_/CLK _1609_/Q vdd gnd DFFSR
XFILL_1__1656_ vdd gnd FILL
XFILL_1__1725_ vdd gnd FILL
XFILL92250x74250 vdd gnd FILL
XFILL_2__1001_ vdd gnd FILL
XFILL_1__1587_ vdd gnd FILL
XFILL_2__978_ vdd gnd FILL
XFILL_2__1765_ vdd gnd FILL
X_984_ _984_/A _991_/B _985_/C vdd gnd AND2X2
XFILL_2__1696_ vdd gnd FILL
XFILL_3__1110_ vdd gnd FILL
XFILL_0__1401_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
XFILL_3__1041_ vdd gnd FILL
XFILL_0__1332_ vdd gnd FILL
XFILL_0__1263_ vdd gnd FILL
XFILL_1__996_ vdd gnd FILL
X_1325_ _1325_/A _1325_/B _1326_/A vdd gnd NOR2X1
XFILL_1__1510_ vdd gnd FILL
X_1256_ _1256_/A _1256_/B _1256_/C _1262_/C vdd gnd AOI21X1
X_1187_ _999_/A _1670_/B _1361_/B vdd gnd NAND2X1
XFILL_2__901_ vdd gnd FILL
XFILL_1__1441_ vdd gnd FILL
XFILL_1__1372_ vdd gnd FILL
XFILL_1__1639_ vdd gnd FILL
XFILL_1__1708_ vdd gnd FILL
XFILL_2__1481_ vdd gnd FILL
XFILL_2__1550_ vdd gnd FILL
X_967_ _967_/A _969_/A vdd gnd INVX1
XFILL_2__1817_ vdd gnd FILL
XFILL_2__1679_ vdd gnd FILL
XFILL_2__1748_ vdd gnd FILL
X_898_ _898_/A _898_/B _915_/B vdd gnd NOR2X1
X_1110_ _1220_/C _1246_/B _1246_/A _1125_/A vdd gnd OAI21X1
X_1041_ _978_/A _988_/B _1048_/C vdd gnd AND2X2
XFILL_0__1177_ vdd gnd FILL
XFILL_3__1024_ vdd gnd FILL
XFILL_0__1246_ vdd gnd FILL
XFILL_0__1315_ vdd gnd FILL
XFILL_3__1788_ vdd gnd FILL
XFILL_1__979_ vdd gnd FILL
X_1308_ _1308_/A _1308_/B _1342_/A _1341_/C vdd gnd AOI21X1
X_1239_ _1329_/A _1307_/A _1248_/B vdd gnd NAND2X1
XFILL_1__1424_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
XFILL_1__1355_ vdd gnd FILL
XFILL_2__1602_ vdd gnd FILL
XFILL_2__1533_ vdd gnd FILL
XFILL_2__1464_ vdd gnd FILL
XFILL_2__1395_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
XFILL_3__1711_ vdd gnd FILL
XFILL_3__1642_ vdd gnd FILL
XFILL_1__902_ vdd gnd FILL
X_1590_ _949_/A _1590_/B _1590_/C _1591_/A vdd gnd OAI21X1
XFILL_0__1795_ vdd gnd FILL
X_1024_ _1491_/A _1496_/A vdd gnd INVX2
XFILL_3__1573_ vdd gnd FILL
XFILL_1__1140_ vdd gnd FILL
X_1788_ _1788_/A _1805_/A _1798_/C vdd gnd NAND2X1
XFILL_1__1071_ vdd gnd FILL
XFILL_0__1229_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_0__920_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_0__1580_ vdd gnd FILL
XFILL_2__1516_ vdd gnd FILL
XFILL_2__1447_ vdd gnd FILL
XFILL_2__1378_ vdd gnd FILL
X_1711_ _988_/B _1713_/B _1712_/C vdd gnd NAND2X1
X_1642_ ABCmd_i[0] _1780_/A _1780_/D vdd gnd NAND2X1
XFILL_0__1014_ vdd gnd FILL
X_1573_ _1586_/C _1573_/B _1573_/C _1581_/C vdd gnd NAND3X1
XFILL_0__1778_ vdd gnd FILL
X_1007_ _978_/B _1121_/B vdd gnd INVX1
XFILL_3__1556_ vdd gnd FILL
XFILL_3__1487_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_1__1123_ vdd gnd FILL
XFILL_2__1163_ vdd gnd FILL
XFILL_2__1232_ vdd gnd FILL
XFILL_2__1301_ vdd gnd FILL
XFILL_0__903_ vdd gnd FILL
XFILL_2__1094_ vdd gnd FILL
XFILL_0__1701_ vdd gnd FILL
XFILL_3__976_ vdd gnd FILL
XFILL_0__1563_ vdd gnd FILL
XFILL_0__1494_ vdd gnd FILL
XFILL_1__1810_ vdd gnd FILL
X_1625_ _1625_/D vdd _1631_/R _1631_/CLK _999_/A vdd gnd DFFSR
XFILL_2_BUFX2_insert33 vdd gnd FILL
XFILL_2_BUFX2_insert22 vdd gnd FILL
X_1556_ _1556_/A _911_/A _1556_/C _1556_/D _1622_/D vdd gnd AOI22X1
XFILL_1__1672_ vdd gnd FILL
XFILL_1__1741_ vdd gnd FILL
XFILL_3__1608_ vdd gnd FILL
XFILL92850x11850 vdd gnd FILL
XFILL_3__1539_ vdd gnd FILL
X_1487_ _1822_/A _1533_/A vdd gnd INVX1
XFILL_2__994_ vdd gnd FILL
XFILL_1__1037_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_2__1781_ vdd gnd FILL
XFILL_2__1146_ vdd gnd FILL
XFILL_2__1215_ vdd gnd FILL
XFILL_2__1077_ vdd gnd FILL
X_1410_ _1413_/A _1413_/B _1471_/C _1411_/B vdd gnd OAI21X1
XFILL_3__959_ vdd gnd FILL
X_1272_ ABCmd_i[7] _1741_/A _1273_/A vdd gnd NOR2X1
X_1341_ _1341_/A _1400_/B _1341_/C _1343_/A vdd gnd NAND3X1
XFILL_3__1324_ vdd gnd FILL
XFILL_3__1255_ vdd gnd FILL
XFILL_0__1546_ vdd gnd FILL
XFILL_0__1477_ vdd gnd FILL
XFILL_3__1186_ vdd gnd FILL
X_1608_ _949_/A _918_/C _1608_/C _1632_/D vdd gnd OAI21X1
X_1539_ _1567_/B _1539_/B _1539_/C _1565_/A vdd gnd OAI21X1
XFILL92850x23550 vdd gnd FILL
XFILL_1__1655_ vdd gnd FILL
XFILL_1__1724_ vdd gnd FILL
XFILL_1__1586_ vdd gnd FILL
XFILL_2__1000_ vdd gnd FILL
XFILL_2__977_ vdd gnd FILL
X_983_ _983_/A _983_/B _983_/C _994_/C vdd gnd OAI21X1
XFILL_2__1695_ vdd gnd FILL
XFILL_2__1764_ vdd gnd FILL
XFILL_0__1400_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
XFILL_0__1262_ vdd gnd FILL
XFILL_2__1129_ vdd gnd FILL
XFILL_1__995_ vdd gnd FILL
X_1186_ _1190_/C _1186_/B _1429_/A vdd gnd OR2X2
X_1324_ _1324_/A _1324_/B _1379_/C _1326_/B vdd gnd NAND3X1
X_1255_ _1350_/A _1350_/B _1350_/C _1367_/A vdd gnd NAND3X1
XFILL_1__1440_ vdd gnd FILL
XFILL_3__1169_ vdd gnd FILL
XFILL_0__1529_ vdd gnd FILL
XFILL_2__900_ vdd gnd FILL
XFILL_1__1371_ vdd gnd FILL
XFILL_3__1307_ vdd gnd FILL
XFILL_3__1238_ vdd gnd FILL
XFILL92850x35250 vdd gnd FILL
XFILL_1__1638_ vdd gnd FILL
XFILL_1__1707_ vdd gnd FILL
XFILL_2__1480_ vdd gnd FILL
XFILL_1__1569_ vdd gnd FILL
XFILL_2__1816_ vdd gnd FILL
X_966_ _972_/A _992_/A _983_/C vdd gnd OR2X2
XFILL_2__1678_ vdd gnd FILL
XFILL_2__1747_ vdd gnd FILL
X_897_ _918_/C _921_/C vdd gnd INVX1
X_1040_ _976_/A _962_/B _1047_/C vdd gnd AND2X2
XFILL_0__1314_ vdd gnd FILL
XFILL_0__1176_ vdd gnd FILL
XFILL_0__1245_ vdd gnd FILL
X_1169_ _1186_/B _1184_/A _1169_/C _1172_/C vdd gnd OAI21X1
XFILL_1__978_ vdd gnd FILL
X_1307_ _1307_/A _1307_/B _1342_/A vdd gnd NOR2X1
XFILL_1__1423_ vdd gnd FILL
X_1238_ _1387_/A _1387_/B _1307_/A vdd gnd XNOR2X1
XFILL_1__1285_ vdd gnd FILL
XFILL_1__1354_ vdd gnd FILL
XFILL_2__1601_ vdd gnd FILL
XFILL_2__1532_ vdd gnd FILL
XFILL_3_CLKBUF1_insert10 vdd gnd FILL
XFILL_2__1463_ vdd gnd FILL
XFILL_2__1394_ vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_1__901_ vdd gnd FILL
XFILL_0__1794_ vdd gnd FILL
X_1023_ _991_/A _1026_/A vdd gnd INVX1
X_949_ _949_/A _949_/B _949_/C _949_/Y vdd gnd OAI21X1
XFILL_1__1070_ vdd gnd FILL
XFILL_3__1006_ vdd gnd FILL
XFILL_0__1228_ vdd gnd FILL
X_1787_ _1804_/A _1799_/B _1811_/C vdd gnd NAND2X1
XFILL_0__1159_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_3__992_ vdd gnd FILL
XFILL_2__1446_ vdd gnd FILL
XFILL_2__1515_ vdd gnd FILL
XFILL_2__1377_ vdd gnd FILL
XFILL_0__1013_ vdd gnd FILL
X_1710_ _1778_/A _1716_/B _1713_/B vdd gnd AND2X2
X_1641_ ABCmd_i[1] _1780_/A vdd gnd INVX2
XFILL_0__979_ vdd gnd FILL
X_1572_ _1572_/A _1572_/B _1572_/C _1573_/C vdd gnd OAI21X1
XFILL_0__1777_ vdd gnd FILL
X_1006_ _953_/B _1211_/A _955_/A _1009_/B vdd gnd OAI21X1
XFILL_1__1053_ vdd gnd FILL
XFILL_1__1122_ vdd gnd FILL
XFILL_2__1300_ vdd gnd FILL
XFILL_0__902_ vdd gnd FILL
XFILL_2__1093_ vdd gnd FILL
XFILL_2__1231_ vdd gnd FILL
XFILL_2__1162_ vdd gnd FILL
XFILL_0__1700_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL_3__1340_ vdd gnd FILL
XFILL_0__1562_ vdd gnd FILL
XFILL_3__1271_ vdd gnd FILL
XFILL_0__1493_ vdd gnd FILL
XFILL_1__1740_ vdd gnd FILL
XFILL_2_BUFX2_insert34 vdd gnd FILL
X_1555_ _1555_/A _1555_/B _911_/A _1556_/D vdd gnd AOI21X1
XFILL_2_BUFX2_insert23 vdd gnd FILL
X_1624_ _1624_/D vdd _1624_/R _1624_/CLK _1825_/A vdd gnd DFFSR
XFILL_1__1671_ vdd gnd FILL
X_1486_ _1486_/A _911_/A _1486_/C _1486_/D _1620_/D vdd gnd AOI22X1
XFILL_2__993_ vdd gnd FILL
XFILL_1__1036_ vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_2__1780_ vdd gnd FILL
XFILL_2__1145_ vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
XFILL_2__1214_ vdd gnd FILL
X_1340_ _1405_/C _1375_/B _1375_/A _1347_/A vdd gnd AOI21X1
X_1271_ _1515_/A _1422_/A _1274_/B vdd gnd XOR2X1
XFILL_0__1545_ vdd gnd FILL
XFILL_0__1476_ vdd gnd FILL
XFILL93150x70350 vdd gnd FILL
XFILL_1__1723_ vdd gnd FILL
X_1607_ _1781_/A _918_/C _1608_/C vdd gnd NAND2X1
X_1469_ _1510_/B _1473_/A _1470_/C vdd gnd NAND2X1
X_1538_ _1538_/A _1538_/B _1538_/C _1562_/A vdd gnd AOI21X1
XFILL_1__1654_ vdd gnd FILL
XFILL_1__1585_ vdd gnd FILL
XFILL_2__976_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
X_982_ _982_/A _982_/B _982_/C _982_/Y vdd gnd OAI21X1
XFILL_2__1763_ vdd gnd FILL
XFILL_2__1694_ vdd gnd FILL
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1261_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_2__1059_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
XFILL_1__994_ vdd gnd FILL
X_1323_ _1379_/A _1323_/B _1323_/C _1326_/C vdd gnd NAND3X1
X_1185_ _960_/A _1361_/A _1185_/C _1190_/C vdd gnd OAI21X1
X_1254_ _1339_/B _1299_/C _1339_/A _1350_/B vdd gnd NAND3X1
XFILL_1__1370_ vdd gnd FILL
XFILL93150x82050 vdd gnd FILL
XFILL_0__1528_ vdd gnd FILL
XFILL_0__1459_ vdd gnd FILL
XFILL_1__1706_ vdd gnd FILL
XFILL_1__1637_ vdd gnd FILL
XFILL_1__1499_ vdd gnd FILL
XFILL_1__1568_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
XFILL_2__1815_ vdd gnd FILL
X_965_ _986_/A _986_/D _992_/A vdd gnd NAND2X1
XFILL_2__1677_ vdd gnd FILL
XFILL_2__1746_ vdd gnd FILL
X_896_ _898_/B _896_/B _896_/Y vdd gnd NAND2X1
XFILL_3__1022_ vdd gnd FILL
XFILL_0__1313_ vdd gnd FILL
XFILL_0__1244_ vdd gnd FILL
XFILL_0__1175_ vdd gnd FILL
XFILL_3__1786_ vdd gnd FILL
XFILL_1__977_ vdd gnd FILL
X_1306_ _1373_/B _1373_/A _1405_/A vdd gnd XNOR2X1
X_1168_ _1679_/A _962_/B _964_/A _978_/B _1184_/A vdd gnd AOI22X1
X_1237_ _1237_/A _1237_/B _1237_/C _1329_/A vdd gnd OAI21X1
X_1099_ _1212_/A _1099_/B _1099_/C _1105_/B vdd gnd NAND3X1
XFILL_1__1353_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
XFILL_1__1284_ vdd gnd FILL
XFILL_2__1600_ vdd gnd FILL
XFILL_2__1531_ vdd gnd FILL
XFILL_2__1462_ vdd gnd FILL
XFILL91950x11850 vdd gnd FILL
XFILL_2__1393_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
XFILL_0__1793_ vdd gnd FILL
XFILL_2__1729_ vdd gnd FILL
XFILL_1__900_ vdd gnd FILL
X_948_ _948_/A _949_/B _949_/C vdd gnd NAND2X1
XFILL_3__1571_ vdd gnd FILL
X_1022_ _985_/C _1325_/B _1088_/A vdd gnd NAND2X1
XFILL_0__1227_ vdd gnd FILL
X_1786_ _1809_/A _1809_/C _1803_/C _1804_/A vdd gnd OAI21X1
XFILL_0__1158_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
XFILL_3__1769_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_2__1514_ vdd gnd FILL
XFILL_2__1445_ vdd gnd FILL
XFILL_2__1376_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
X_1640_ _1684_/D _1661_/A vdd gnd INVX1
XFILL_0__1012_ vdd gnd FILL
X_1571_ _1583_/C _1572_/C vdd gnd INVX1
XFILL_0__1776_ vdd gnd FILL
XFILL_3__1554_ vdd gnd FILL
XFILL_3__1485_ vdd gnd FILL
X_1005_ _1005_/A _1005_/B _1005_/C _1063_/C vdd gnd NAND3X1
XFILL_1__1121_ vdd gnd FILL
XFILL_1__1052_ vdd gnd FILL
X_1769_ _1769_/A _1769_/B _1769_/C _1770_/B vdd gnd AOI21X1
XFILL_2__1230_ vdd gnd FILL
XFILL_0__901_ vdd gnd FILL
XFILL_2__1092_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_2__1161_ vdd gnd FILL
XFILL91950x35250 vdd gnd FILL
XFILL_2__1359_ vdd gnd FILL
XFILL_2__1428_ vdd gnd FILL
XFILL_0__1561_ vdd gnd FILL
XFILL_0__1492_ vdd gnd FILL
X_1554_ _949_/A _1554_/B _915_/A _1555_/B vdd gnd AOI21X1
XFILL_2_BUFX2_insert35 vdd gnd FILL
XFILL_2_BUFX2_insert24 vdd gnd FILL
XFILL_2_BUFX2_insert13 vdd gnd FILL
X_1485_ _1485_/A _899_/A _911_/A _1486_/D vdd gnd AOI21X1
X_1623_ _1623_/D vdd _1624_/R _1624_/CLK _1824_/A vdd gnd DFFSR
.ends

