VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_wrapper
  CLASS BLOCK ;
  FOREIGN ALU_wrapper ;
  ORIGIN 6.000 6.000 ;
  SIZE 948.000 BY 951.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 936.450 899.700 945.450 938.700 ;
        RECT 0.600 897.300 945.450 899.700 ;
        RECT 936.450 821.700 945.450 897.300 ;
        RECT 0.600 819.300 945.450 821.700 ;
        RECT 936.450 743.700 945.450 819.300 ;
        RECT 0.600 741.300 945.450 743.700 ;
        RECT 936.450 665.700 945.450 741.300 ;
        RECT 0.600 663.300 945.450 665.700 ;
        RECT 936.450 587.700 945.450 663.300 ;
        RECT 0.600 585.300 945.450 587.700 ;
        RECT 936.450 509.700 945.450 585.300 ;
        RECT 0.600 507.300 945.450 509.700 ;
        RECT 936.450 431.700 945.450 507.300 ;
        RECT 0.600 429.300 945.450 431.700 ;
        RECT 936.450 353.700 945.450 429.300 ;
        RECT 0.600 351.300 945.450 353.700 ;
        RECT 936.450 275.700 945.450 351.300 ;
        RECT 0.600 273.300 945.450 275.700 ;
        RECT 936.450 197.700 945.450 273.300 ;
        RECT 0.600 195.300 945.450 197.700 ;
        RECT 936.450 119.700 945.450 195.300 ;
        RECT 0.600 117.300 945.450 119.700 ;
        RECT 936.450 41.700 945.450 117.300 ;
        RECT 0.600 39.300 945.450 41.700 ;
        RECT 936.450 0.300 945.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 936.300 935.400 938.700 ;
        RECT -9.450 860.700 -0.450 936.300 ;
        RECT -9.450 858.300 935.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT -9.450 780.300 935.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT -9.450 702.300 935.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 190.950 700.950 193.050 702.300 ;
        RECT 298.950 700.950 301.050 702.300 ;
        RECT 511.950 700.950 514.050 702.300 ;
        RECT -9.450 624.300 935.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 238.950 622.950 241.050 624.300 ;
        RECT 259.950 622.950 262.050 624.300 ;
        RECT 430.950 622.950 433.050 624.300 ;
        RECT 529.950 622.950 532.050 624.300 ;
        RECT 553.950 622.800 556.050 624.300 ;
        RECT 429.000 606.450 433.050 607.050 ;
        RECT 428.550 604.950 433.050 606.450 ;
        RECT 553.950 606.450 558.000 607.050 ;
        RECT 553.950 604.950 558.450 606.450 ;
        RECT 428.550 601.050 429.450 604.950 ;
        RECT 557.550 601.050 558.450 604.950 ;
        RECT 428.550 599.550 433.050 601.050 ;
        RECT 557.550 599.550 562.050 601.050 ;
        RECT 429.000 598.950 433.050 599.550 ;
        RECT 558.000 598.950 562.050 599.550 ;
        RECT -9.450 546.300 935.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 73.950 544.950 76.050 546.300 ;
        RECT 292.950 544.950 295.050 546.300 ;
        RECT 589.950 544.950 592.050 546.300 ;
        RECT -9.450 468.300 935.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 118.950 466.950 121.050 468.300 ;
        RECT 410.550 466.050 411.450 468.300 ;
        RECT 496.950 466.950 499.050 468.300 ;
        RECT 520.950 466.950 523.050 468.300 ;
        RECT 406.950 464.550 411.450 466.050 ;
        RECT 406.950 463.950 411.000 464.550 ;
        RECT 118.950 392.700 121.500 394.050 ;
        RECT -9.450 390.300 935.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 49.950 388.950 52.050 390.300 ;
        RECT 166.950 388.950 169.050 390.300 ;
        RECT 244.950 388.950 247.050 390.300 ;
        RECT 304.950 388.950 307.050 390.300 ;
        RECT 355.950 388.950 358.050 390.300 ;
        RECT -9.450 312.300 935.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 16.950 310.950 19.050 312.300 ;
        RECT 160.950 310.950 163.050 312.300 ;
        RECT -9.450 234.300 935.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 80.550 232.050 81.450 234.300 ;
        RECT 187.950 232.950 190.050 234.300 ;
        RECT 76.950 230.550 81.450 232.050 ;
        RECT 76.950 229.950 81.000 230.550 ;
        RECT -9.450 156.300 935.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT -9.450 78.300 935.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 935.400 2.700 ;
      LAYER metal2 ;
        RECT 190.950 697.950 193.050 703.050 ;
        RECT 298.950 700.950 301.050 703.050 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 223.950 697.950 226.050 700.050 ;
        RECT 221.400 681.450 222.600 682.650 ;
        RECT 224.400 681.450 225.450 697.950 ;
        RECT 299.400 685.050 300.450 700.950 ;
        RECT 298.950 682.950 301.050 685.050 ;
        RECT 329.400 681.900 330.600 682.650 ;
        RECT 221.400 680.400 225.450 681.450 ;
        RECT 328.950 679.800 331.050 681.900 ;
        RECT 512.400 676.050 513.450 700.950 ;
        RECT 505.950 673.950 508.050 676.050 ;
        RECT 511.950 673.950 514.050 676.050 ;
        RECT 506.400 648.600 507.450 673.950 ;
        RECT 257.400 648.450 258.600 648.600 ;
        RECT 257.400 647.400 261.450 648.450 ;
        RECT 257.400 646.350 258.600 647.400 ;
        RECT 260.400 625.050 261.450 647.400 ;
        RECT 506.400 646.350 507.600 648.600 ;
        RECT 238.950 622.950 241.050 625.050 ;
        RECT 259.950 622.950 262.050 625.050 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 529.950 622.950 532.050 625.050 ;
        RECT 239.400 570.600 240.450 622.950 ;
        RECT 431.400 607.050 432.450 622.950 ;
        RECT 430.950 604.950 433.050 607.050 ;
        RECT 518.400 603.900 519.600 604.650 ;
        RECT 530.400 604.050 531.450 622.950 ;
        RECT 553.950 622.800 556.050 624.900 ;
        RECT 554.400 607.050 555.450 622.800 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 517.950 601.800 520.050 603.900 ;
        RECT 529.950 601.950 532.050 604.050 ;
        RECT 581.400 602.400 582.600 604.650 ;
        RECT 430.950 597.450 433.050 601.050 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 430.950 597.000 435.450 597.450 ;
        RECT 431.400 596.400 435.450 597.000 ;
        RECT 434.400 570.600 435.450 596.400 ;
        RECT 560.400 583.050 561.450 598.950 ;
        RECT 581.400 591.450 582.450 602.400 ;
        RECT 578.400 590.400 582.450 591.450 ;
        RECT 578.400 583.050 579.450 590.400 ;
        RECT 559.950 580.950 562.050 583.050 ;
        RECT 577.950 580.950 580.050 583.050 ;
        RECT 239.400 568.350 240.600 570.600 ;
        RECT 434.400 568.350 435.600 570.600 ;
        RECT 73.950 544.950 76.050 547.050 ;
        RECT 11.400 524.400 12.600 526.650 ;
        RECT 11.400 507.450 12.450 524.400 ;
        RECT 11.400 506.400 15.450 507.450 ;
        RECT 14.400 502.050 15.450 506.400 ;
        RECT 74.400 502.050 75.450 544.950 ;
        RECT 292.950 541.950 295.050 547.050 ;
        RECT 589.950 544.950 592.050 547.050 ;
        RECT 316.950 541.950 319.050 544.050 ;
        RECT 317.400 532.050 318.450 541.950 ;
        RECT 590.400 538.050 591.450 544.950 ;
        RECT 529.950 534.450 532.050 538.050 ;
        RECT 589.950 535.950 592.050 538.050 ;
        RECT 527.400 534.000 532.050 534.450 ;
        RECT 527.400 533.400 531.450 534.000 ;
        RECT 316.950 529.950 319.050 532.050 ;
        RECT 334.950 529.950 337.050 532.050 ;
        RECT 320.400 525.900 321.600 526.650 ;
        RECT 335.400 526.050 336.450 529.950 ;
        RECT 319.950 523.800 322.050 525.900 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 512.400 525.900 513.600 526.650 ;
        RECT 527.400 526.050 528.450 533.400 ;
        RECT 511.950 523.800 514.050 525.900 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 13.950 499.950 16.050 502.050 ;
        RECT 73.950 499.950 76.050 502.050 ;
        RECT 74.400 492.450 75.450 499.950 ;
        RECT 71.400 491.400 75.450 492.450 ;
        RECT 118.950 492.600 123.000 493.050 ;
        RECT 26.400 486.000 27.600 487.650 ;
        RECT 25.950 481.950 28.050 486.000 ;
        RECT 71.400 484.050 72.450 491.400 ;
        RECT 118.950 490.950 123.600 492.600 ;
        RECT 499.950 491.100 502.050 493.200 ;
        RECT 122.400 490.350 123.600 490.950 ;
        RECT 500.400 490.350 501.600 491.100 ;
        RECT 118.950 484.950 121.050 487.050 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 119.400 469.050 120.450 484.950 ;
        RECT 520.950 484.650 523.050 486.750 ;
        RECT 521.400 469.050 522.450 484.650 ;
        RECT 118.950 466.950 121.050 469.050 ;
        RECT 496.950 466.950 499.050 469.050 ;
        RECT 520.950 466.950 523.050 469.050 ;
        RECT 406.950 463.950 409.050 466.050 ;
        RECT 77.400 446.400 78.600 448.650 ;
        RECT 140.400 446.400 141.600 448.650 ;
        RECT 257.400 446.400 258.600 448.650 ;
        RECT 278.400 446.400 279.600 448.650 ;
        RECT 347.400 446.400 348.600 448.650 ;
        RECT 77.400 421.050 78.450 446.400 ;
        RECT 140.400 444.450 141.450 446.400 ;
        RECT 137.400 443.400 141.450 444.450 ;
        RECT 137.400 424.050 138.450 443.400 ;
        RECT 118.950 421.950 121.050 424.050 ;
        RECT 136.950 421.950 139.050 424.050 ;
        RECT 64.950 418.950 67.050 421.050 ;
        RECT 76.950 418.950 79.050 421.050 ;
        RECT 65.400 394.050 66.450 418.950 ;
        RECT 119.400 394.050 120.450 421.950 ;
        RECT 49.950 388.950 52.050 394.050 ;
        RECT 64.950 391.950 67.050 394.050 ;
        RECT 118.950 391.950 121.050 394.050 ;
        RECT 257.400 391.050 258.450 446.400 ;
        RECT 278.400 418.050 279.450 446.400 ;
        RECT 347.400 442.050 348.450 446.400 ;
        RECT 407.400 442.050 408.450 463.950 ;
        RECT 482.400 447.900 483.600 448.650 ;
        RECT 497.400 448.050 498.450 466.950 ;
        RECT 481.950 445.800 484.050 447.900 ;
        RECT 496.950 445.950 499.050 448.050 ;
        RECT 346.950 439.950 349.050 442.050 ;
        RECT 406.950 439.950 409.050 442.050 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 296.400 397.050 297.450 415.950 ;
        RECT 337.950 414.000 340.050 418.050 ;
        RECT 338.400 412.350 339.600 414.000 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 353.400 405.450 354.450 412.950 ;
        RECT 353.400 404.400 357.450 405.450 ;
        RECT 295.950 394.950 298.050 397.050 ;
        RECT 304.950 394.950 307.050 397.050 ;
        RECT 305.400 391.050 306.450 394.950 ;
        RECT 356.400 391.050 357.450 404.400 ;
        RECT 166.950 388.950 169.050 391.050 ;
        RECT 244.950 388.950 250.050 391.050 ;
        RECT 256.950 388.950 259.050 391.050 ;
        RECT 304.950 388.950 307.050 391.050 ;
        RECT 355.950 388.950 358.050 391.050 ;
        RECT 167.400 373.050 168.450 388.950 ;
        RECT 166.950 370.950 169.050 373.050 ;
        RECT 125.400 369.900 126.600 370.650 ;
        RECT 124.950 367.800 127.050 369.900 ;
        RECT 116.400 336.450 117.600 336.600 ;
        RECT 113.400 335.400 117.600 336.450 ;
        RECT 113.400 316.050 114.450 335.400 ;
        RECT 116.400 334.350 117.600 335.400 ;
        RECT 112.950 313.950 115.050 316.050 ;
        RECT 4.950 307.950 7.050 310.050 ;
        RECT 16.950 307.950 19.050 313.050 ;
        RECT 5.400 283.050 6.450 307.950 ;
        RECT 113.400 291.450 114.450 313.950 ;
        RECT 160.950 310.950 163.050 316.050 ;
        RECT 116.400 291.450 117.600 292.650 ;
        RECT 113.400 290.400 117.600 291.450 ;
        RECT 4.950 280.950 7.050 283.050 ;
        RECT 58.950 280.950 61.050 283.050 ;
        RECT 59.400 258.600 60.450 280.950 ;
        RECT 59.400 256.350 60.600 258.600 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 76.950 229.950 79.050 232.050 ;
        RECT 59.400 213.900 60.600 214.650 ;
        RECT 77.400 214.050 78.450 229.950 ;
        RECT 58.950 211.800 61.050 213.900 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 146.400 213.900 147.600 214.650 ;
        RECT 188.400 214.050 189.450 232.950 ;
        RECT 145.950 211.800 148.050 213.900 ;
        RECT 187.950 211.950 190.050 214.050 ;
      LAYER metal3 ;
        RECT 190.950 699.600 193.050 700.050 ;
        RECT 223.950 699.600 226.050 700.050 ;
        RECT 190.950 698.400 226.050 699.600 ;
        RECT 190.950 697.950 193.050 698.400 ;
        RECT 223.950 697.950 226.050 698.400 ;
        RECT 298.950 681.600 301.050 685.050 ;
        RECT 328.950 681.600 331.050 681.900 ;
        RECT 298.950 681.000 331.050 681.600 ;
        RECT 299.400 680.400 331.050 681.000 ;
        RECT 328.950 679.800 331.050 680.400 ;
        RECT 505.950 675.600 508.050 676.050 ;
        RECT 511.950 675.600 514.050 676.050 ;
        RECT 505.950 674.400 514.050 675.600 ;
        RECT 505.950 673.950 508.050 674.400 ;
        RECT 511.950 673.950 514.050 674.400 ;
        RECT 517.950 603.600 520.050 603.900 ;
        RECT 529.950 603.600 532.050 604.050 ;
        RECT 517.950 602.400 532.050 603.600 ;
        RECT 517.950 601.800 520.050 602.400 ;
        RECT 529.950 601.950 532.050 602.400 ;
        RECT 559.950 582.600 562.050 583.050 ;
        RECT 577.950 582.600 580.050 583.050 ;
        RECT 559.950 581.400 580.050 582.600 ;
        RECT 559.950 580.950 562.050 581.400 ;
        RECT 577.950 580.950 580.050 581.400 ;
        RECT 292.950 543.600 295.050 544.050 ;
        RECT 316.950 543.600 319.050 544.050 ;
        RECT 292.950 542.400 319.050 543.600 ;
        RECT 292.950 541.950 295.050 542.400 ;
        RECT 316.950 541.950 319.050 542.400 ;
        RECT 529.950 537.600 532.050 538.050 ;
        RECT 589.950 537.600 592.050 538.050 ;
        RECT 529.950 536.400 592.050 537.600 ;
        RECT 529.950 535.950 532.050 536.400 ;
        RECT 589.950 535.950 592.050 536.400 ;
        RECT 316.950 531.600 319.050 532.050 ;
        RECT 334.950 531.600 337.050 532.050 ;
        RECT 316.950 530.400 337.050 531.600 ;
        RECT 316.950 529.950 319.050 530.400 ;
        RECT 334.950 529.950 337.050 530.400 ;
        RECT 319.950 525.600 322.050 525.900 ;
        RECT 334.950 525.600 337.050 526.050 ;
        RECT 319.950 524.400 337.050 525.600 ;
        RECT 319.950 523.800 322.050 524.400 ;
        RECT 334.950 523.950 337.050 524.400 ;
        RECT 511.950 525.600 514.050 525.900 ;
        RECT 526.950 525.600 529.050 526.050 ;
        RECT 511.950 524.400 529.050 525.600 ;
        RECT 511.950 523.800 514.050 524.400 ;
        RECT 526.950 523.950 529.050 524.400 ;
        RECT 13.950 501.600 16.050 502.050 ;
        RECT 73.950 501.600 76.050 502.050 ;
        RECT 13.950 500.400 76.050 501.600 ;
        RECT 13.950 499.950 16.050 500.400 ;
        RECT 73.950 499.950 76.050 500.400 ;
        RECT 118.950 490.950 121.050 493.050 ;
        RECT 499.950 492.600 502.050 493.200 ;
        RECT 499.950 491.400 519.600 492.600 ;
        RECT 499.950 491.100 502.050 491.400 ;
        RECT 119.400 487.050 120.600 490.950 ;
        RECT 518.400 487.050 519.600 491.400 ;
        RECT 118.950 484.950 121.050 487.050 ;
        RECT 518.400 486.750 522.000 487.050 ;
        RECT 518.400 485.400 523.050 486.750 ;
        RECT 519.000 484.950 523.050 485.400 ;
        RECT 520.950 484.650 523.050 484.950 ;
        RECT 25.950 483.600 28.050 484.050 ;
        RECT 70.950 483.600 73.050 484.050 ;
        RECT 25.950 482.400 73.050 483.600 ;
        RECT 25.950 481.950 28.050 482.400 ;
        RECT 70.950 481.950 73.050 482.400 ;
        RECT 481.950 447.600 484.050 447.900 ;
        RECT 496.950 447.600 499.050 448.050 ;
        RECT 481.950 446.400 499.050 447.600 ;
        RECT 481.950 445.800 484.050 446.400 ;
        RECT 496.950 445.950 499.050 446.400 ;
        RECT 346.950 441.600 349.050 442.050 ;
        RECT 406.950 441.600 409.050 442.050 ;
        RECT 346.950 440.400 409.050 441.600 ;
        RECT 346.950 439.950 349.050 440.400 ;
        RECT 406.950 439.950 409.050 440.400 ;
        RECT 118.950 423.600 121.050 424.050 ;
        RECT 136.950 423.600 139.050 424.050 ;
        RECT 118.950 422.400 139.050 423.600 ;
        RECT 118.950 421.950 121.050 422.400 ;
        RECT 136.950 421.950 139.050 422.400 ;
        RECT 64.950 420.600 67.050 421.050 ;
        RECT 76.950 420.600 79.050 421.050 ;
        RECT 64.950 419.400 79.050 420.600 ;
        RECT 64.950 418.950 67.050 419.400 ;
        RECT 76.950 418.950 79.050 419.400 ;
        RECT 277.950 417.600 280.050 418.050 ;
        RECT 295.950 417.600 298.050 418.050 ;
        RECT 277.950 416.400 298.050 417.600 ;
        RECT 277.950 415.950 280.050 416.400 ;
        RECT 295.950 415.950 298.050 416.400 ;
        RECT 337.950 417.600 340.050 418.050 ;
        RECT 337.950 417.000 354.600 417.600 ;
        RECT 337.950 416.400 355.050 417.000 ;
        RECT 337.950 415.950 340.050 416.400 ;
        RECT 352.950 412.950 355.050 416.400 ;
        RECT 295.950 396.600 298.050 397.050 ;
        RECT 304.950 396.600 307.050 397.050 ;
        RECT 295.950 395.400 307.050 396.600 ;
        RECT 295.950 394.950 298.050 395.400 ;
        RECT 304.950 394.950 307.050 395.400 ;
        RECT 49.950 393.600 52.050 394.050 ;
        RECT 64.950 393.600 67.050 394.050 ;
        RECT 49.950 392.400 67.050 393.600 ;
        RECT 49.950 391.950 52.050 392.400 ;
        RECT 64.950 391.950 67.050 392.400 ;
        RECT 247.950 390.600 250.050 391.050 ;
        RECT 256.950 390.600 259.050 391.050 ;
        RECT 247.950 389.400 259.050 390.600 ;
        RECT 247.950 388.950 250.050 389.400 ;
        RECT 256.950 388.950 259.050 389.400 ;
        RECT 124.950 369.600 127.050 369.900 ;
        RECT 166.950 369.600 169.050 373.050 ;
        RECT 124.950 369.000 169.050 369.600 ;
        RECT 124.950 368.400 168.600 369.000 ;
        RECT 124.950 367.800 127.050 368.400 ;
        RECT 112.950 315.600 115.050 316.050 ;
        RECT 160.950 315.600 163.050 316.050 ;
        RECT 112.950 314.400 163.050 315.600 ;
        RECT 112.950 313.950 115.050 314.400 ;
        RECT 160.950 313.950 163.050 314.400 ;
        RECT 4.950 309.600 7.050 310.050 ;
        RECT 16.950 309.600 19.050 310.050 ;
        RECT 4.950 308.400 19.050 309.600 ;
        RECT 4.950 307.950 7.050 308.400 ;
        RECT 16.950 307.950 19.050 308.400 ;
        RECT 4.950 282.600 7.050 283.050 ;
        RECT 58.950 282.600 61.050 283.050 ;
        RECT 4.950 281.400 61.050 282.600 ;
        RECT 4.950 280.950 7.050 281.400 ;
        RECT 58.950 280.950 61.050 281.400 ;
        RECT 58.950 213.600 61.050 213.900 ;
        RECT 76.950 213.600 79.050 214.050 ;
        RECT 58.950 212.400 79.050 213.600 ;
        RECT 58.950 211.800 61.050 212.400 ;
        RECT 76.950 211.950 79.050 212.400 ;
        RECT 145.950 213.600 148.050 213.900 ;
        RECT 187.950 213.600 190.050 214.050 ;
        RECT 145.950 212.400 190.050 213.600 ;
        RECT 145.950 211.800 148.050 212.400 ;
        RECT 187.950 211.950 190.050 212.400 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal1 ;
        RECT 256.950 600.450 259.050 601.050 ;
        RECT 256.950 599.550 264.450 600.450 ;
        RECT 256.950 598.950 259.050 599.550 ;
        RECT 263.550 595.050 264.450 599.550 ;
        RECT 262.950 592.950 265.050 595.050 ;
        RECT 349.950 189.450 352.050 190.050 ;
        RECT 358.950 189.450 361.050 190.050 ;
        RECT 349.950 188.550 361.050 189.450 ;
        RECT 349.950 187.950 352.050 188.550 ;
        RECT 358.950 187.950 361.050 188.550 ;
      LAYER metal2 ;
        RECT 140.400 937.050 141.450 945.450 ;
        RECT 139.950 934.950 142.050 937.050 ;
        RECT 283.950 934.950 286.050 937.050 ;
        RECT 284.400 912.450 285.450 934.950 ;
        RECT 281.400 911.400 285.450 912.450 ;
        RECT 281.400 834.450 282.450 911.400 ;
        RECT 278.400 833.400 282.450 834.450 ;
        RECT 278.400 822.450 279.450 833.400 ;
        RECT 275.400 821.400 279.450 822.450 ;
        RECT 275.400 793.050 276.450 821.400 ;
        RECT 268.950 790.950 271.050 793.050 ;
        RECT 274.950 790.950 277.050 793.050 ;
        RECT 269.400 754.050 270.450 790.950 ;
        RECT 262.950 751.950 265.050 754.050 ;
        RECT 268.950 751.950 271.050 754.050 ;
        RECT 4.950 728.100 7.050 730.200 ;
        RECT 10.950 728.100 13.050 730.200 ;
        RECT 5.400 685.050 6.450 728.100 ;
        RECT 11.400 727.350 12.600 728.100 ;
        RECT 163.950 727.950 166.050 730.050 ;
        RECT 169.950 728.100 172.050 730.200 ;
        RECT 164.400 703.050 165.450 727.950 ;
        RECT 170.400 727.350 171.600 728.100 ;
        RECT 263.400 703.050 264.450 751.950 ;
        RECT 163.950 700.950 166.050 703.050 ;
        RECT 262.950 700.950 265.050 703.050 ;
        RECT 164.400 688.200 165.450 700.950 ;
        RECT 385.950 688.950 388.050 691.050 ;
        RECT 418.950 688.950 421.050 691.050 ;
        RECT 517.950 688.950 520.050 691.050 ;
        RECT 538.950 688.950 541.050 691.050 ;
        RECT 130.950 685.950 133.050 688.050 ;
        RECT 163.950 686.100 166.050 688.200 ;
        RECT 172.950 685.950 175.050 688.050 ;
        RECT 4.950 682.950 7.050 685.050 ;
        RECT 13.950 683.100 16.050 685.200 ;
        RECT 25.950 683.100 28.050 685.200 ;
        RECT 14.400 682.350 15.600 683.100 ;
        RECT 26.400 670.050 27.450 683.100 ;
        RECT 59.400 677.400 60.600 679.650 ;
        RECT 59.400 670.050 60.450 677.400 ;
        RECT 131.400 670.050 132.450 685.950 ;
        RECT 161.400 677.400 162.600 679.650 ;
        RECT 161.400 670.050 162.450 677.400 ;
        RECT 173.400 670.050 174.450 685.950 ;
        RECT 25.950 667.950 28.050 670.050 ;
        RECT 58.950 667.950 61.050 670.050 ;
        RECT 130.950 667.950 133.050 670.050 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 172.950 669.450 175.050 670.050 ;
        RECT 170.400 668.400 175.050 669.450 ;
        RECT 170.400 640.050 171.450 668.400 ;
        RECT 172.950 667.950 175.050 668.400 ;
        RECT 386.400 655.050 387.450 688.950 ;
        RECT 419.400 684.600 420.450 688.950 ;
        RECT 419.400 682.350 420.600 684.600 ;
        RECT 518.400 684.450 519.450 688.950 ;
        RECT 521.400 684.450 522.600 684.600 ;
        RECT 518.400 683.400 522.600 684.450 ;
        RECT 521.400 682.350 522.600 683.400 ;
        RECT 539.400 673.050 540.450 688.950 ;
        RECT 538.950 670.950 541.050 673.050 ;
        RECT 556.950 670.950 559.050 673.050 ;
        RECT 343.950 652.950 346.050 655.050 ;
        RECT 385.950 652.950 388.050 655.050 ;
        RECT 344.400 649.050 345.450 652.950 ;
        RECT 557.400 649.050 558.450 670.950 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 556.950 646.950 559.050 649.050 ;
        RECT 206.400 645.900 207.600 646.650 ;
        RECT 335.400 645.900 336.600 646.650 ;
        RECT 193.950 643.800 196.050 645.900 ;
        RECT 205.950 643.800 208.050 645.900 ;
        RECT 334.950 643.800 337.050 645.900 ;
        RECT 586.950 643.950 589.050 646.050 ;
        RECT 194.400 640.050 195.450 643.800 ;
        RECT 169.950 637.950 172.050 640.050 ;
        RECT 193.950 637.950 196.050 640.050 ;
        RECT 206.400 631.050 207.450 643.800 ;
        RECT 205.950 628.950 208.050 631.050 ;
        RECT 253.950 628.950 256.050 631.050 ;
        RECT 254.400 625.050 255.450 628.950 ;
        RECT 335.400 625.050 336.450 643.800 ;
        RECT 587.400 625.050 588.450 643.950 ;
        RECT 694.950 631.950 697.050 634.050 ;
        RECT 709.950 631.950 712.050 634.050 ;
        RECT 695.400 625.050 696.450 631.950 ;
        RECT 253.950 622.950 256.050 625.050 ;
        RECT 334.950 622.950 337.050 625.050 ;
        RECT 586.950 622.950 589.050 625.050 ;
        RECT 694.950 622.950 697.050 625.050 ;
        RECT 254.400 606.450 255.450 622.950 ;
        RECT 710.400 607.200 711.450 631.950 ;
        RECT 254.400 605.400 258.450 606.450 ;
        RECT 257.400 601.050 258.450 605.400 ;
        RECT 703.950 604.950 706.050 607.050 ;
        RECT 709.950 605.100 712.050 607.200 ;
        RECT 256.950 598.950 259.050 601.050 ;
        RECT 262.950 592.950 265.050 595.050 ;
        RECT 263.400 586.050 264.450 592.950 ;
        RECT 262.950 583.950 265.050 586.050 ;
        RECT 283.800 583.950 285.900 586.050 ;
        RECT 284.400 579.450 285.450 583.950 ;
        RECT 284.400 578.400 288.450 579.450 ;
        RECT 287.400 550.050 288.450 578.400 ;
        RECT 274.950 547.950 277.050 550.050 ;
        RECT 286.950 547.950 289.050 550.050 ;
        RECT 704.400 549.450 705.450 604.950 ;
        RECT 710.400 604.350 711.600 605.100 ;
        RECT 704.400 548.400 708.450 549.450 ;
        RECT 275.400 460.050 276.450 547.950 ;
        RECT 707.400 528.600 708.450 548.400 ;
        RECT 707.400 526.350 708.600 528.600 ;
        RECT 253.950 457.950 256.050 460.050 ;
        RECT 274.950 457.950 277.050 460.050 ;
        RECT 254.400 424.050 255.450 457.950 ;
        RECT 220.950 421.950 223.050 424.050 ;
        RECT 253.950 421.950 256.050 424.050 ;
        RECT 298.950 421.950 301.050 424.050 ;
        RECT 194.400 410.400 195.600 412.650 ;
        RECT 194.400 406.050 195.450 410.400 ;
        RECT 221.400 406.050 222.450 421.950 ;
        RECT 193.950 403.950 196.050 406.050 ;
        RECT 220.950 403.950 223.050 406.050 ;
        RECT 299.400 373.050 300.450 421.950 ;
        RECT 298.950 370.950 301.050 373.050 ;
        RECT 331.950 361.950 334.050 364.050 ;
        RECT 332.400 346.050 333.450 361.950 ;
        RECT 332.400 344.400 337.050 346.050 ;
        RECT 333.000 343.950 337.050 344.400 ;
        RECT 394.800 343.950 396.900 346.050 ;
        RECT 395.400 340.050 396.450 343.950 ;
        RECT 394.950 337.950 397.050 340.050 ;
        RECT 394.950 331.950 397.050 334.050 ;
        RECT 395.400 301.050 396.450 331.950 ;
        RECT 394.950 298.950 397.050 301.050 ;
        RECT 409.950 298.950 412.050 301.050 ;
        RECT 410.400 261.450 411.450 298.950 ;
        RECT 407.400 260.400 411.450 261.450 ;
        RECT 407.400 255.900 408.450 260.400 ;
        RECT 413.400 255.900 414.600 256.650 ;
        RECT 406.950 253.800 409.050 255.900 ;
        RECT 412.950 253.800 415.050 255.900 ;
        RECT 407.400 229.050 408.450 253.800 ;
        RECT 349.950 226.950 352.050 229.050 ;
        RECT 355.950 226.950 358.050 229.050 ;
        RECT 406.950 226.950 409.050 229.050 ;
        RECT 350.400 190.050 351.450 226.950 ;
        RECT 356.400 216.600 357.450 226.950 ;
        RECT 356.400 214.350 357.600 216.600 ;
        RECT 349.950 187.950 352.050 190.050 ;
        RECT 358.950 187.950 361.050 190.050 ;
        RECT 317.400 176.400 318.600 178.650 ;
        RECT 317.400 160.050 318.450 176.400 ;
        RECT 359.400 160.050 360.450 187.950 ;
        RECT 52.950 157.950 55.050 160.050 ;
        RECT 316.950 157.950 319.050 160.050 ;
        RECT 358.950 157.950 361.050 160.050 ;
        RECT 53.400 138.600 54.450 157.950 ;
        RECT 53.400 136.350 54.600 138.600 ;
      LAYER metal3 ;
        RECT 139.950 936.600 142.050 937.050 ;
        RECT 283.950 936.600 286.050 937.050 ;
        RECT 139.950 935.400 286.050 936.600 ;
        RECT 139.950 934.950 142.050 935.400 ;
        RECT 283.950 934.950 286.050 935.400 ;
        RECT 268.950 792.600 271.050 793.050 ;
        RECT 274.950 792.600 277.050 793.050 ;
        RECT 268.950 791.400 277.050 792.600 ;
        RECT 268.950 790.950 271.050 791.400 ;
        RECT 274.950 790.950 277.050 791.400 ;
        RECT 262.950 753.600 265.050 754.050 ;
        RECT 268.950 753.600 271.050 754.050 ;
        RECT 262.950 752.400 271.050 753.600 ;
        RECT 262.950 751.950 265.050 752.400 ;
        RECT 268.950 751.950 271.050 752.400 ;
        RECT 4.950 729.750 7.050 730.200 ;
        RECT 10.950 729.750 13.050 730.200 ;
        RECT 4.950 728.550 13.050 729.750 ;
        RECT 4.950 728.100 7.050 728.550 ;
        RECT 10.950 728.100 13.050 728.550 ;
        RECT 163.950 729.600 166.050 730.050 ;
        RECT 169.950 729.600 172.050 730.200 ;
        RECT 163.950 728.400 172.050 729.600 ;
        RECT 163.950 727.950 166.050 728.400 ;
        RECT 169.950 728.100 172.050 728.400 ;
        RECT 163.950 702.600 166.050 703.050 ;
        RECT 262.950 702.600 265.050 703.050 ;
        RECT 163.950 701.400 265.050 702.600 ;
        RECT 163.950 700.950 166.050 701.400 ;
        RECT 262.950 700.950 265.050 701.400 ;
        RECT 385.950 690.600 388.050 691.050 ;
        RECT 418.950 690.600 421.050 691.050 ;
        RECT 517.950 690.600 520.050 691.050 ;
        RECT 538.950 690.600 541.050 691.050 ;
        RECT 385.950 689.400 541.050 690.600 ;
        RECT 385.950 688.950 388.050 689.400 ;
        RECT 418.950 688.950 421.050 689.400 ;
        RECT 517.950 688.950 520.050 689.400 ;
        RECT 538.950 688.950 541.050 689.400 ;
        RECT 130.950 687.600 133.050 688.050 ;
        RECT 163.950 687.600 166.050 688.200 ;
        RECT 172.950 687.600 175.050 688.050 ;
        RECT 130.950 686.400 175.050 687.600 ;
        RECT 130.950 685.950 133.050 686.400 ;
        RECT 163.950 686.100 166.050 686.400 ;
        RECT 172.950 685.950 175.050 686.400 ;
        RECT 4.950 684.600 7.050 685.050 ;
        RECT 13.950 684.750 16.050 685.200 ;
        RECT 25.950 684.750 28.050 685.200 ;
        RECT 13.950 684.600 28.050 684.750 ;
        RECT 4.950 683.550 28.050 684.600 ;
        RECT 4.950 683.400 16.050 683.550 ;
        RECT 4.950 682.950 7.050 683.400 ;
        RECT 13.950 683.100 16.050 683.400 ;
        RECT 25.950 683.100 28.050 683.550 ;
        RECT 538.950 672.600 541.050 673.050 ;
        RECT 556.950 672.600 559.050 673.050 ;
        RECT 538.950 671.400 559.050 672.600 ;
        RECT 538.950 670.950 541.050 671.400 ;
        RECT 556.950 670.950 559.050 671.400 ;
        RECT 25.950 669.600 28.050 670.050 ;
        RECT 58.950 669.600 61.050 670.050 ;
        RECT 130.950 669.600 133.050 670.050 ;
        RECT 25.950 668.400 133.050 669.600 ;
        RECT 25.950 667.950 28.050 668.400 ;
        RECT 58.950 667.950 61.050 668.400 ;
        RECT 130.950 667.950 133.050 668.400 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 172.950 669.600 175.050 670.050 ;
        RECT 160.950 668.400 175.050 669.600 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 172.950 667.950 175.050 668.400 ;
        RECT 343.950 654.600 346.050 655.050 ;
        RECT 385.950 654.600 388.050 655.050 ;
        RECT 343.950 653.400 388.050 654.600 ;
        RECT 343.950 652.950 346.050 653.400 ;
        RECT 385.950 652.950 388.050 653.400 ;
        RECT 343.950 648.600 346.050 649.050 ;
        RECT 335.400 647.400 346.050 648.600 ;
        RECT 335.400 645.900 336.600 647.400 ;
        RECT 343.950 646.950 346.050 647.400 ;
        RECT 556.950 648.600 559.050 649.050 ;
        RECT 556.950 647.400 585.600 648.600 ;
        RECT 556.950 646.950 559.050 647.400 ;
        RECT 584.400 646.050 585.600 647.400 ;
        RECT 193.950 645.450 196.050 645.900 ;
        RECT 205.950 645.450 208.050 645.900 ;
        RECT 193.950 644.250 208.050 645.450 ;
        RECT 193.950 643.800 196.050 644.250 ;
        RECT 205.950 643.800 208.050 644.250 ;
        RECT 334.950 643.800 337.050 645.900 ;
        RECT 584.400 644.400 589.050 646.050 ;
        RECT 585.000 643.950 589.050 644.400 ;
        RECT 169.950 639.600 172.050 640.050 ;
        RECT 193.950 639.600 196.050 640.050 ;
        RECT 169.950 638.400 196.050 639.600 ;
        RECT 169.950 637.950 172.050 638.400 ;
        RECT 193.950 637.950 196.050 638.400 ;
        RECT 694.950 633.600 697.050 634.050 ;
        RECT 709.950 633.600 712.050 634.050 ;
        RECT 694.950 632.400 712.050 633.600 ;
        RECT 694.950 631.950 697.050 632.400 ;
        RECT 709.950 631.950 712.050 632.400 ;
        RECT 205.950 630.600 208.050 631.050 ;
        RECT 253.950 630.600 256.050 631.050 ;
        RECT 205.950 629.400 256.050 630.600 ;
        RECT 205.950 628.950 208.050 629.400 ;
        RECT 253.950 628.950 256.050 629.400 ;
        RECT 253.950 624.600 256.050 625.050 ;
        RECT 334.950 624.600 337.050 625.050 ;
        RECT 253.950 623.400 337.050 624.600 ;
        RECT 253.950 622.950 256.050 623.400 ;
        RECT 334.950 622.950 337.050 623.400 ;
        RECT 586.950 624.600 589.050 625.050 ;
        RECT 694.950 624.600 697.050 625.050 ;
        RECT 586.950 623.400 697.050 624.600 ;
        RECT 586.950 622.950 589.050 623.400 ;
        RECT 694.950 622.950 697.050 623.400 ;
        RECT 703.950 606.600 706.050 607.050 ;
        RECT 709.950 606.600 712.050 607.200 ;
        RECT 703.950 605.400 712.050 606.600 ;
        RECT 703.950 604.950 706.050 605.400 ;
        RECT 709.950 605.100 712.050 605.400 ;
        RECT 262.950 585.600 265.050 586.050 ;
        RECT 283.800 585.600 285.900 586.050 ;
        RECT 262.950 584.400 285.900 585.600 ;
        RECT 262.950 583.950 265.050 584.400 ;
        RECT 283.800 583.950 285.900 584.400 ;
        RECT 274.950 549.600 277.050 550.050 ;
        RECT 286.950 549.600 289.050 550.050 ;
        RECT 274.950 548.400 289.050 549.600 ;
        RECT 274.950 547.950 277.050 548.400 ;
        RECT 286.950 547.950 289.050 548.400 ;
        RECT 253.950 459.600 256.050 460.050 ;
        RECT 274.950 459.600 277.050 460.050 ;
        RECT 253.950 458.400 277.050 459.600 ;
        RECT 253.950 457.950 256.050 458.400 ;
        RECT 274.950 457.950 277.050 458.400 ;
        RECT 220.950 423.600 223.050 424.050 ;
        RECT 253.950 423.600 256.050 424.050 ;
        RECT 298.950 423.600 301.050 424.050 ;
        RECT 220.950 422.400 301.050 423.600 ;
        RECT 220.950 421.950 223.050 422.400 ;
        RECT 253.950 421.950 256.050 422.400 ;
        RECT 298.950 421.950 301.050 422.400 ;
        RECT 193.950 405.600 196.050 406.050 ;
        RECT 220.950 405.600 223.050 406.050 ;
        RECT 193.950 404.400 223.050 405.600 ;
        RECT 193.950 403.950 196.050 404.400 ;
        RECT 220.950 403.950 223.050 404.400 ;
        RECT 298.950 369.600 301.050 373.050 ;
        RECT 298.950 369.000 333.600 369.600 ;
        RECT 299.400 368.400 333.600 369.000 ;
        RECT 332.400 364.050 333.600 368.400 ;
        RECT 331.950 361.950 334.050 364.050 ;
        RECT 334.950 345.600 337.050 346.050 ;
        RECT 394.800 345.600 396.900 346.050 ;
        RECT 334.950 344.400 396.900 345.600 ;
        RECT 334.950 343.950 337.050 344.400 ;
        RECT 394.800 343.950 396.900 344.400 ;
        RECT 394.950 337.950 397.050 340.050 ;
        RECT 395.400 334.050 396.600 337.950 ;
        RECT 394.950 331.950 397.050 334.050 ;
        RECT 394.950 300.600 397.050 301.050 ;
        RECT 409.950 300.600 412.050 301.050 ;
        RECT 394.950 299.400 412.050 300.600 ;
        RECT 394.950 298.950 397.050 299.400 ;
        RECT 409.950 298.950 412.050 299.400 ;
        RECT 406.950 255.450 409.050 255.900 ;
        RECT 412.950 255.450 415.050 255.900 ;
        RECT 406.950 254.250 415.050 255.450 ;
        RECT 406.950 253.800 409.050 254.250 ;
        RECT 412.950 253.800 415.050 254.250 ;
        RECT 349.950 228.600 352.050 229.050 ;
        RECT 355.950 228.600 358.050 229.050 ;
        RECT 406.950 228.600 409.050 229.050 ;
        RECT 349.950 227.400 409.050 228.600 ;
        RECT 349.950 226.950 352.050 227.400 ;
        RECT 355.950 226.950 358.050 227.400 ;
        RECT 406.950 226.950 409.050 227.400 ;
        RECT 52.950 159.600 55.050 160.050 ;
        RECT 316.950 159.600 319.050 160.050 ;
        RECT 358.950 159.600 361.050 160.050 ;
        RECT 52.950 158.400 361.050 159.600 ;
        RECT 52.950 157.950 55.050 158.400 ;
        RECT 316.950 157.950 319.050 158.400 ;
        RECT 358.950 157.950 361.050 158.400 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal2 ;
        RECT 146.400 865.050 147.450 945.450 ;
        RECT 85.950 862.950 88.050 865.050 ;
        RECT 145.950 862.950 148.050 865.050 ;
        RECT 86.400 841.200 87.450 862.950 ;
        RECT 146.400 850.050 147.450 862.950 ;
        RECT 145.950 847.950 148.050 850.050 ;
        RECT 178.950 847.950 181.050 850.050 ;
        RECT 85.950 839.100 88.050 841.200 ;
        RECT 179.400 841.050 180.450 847.950 ;
        RECT 86.400 838.350 87.600 839.100 ;
        RECT 178.950 838.950 181.050 841.050 ;
        RECT 184.950 839.100 187.050 841.200 ;
        RECT 88.950 832.950 91.050 835.050 ;
        RECT 44.400 800.400 45.600 802.650 ;
        RECT 44.400 796.050 45.450 800.400 ;
        RECT 89.400 796.050 90.450 832.950 ;
        RECT 179.400 807.600 180.450 838.950 ;
        RECT 185.400 838.350 186.600 839.100 ;
        RECT 179.400 805.350 180.600 807.600 ;
        RECT 43.950 793.950 46.050 796.050 ;
        RECT 88.950 793.950 91.050 796.050 ;
        RECT 89.400 772.050 90.450 793.950 ;
        RECT 88.950 769.950 91.050 772.050 ;
        RECT 145.950 769.950 148.050 772.050 ;
        RECT 146.400 739.050 147.450 769.950 ;
        RECT 136.950 736.800 139.050 738.900 ;
        RECT 145.950 736.950 148.050 739.050 ;
        RECT 137.400 684.450 138.450 736.800 ;
        RECT 134.400 683.400 138.450 684.450 ;
        RECT 134.400 673.050 135.450 683.400 ;
        RECT 133.950 670.950 136.050 673.050 ;
        RECT 220.950 667.950 223.050 670.050 ;
        RECT 221.400 651.600 222.450 667.950 ;
        RECT 221.400 649.350 222.600 651.600 ;
      LAYER metal3 ;
        RECT 85.950 864.600 88.050 865.050 ;
        RECT 145.950 864.600 148.050 865.050 ;
        RECT 85.950 863.400 148.050 864.600 ;
        RECT 85.950 862.950 88.050 863.400 ;
        RECT 145.950 862.950 148.050 863.400 ;
        RECT 145.950 849.600 148.050 850.050 ;
        RECT 178.950 849.600 181.050 850.050 ;
        RECT 145.950 848.400 181.050 849.600 ;
        RECT 145.950 847.950 148.050 848.400 ;
        RECT 178.950 847.950 181.050 848.400 ;
        RECT 85.950 839.100 88.050 841.200 ;
        RECT 178.950 840.600 181.050 841.050 ;
        RECT 184.950 840.600 187.050 841.200 ;
        RECT 178.950 839.400 187.050 840.600 ;
        RECT 86.400 837.600 87.600 839.100 ;
        RECT 178.950 838.950 181.050 839.400 ;
        RECT 184.950 839.100 187.050 839.400 ;
        RECT 86.400 837.000 90.600 837.600 ;
        RECT 86.400 836.400 91.050 837.000 ;
        RECT 88.950 832.950 91.050 836.400 ;
        RECT 43.950 795.600 46.050 796.050 ;
        RECT 88.950 795.600 91.050 796.050 ;
        RECT 43.950 794.400 91.050 795.600 ;
        RECT 43.950 793.950 46.050 794.400 ;
        RECT 88.950 793.950 91.050 794.400 ;
        RECT 88.950 771.600 91.050 772.050 ;
        RECT 145.950 771.600 148.050 772.050 ;
        RECT 88.950 770.400 148.050 771.600 ;
        RECT 88.950 769.950 91.050 770.400 ;
        RECT 145.950 769.950 148.050 770.400 ;
        RECT 136.950 738.600 139.050 738.900 ;
        RECT 145.950 738.600 148.050 739.050 ;
        RECT 136.950 737.400 148.050 738.600 ;
        RECT 136.950 736.800 139.050 737.400 ;
        RECT 145.950 736.950 148.050 737.400 ;
        RECT 133.950 672.600 136.050 673.050 ;
        RECT 133.950 671.400 192.600 672.600 ;
        RECT 133.950 670.950 136.050 671.400 ;
        RECT 191.400 669.600 192.600 671.400 ;
        RECT 220.950 669.600 223.050 670.050 ;
        RECT 191.400 668.400 223.050 669.600 ;
        RECT 220.950 667.950 223.050 668.400 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal1 ;
        RECT 592.950 885.450 595.050 886.050 ;
        RECT 598.950 885.450 601.050 886.050 ;
        RECT 592.950 884.550 601.050 885.450 ;
        RECT 592.950 883.950 595.050 884.550 ;
        RECT 598.950 883.950 601.050 884.550 ;
        RECT 469.950 765.450 472.050 766.050 ;
        RECT 481.950 765.450 484.050 766.050 ;
        RECT 469.950 764.550 484.050 765.450 ;
        RECT 469.950 763.950 472.050 764.550 ;
        RECT 481.950 763.950 484.050 764.550 ;
        RECT 457.950 721.950 460.050 724.050 ;
        RECT 458.550 718.050 459.450 721.950 ;
        RECT 457.950 715.950 460.050 718.050 ;
      LAYER metal2 ;
        RECT 596.400 924.450 597.450 945.450 ;
        RECT 593.400 923.400 597.450 924.450 ;
        RECT 593.400 913.050 594.450 923.400 ;
        RECT 592.950 910.950 595.050 913.050 ;
        RECT 599.400 912.900 600.600 913.650 ;
        RECT 598.950 910.800 601.050 912.900 ;
        RECT 599.400 886.050 600.450 910.800 ;
        RECT 592.950 883.950 595.050 886.050 ;
        RECT 598.950 883.950 601.050 886.050 ;
        RECT 563.400 878.400 564.600 880.650 ;
        RECT 563.400 853.050 564.450 878.400 ;
        RECT 593.400 853.050 594.450 883.950 ;
        RECT 460.950 850.950 463.050 853.050 ;
        RECT 514.950 850.950 517.050 853.050 ;
        RECT 562.950 850.950 565.050 853.050 ;
        RECT 592.950 850.950 595.050 853.050 ;
        RECT 461.400 840.600 462.450 850.950 ;
        RECT 461.400 838.350 462.600 840.600 ;
        RECT 515.400 829.050 516.450 850.950 ;
        RECT 502.950 826.950 505.050 829.050 ;
        RECT 514.950 826.950 517.050 829.050 ;
        RECT 503.400 778.050 504.450 826.950 ;
        RECT 563.400 801.900 564.600 802.650 ;
        RECT 547.950 799.800 550.050 801.900 ;
        RECT 562.950 799.800 565.050 801.900 ;
        RECT 599.400 800.400 600.600 802.650 ;
        RECT 548.400 793.050 549.450 799.800 ;
        RECT 563.400 796.050 564.450 799.800 ;
        RECT 599.400 796.050 600.450 800.400 ;
        RECT 562.950 793.950 565.050 796.050 ;
        RECT 598.950 793.950 601.050 796.050 ;
        RECT 538.950 790.950 541.050 793.050 ;
        RECT 547.950 790.950 550.050 793.050 ;
        RECT 481.950 775.950 484.050 778.050 ;
        RECT 502.950 775.950 505.050 778.050 ;
        RECT 514.950 775.950 517.050 778.050 ;
        RECT 482.400 766.050 483.450 775.950 ;
        RECT 469.950 763.950 472.050 766.050 ;
        RECT 481.950 763.950 484.050 766.050 ;
        RECT 503.400 765.450 504.450 775.950 ;
        RECT 515.400 772.050 516.450 775.950 ;
        RECT 539.400 772.050 540.450 790.950 ;
        RECT 514.950 769.950 517.050 772.050 ;
        RECT 538.950 769.950 541.050 772.050 ;
        RECT 500.400 764.400 504.450 765.450 ;
        RECT 470.400 736.050 471.450 763.950 ;
        RECT 500.400 762.600 501.450 764.400 ;
        RECT 539.400 762.600 540.450 769.950 ;
        RECT 500.400 760.350 501.600 762.600 ;
        RECT 539.400 760.350 540.600 762.600 ;
        RECT 457.950 733.950 460.050 736.050 ;
        RECT 469.950 733.950 472.050 736.050 ;
        RECT 398.400 722.400 399.600 724.650 ;
        RECT 458.400 724.050 459.450 733.950 ;
        RECT 398.400 718.050 399.450 722.400 ;
        RECT 457.950 721.950 460.050 724.050 ;
        RECT 397.950 715.950 400.050 718.050 ;
        RECT 403.950 715.950 406.050 718.050 ;
        RECT 404.400 697.050 405.450 715.950 ;
        RECT 457.950 714.450 460.050 718.050 ;
        RECT 457.950 714.000 462.450 714.450 ;
        RECT 458.400 713.400 462.450 714.000 ;
        RECT 370.950 694.950 373.050 697.050 ;
        RECT 403.950 694.950 406.050 697.050 ;
        RECT 371.400 687.450 372.450 694.950 ;
        RECT 404.400 688.050 405.450 694.950 ;
        RECT 461.400 688.050 462.450 713.400 ;
        RECT 368.400 686.400 372.450 687.450 ;
        RECT 368.400 666.450 369.450 686.400 ;
        RECT 403.950 684.000 406.050 688.050 ;
        RECT 460.950 685.950 463.050 688.050 ;
        RECT 404.400 682.350 405.600 684.000 ;
        RECT 365.400 665.400 369.450 666.450 ;
        RECT 365.400 658.050 366.450 665.400 ;
        RECT 364.950 655.950 367.050 658.050 ;
        RECT 370.950 655.950 373.050 658.050 ;
        RECT 371.400 652.200 372.450 655.950 ;
        RECT 370.950 650.100 373.050 652.200 ;
        RECT 371.400 649.350 372.600 650.100 ;
        RECT 359.400 645.900 360.600 646.650 ;
        RECT 358.950 643.800 361.050 645.900 ;
      LAYER metal3 ;
        RECT 592.950 912.600 595.050 913.050 ;
        RECT 598.950 912.600 601.050 912.900 ;
        RECT 592.950 911.400 601.050 912.600 ;
        RECT 592.950 910.950 595.050 911.400 ;
        RECT 598.950 910.800 601.050 911.400 ;
        RECT 460.950 852.600 463.050 853.050 ;
        RECT 514.950 852.600 517.050 853.050 ;
        RECT 562.950 852.600 565.050 853.050 ;
        RECT 592.950 852.600 595.050 853.050 ;
        RECT 460.950 851.400 595.050 852.600 ;
        RECT 460.950 850.950 463.050 851.400 ;
        RECT 514.950 850.950 517.050 851.400 ;
        RECT 562.950 850.950 565.050 851.400 ;
        RECT 592.950 850.950 595.050 851.400 ;
        RECT 502.950 828.600 505.050 829.050 ;
        RECT 514.950 828.600 517.050 829.050 ;
        RECT 502.950 827.400 517.050 828.600 ;
        RECT 502.950 826.950 505.050 827.400 ;
        RECT 514.950 826.950 517.050 827.400 ;
        RECT 547.950 801.450 550.050 801.900 ;
        RECT 562.950 801.450 565.050 801.900 ;
        RECT 547.950 800.250 565.050 801.450 ;
        RECT 547.950 799.800 550.050 800.250 ;
        RECT 562.950 799.800 565.050 800.250 ;
        RECT 562.950 795.600 565.050 796.050 ;
        RECT 598.950 795.600 601.050 796.050 ;
        RECT 562.950 794.400 601.050 795.600 ;
        RECT 562.950 793.950 565.050 794.400 ;
        RECT 598.950 793.950 601.050 794.400 ;
        RECT 538.950 792.600 541.050 793.050 ;
        RECT 547.950 792.600 550.050 793.050 ;
        RECT 538.950 791.400 550.050 792.600 ;
        RECT 538.950 790.950 541.050 791.400 ;
        RECT 547.950 790.950 550.050 791.400 ;
        RECT 481.950 777.600 484.050 778.050 ;
        RECT 502.950 777.600 505.050 778.050 ;
        RECT 514.950 777.600 517.050 778.050 ;
        RECT 481.950 776.400 517.050 777.600 ;
        RECT 481.950 775.950 484.050 776.400 ;
        RECT 502.950 775.950 505.050 776.400 ;
        RECT 514.950 775.950 517.050 776.400 ;
        RECT 514.950 771.600 517.050 772.050 ;
        RECT 538.950 771.600 541.050 772.050 ;
        RECT 514.950 770.400 541.050 771.600 ;
        RECT 514.950 769.950 517.050 770.400 ;
        RECT 538.950 769.950 541.050 770.400 ;
        RECT 457.950 735.600 460.050 736.050 ;
        RECT 469.950 735.600 472.050 736.050 ;
        RECT 457.950 734.400 472.050 735.600 ;
        RECT 457.950 733.950 460.050 734.400 ;
        RECT 469.950 733.950 472.050 734.400 ;
        RECT 397.950 717.600 400.050 718.050 ;
        RECT 403.950 717.600 406.050 718.050 ;
        RECT 397.950 716.400 406.050 717.600 ;
        RECT 397.950 715.950 400.050 716.400 ;
        RECT 403.950 715.950 406.050 716.400 ;
        RECT 370.950 696.600 373.050 697.050 ;
        RECT 403.950 696.600 406.050 697.050 ;
        RECT 370.950 695.400 406.050 696.600 ;
        RECT 370.950 694.950 373.050 695.400 ;
        RECT 403.950 694.950 406.050 695.400 ;
        RECT 403.950 687.600 406.050 688.050 ;
        RECT 460.950 687.600 463.050 688.050 ;
        RECT 403.950 686.400 463.050 687.600 ;
        RECT 403.950 685.950 406.050 686.400 ;
        RECT 460.950 685.950 463.050 686.400 ;
        RECT 364.950 657.600 367.050 658.050 ;
        RECT 370.950 657.600 373.050 658.050 ;
        RECT 364.950 656.400 373.050 657.600 ;
        RECT 364.950 655.950 367.050 656.400 ;
        RECT 370.950 655.950 373.050 656.400 ;
        RECT 370.950 651.600 373.050 652.200 ;
        RECT 359.400 650.400 373.050 651.600 ;
        RECT 359.400 645.900 360.600 650.400 ;
        RECT 370.950 650.100 373.050 650.400 ;
        RECT 358.950 643.800 361.050 645.900 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal1 ;
        RECT 565.950 807.450 570.000 808.050 ;
        RECT 565.950 805.950 570.450 807.450 ;
        RECT 569.550 802.050 570.450 805.950 ;
        RECT 565.950 800.550 570.450 802.050 ;
        RECT 565.950 799.950 570.000 800.550 ;
        RECT 558.000 729.450 562.050 730.050 ;
        RECT 557.550 727.950 562.050 729.450 ;
        RECT 557.550 724.050 558.450 727.950 ;
        RECT 553.950 722.550 558.450 724.050 ;
        RECT 553.950 721.950 558.000 722.550 ;
      LAYER metal2 ;
        RECT 614.400 944.400 618.450 945.450 ;
        RECT 617.400 925.050 618.450 944.400 ;
        RECT 550.950 922.950 553.050 925.050 ;
        RECT 616.950 922.950 619.050 925.050 ;
        RECT 551.400 847.050 552.450 922.950 ;
        RECT 617.400 918.600 618.450 922.950 ;
        RECT 617.400 916.350 618.600 918.600 ;
        RECT 550.950 844.950 553.050 847.050 ;
        RECT 565.950 844.800 568.050 846.900 ;
        RECT 566.400 808.050 567.450 844.800 ;
        RECT 565.950 805.950 568.050 808.050 ;
        RECT 557.400 800.400 558.600 802.650 ;
        RECT 557.400 793.050 558.450 800.400 ;
        RECT 565.950 799.950 568.050 802.050 ;
        RECT 566.400 793.050 567.450 799.950 ;
        RECT 556.950 790.950 559.050 793.050 ;
        RECT 565.950 790.950 568.050 793.050 ;
        RECT 557.400 787.050 558.450 790.950 ;
        RECT 547.950 784.950 550.050 787.050 ;
        RECT 556.950 784.950 559.050 787.050 ;
        RECT 548.400 763.050 549.450 784.950 ;
        RECT 547.800 760.950 549.900 763.050 ;
        RECT 556.950 754.950 559.050 757.050 ;
        RECT 557.400 735.450 558.450 754.950 ;
        RECT 557.400 734.400 561.450 735.450 ;
        RECT 560.400 730.050 561.450 734.400 ;
        RECT 559.950 727.950 562.050 730.050 ;
        RECT 553.950 721.950 556.050 724.050 ;
        RECT 554.400 661.050 555.450 721.950 ;
        RECT 448.950 658.950 451.050 661.050 ;
        RECT 553.950 658.950 556.050 661.050 ;
        RECT 449.400 651.600 450.450 658.950 ;
        RECT 449.400 649.350 450.600 651.600 ;
      LAYER metal3 ;
        RECT 550.950 924.600 553.050 925.050 ;
        RECT 616.950 924.600 619.050 925.050 ;
        RECT 550.950 923.400 619.050 924.600 ;
        RECT 550.950 922.950 553.050 923.400 ;
        RECT 616.950 922.950 619.050 923.400 ;
        RECT 550.950 846.600 553.050 847.050 ;
        RECT 565.950 846.600 568.050 846.900 ;
        RECT 550.950 845.400 568.050 846.600 ;
        RECT 550.950 844.950 553.050 845.400 ;
        RECT 565.950 844.800 568.050 845.400 ;
        RECT 556.950 792.600 559.050 793.050 ;
        RECT 565.950 792.600 568.050 793.050 ;
        RECT 556.950 791.400 568.050 792.600 ;
        RECT 556.950 790.950 559.050 791.400 ;
        RECT 565.950 790.950 568.050 791.400 ;
        RECT 547.950 786.600 550.050 787.050 ;
        RECT 556.950 786.600 559.050 787.050 ;
        RECT 547.950 785.400 559.050 786.600 ;
        RECT 547.950 784.950 550.050 785.400 ;
        RECT 556.950 784.950 559.050 785.400 ;
        RECT 547.800 762.000 549.900 763.050 ;
        RECT 547.800 760.950 550.050 762.000 ;
        RECT 547.950 759.600 550.050 760.950 ;
        RECT 547.950 759.000 558.600 759.600 ;
        RECT 548.400 758.400 559.050 759.000 ;
        RECT 556.950 754.950 559.050 758.400 ;
        RECT 448.950 660.600 451.050 661.050 ;
        RECT 553.950 660.600 556.050 661.050 ;
        RECT 448.950 659.400 556.050 660.600 ;
        RECT 448.950 658.950 451.050 659.400 ;
        RECT 553.950 658.950 556.050 659.400 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal2 ;
        RECT 659.400 944.400 663.450 945.450 ;
        RECT 662.400 918.600 663.450 944.400 ;
        RECT 662.400 918.450 663.600 918.600 ;
        RECT 662.400 917.400 666.450 918.450 ;
        RECT 662.400 916.350 663.600 917.400 ;
        RECT 665.400 889.050 666.450 917.400 ;
        RECT 658.950 886.950 661.050 889.050 ;
        RECT 664.800 886.950 666.900 889.050 ;
        RECT 659.400 847.050 660.450 886.950 ;
        RECT 658.950 844.950 661.050 847.050 ;
        RECT 667.950 844.950 670.050 847.050 ;
        RECT 668.400 811.050 669.450 844.950 ;
        RECT 661.950 807.000 664.050 811.050 ;
        RECT 667.950 808.950 670.050 811.050 ;
        RECT 662.400 805.350 663.600 807.000 ;
      LAYER metal3 ;
        RECT 658.950 888.600 661.050 889.050 ;
        RECT 664.800 888.600 666.900 889.050 ;
        RECT 658.950 887.400 666.900 888.600 ;
        RECT 658.950 886.950 661.050 887.400 ;
        RECT 664.800 886.950 666.900 887.400 ;
        RECT 658.950 846.600 661.050 847.050 ;
        RECT 667.950 846.600 670.050 847.050 ;
        RECT 658.950 845.400 670.050 846.600 ;
        RECT 658.950 844.950 661.050 845.400 ;
        RECT 667.950 844.950 670.050 845.400 ;
        RECT 661.950 810.600 664.050 811.050 ;
        RECT 667.950 810.600 670.050 811.050 ;
        RECT 661.950 809.400 670.050 810.600 ;
        RECT 661.950 808.950 664.050 809.400 ;
        RECT 667.950 808.950 670.050 809.400 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal1 ;
        RECT 505.950 903.450 508.050 904.050 ;
        RECT 511.950 903.450 514.050 904.050 ;
        RECT 505.950 902.550 514.050 903.450 ;
        RECT 505.950 901.950 508.050 902.550 ;
        RECT 511.950 901.950 514.050 902.550 ;
      LAYER metal2 ;
        RECT 934.950 931.950 937.050 934.050 ;
        RECT 532.950 928.950 535.050 931.050 ;
        RECT 691.950 928.950 694.050 931.050 ;
        RECT 265.950 907.950 268.050 910.050 ;
        RECT 304.950 907.950 307.050 910.050 ;
        RECT 266.400 886.200 267.450 907.950 ;
        RECT 305.400 895.050 306.450 907.950 ;
        RECT 504.000 903.450 508.050 904.050 ;
        RECT 503.400 901.950 508.050 903.450 ;
        RECT 304.950 892.950 307.050 895.050 ;
        RECT 403.950 892.950 406.050 895.050 ;
        RECT 404.400 886.200 405.450 892.950 ;
        RECT 253.950 884.100 256.050 886.200 ;
        RECT 265.950 884.100 268.050 886.200 ;
        RECT 403.950 884.100 406.050 886.200 ;
        RECT 254.400 883.350 255.600 884.100 ;
        RECT 266.400 883.350 267.600 884.100 ;
        RECT 404.400 883.350 405.600 884.100 ;
        RECT 503.400 883.050 504.450 901.950 ;
        RECT 511.950 898.950 514.050 904.050 ;
        RECT 533.400 901.050 534.450 928.950 ;
        RECT 532.950 898.950 535.050 901.050 ;
        RECT 689.400 885.450 690.600 885.600 ;
        RECT 692.400 885.450 693.450 928.950 ;
        RECT 689.400 884.400 693.450 885.450 ;
        RECT 689.400 883.350 690.600 884.400 ;
        RECT 502.950 880.950 505.050 883.050 ;
        RECT 935.400 880.050 936.450 931.950 ;
        RECT 934.950 877.950 937.050 880.050 ;
      LAYER metal3 ;
        RECT 934.950 933.600 937.050 934.050 ;
        RECT 692.400 932.400 937.050 933.600 ;
        RECT 692.400 931.050 693.600 932.400 ;
        RECT 934.950 931.950 937.050 932.400 ;
        RECT 532.950 930.600 535.050 931.050 ;
        RECT 691.950 930.600 694.050 931.050 ;
        RECT 532.950 929.400 694.050 930.600 ;
        RECT 532.950 928.950 535.050 929.400 ;
        RECT 691.950 928.950 694.050 929.400 ;
        RECT 265.950 909.600 268.050 910.050 ;
        RECT 304.950 909.600 307.050 910.050 ;
        RECT 265.950 908.400 307.050 909.600 ;
        RECT 265.950 907.950 268.050 908.400 ;
        RECT 304.950 907.950 307.050 908.400 ;
        RECT 511.950 900.600 514.050 901.050 ;
        RECT 532.950 900.600 535.050 901.050 ;
        RECT 511.950 899.400 535.050 900.600 ;
        RECT 511.950 898.950 514.050 899.400 ;
        RECT 532.950 898.950 535.050 899.400 ;
        RECT 304.950 894.600 307.050 895.050 ;
        RECT 403.950 894.600 406.050 895.050 ;
        RECT 304.950 893.400 406.050 894.600 ;
        RECT 304.950 892.950 307.050 893.400 ;
        RECT 403.950 892.950 406.050 893.400 ;
        RECT 253.950 885.600 256.050 886.200 ;
        RECT 265.950 885.600 268.050 886.200 ;
        RECT 253.950 884.400 268.050 885.600 ;
        RECT 253.950 884.100 256.050 884.400 ;
        RECT 265.950 884.100 268.050 884.400 ;
        RECT 403.950 885.600 406.050 886.200 ;
        RECT 403.950 884.400 420.600 885.600 ;
        RECT 403.950 884.100 406.050 884.400 ;
        RECT 419.400 882.600 420.600 884.400 ;
        RECT 502.950 882.600 505.050 883.050 ;
        RECT 419.400 881.400 505.050 882.600 ;
        RECT 502.950 880.950 505.050 881.400 ;
        RECT 934.950 879.600 937.050 880.050 ;
        RECT 934.950 878.400 942.600 879.600 ;
        RECT 934.950 877.950 937.050 878.400 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal2 ;
        RECT 934.950 844.950 937.050 847.050 ;
        RECT 665.400 833.400 666.600 835.650 ;
        RECT 665.400 826.050 666.450 833.400 ;
        RECT 655.950 823.950 658.050 826.050 ;
        RECT 664.950 823.950 667.050 826.050 ;
        RECT 656.400 793.050 657.450 823.950 ;
        RECT 935.400 817.050 936.450 844.950 ;
        RECT 934.950 814.950 937.050 817.050 ;
        RECT 853.950 811.950 856.050 814.050 ;
        RECT 683.400 800.400 684.600 802.650 ;
        RECT 683.400 793.050 684.450 800.400 ;
        RECT 854.400 799.050 855.450 811.950 ;
        RECT 814.950 796.950 817.050 799.050 ;
        RECT 853.800 796.950 855.900 799.050 ;
        RECT 637.950 790.950 640.050 793.050 ;
        RECT 655.950 790.950 658.050 793.050 ;
        RECT 682.950 790.950 685.050 793.050 ;
        RECT 638.400 775.050 639.450 790.950 ;
        RECT 760.950 787.950 763.050 790.050 ;
        RECT 761.400 784.050 762.450 787.950 ;
        RECT 815.400 784.050 816.450 796.950 ;
        RECT 760.950 781.950 763.050 784.050 ;
        RECT 814.950 781.950 817.050 784.050 ;
        RECT 592.950 772.950 595.050 775.050 ;
        RECT 637.950 772.950 640.050 775.050 ;
        RECT 593.400 754.050 594.450 772.950 ;
        RECT 571.950 751.800 574.050 753.900 ;
        RECT 592.950 751.950 595.050 754.050 ;
        RECT 572.400 730.200 573.450 751.800 ;
        RECT 565.950 728.100 568.050 730.200 ;
        RECT 571.950 728.100 574.050 730.200 ;
        RECT 566.400 727.350 567.600 728.100 ;
        RECT 551.400 723.900 552.600 724.650 ;
        RECT 572.400 724.050 573.450 728.100 ;
        RECT 550.950 721.800 553.050 723.900 ;
        RECT 571.950 721.950 574.050 724.050 ;
      LAYER metal3 ;
        RECT 934.950 846.600 937.050 847.050 ;
        RECT 934.950 845.400 942.600 846.600 ;
        RECT 934.950 844.950 937.050 845.400 ;
        RECT 655.950 825.600 658.050 826.050 ;
        RECT 664.950 825.600 667.050 826.050 ;
        RECT 655.950 824.400 667.050 825.600 ;
        RECT 655.950 823.950 658.050 824.400 ;
        RECT 664.950 823.950 667.050 824.400 ;
        RECT 934.950 816.600 937.050 817.050 ;
        RECT 908.400 815.400 937.050 816.600 ;
        RECT 853.950 813.600 856.050 814.050 ;
        RECT 908.400 813.600 909.600 815.400 ;
        RECT 934.950 814.950 937.050 815.400 ;
        RECT 853.950 812.400 909.600 813.600 ;
        RECT 853.950 811.950 856.050 812.400 ;
        RECT 814.950 798.600 817.050 799.050 ;
        RECT 853.800 798.600 855.900 799.050 ;
        RECT 814.950 797.400 855.900 798.600 ;
        RECT 814.950 796.950 817.050 797.400 ;
        RECT 853.800 796.950 855.900 797.400 ;
        RECT 637.950 792.600 640.050 793.050 ;
        RECT 655.950 792.600 658.050 793.050 ;
        RECT 682.950 792.600 685.050 793.050 ;
        RECT 637.950 791.400 685.050 792.600 ;
        RECT 637.950 790.950 640.050 791.400 ;
        RECT 655.950 790.950 658.050 791.400 ;
        RECT 682.950 790.950 685.050 791.400 ;
        RECT 683.400 789.600 684.600 790.950 ;
        RECT 760.950 789.600 763.050 790.050 ;
        RECT 683.400 788.400 763.050 789.600 ;
        RECT 760.950 787.950 763.050 788.400 ;
        RECT 760.950 783.600 763.050 784.050 ;
        RECT 814.950 783.600 817.050 784.050 ;
        RECT 760.950 782.400 817.050 783.600 ;
        RECT 760.950 781.950 763.050 782.400 ;
        RECT 814.950 781.950 817.050 782.400 ;
        RECT 592.950 774.600 595.050 775.050 ;
        RECT 637.950 774.600 640.050 775.050 ;
        RECT 592.950 773.400 640.050 774.600 ;
        RECT 592.950 772.950 595.050 773.400 ;
        RECT 637.950 772.950 640.050 773.400 ;
        RECT 571.950 753.600 574.050 753.900 ;
        RECT 592.950 753.600 595.050 754.050 ;
        RECT 571.950 752.400 595.050 753.600 ;
        RECT 571.950 751.800 574.050 752.400 ;
        RECT 592.950 751.950 595.050 752.400 ;
        RECT 565.950 729.750 568.050 730.200 ;
        RECT 571.950 729.750 574.050 730.200 ;
        RECT 565.950 728.550 574.050 729.750 ;
        RECT 565.950 728.100 568.050 728.550 ;
        RECT 571.950 728.100 574.050 728.550 ;
        RECT 550.950 723.600 553.050 723.900 ;
        RECT 571.950 723.600 574.050 724.050 ;
        RECT 550.950 722.400 574.050 723.600 ;
        RECT 550.950 721.800 553.050 722.400 ;
        RECT 571.950 721.950 574.050 722.400 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal2 ;
        RECT 652.950 868.950 655.050 871.050 ;
        RECT 820.950 868.950 823.050 871.050 ;
        RECT 653.400 840.600 654.450 868.950 ;
        RECT 821.400 853.050 822.450 868.950 ;
        RECT 821.400 851.400 826.050 853.050 ;
        RECT 822.000 850.950 826.050 851.400 ;
        RECT 880.950 850.950 883.050 853.050 ;
        RECT 881.400 841.050 882.450 850.950 ;
        RECT 653.400 840.450 654.600 840.600 ;
        RECT 650.400 839.400 654.600 840.450 ;
        RECT 521.400 833.400 522.600 835.650 ;
        RECT 605.400 833.400 606.600 835.650 ;
        RECT 521.400 829.050 522.450 833.400 ;
        RECT 605.400 831.450 606.450 833.400 ;
        RECT 650.400 832.050 651.450 839.400 ;
        RECT 653.400 838.350 654.600 839.400 ;
        RECT 880.950 838.950 883.050 841.050 ;
        RECT 602.400 830.400 606.450 831.450 ;
        RECT 520.950 826.950 523.050 829.050 ;
        RECT 553.950 826.950 556.050 829.050 ;
        RECT 554.400 820.050 555.450 826.950 ;
        RECT 602.400 820.050 603.450 830.400 ;
        RECT 622.950 829.950 625.050 832.050 ;
        RECT 649.950 829.950 652.050 832.050 ;
        RECT 623.400 820.050 624.450 829.950 ;
        RECT 553.950 817.950 556.050 820.050 ;
        RECT 601.950 817.950 604.050 820.050 ;
        RECT 607.950 817.950 610.050 820.050 ;
        RECT 622.950 817.950 625.050 820.050 ;
        RECT 608.400 762.450 609.450 817.950 ;
        RECT 610.950 762.450 613.050 763.200 ;
        RECT 608.400 761.400 613.050 762.450 ;
        RECT 610.950 761.100 613.050 761.400 ;
        RECT 619.950 761.100 622.050 763.200 ;
        RECT 581.400 755.400 582.600 757.650 ;
        RECT 581.400 744.450 582.450 755.400 ;
        RECT 578.400 743.400 582.450 744.450 ;
        RECT 578.400 736.050 579.450 743.400 ;
        RECT 611.400 736.050 612.450 761.100 ;
        RECT 620.400 760.350 621.600 761.100 ;
        RECT 577.950 733.950 580.050 736.050 ;
        RECT 610.800 733.950 612.900 736.050 ;
        RECT 491.400 722.400 492.600 724.650 ;
        RECT 491.400 709.050 492.450 722.400 ;
        RECT 578.400 709.050 579.450 733.950 ;
        RECT 490.950 706.950 493.050 709.050 ;
        RECT 577.950 706.950 580.050 709.050 ;
        RECT 482.400 678.000 483.600 679.650 ;
        RECT 481.950 673.950 484.050 678.000 ;
        RECT 491.400 676.050 492.450 706.950 ;
        RECT 490.950 673.950 493.050 676.050 ;
      LAYER metal3 ;
        RECT 652.950 870.600 655.050 871.050 ;
        RECT 820.950 870.600 823.050 871.050 ;
        RECT 652.950 869.400 823.050 870.600 ;
        RECT 652.950 868.950 655.050 869.400 ;
        RECT 820.950 868.950 823.050 869.400 ;
        RECT 823.950 852.600 826.050 853.050 ;
        RECT 880.950 852.600 883.050 853.050 ;
        RECT 823.950 851.400 883.050 852.600 ;
        RECT 823.950 850.950 826.050 851.400 ;
        RECT 880.950 850.950 883.050 851.400 ;
        RECT 880.950 840.600 883.050 841.050 ;
        RECT 880.950 839.400 942.600 840.600 ;
        RECT 880.950 838.950 883.050 839.400 ;
        RECT 622.950 831.600 625.050 832.050 ;
        RECT 649.950 831.600 652.050 832.050 ;
        RECT 622.950 830.400 652.050 831.600 ;
        RECT 622.950 829.950 625.050 830.400 ;
        RECT 649.950 829.950 652.050 830.400 ;
        RECT 520.950 828.600 523.050 829.050 ;
        RECT 553.950 828.600 556.050 829.050 ;
        RECT 520.950 827.400 556.050 828.600 ;
        RECT 520.950 826.950 523.050 827.400 ;
        RECT 553.950 826.950 556.050 827.400 ;
        RECT 553.950 819.600 556.050 820.050 ;
        RECT 601.950 819.600 604.050 820.050 ;
        RECT 607.950 819.600 610.050 820.050 ;
        RECT 622.950 819.600 625.050 820.050 ;
        RECT 553.950 818.400 625.050 819.600 ;
        RECT 553.950 817.950 556.050 818.400 ;
        RECT 601.950 817.950 604.050 818.400 ;
        RECT 607.950 817.950 610.050 818.400 ;
        RECT 622.950 817.950 625.050 818.400 ;
        RECT 610.950 762.750 613.050 763.200 ;
        RECT 619.950 762.750 622.050 763.200 ;
        RECT 610.950 761.550 622.050 762.750 ;
        RECT 610.950 761.100 613.050 761.550 ;
        RECT 619.950 761.100 622.050 761.550 ;
        RECT 577.950 735.600 580.050 736.050 ;
        RECT 610.800 735.600 612.900 736.050 ;
        RECT 577.950 734.400 612.900 735.600 ;
        RECT 577.950 733.950 580.050 734.400 ;
        RECT 610.800 733.950 612.900 734.400 ;
        RECT 490.950 708.600 493.050 709.050 ;
        RECT 577.950 708.600 580.050 709.050 ;
        RECT 490.950 707.400 580.050 708.600 ;
        RECT 490.950 706.950 493.050 707.400 ;
        RECT 577.950 706.950 580.050 707.400 ;
        RECT 481.950 675.600 484.050 676.050 ;
        RECT 490.950 675.600 493.050 676.050 ;
        RECT 481.950 674.400 493.050 675.600 ;
        RECT 481.950 673.950 484.050 674.400 ;
        RECT 490.950 673.950 493.050 674.400 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal2 ;
        RECT 17.400 98.400 18.600 100.650 ;
        RECT 17.400 67.050 18.450 98.400 ;
        RECT 7.950 64.950 10.050 67.050 ;
        RECT 16.950 64.950 19.050 67.050 ;
        RECT 8.400 -2.550 9.450 64.950 ;
        RECT 8.400 -3.600 12.450 -2.550 ;
      LAYER metal3 ;
        RECT 7.950 66.600 10.050 67.050 ;
        RECT 16.950 66.600 19.050 67.050 ;
        RECT 7.950 65.400 19.050 66.600 ;
        RECT 7.950 64.950 10.050 65.400 ;
        RECT 16.950 64.950 19.050 65.400 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal2 ;
        RECT 20.400 20.400 21.600 22.650 ;
        RECT 20.400 -2.550 21.450 20.400 ;
        RECT 17.400 -3.600 21.450 -2.550 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal2 ;
        RECT 32.400 20.400 33.600 22.650 ;
        RECT 32.400 -2.550 33.450 20.400 ;
        RECT 32.400 -3.600 36.450 -2.550 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal2 ;
        RECT 50.400 20.400 51.600 22.650 ;
        RECT 50.400 -2.550 51.450 20.400 ;
        RECT 50.400 -3.600 54.450 -2.550 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal2 ;
        RECT 95.400 20.400 96.600 22.650 ;
        RECT 95.400 -2.550 96.450 20.400 ;
        RECT 92.400 -3.600 96.450 -2.550 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal2 ;
        RECT 11.400 567.900 12.600 568.650 ;
        RECT 10.950 565.800 13.050 567.900 ;
      LAYER metal3 ;
        RECT 10.950 567.600 13.050 567.900 ;
        RECT -3.600 566.400 13.050 567.600 ;
        RECT 10.950 565.800 13.050 566.400 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal2 ;
        RECT 32.400 411.000 33.600 412.650 ;
        RECT 31.950 406.950 34.050 411.000 ;
      LAYER metal3 ;
        RECT -3.600 414.600 -2.400 417.600 ;
        RECT -6.600 413.400 -2.400 414.600 ;
        RECT -6.600 408.600 -5.400 413.400 ;
        RECT 31.950 408.600 34.050 409.050 ;
        RECT -6.600 407.400 34.050 408.600 ;
        RECT 31.950 406.950 34.050 407.400 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal2 ;
        RECT 11.400 411.900 12.600 412.650 ;
        RECT 10.950 409.800 13.050 411.900 ;
      LAYER metal3 ;
        RECT 10.950 411.600 13.050 411.900 ;
        RECT -3.600 410.400 13.050 411.600 ;
        RECT 10.950 409.800 13.050 410.400 ;
    END
  END ACC_o[0]
  PIN Done_o
    PORT
      LAYER metal1 ;
        RECT 180.000 105.450 184.050 106.050 ;
        RECT 179.550 103.950 184.050 105.450 ;
        RECT 179.550 100.050 180.450 103.950 ;
        RECT 175.950 98.550 180.450 100.050 ;
        RECT 175.950 97.950 180.000 98.550 ;
      LAYER metal2 ;
        RECT 176.400 216.450 177.600 216.600 ;
        RECT 176.400 215.400 180.450 216.450 ;
        RECT 176.400 214.350 177.600 215.400 ;
        RECT 179.400 187.050 180.450 215.400 ;
        RECT 172.950 184.950 175.050 187.050 ;
        RECT 178.950 184.950 181.050 187.050 ;
        RECT 173.400 145.050 174.450 184.950 ;
        RECT 172.950 142.950 175.050 145.050 ;
        RECT 184.950 142.950 187.050 145.050 ;
        RECT 185.400 114.450 186.450 142.950 ;
        RECT 182.400 113.400 186.450 114.450 ;
        RECT 182.400 106.050 183.450 113.400 ;
        RECT 181.950 103.950 184.050 106.050 ;
        RECT 175.950 97.950 178.050 100.050 ;
        RECT 176.400 67.050 177.450 97.950 ;
        RECT 169.950 64.950 172.050 67.050 ;
        RECT 175.950 64.950 178.050 67.050 ;
        RECT 170.400 27.450 171.450 64.950 ;
        RECT 167.400 26.400 171.450 27.450 ;
        RECT 167.400 4.050 168.450 26.400 ;
        RECT 166.950 1.950 169.050 4.050 ;
        RECT 172.950 1.950 175.050 4.050 ;
        RECT 173.400 -3.600 174.450 1.950 ;
      LAYER metal3 ;
        RECT 172.950 186.600 175.050 187.050 ;
        RECT 178.950 186.600 181.050 187.050 ;
        RECT 172.950 185.400 181.050 186.600 ;
        RECT 172.950 184.950 175.050 185.400 ;
        RECT 178.950 184.950 181.050 185.400 ;
        RECT 172.950 144.600 175.050 145.050 ;
        RECT 184.950 144.600 187.050 145.050 ;
        RECT 172.950 143.400 187.050 144.600 ;
        RECT 172.950 142.950 175.050 143.400 ;
        RECT 184.950 142.950 187.050 143.400 ;
        RECT 169.950 66.600 172.050 67.050 ;
        RECT 175.950 66.600 178.050 67.050 ;
        RECT 169.950 65.400 178.050 66.600 ;
        RECT 169.950 64.950 172.050 65.400 ;
        RECT 175.950 64.950 178.050 65.400 ;
        RECT 166.950 3.600 169.050 4.050 ;
        RECT 172.950 3.600 175.050 4.050 ;
        RECT 166.950 2.400 175.050 3.600 ;
        RECT 166.950 1.950 169.050 2.400 ;
        RECT 172.950 1.950 175.050 2.400 ;
    END
  END Done_o
  PIN LoadA_i
    PORT
      LAYER metal1 ;
        RECT 64.950 886.950 67.050 889.050 ;
        RECT 65.550 880.050 66.450 886.950 ;
        RECT 61.950 878.550 66.450 880.050 ;
        RECT 61.950 877.950 66.000 878.550 ;
      LAYER metal2 ;
        RECT 65.400 944.400 69.450 945.450 ;
        RECT 65.400 919.050 66.450 944.400 ;
        RECT 64.800 916.950 66.900 919.050 ;
        RECT 64.800 910.950 66.900 913.050 ;
        RECT 65.400 889.050 66.450 910.950 ;
        RECT 64.950 886.950 67.050 889.050 ;
        RECT 61.950 877.950 64.050 880.050 ;
        RECT 62.400 868.050 63.450 877.950 ;
        RECT 49.950 865.950 52.050 868.050 ;
        RECT 61.950 865.950 64.050 868.050 ;
        RECT 50.400 834.450 51.450 865.950 ;
        RECT 50.400 833.400 54.450 834.450 ;
        RECT 53.400 808.050 54.450 833.400 ;
        RECT 52.950 805.950 55.050 808.050 ;
        RECT 52.950 799.950 55.050 802.050 ;
        RECT 53.400 775.050 54.450 799.950 ;
        RECT 52.950 772.950 55.050 775.050 ;
        RECT 76.800 772.950 78.900 775.050 ;
        RECT 77.400 763.050 78.450 772.950 ;
        RECT 76.950 760.950 79.050 763.050 ;
        RECT 40.950 751.950 43.050 754.050 ;
        RECT 41.400 721.050 42.450 751.950 ;
        RECT 31.950 718.950 34.050 721.050 ;
        RECT 40.950 718.950 43.050 721.050 ;
        RECT 32.400 678.450 33.450 718.950 ;
        RECT 38.400 678.450 39.600 679.650 ;
        RECT 32.400 677.400 39.600 678.450 ;
        RECT 35.400 655.050 36.450 677.400 ;
        RECT 91.950 655.950 94.050 658.050 ;
        RECT 34.950 652.950 37.050 655.050 ;
        RECT 35.400 651.600 36.450 652.950 ;
        RECT 92.400 651.600 93.450 655.950 ;
        RECT 35.400 649.350 36.600 651.600 ;
        RECT 92.400 649.350 93.600 651.600 ;
      LAYER metal3 ;
        RECT 64.800 916.950 66.900 919.050 ;
        RECT 65.250 913.050 66.450 916.950 ;
        RECT 64.800 910.950 66.900 913.050 ;
        RECT 49.950 867.600 52.050 868.050 ;
        RECT 61.950 867.600 64.050 868.050 ;
        RECT 49.950 866.400 64.050 867.600 ;
        RECT 49.950 865.950 52.050 866.400 ;
        RECT 61.950 865.950 64.050 866.400 ;
        RECT 52.950 805.950 55.050 808.050 ;
        RECT 53.400 802.050 54.600 805.950 ;
        RECT 52.950 799.950 55.050 802.050 ;
        RECT 52.950 774.600 55.050 775.050 ;
        RECT 76.800 774.600 78.900 775.050 ;
        RECT 52.950 773.400 78.900 774.600 ;
        RECT 52.950 772.950 55.050 773.400 ;
        RECT 76.800 772.950 78.900 773.400 ;
        RECT 76.950 762.600 79.050 763.050 ;
        RECT 65.400 761.400 79.050 762.600 ;
        RECT 40.950 753.600 43.050 754.050 ;
        RECT 65.400 753.600 66.600 761.400 ;
        RECT 76.950 760.950 79.050 761.400 ;
        RECT 40.950 752.400 66.600 753.600 ;
        RECT 40.950 751.950 43.050 752.400 ;
        RECT 31.950 720.600 34.050 721.050 ;
        RECT 40.950 720.600 43.050 721.050 ;
        RECT 31.950 719.400 43.050 720.600 ;
        RECT 31.950 718.950 34.050 719.400 ;
        RECT 40.950 718.950 43.050 719.400 ;
        RECT 91.950 657.600 94.050 658.050 ;
        RECT 71.400 656.400 94.050 657.600 ;
        RECT 34.950 654.600 37.050 655.050 ;
        RECT 71.400 654.600 72.600 656.400 ;
        RECT 91.950 655.950 94.050 656.400 ;
        RECT 34.950 653.400 72.600 654.600 ;
        RECT 34.950 652.950 37.050 653.400 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal1 ;
        RECT 85.950 885.450 90.000 886.050 ;
        RECT 85.950 883.950 90.450 885.450 ;
        RECT 89.550 880.050 90.450 883.950 ;
        RECT 85.950 878.550 90.450 880.050 ;
        RECT 85.950 877.950 90.000 878.550 ;
      LAYER metal2 ;
        RECT 74.400 944.400 78.450 945.450 ;
        RECT 77.400 919.050 78.450 944.400 ;
        RECT 76.950 916.950 79.050 919.050 ;
        RECT 82.950 909.450 85.050 913.050 ;
        RECT 82.950 909.000 87.450 909.450 ;
        RECT 83.400 908.400 87.450 909.000 ;
        RECT 86.400 886.050 87.450 908.400 ;
        RECT 85.950 883.950 88.050 886.050 ;
        RECT 85.950 877.950 88.050 880.050 ;
        RECT 86.400 873.450 87.450 877.950 ;
        RECT 86.400 872.400 90.450 873.450 ;
        RECT 89.400 844.050 90.450 872.400 ;
        RECT 88.950 841.950 91.050 844.050 ;
        RECT 85.950 829.950 88.050 832.050 ;
        RECT 86.400 808.050 87.450 829.950 ;
        RECT 85.950 805.950 88.050 808.050 ;
        RECT 82.950 796.950 85.050 799.050 ;
        RECT 83.400 766.050 84.450 796.950 ;
        RECT 82.950 763.950 85.050 766.050 ;
        RECT 91.950 751.950 94.050 754.050 ;
        RECT 92.400 729.450 93.450 751.950 ;
        RECT 92.400 728.400 96.450 729.450 ;
        RECT 95.400 706.050 96.450 728.400 ;
        RECT 40.950 703.950 43.050 706.050 ;
        RECT 94.950 703.950 97.050 706.050 ;
        RECT 41.400 685.200 42.450 703.950 ;
        RECT 40.950 683.100 43.050 685.200 ;
        RECT 41.400 682.350 42.600 683.100 ;
        RECT 40.950 673.950 43.050 676.050 ;
        RECT 41.400 657.450 42.450 673.950 ;
        RECT 41.400 656.400 45.450 657.450 ;
        RECT 44.400 613.050 45.450 656.400 ;
        RECT 43.950 610.950 46.050 613.050 ;
        RECT 79.950 610.950 82.050 613.050 ;
        RECT 100.950 610.950 103.050 613.050 ;
        RECT 80.400 606.600 81.450 610.950 ;
        RECT 101.400 607.050 102.450 610.950 ;
        RECT 80.400 604.350 81.600 606.600 ;
        RECT 100.950 604.950 103.050 607.050 ;
        RECT 104.400 601.050 105.600 601.650 ;
        RECT 100.950 599.400 105.600 601.050 ;
        RECT 100.950 598.950 105.000 599.400 ;
        RECT 98.400 573.450 99.600 573.600 ;
        RECT 101.400 573.450 102.450 598.950 ;
        RECT 98.400 572.400 102.450 573.450 ;
        RECT 98.400 571.350 99.600 572.400 ;
      LAYER metal3 ;
        RECT 76.950 918.600 81.000 919.050 ;
        RECT 76.950 916.950 81.600 918.600 ;
        RECT 80.400 915.600 81.600 916.950 ;
        RECT 80.400 915.000 84.600 915.600 ;
        RECT 80.400 914.400 85.050 915.000 ;
        RECT 82.950 910.950 85.050 914.400 ;
        RECT 88.950 843.600 93.000 844.050 ;
        RECT 88.950 841.950 93.600 843.600 ;
        RECT 85.950 831.600 88.050 832.050 ;
        RECT 92.400 831.600 93.600 841.950 ;
        RECT 85.950 830.400 93.600 831.600 ;
        RECT 85.950 829.950 88.050 830.400 ;
        RECT 85.950 805.950 88.050 808.050 ;
        RECT 86.400 799.050 87.600 805.950 ;
        RECT 82.950 797.400 87.600 799.050 ;
        RECT 82.950 796.950 87.000 797.400 ;
        RECT 82.950 765.600 87.000 766.050 ;
        RECT 82.950 763.950 87.600 765.600 ;
        RECT 86.400 762.600 87.600 763.950 ;
        RECT 86.400 761.400 90.600 762.600 ;
        RECT 89.400 754.050 90.600 761.400 ;
        RECT 89.400 752.400 94.050 754.050 ;
        RECT 90.000 751.950 94.050 752.400 ;
        RECT 40.950 705.600 43.050 706.050 ;
        RECT 94.950 705.600 97.050 706.050 ;
        RECT 40.950 704.400 97.050 705.600 ;
        RECT 40.950 703.950 43.050 704.400 ;
        RECT 94.950 703.950 97.050 704.400 ;
        RECT 40.950 683.100 43.050 685.200 ;
        RECT 41.400 676.050 42.600 683.100 ;
        RECT 40.950 673.950 43.050 676.050 ;
        RECT 43.950 612.600 46.050 613.050 ;
        RECT 79.950 612.600 82.050 613.050 ;
        RECT 100.950 612.600 103.050 613.050 ;
        RECT 43.950 611.400 103.050 612.600 ;
        RECT 43.950 610.950 46.050 611.400 ;
        RECT 79.950 610.950 82.050 611.400 ;
        RECT 100.950 610.950 103.050 611.400 ;
        RECT 100.950 604.950 103.050 607.050 ;
        RECT 101.400 601.050 102.600 604.950 ;
        RECT 100.950 598.950 103.050 601.050 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal1 ;
        RECT 52.950 720.450 55.050 721.050 ;
        RECT 61.950 720.450 64.050 721.050 ;
        RECT 52.950 719.550 64.050 720.450 ;
        RECT 52.950 718.950 55.050 719.550 ;
        RECT 61.950 718.950 64.050 719.550 ;
        RECT 73.950 642.450 76.050 643.050 ;
        RECT 79.950 642.450 82.050 643.050 ;
        RECT 73.950 641.550 82.050 642.450 ;
        RECT 73.950 640.950 76.050 641.550 ;
        RECT 79.950 640.950 82.050 641.550 ;
      LAYER metal2 ;
        RECT 80.400 910.050 81.450 945.450 ;
        RECT 67.950 907.950 70.050 910.050 ;
        RECT 79.950 907.950 82.050 910.050 ;
        RECT 68.400 879.450 69.450 907.950 ;
        RECT 68.400 878.400 72.450 879.450 ;
        RECT 71.400 834.450 72.450 878.400 ;
        RECT 68.400 833.400 72.450 834.450 ;
        RECT 68.400 801.450 69.450 833.400 ;
        RECT 68.400 800.400 72.450 801.450 ;
        RECT 71.400 745.050 72.450 800.400 ;
        RECT 64.950 742.950 67.050 745.050 ;
        RECT 70.950 742.950 73.050 745.050 ;
        RECT 65.400 732.450 66.450 742.950 ;
        RECT 62.400 731.400 66.450 732.450 ;
        RECT 62.400 721.050 63.450 731.400 ;
        RECT 52.950 718.950 55.050 721.050 ;
        RECT 61.950 718.950 64.050 721.050 ;
        RECT 53.400 679.050 54.450 718.950 ;
        RECT 52.950 676.950 55.050 679.050 ;
        RECT 73.950 676.950 76.050 679.050 ;
        RECT 74.400 652.200 75.450 676.950 ;
        RECT 73.950 650.100 76.050 652.200 ;
        RECT 79.950 650.100 82.050 652.200 ;
        RECT 74.400 649.350 75.600 650.100 ;
        RECT 80.400 643.050 81.450 650.100 ;
        RECT 73.950 640.950 76.050 643.050 ;
        RECT 79.950 640.950 82.050 643.050 ;
        RECT 68.400 600.900 69.600 601.650 ;
        RECT 74.400 601.050 75.450 640.950 ;
        RECT 67.950 598.800 70.050 600.900 ;
        RECT 73.950 598.950 76.050 601.050 ;
      LAYER metal3 ;
        RECT 67.950 909.600 70.050 910.050 ;
        RECT 79.950 909.600 82.050 910.050 ;
        RECT 67.950 908.400 82.050 909.600 ;
        RECT 67.950 907.950 70.050 908.400 ;
        RECT 79.950 907.950 82.050 908.400 ;
        RECT 64.950 744.600 67.050 745.050 ;
        RECT 70.950 744.600 73.050 745.050 ;
        RECT 64.950 743.400 73.050 744.600 ;
        RECT 64.950 742.950 67.050 743.400 ;
        RECT 70.950 742.950 73.050 743.400 ;
        RECT 52.950 678.600 55.050 679.050 ;
        RECT 73.950 678.600 76.050 679.050 ;
        RECT 52.950 677.400 76.050 678.600 ;
        RECT 52.950 676.950 55.050 677.400 ;
        RECT 73.950 676.950 76.050 677.400 ;
        RECT 73.950 651.750 76.050 652.200 ;
        RECT 79.950 651.750 82.050 652.200 ;
        RECT 73.950 650.550 82.050 651.750 ;
        RECT 73.950 650.100 76.050 650.550 ;
        RECT 79.950 650.100 82.050 650.550 ;
        RECT 67.950 600.600 70.050 600.900 ;
        RECT 73.950 600.600 76.050 601.050 ;
        RECT 67.950 599.400 76.050 600.600 ;
        RECT 67.950 598.800 70.050 599.400 ;
        RECT 73.950 598.950 76.050 599.400 ;
    END
  END LoadCmd_i
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 310.950 426.450 313.050 427.050 ;
        RECT 319.950 426.450 322.050 427.050 ;
        RECT 310.950 425.550 322.050 426.450 ;
        RECT 310.950 424.950 313.050 425.550 ;
        RECT 319.950 424.950 322.050 425.550 ;
      LAYER metal2 ;
        RECT 317.400 489.000 318.600 490.650 ;
        RECT 316.950 484.950 319.050 489.000 ;
        RECT 338.400 488.400 339.600 490.650 ;
        RECT 338.400 487.050 339.450 488.400 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 338.400 454.050 339.450 484.950 ;
        RECT 337.950 451.950 340.050 454.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 320.400 427.050 321.450 445.950 ;
        RECT 310.950 424.950 313.050 427.050 ;
        RECT 319.950 424.950 322.050 427.050 ;
        RECT 227.400 410.400 228.600 412.650 ;
        RECT 227.400 400.050 228.450 410.400 ;
        RECT 19.950 397.950 22.050 400.050 ;
        RECT 226.950 397.950 229.050 400.050 ;
        RECT 16.950 372.450 19.050 373.200 ;
        RECT 20.400 372.450 21.450 397.950 ;
        RECT 227.400 394.050 228.450 397.950 ;
        RECT 311.400 394.050 312.450 424.950 ;
        RECT 226.950 391.950 229.050 394.050 ;
        RECT 310.950 391.950 313.050 394.050 ;
        RECT 16.950 371.400 21.450 372.450 ;
        RECT 16.950 371.100 19.050 371.400 ;
        RECT 17.400 370.350 18.600 371.100 ;
        RECT 17.400 333.450 18.600 334.650 ;
        RECT 20.400 333.450 21.450 371.400 ;
        RECT 17.400 332.400 21.450 333.450 ;
      LAYER metal3 ;
        RECT 316.950 486.600 319.050 487.050 ;
        RECT 337.950 486.600 340.050 487.050 ;
        RECT 316.950 485.400 340.050 486.600 ;
        RECT 316.950 484.950 319.050 485.400 ;
        RECT 337.950 484.950 340.050 485.400 ;
        RECT 337.950 453.600 340.050 454.050 ;
        RECT 329.400 452.400 340.050 453.600 ;
        RECT 319.950 447.600 322.050 448.050 ;
        RECT 329.400 447.600 330.600 452.400 ;
        RECT 337.950 451.950 340.050 452.400 ;
        RECT 319.950 446.400 330.600 447.600 ;
        RECT 319.950 445.950 322.050 446.400 ;
        RECT 19.950 399.600 22.050 400.050 ;
        RECT 226.950 399.600 229.050 400.050 ;
        RECT 19.950 398.400 229.050 399.600 ;
        RECT 19.950 397.950 22.050 398.400 ;
        RECT 226.950 397.950 229.050 398.400 ;
        RECT 226.950 393.600 229.050 394.050 ;
        RECT 310.950 393.600 313.050 394.050 ;
        RECT 226.950 392.400 313.050 393.600 ;
        RECT 226.950 391.950 229.050 392.400 ;
        RECT 310.950 391.950 313.050 392.400 ;
        RECT 16.950 372.600 19.050 373.200 ;
        RECT -3.600 371.400 19.050 372.600 ;
        RECT 16.950 371.100 19.050 371.400 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 4.950 601.950 7.050 604.050 ;
        RECT 5.400 598.050 6.450 601.950 ;
        RECT 17.400 600.000 18.600 601.650 ;
        RECT 4.950 595.950 7.050 598.050 ;
        RECT 16.950 595.950 19.050 600.000 ;
      LAYER metal3 ;
        RECT -3.600 603.600 -2.400 606.600 ;
        RECT 4.950 603.600 7.050 604.050 ;
        RECT -3.600 602.400 7.050 603.600 ;
        RECT 4.950 601.950 7.050 602.400 ;
        RECT 4.950 597.600 7.050 598.050 ;
        RECT 16.950 597.600 19.050 598.050 ;
        RECT 4.950 596.400 19.050 597.600 ;
        RECT 4.950 595.950 7.050 596.400 ;
        RECT 16.950 595.950 19.050 596.400 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 14.100 929.400 15.900 935.400 ;
        RECT 17.100 930.000 18.900 936.000 ;
        RECT 15.000 929.100 15.900 929.400 ;
        RECT 20.100 929.400 21.900 935.400 ;
        RECT 23.100 929.400 24.900 936.000 ;
        RECT 35.100 929.400 36.900 936.000 ;
        RECT 38.100 929.400 39.900 935.400 ;
        RECT 41.100 929.400 42.900 936.000 ;
        RECT 53.100 929.400 54.900 935.400 ;
        RECT 56.100 929.400 57.900 936.000 ;
        RECT 68.100 929.400 69.900 936.000 ;
        RECT 71.100 929.400 72.900 935.400 ;
        RECT 74.100 929.400 75.900 936.000 ;
        RECT 86.100 929.400 87.900 936.000 ;
        RECT 89.100 929.400 90.900 935.400 ;
        RECT 92.100 929.400 93.900 936.000 ;
        RECT 107.100 929.400 108.900 935.400 ;
        RECT 110.100 930.000 111.900 936.000 ;
        RECT 20.100 929.100 21.600 929.400 ;
        RECT 15.000 928.200 21.600 929.100 ;
        RECT 15.000 916.050 15.900 928.200 ;
        RECT 20.100 916.050 21.900 917.850 ;
        RECT 38.100 916.050 39.300 929.400 ;
        RECT 48.000 918.450 52.050 919.050 ;
        RECT 47.550 916.950 52.050 918.450 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 19.950 913.950 22.050 916.050 ;
        RECT 22.950 913.950 25.050 916.050 ;
        RECT 34.950 913.950 37.050 916.050 ;
        RECT 37.950 913.950 40.050 916.050 ;
        RECT 40.950 913.950 43.050 916.050 ;
        RECT 15.000 910.200 15.900 913.950 ;
        RECT 17.100 912.150 18.900 913.950 ;
        RECT 23.100 912.150 24.900 913.950 ;
        RECT 35.250 912.150 37.050 913.950 ;
        RECT 15.000 909.000 18.300 910.200 ;
        RECT 16.500 900.600 18.300 909.000 ;
        RECT 23.100 900.000 24.900 909.600 ;
        RECT 38.100 908.700 39.300 913.950 ;
        RECT 41.100 912.150 42.900 913.950 ;
        RECT 47.550 913.050 48.450 916.950 ;
        RECT 53.700 916.050 54.900 929.400 ;
        RECT 56.100 916.050 57.900 917.850 ;
        RECT 71.100 916.050 72.300 929.400 ;
        RECT 89.700 916.050 90.900 929.400 ;
        RECT 108.000 929.100 108.900 929.400 ;
        RECT 113.100 929.400 114.900 935.400 ;
        RECT 116.100 929.400 117.900 936.000 ;
        RECT 113.100 929.100 114.600 929.400 ;
        RECT 108.000 928.200 114.600 929.100 ;
        RECT 108.000 916.050 108.900 928.200 ;
        RECT 131.400 923.400 133.200 936.000 ;
        RECT 136.500 924.900 138.300 935.400 ;
        RECT 139.500 929.400 141.300 936.000 ;
        RECT 155.700 929.400 157.500 936.000 ;
        RECT 139.200 926.100 141.000 927.900 ;
        RECT 156.000 926.100 157.800 927.900 ;
        RECT 158.700 924.900 160.500 935.400 ;
        RECT 136.500 923.400 138.900 924.900 ;
        RECT 115.950 921.450 118.050 922.050 ;
        RECT 121.950 921.450 124.050 922.050 ;
        RECT 115.950 920.550 124.050 921.450 ;
        RECT 115.950 919.950 118.050 920.550 ;
        RECT 121.950 919.950 124.050 920.550 ;
        RECT 113.100 916.050 114.900 917.850 ;
        RECT 131.100 916.050 132.900 917.850 ;
        RECT 137.700 916.050 138.900 923.400 ;
        RECT 158.100 923.400 160.500 924.900 ;
        RECT 163.800 923.400 165.600 936.000 ;
        RECT 176.700 929.400 178.500 936.000 ;
        RECT 177.000 926.100 178.800 927.900 ;
        RECT 179.700 924.900 181.500 935.400 ;
        RECT 179.100 923.400 181.500 924.900 ;
        RECT 184.800 923.400 186.600 936.000 ;
        RECT 197.100 924.300 198.900 935.400 ;
        RECT 200.100 925.500 201.900 936.000 ;
        RECT 197.100 923.400 201.600 924.300 ;
        RECT 204.600 923.400 206.400 935.400 ;
        RECT 209.100 925.500 210.900 936.000 ;
        RECT 212.100 924.600 213.900 935.400 ;
        RECT 158.100 916.050 159.300 923.400 ;
        RECT 164.100 916.050 165.900 917.850 ;
        RECT 179.100 916.050 180.300 923.400 ;
        RECT 199.500 921.300 201.600 923.400 ;
        RECT 205.200 922.050 206.400 923.400 ;
        RECT 209.100 923.400 213.900 924.600 ;
        RECT 227.100 923.400 228.900 936.000 ;
        RECT 232.200 924.600 234.000 935.400 ;
        RECT 248.100 929.400 249.900 936.000 ;
        RECT 251.100 929.400 252.900 935.400 ;
        RECT 254.100 929.400 255.900 936.000 ;
        RECT 269.100 929.400 270.900 936.000 ;
        RECT 272.100 929.400 273.900 935.400 ;
        RECT 275.100 930.000 276.900 936.000 ;
        RECT 230.400 923.400 234.000 924.600 ;
        RECT 209.100 922.500 211.200 923.400 ;
        RECT 205.200 921.000 206.700 922.050 ;
        RECT 202.800 919.500 204.900 919.800 ;
        RECT 185.100 916.050 186.900 917.850 ;
        RECT 201.000 917.700 204.900 919.500 ;
        RECT 205.800 919.050 206.700 921.000 ;
        RECT 205.800 916.950 207.900 919.050 ;
        RECT 205.800 916.800 207.300 916.950 ;
        RECT 202.200 916.050 204.000 916.500 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 55.950 913.950 58.050 916.050 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 73.950 913.950 76.050 916.050 ;
        RECT 85.950 913.950 88.050 916.050 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 106.950 913.950 109.050 916.050 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 130.950 913.950 133.050 916.050 ;
        RECT 133.950 913.950 136.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 154.950 913.950 157.050 916.050 ;
        RECT 157.950 913.950 160.050 916.050 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 175.950 913.950 178.050 916.050 ;
        RECT 178.950 913.950 181.050 916.050 ;
        RECT 181.950 913.950 184.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 197.100 914.700 204.000 916.050 ;
        RECT 204.900 915.900 207.300 916.800 ;
        RECT 211.800 916.050 213.600 917.850 ;
        RECT 227.250 916.050 229.050 917.850 ;
        RECT 230.400 916.050 231.300 923.400 ;
        RECT 233.100 916.050 234.900 917.850 ;
        RECT 251.100 916.050 252.300 929.400 ;
        RECT 272.400 929.100 273.900 929.400 ;
        RECT 278.100 929.400 279.900 935.400 ;
        RECT 290.100 929.400 291.900 936.000 ;
        RECT 293.100 929.400 294.900 935.400 ;
        RECT 305.100 929.400 306.900 935.400 ;
        RECT 308.100 930.000 309.900 936.000 ;
        RECT 278.100 929.100 279.000 929.400 ;
        RECT 272.400 928.200 279.000 929.100 ;
        RECT 272.100 916.050 273.900 917.850 ;
        RECT 278.100 916.050 279.000 928.200 ;
        RECT 290.100 916.050 291.900 917.850 ;
        RECT 293.100 916.050 294.300 929.400 ;
        RECT 306.000 929.100 306.900 929.400 ;
        RECT 311.100 929.400 312.900 935.400 ;
        RECT 314.100 929.400 315.900 936.000 ;
        RECT 329.100 929.400 330.900 936.000 ;
        RECT 332.100 929.400 333.900 935.400 ;
        RECT 335.100 929.400 336.900 936.000 ;
        RECT 347.700 929.400 349.500 936.000 ;
        RECT 311.100 929.100 312.600 929.400 ;
        RECT 306.000 928.200 312.600 929.100 ;
        RECT 306.000 916.050 306.900 928.200 ;
        RECT 307.950 921.450 310.050 922.050 ;
        RECT 328.950 921.450 331.050 922.050 ;
        RECT 307.950 920.550 331.050 921.450 ;
        RECT 307.950 919.950 310.050 920.550 ;
        RECT 328.950 919.950 331.050 920.550 ;
        RECT 311.100 916.050 312.900 917.850 ;
        RECT 332.700 916.050 333.900 929.400 ;
        RECT 348.000 926.100 349.800 927.900 ;
        RECT 350.700 924.900 352.500 935.400 ;
        RECT 350.100 923.400 352.500 924.900 ;
        RECT 355.800 923.400 357.600 936.000 ;
        RECT 368.100 929.400 369.900 936.000 ;
        RECT 371.100 929.400 372.900 935.400 ;
        RECT 374.100 929.400 375.900 936.000 ;
        RECT 386.700 929.400 388.500 936.000 ;
        RECT 350.100 916.050 351.300 923.400 ;
        RECT 356.100 916.050 357.900 917.850 ;
        RECT 371.100 916.050 372.300 929.400 ;
        RECT 387.000 926.100 388.800 927.900 ;
        RECT 389.700 924.900 391.500 935.400 ;
        RECT 389.100 923.400 391.500 924.900 ;
        RECT 394.800 923.400 396.600 936.000 ;
        RECT 410.100 923.400 411.900 936.000 ;
        RECT 415.200 924.600 417.000 935.400 ;
        RECT 431.700 929.400 433.500 936.000 ;
        RECT 421.950 925.950 427.050 928.050 ;
        RECT 432.000 926.100 433.800 927.900 ;
        RECT 434.700 924.900 436.500 935.400 ;
        RECT 413.400 923.400 417.000 924.600 ;
        RECT 434.100 923.400 436.500 924.900 ;
        RECT 439.800 923.400 441.600 936.000 ;
        RECT 452.100 929.400 453.900 936.000 ;
        RECT 455.100 929.400 456.900 935.400 ;
        RECT 458.100 929.400 459.900 936.000 ;
        RECT 389.100 916.050 390.300 923.400 ;
        RECT 391.950 921.450 394.050 922.050 ;
        RECT 400.950 921.450 403.050 922.050 ;
        RECT 391.950 920.550 403.050 921.450 ;
        RECT 391.950 919.950 394.050 920.550 ;
        RECT 400.950 919.950 403.050 920.550 ;
        RECT 395.100 916.050 396.900 917.850 ;
        RECT 410.250 916.050 412.050 917.850 ;
        RECT 413.400 916.050 414.300 923.400 ;
        RECT 416.100 916.050 417.900 917.850 ;
        RECT 434.100 916.050 435.300 923.400 ;
        RECT 447.000 918.450 451.050 919.050 ;
        RECT 440.100 916.050 441.900 917.850 ;
        RECT 446.550 916.950 451.050 918.450 ;
        RECT 197.100 913.950 199.200 914.700 ;
        RECT 43.950 911.550 48.450 913.050 ;
        RECT 43.950 910.950 48.000 911.550 ;
        RECT 38.100 907.800 42.300 908.700 ;
        RECT 35.400 900.000 37.200 906.600 ;
        RECT 40.500 900.600 42.300 907.800 ;
        RECT 53.700 903.600 54.900 913.950 ;
        RECT 68.250 912.150 70.050 913.950 ;
        RECT 55.950 909.450 58.050 910.050 ;
        RECT 61.950 909.450 64.050 910.050 ;
        RECT 55.950 908.550 64.050 909.450 ;
        RECT 55.950 907.950 58.050 908.550 ;
        RECT 61.950 907.950 64.050 908.550 ;
        RECT 71.100 908.700 72.300 913.950 ;
        RECT 74.100 912.150 75.900 913.950 ;
        RECT 86.100 912.150 87.900 913.950 ;
        RECT 89.700 908.700 90.900 913.950 ;
        RECT 91.950 912.150 93.750 913.950 ;
        RECT 108.000 910.200 108.900 913.950 ;
        RECT 110.100 912.150 111.900 913.950 ;
        RECT 116.100 912.150 117.900 913.950 ;
        RECT 134.100 912.150 135.900 913.950 ;
        RECT 108.000 909.000 111.300 910.200 ;
        RECT 137.700 909.600 138.900 913.950 ;
        RECT 140.100 912.150 141.900 913.950 ;
        RECT 155.100 912.150 156.900 913.950 ;
        RECT 158.100 909.600 159.300 913.950 ;
        RECT 161.100 912.150 162.900 913.950 ;
        RECT 176.100 912.150 177.900 913.950 ;
        RECT 179.100 909.600 180.300 913.950 ;
        RECT 182.100 912.150 183.900 913.950 ;
        RECT 197.400 912.150 199.200 913.950 ;
        RECT 202.200 911.400 204.000 913.200 ;
        RECT 71.100 907.800 75.300 908.700 ;
        RECT 53.100 900.600 54.900 903.600 ;
        RECT 56.100 900.000 57.900 903.600 ;
        RECT 68.400 900.000 70.200 906.600 ;
        RECT 73.500 900.600 75.300 907.800 ;
        RECT 86.700 907.800 90.900 908.700 ;
        RECT 86.700 900.600 88.500 907.800 ;
        RECT 91.800 900.000 93.600 906.600 ;
        RECT 109.500 900.600 111.300 909.000 ;
        RECT 116.100 900.000 117.900 909.600 ;
        RECT 137.700 908.700 141.300 909.600 ;
        RECT 131.100 905.700 138.900 907.050 ;
        RECT 131.100 900.600 132.900 905.700 ;
        RECT 134.100 900.000 135.900 904.800 ;
        RECT 137.100 900.600 138.900 905.700 ;
        RECT 140.100 906.600 141.300 908.700 ;
        RECT 155.700 908.700 159.300 909.600 ;
        RECT 176.700 908.700 180.300 909.600 ;
        RECT 201.900 909.300 204.000 911.400 ;
        RECT 155.700 906.600 156.900 908.700 ;
        RECT 140.100 900.600 141.900 906.600 ;
        RECT 155.100 900.600 156.900 906.600 ;
        RECT 158.100 905.700 165.900 907.050 ;
        RECT 176.700 906.600 177.900 908.700 ;
        RECT 197.700 908.400 204.000 909.300 ;
        RECT 204.900 910.200 206.100 915.900 ;
        RECT 207.300 913.200 209.100 915.000 ;
        RECT 211.800 913.950 213.900 916.050 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 289.950 913.950 292.050 916.050 ;
        RECT 292.950 913.950 295.050 916.050 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 307.950 913.950 310.050 916.050 ;
        RECT 310.950 913.950 313.050 916.050 ;
        RECT 313.950 913.950 316.050 916.050 ;
        RECT 328.950 913.950 331.050 916.050 ;
        RECT 331.950 913.950 334.050 916.050 ;
        RECT 334.950 913.950 337.050 916.050 ;
        RECT 346.950 913.950 349.050 916.050 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 355.950 913.950 358.050 916.050 ;
        RECT 367.950 913.950 370.050 916.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 373.950 913.950 376.050 916.050 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 388.950 913.950 391.050 916.050 ;
        RECT 391.950 913.950 394.050 916.050 ;
        RECT 394.950 913.950 397.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 412.950 913.950 415.050 916.050 ;
        RECT 415.950 913.950 418.050 916.050 ;
        RECT 430.950 913.950 433.050 916.050 ;
        RECT 433.950 913.950 436.050 916.050 ;
        RECT 436.950 913.950 439.050 916.050 ;
        RECT 439.950 913.950 442.050 916.050 ;
        RECT 207.000 911.100 209.100 913.200 ;
        RECT 158.100 900.600 159.900 905.700 ;
        RECT 161.100 900.000 162.900 904.800 ;
        RECT 164.100 900.600 165.900 905.700 ;
        RECT 176.100 900.600 177.900 906.600 ;
        RECT 179.100 905.700 186.900 907.050 ;
        RECT 197.700 906.600 198.900 908.400 ;
        RECT 204.900 908.100 207.900 910.200 ;
        RECT 204.900 906.600 206.100 908.100 ;
        RECT 209.100 907.500 211.200 908.700 ;
        RECT 209.100 906.600 213.900 907.500 ;
        RECT 179.100 900.600 180.900 905.700 ;
        RECT 182.100 900.000 183.900 904.800 ;
        RECT 185.100 900.600 186.900 905.700 ;
        RECT 197.100 900.600 198.900 906.600 ;
        RECT 200.100 900.000 201.900 905.700 ;
        RECT 204.600 900.600 206.400 906.600 ;
        RECT 209.100 900.000 210.900 905.700 ;
        RECT 212.100 900.600 213.900 906.600 ;
        RECT 230.400 903.600 231.300 913.950 ;
        RECT 248.250 912.150 250.050 913.950 ;
        RECT 251.100 908.700 252.300 913.950 ;
        RECT 254.100 912.150 255.900 913.950 ;
        RECT 269.100 912.150 270.900 913.950 ;
        RECT 275.100 912.150 276.900 913.950 ;
        RECT 278.100 910.200 279.000 913.950 ;
        RECT 251.100 907.800 255.300 908.700 ;
        RECT 227.100 900.000 228.900 903.600 ;
        RECT 230.100 900.600 231.900 903.600 ;
        RECT 233.100 900.000 234.900 903.600 ;
        RECT 248.400 900.000 250.200 906.600 ;
        RECT 253.500 900.600 255.300 907.800 ;
        RECT 269.100 900.000 270.900 909.600 ;
        RECT 275.700 909.000 279.000 910.200 ;
        RECT 275.700 900.600 277.500 909.000 ;
        RECT 293.100 903.600 294.300 913.950 ;
        RECT 301.950 912.450 304.050 913.050 ;
        RECT 296.550 912.000 304.050 912.450 ;
        RECT 295.950 911.550 304.050 912.000 ;
        RECT 295.950 907.950 298.050 911.550 ;
        RECT 301.950 910.950 304.050 911.550 ;
        RECT 306.000 910.200 306.900 913.950 ;
        RECT 308.100 912.150 309.900 913.950 ;
        RECT 314.100 912.150 315.900 913.950 ;
        RECT 329.100 912.150 330.900 913.950 ;
        RECT 306.000 909.000 309.300 910.200 ;
        RECT 290.100 900.000 291.900 903.600 ;
        RECT 293.100 900.600 294.900 903.600 ;
        RECT 307.500 900.600 309.300 909.000 ;
        RECT 314.100 900.000 315.900 909.600 ;
        RECT 332.700 908.700 333.900 913.950 ;
        RECT 334.950 912.150 336.750 913.950 ;
        RECT 347.100 912.150 348.900 913.950 ;
        RECT 350.100 909.600 351.300 913.950 ;
        RECT 353.100 912.150 354.900 913.950 ;
        RECT 368.250 912.150 370.050 913.950 ;
        RECT 329.700 907.800 333.900 908.700 ;
        RECT 347.700 908.700 351.300 909.600 ;
        RECT 371.100 908.700 372.300 913.950 ;
        RECT 374.100 912.150 375.900 913.950 ;
        RECT 386.100 912.150 387.900 913.950 ;
        RECT 389.100 909.600 390.300 913.950 ;
        RECT 392.100 912.150 393.900 913.950 ;
        RECT 386.700 908.700 390.300 909.600 ;
        RECT 329.700 900.600 331.500 907.800 ;
        RECT 347.700 906.600 348.900 908.700 ;
        RECT 371.100 907.800 375.300 908.700 ;
        RECT 334.800 900.000 336.600 906.600 ;
        RECT 347.100 900.600 348.900 906.600 ;
        RECT 350.100 905.700 357.900 907.050 ;
        RECT 350.100 900.600 351.900 905.700 ;
        RECT 353.100 900.000 354.900 904.800 ;
        RECT 356.100 900.600 357.900 905.700 ;
        RECT 368.400 900.000 370.200 906.600 ;
        RECT 373.500 900.600 375.300 907.800 ;
        RECT 386.700 906.600 387.900 908.700 ;
        RECT 386.100 900.600 387.900 906.600 ;
        RECT 389.100 905.700 396.900 907.050 ;
        RECT 389.100 900.600 390.900 905.700 ;
        RECT 392.100 900.000 393.900 904.800 ;
        RECT 395.100 900.600 396.900 905.700 ;
        RECT 413.400 903.600 414.300 913.950 ;
        RECT 431.100 912.150 432.900 913.950 ;
        RECT 434.100 909.600 435.300 913.950 ;
        RECT 437.100 912.150 438.900 913.950 ;
        RECT 446.550 913.050 447.450 916.950 ;
        RECT 455.100 916.050 456.300 929.400 ;
        RECT 470.400 923.400 472.200 936.000 ;
        RECT 475.500 924.900 477.300 935.400 ;
        RECT 478.500 929.400 480.300 936.000 ;
        RECT 478.200 926.100 480.000 927.900 ;
        RECT 475.500 923.400 477.900 924.900 ;
        RECT 494.400 923.400 496.200 936.000 ;
        RECT 499.500 924.900 501.300 935.400 ;
        RECT 502.500 929.400 504.300 936.000 ;
        RECT 515.700 929.400 517.500 936.000 ;
        RECT 502.200 926.100 504.000 927.900 ;
        RECT 516.000 926.100 517.800 927.900 ;
        RECT 518.700 924.900 520.500 935.400 ;
        RECT 499.500 923.400 501.900 924.900 ;
        RECT 470.100 916.050 471.900 917.850 ;
        RECT 476.700 916.050 477.900 923.400 ;
        RECT 494.100 916.050 495.900 917.850 ;
        RECT 500.700 916.050 501.900 923.400 ;
        RECT 518.100 923.400 520.500 924.900 ;
        RECT 523.800 923.400 525.600 936.000 ;
        RECT 539.100 923.400 540.900 936.000 ;
        RECT 544.200 924.600 546.000 935.400 ;
        RECT 557.100 929.400 558.900 935.400 ;
        RECT 560.100 929.400 561.900 936.000 ;
        RECT 542.400 923.400 546.000 924.600 ;
        RECT 518.100 916.050 519.300 923.400 ;
        RECT 524.100 916.050 525.900 917.850 ;
        RECT 539.250 916.050 541.050 917.850 ;
        RECT 542.400 916.050 543.300 923.400 ;
        RECT 545.100 916.050 546.900 917.850 ;
        RECT 557.700 916.050 558.900 929.400 ;
        RECT 572.100 924.600 573.900 935.400 ;
        RECT 575.100 925.500 576.900 936.000 ;
        RECT 578.100 934.500 585.900 935.400 ;
        RECT 578.100 924.600 579.900 934.500 ;
        RECT 572.100 923.700 579.900 924.600 ;
        RECT 581.100 922.500 582.900 933.600 ;
        RECT 584.100 923.400 585.900 934.500 ;
        RECT 599.100 923.400 600.900 936.000 ;
        RECT 604.200 924.600 606.000 935.400 ;
        RECT 617.700 929.400 619.500 936.000 ;
        RECT 618.000 926.100 619.800 927.900 ;
        RECT 620.700 924.900 622.500 935.400 ;
        RECT 602.400 923.400 606.000 924.600 ;
        RECT 620.100 923.400 622.500 924.900 ;
        RECT 625.800 923.400 627.600 936.000 ;
        RECT 638.100 929.400 639.900 935.400 ;
        RECT 641.100 929.400 642.900 936.000 ;
        RECT 578.100 921.600 582.900 922.500 ;
        RECT 560.100 916.050 561.900 917.850 ;
        RECT 575.250 916.050 577.050 917.850 ;
        RECT 578.100 916.050 579.000 921.600 ;
        RECT 581.100 916.050 582.900 917.850 ;
        RECT 599.250 916.050 601.050 917.850 ;
        RECT 602.400 916.050 603.300 923.400 ;
        RECT 605.100 916.050 606.900 917.850 ;
        RECT 620.100 916.050 621.300 923.400 ;
        RECT 626.100 916.050 627.900 917.850 ;
        RECT 638.700 916.050 639.900 929.400 ;
        RECT 656.100 923.400 657.900 936.000 ;
        RECT 659.100 923.400 660.900 935.400 ;
        RECT 662.100 923.400 663.900 936.000 ;
        RECT 674.100 923.400 675.900 935.400 ;
        RECT 677.100 924.300 678.900 935.400 ;
        RECT 680.100 925.200 681.900 936.000 ;
        RECT 683.100 924.300 684.900 935.400 ;
        RECT 698.700 929.400 700.500 936.000 ;
        RECT 699.000 926.100 700.800 927.900 ;
        RECT 701.700 924.900 703.500 935.400 ;
        RECT 677.100 923.400 684.900 924.300 ;
        RECT 701.100 923.400 703.500 924.900 ;
        RECT 706.800 923.400 708.600 936.000 ;
        RECT 719.100 923.400 720.900 935.400 ;
        RECT 722.100 924.000 723.900 936.000 ;
        RECT 725.100 929.400 726.900 935.400 ;
        RECT 728.100 929.400 729.900 936.000 ;
        RECT 641.100 916.050 642.900 917.850 ;
        RECT 659.550 916.050 660.600 923.400 ;
        RECT 674.400 916.050 675.300 923.400 ;
        RECT 679.950 916.050 681.750 917.850 ;
        RECT 701.100 916.050 702.300 923.400 ;
        RECT 707.100 916.050 708.900 917.850 ;
        RECT 719.700 916.050 720.600 923.400 ;
        RECT 723.000 916.050 724.800 917.850 ;
        RECT 451.950 913.950 454.050 916.050 ;
        RECT 454.950 913.950 457.050 916.050 ;
        RECT 457.950 913.950 460.050 916.050 ;
        RECT 469.950 913.950 472.050 916.050 ;
        RECT 472.950 913.950 475.050 916.050 ;
        RECT 475.950 913.950 478.050 916.050 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 493.950 913.950 496.050 916.050 ;
        RECT 496.950 913.950 499.050 916.050 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 514.950 913.950 517.050 916.050 ;
        RECT 517.950 913.950 520.050 916.050 ;
        RECT 520.950 913.950 523.050 916.050 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 538.950 913.950 541.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 556.950 913.950 559.050 916.050 ;
        RECT 559.950 913.950 562.050 916.050 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 574.950 913.950 577.050 916.050 ;
        RECT 577.950 913.950 580.050 916.050 ;
        RECT 580.950 913.950 583.050 916.050 ;
        RECT 583.950 913.950 586.050 916.050 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 601.950 913.950 604.050 916.050 ;
        RECT 604.950 913.950 607.050 916.050 ;
        RECT 616.950 913.950 619.050 916.050 ;
        RECT 619.950 913.950 622.050 916.050 ;
        RECT 622.950 913.950 625.050 916.050 ;
        RECT 625.950 913.950 628.050 916.050 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 640.950 913.950 643.050 916.050 ;
        RECT 656.400 913.950 660.600 916.050 ;
        RECT 661.500 913.950 663.600 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 676.950 913.950 679.050 916.050 ;
        RECT 679.950 913.950 682.050 916.050 ;
        RECT 682.950 913.950 685.050 916.050 ;
        RECT 697.950 913.950 700.050 916.050 ;
        RECT 700.950 913.950 703.050 916.050 ;
        RECT 703.950 913.950 706.050 916.050 ;
        RECT 706.950 913.950 709.050 916.050 ;
        RECT 719.100 913.950 721.200 916.050 ;
        RECT 722.400 913.950 724.500 916.050 ;
        RECT 442.950 911.550 447.450 913.050 ;
        RECT 452.250 912.150 454.050 913.950 ;
        RECT 442.950 910.950 447.000 911.550 ;
        RECT 431.700 908.700 435.300 909.600 ;
        RECT 455.100 908.700 456.300 913.950 ;
        RECT 458.100 912.150 459.900 913.950 ;
        RECT 473.100 912.150 474.900 913.950 ;
        RECT 476.700 909.600 477.900 913.950 ;
        RECT 479.100 912.150 480.900 913.950 ;
        RECT 497.100 912.150 498.900 913.950 ;
        RECT 500.700 909.600 501.900 913.950 ;
        RECT 503.100 912.150 504.900 913.950 ;
        RECT 515.100 912.150 516.900 913.950 ;
        RECT 518.100 909.600 519.300 913.950 ;
        RECT 521.100 912.150 522.900 913.950 ;
        RECT 476.700 908.700 480.300 909.600 ;
        RECT 500.700 908.700 504.300 909.600 ;
        RECT 431.700 906.600 432.900 908.700 ;
        RECT 455.100 907.800 459.300 908.700 ;
        RECT 410.100 900.000 411.900 903.600 ;
        RECT 413.100 900.600 414.900 903.600 ;
        RECT 416.100 900.000 417.900 903.600 ;
        RECT 431.100 900.600 432.900 906.600 ;
        RECT 434.100 905.700 441.900 907.050 ;
        RECT 434.100 900.600 435.900 905.700 ;
        RECT 437.100 900.000 438.900 904.800 ;
        RECT 440.100 900.600 441.900 905.700 ;
        RECT 452.400 900.000 454.200 906.600 ;
        RECT 457.500 900.600 459.300 907.800 ;
        RECT 470.100 905.700 477.900 907.050 ;
        RECT 470.100 900.600 471.900 905.700 ;
        RECT 473.100 900.000 474.900 904.800 ;
        RECT 476.100 900.600 477.900 905.700 ;
        RECT 479.100 906.600 480.300 908.700 ;
        RECT 479.100 900.600 480.900 906.600 ;
        RECT 494.100 905.700 501.900 907.050 ;
        RECT 494.100 900.600 495.900 905.700 ;
        RECT 497.100 900.000 498.900 904.800 ;
        RECT 500.100 900.600 501.900 905.700 ;
        RECT 503.100 906.600 504.300 908.700 ;
        RECT 515.700 908.700 519.300 909.600 ;
        RECT 515.700 906.600 516.900 908.700 ;
        RECT 503.100 900.600 504.900 906.600 ;
        RECT 515.100 900.600 516.900 906.600 ;
        RECT 518.100 905.700 525.900 907.050 ;
        RECT 518.100 900.600 519.900 905.700 ;
        RECT 521.100 900.000 522.900 904.800 ;
        RECT 524.100 900.600 525.900 905.700 ;
        RECT 542.400 903.600 543.300 913.950 ;
        RECT 557.700 903.600 558.900 913.950 ;
        RECT 572.250 912.150 574.050 913.950 ;
        RECT 559.950 909.450 562.050 910.050 ;
        RECT 574.950 909.450 577.050 909.750 ;
        RECT 559.950 908.550 577.050 909.450 ;
        RECT 559.950 907.950 562.050 908.550 ;
        RECT 574.950 907.650 577.050 908.550 ;
        RECT 578.100 906.600 579.300 913.950 ;
        RECT 584.100 912.150 585.900 913.950 ;
        RECT 580.950 909.450 583.050 910.050 ;
        RECT 589.950 909.450 592.050 910.050 ;
        RECT 580.950 908.550 592.050 909.450 ;
        RECT 580.950 907.950 583.050 908.550 ;
        RECT 589.950 907.950 592.050 908.550 ;
        RECT 539.100 900.000 540.900 903.600 ;
        RECT 542.100 900.600 543.900 903.600 ;
        RECT 545.100 900.000 546.900 903.600 ;
        RECT 557.100 900.600 558.900 903.600 ;
        RECT 560.100 900.000 561.900 903.600 ;
        RECT 572.700 900.000 574.500 906.600 ;
        RECT 577.200 900.600 579.000 906.600 ;
        RECT 581.700 900.000 583.500 906.600 ;
        RECT 602.400 903.600 603.300 913.950 ;
        RECT 617.100 912.150 618.900 913.950 ;
        RECT 620.100 909.600 621.300 913.950 ;
        RECT 623.100 912.150 624.900 913.950 ;
        RECT 617.700 908.700 621.300 909.600 ;
        RECT 617.700 906.600 618.900 908.700 ;
        RECT 599.100 900.000 600.900 903.600 ;
        RECT 602.100 900.600 603.900 903.600 ;
        RECT 605.100 900.000 606.900 903.600 ;
        RECT 617.100 900.600 618.900 906.600 ;
        RECT 620.100 905.700 627.900 907.050 ;
        RECT 620.100 900.600 621.900 905.700 ;
        RECT 623.100 900.000 624.900 904.800 ;
        RECT 626.100 900.600 627.900 905.700 ;
        RECT 638.700 903.600 639.900 913.950 ;
        RECT 659.550 906.600 660.600 913.950 ;
        RECT 661.800 912.150 663.600 913.950 ;
        RECT 674.400 906.600 675.300 913.950 ;
        RECT 676.950 912.150 678.750 913.950 ;
        RECT 683.100 912.150 684.900 913.950 ;
        RECT 698.100 912.150 699.900 913.950 ;
        RECT 701.100 909.600 702.300 913.950 ;
        RECT 704.100 912.150 705.900 913.950 ;
        RECT 698.700 908.700 702.300 909.600 ;
        RECT 698.700 906.600 699.900 908.700 ;
        RECT 638.100 900.600 639.900 903.600 ;
        RECT 641.100 900.000 642.900 903.600 ;
        RECT 656.100 900.000 657.900 906.600 ;
        RECT 659.100 900.600 660.900 906.600 ;
        RECT 662.100 900.000 663.900 906.600 ;
        RECT 674.400 905.400 679.500 906.600 ;
        RECT 674.700 900.000 676.500 903.600 ;
        RECT 677.700 900.600 679.500 905.400 ;
        RECT 682.200 900.000 684.000 906.600 ;
        RECT 698.100 900.600 699.900 906.600 ;
        RECT 701.100 905.700 708.900 907.050 ;
        RECT 701.100 900.600 702.900 905.700 ;
        RECT 704.100 900.000 705.900 904.800 ;
        RECT 707.100 900.600 708.900 905.700 ;
        RECT 719.700 906.600 720.600 913.950 ;
        RECT 726.000 909.300 726.900 929.400 ;
        RECT 740.100 923.400 741.900 935.400 ;
        RECT 744.600 923.400 746.400 936.000 ;
        RECT 747.600 924.900 749.400 935.400 ;
        RECT 764.700 929.400 766.500 936.000 ;
        RECT 765.000 926.100 766.800 927.900 ;
        RECT 767.700 924.900 769.500 935.400 ;
        RECT 747.600 923.400 750.000 924.900 ;
        RECT 740.100 921.900 741.300 923.400 ;
        RECT 740.100 920.700 747.900 921.900 ;
        RECT 746.100 920.100 747.900 920.700 ;
        RECT 744.000 916.050 745.800 917.850 ;
        RECT 727.800 913.950 729.900 916.050 ;
        RECT 740.100 913.950 742.200 916.050 ;
        RECT 743.400 913.950 745.500 916.050 ;
        RECT 727.950 912.150 729.750 913.950 ;
        RECT 740.400 912.150 742.200 913.950 ;
        RECT 746.700 909.600 747.600 920.100 ;
        RECT 748.800 916.050 750.000 923.400 ;
        RECT 767.100 923.400 769.500 924.900 ;
        RECT 772.800 923.400 774.600 936.000 ;
        RECT 785.100 929.400 786.900 935.400 ;
        RECT 788.100 930.000 789.900 936.000 ;
        RECT 786.000 929.100 786.900 929.400 ;
        RECT 791.100 929.400 792.900 935.400 ;
        RECT 794.100 929.400 795.900 936.000 ;
        RECT 809.100 929.400 810.900 935.400 ;
        RECT 812.100 929.400 813.900 936.000 ;
        RECT 824.100 929.400 825.900 936.000 ;
        RECT 827.100 929.400 828.900 935.400 ;
        RECT 830.100 930.000 831.900 936.000 ;
        RECT 791.100 929.100 792.600 929.400 ;
        RECT 786.000 928.200 792.600 929.100 ;
        RECT 767.100 916.050 768.300 923.400 ;
        RECT 773.100 916.050 774.900 917.850 ;
        RECT 786.000 916.050 786.900 928.200 ;
        RECT 796.950 918.450 799.050 919.050 ;
        RECT 802.950 918.450 805.050 919.050 ;
        RECT 791.100 916.050 792.900 917.850 ;
        RECT 796.950 917.550 805.050 918.450 ;
        RECT 796.950 916.950 799.050 917.550 ;
        RECT 802.950 916.950 805.050 917.550 ;
        RECT 809.700 916.050 810.900 929.400 ;
        RECT 827.400 929.100 828.900 929.400 ;
        RECT 833.100 929.400 834.900 935.400 ;
        RECT 833.100 929.100 834.000 929.400 ;
        RECT 827.400 928.200 834.000 929.100 ;
        RECT 812.100 916.050 813.900 917.850 ;
        RECT 827.100 916.050 828.900 917.850 ;
        RECT 833.100 916.050 834.000 928.200 ;
        RECT 845.100 924.300 846.900 935.400 ;
        RECT 848.100 925.200 849.900 936.000 ;
        RECT 851.100 924.300 852.900 935.400 ;
        RECT 845.100 923.400 852.900 924.300 ;
        RECT 854.100 923.400 855.900 935.400 ;
        RECT 869.700 929.400 871.500 936.000 ;
        RECT 870.000 926.100 871.800 927.900 ;
        RECT 872.700 924.900 874.500 935.400 ;
        RECT 872.100 923.400 874.500 924.900 ;
        RECT 877.800 923.400 879.600 936.000 ;
        RECT 890.400 923.400 892.200 936.000 ;
        RECT 895.500 924.900 897.300 935.400 ;
        RECT 898.500 929.400 900.300 936.000 ;
        RECT 914.100 929.400 915.900 936.000 ;
        RECT 917.100 929.400 918.900 935.400 ;
        RECT 898.200 926.100 900.000 927.900 ;
        RECT 895.500 923.400 897.900 924.900 ;
        RECT 848.250 916.050 850.050 917.850 ;
        RECT 854.700 916.050 855.600 923.400 ;
        RECT 872.100 916.050 873.300 923.400 ;
        RECT 878.100 916.050 879.900 917.850 ;
        RECT 890.100 916.050 891.900 917.850 ;
        RECT 896.700 916.050 897.900 923.400 ;
        RECT 914.100 916.050 915.900 917.850 ;
        RECT 917.100 916.050 918.300 929.400 ;
        RECT 748.800 913.950 750.900 916.050 ;
        RECT 763.950 913.950 766.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 769.950 913.950 772.050 916.050 ;
        RECT 772.950 913.950 775.050 916.050 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 793.950 913.950 796.050 916.050 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 826.950 913.950 829.050 916.050 ;
        RECT 829.950 913.950 832.050 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 844.950 913.950 847.050 916.050 ;
        RECT 847.950 913.950 850.050 916.050 ;
        RECT 850.950 913.950 853.050 916.050 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 868.950 913.950 871.050 916.050 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 892.950 913.950 895.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 913.950 913.950 916.050 916.050 ;
        RECT 916.950 913.950 919.050 916.050 ;
        RECT 721.500 908.400 729.900 909.300 ;
        RECT 746.700 908.700 748.800 909.600 ;
        RECT 721.500 907.500 723.300 908.400 ;
        RECT 719.700 904.800 722.400 906.600 ;
        RECT 720.600 900.600 722.400 904.800 ;
        RECT 723.600 900.000 725.400 906.600 ;
        RECT 728.100 900.600 729.900 908.400 ;
        RECT 743.400 907.800 748.800 908.700 ;
        RECT 743.400 903.600 744.300 907.800 ;
        RECT 750.000 906.600 750.900 913.950 ;
        RECT 764.100 912.150 765.900 913.950 ;
        RECT 767.100 909.600 768.300 913.950 ;
        RECT 770.100 912.150 771.900 913.950 ;
        RECT 764.700 908.700 768.300 909.600 ;
        RECT 786.000 910.200 786.900 913.950 ;
        RECT 788.100 912.150 789.900 913.950 ;
        RECT 794.100 912.150 795.900 913.950 ;
        RECT 786.000 909.000 789.300 910.200 ;
        RECT 764.700 906.600 765.900 908.700 ;
        RECT 740.100 900.600 741.900 903.600 ;
        RECT 743.100 900.600 744.900 903.600 ;
        RECT 740.100 900.000 741.300 900.600 ;
        RECT 746.100 900.000 747.900 906.000 ;
        RECT 749.100 900.600 750.900 906.600 ;
        RECT 764.100 900.600 765.900 906.600 ;
        RECT 767.100 905.700 774.900 907.050 ;
        RECT 767.100 900.600 768.900 905.700 ;
        RECT 770.100 900.000 771.900 904.800 ;
        RECT 773.100 900.600 774.900 905.700 ;
        RECT 787.500 900.600 789.300 909.000 ;
        RECT 794.100 900.000 795.900 909.600 ;
        RECT 809.700 903.600 810.900 913.950 ;
        RECT 824.100 912.150 825.900 913.950 ;
        RECT 830.100 912.150 831.900 913.950 ;
        RECT 833.100 910.200 834.000 913.950 ;
        RECT 845.100 912.150 846.900 913.950 ;
        RECT 851.250 912.150 853.050 913.950 ;
        RECT 809.100 900.600 810.900 903.600 ;
        RECT 812.100 900.000 813.900 903.600 ;
        RECT 824.100 900.000 825.900 909.600 ;
        RECT 830.700 909.000 834.000 910.200 ;
        RECT 835.950 909.450 838.050 910.050 ;
        RECT 847.950 909.450 850.050 910.050 ;
        RECT 830.700 900.600 832.500 909.000 ;
        RECT 835.950 908.550 850.050 909.450 ;
        RECT 835.950 907.950 838.050 908.550 ;
        RECT 847.950 907.950 850.050 908.550 ;
        RECT 854.700 906.600 855.600 913.950 ;
        RECT 869.100 912.150 870.900 913.950 ;
        RECT 872.100 909.600 873.300 913.950 ;
        RECT 875.100 912.150 876.900 913.950 ;
        RECT 893.100 912.150 894.900 913.950 ;
        RECT 869.700 908.700 873.300 909.600 ;
        RECT 896.700 909.600 897.900 913.950 ;
        RECT 899.100 912.150 900.900 913.950 ;
        RECT 896.700 908.700 900.300 909.600 ;
        RECT 869.700 906.600 870.900 908.700 ;
        RECT 846.000 900.000 847.800 906.600 ;
        RECT 850.500 905.400 855.600 906.600 ;
        RECT 850.500 900.600 852.300 905.400 ;
        RECT 853.500 900.000 855.300 903.600 ;
        RECT 869.100 900.600 870.900 906.600 ;
        RECT 872.100 905.700 879.900 907.050 ;
        RECT 872.100 900.600 873.900 905.700 ;
        RECT 875.100 900.000 876.900 904.800 ;
        RECT 878.100 900.600 879.900 905.700 ;
        RECT 890.100 905.700 897.900 907.050 ;
        RECT 890.100 900.600 891.900 905.700 ;
        RECT 893.100 900.000 894.900 904.800 ;
        RECT 896.100 900.600 897.900 905.700 ;
        RECT 899.100 906.600 900.300 908.700 ;
        RECT 899.100 900.600 900.900 906.600 ;
        RECT 917.100 903.600 918.300 913.950 ;
        RECT 914.100 900.000 915.900 903.600 ;
        RECT 917.100 900.600 918.900 903.600 ;
        RECT 11.700 889.200 13.500 896.400 ;
        RECT 16.800 890.400 18.600 897.000 ;
        RECT 11.700 888.300 15.900 889.200 ;
        RECT 11.100 883.050 12.900 884.850 ;
        RECT 14.700 883.050 15.900 888.300 ;
        RECT 34.500 888.000 36.300 896.400 ;
        RECT 33.000 886.800 36.300 888.000 ;
        RECT 41.100 887.400 42.900 897.000 ;
        RECT 53.700 889.200 55.500 896.400 ;
        RECT 58.800 890.400 60.600 897.000 ;
        RECT 53.700 888.300 57.900 889.200 ;
        RECT 16.950 883.050 18.750 884.850 ;
        RECT 33.000 883.050 33.900 886.800 ;
        RECT 35.100 883.050 36.900 884.850 ;
        RECT 41.100 883.050 42.900 884.850 ;
        RECT 53.100 883.050 54.900 884.850 ;
        RECT 56.700 883.050 57.900 888.300 ;
        RECT 76.500 888.000 78.300 896.400 ;
        RECT 75.000 886.800 78.300 888.000 ;
        RECT 83.100 887.400 84.900 897.000 ;
        RECT 95.100 893.400 96.900 896.400 ;
        RECT 98.100 893.400 99.900 897.000 ;
        RECT 110.100 893.400 111.900 897.000 ;
        RECT 113.100 893.400 114.900 896.400 ;
        RECT 116.100 893.400 117.900 897.000 ;
        RECT 58.950 883.050 60.750 884.850 ;
        RECT 75.000 883.050 75.900 886.800 ;
        RECT 77.100 883.050 78.900 884.850 ;
        RECT 83.100 883.050 84.900 884.850 ;
        RECT 95.700 883.050 96.900 893.400 ;
        RECT 113.700 883.050 114.600 893.400 ;
        RECT 132.000 890.400 133.800 897.000 ;
        RECT 136.500 891.600 138.300 896.400 ;
        RECT 139.500 893.400 141.300 897.000 ;
        RECT 136.500 890.400 141.600 891.600 ;
        RECT 124.950 888.450 127.050 889.050 ;
        RECT 136.950 888.450 139.050 889.050 ;
        RECT 124.950 887.550 139.050 888.450 ;
        RECT 124.950 886.950 127.050 887.550 ;
        RECT 136.950 886.950 139.050 887.550 ;
        RECT 118.950 885.450 123.000 886.050 ;
        RECT 118.950 883.950 123.450 885.450 ;
        RECT 10.950 880.950 13.050 883.050 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 52.950 880.950 55.050 883.050 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 73.950 880.950 76.050 883.050 ;
        RECT 76.950 880.950 79.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 94.950 880.950 97.050 883.050 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 112.950 880.950 115.050 883.050 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 14.700 867.600 15.900 880.950 ;
        RECT 33.000 868.800 33.900 880.950 ;
        RECT 38.100 879.150 39.900 880.950 ;
        RECT 33.000 867.900 39.600 868.800 ;
        RECT 33.000 867.600 33.900 867.900 ;
        RECT 11.100 861.000 12.900 867.600 ;
        RECT 14.100 861.600 15.900 867.600 ;
        RECT 17.100 861.000 18.900 867.600 ;
        RECT 32.100 861.600 33.900 867.600 ;
        RECT 38.100 867.600 39.600 867.900 ;
        RECT 56.700 867.600 57.900 880.950 ;
        RECT 75.000 868.800 75.900 880.950 ;
        RECT 80.100 879.150 81.900 880.950 ;
        RECT 76.950 876.450 79.050 877.050 ;
        RECT 91.950 876.450 94.050 877.050 ;
        RECT 76.950 875.550 94.050 876.450 ;
        RECT 76.950 874.950 79.050 875.550 ;
        RECT 91.950 874.950 94.050 875.550 ;
        RECT 75.000 867.900 81.600 868.800 ;
        RECT 75.000 867.600 75.900 867.900 ;
        RECT 35.100 861.000 36.900 867.000 ;
        RECT 38.100 861.600 39.900 867.600 ;
        RECT 41.100 861.000 42.900 867.600 ;
        RECT 53.100 861.000 54.900 867.600 ;
        RECT 56.100 861.600 57.900 867.600 ;
        RECT 59.100 861.000 60.900 867.600 ;
        RECT 74.100 861.600 75.900 867.600 ;
        RECT 80.100 867.600 81.600 867.900 ;
        RECT 95.700 867.600 96.900 880.950 ;
        RECT 98.100 879.150 99.900 880.950 ;
        RECT 110.100 879.150 111.900 880.950 ;
        RECT 113.700 873.600 114.600 880.950 ;
        RECT 115.950 879.150 117.750 880.950 ;
        RECT 122.550 880.050 123.450 883.950 ;
        RECT 131.100 883.050 132.900 884.850 ;
        RECT 137.250 883.050 139.050 884.850 ;
        RECT 140.700 883.050 141.600 890.400 ;
        RECT 152.100 890.400 153.900 896.400 ;
        RECT 155.100 891.300 156.900 897.000 ;
        RECT 159.600 890.400 161.400 896.400 ;
        RECT 164.100 891.300 165.900 897.000 ;
        RECT 167.100 890.400 168.900 896.400 ;
        RECT 182.700 893.400 184.500 897.000 ;
        RECT 185.700 891.600 187.500 896.400 ;
        RECT 182.400 890.400 187.500 891.600 ;
        RECT 190.200 890.400 192.000 897.000 ;
        RECT 206.700 893.400 208.500 897.000 ;
        RECT 209.700 891.600 211.500 896.400 ;
        RECT 206.400 890.400 211.500 891.600 ;
        RECT 214.200 890.400 216.000 897.000 ;
        RECT 227.100 890.400 228.900 896.400 ;
        RECT 152.100 889.500 156.900 890.400 ;
        RECT 154.800 888.300 156.900 889.500 ;
        RECT 159.900 888.900 161.100 890.400 ;
        RECT 158.100 886.800 161.100 888.900 ;
        RECT 167.100 888.600 168.300 890.400 ;
        RECT 156.900 883.800 159.000 885.900 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 152.100 880.950 154.200 883.050 ;
        RECT 156.900 882.000 158.700 883.800 ;
        RECT 159.900 881.100 161.100 886.800 ;
        RECT 162.000 887.700 168.300 888.600 ;
        RECT 162.000 885.600 164.100 887.700 ;
        RECT 162.000 883.800 163.800 885.600 ;
        RECT 166.800 883.050 168.600 884.850 ;
        RECT 182.400 883.050 183.300 890.400 ;
        RECT 184.950 883.050 186.750 884.850 ;
        RECT 191.100 883.050 192.900 884.850 ;
        RECT 206.400 883.050 207.300 890.400 ;
        RECT 227.700 888.300 228.900 890.400 ;
        RECT 230.100 891.300 231.900 896.400 ;
        RECT 233.100 892.200 234.900 897.000 ;
        RECT 236.100 891.300 237.900 896.400 ;
        RECT 230.100 889.950 237.900 891.300 ;
        RECT 248.100 890.400 249.900 896.400 ;
        RECT 251.100 890.400 252.900 897.000 ;
        RECT 254.100 893.400 255.900 896.400 ;
        RECT 227.700 887.400 231.300 888.300 ;
        RECT 208.950 883.050 210.750 884.850 ;
        RECT 215.100 883.050 216.900 884.850 ;
        RECT 227.100 883.050 228.900 884.850 ;
        RECT 230.100 883.050 231.300 887.400 ;
        RECT 233.100 883.050 234.900 884.850 ;
        RECT 248.100 883.050 249.300 890.400 ;
        RECT 254.700 889.500 255.900 893.400 ;
        RECT 250.200 888.600 255.900 889.500 ;
        RECT 266.100 893.400 267.900 896.400 ;
        RECT 266.100 889.500 267.300 893.400 ;
        RECT 269.100 890.400 270.900 897.000 ;
        RECT 272.100 890.400 273.900 896.400 ;
        RECT 289.500 890.400 291.300 897.000 ;
        RECT 294.000 890.400 295.800 896.400 ;
        RECT 298.500 890.400 300.300 897.000 ;
        RECT 314.100 891.300 315.900 896.400 ;
        RECT 317.100 892.200 318.900 897.000 ;
        RECT 320.100 891.300 321.900 896.400 ;
        RECT 266.100 888.600 271.800 889.500 ;
        RECT 250.200 887.700 252.000 888.600 ;
        RECT 166.800 882.300 168.900 883.050 ;
        RECT 118.950 878.550 123.450 880.050 ;
        RECT 134.250 879.150 136.050 880.950 ;
        RECT 118.950 877.950 123.000 878.550 ;
        RECT 140.700 873.600 141.600 880.950 ;
        RECT 152.400 879.150 154.200 880.950 ;
        RECT 158.700 880.200 161.100 881.100 ;
        RECT 162.000 880.950 168.900 882.300 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 187.950 880.950 190.050 883.050 ;
        RECT 190.950 880.950 193.050 883.050 ;
        RECT 205.950 880.950 208.050 883.050 ;
        RECT 208.950 880.950 211.050 883.050 ;
        RECT 211.950 880.950 214.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 226.950 880.950 229.050 883.050 ;
        RECT 229.950 880.950 232.050 883.050 ;
        RECT 232.950 880.950 235.050 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 248.100 880.950 250.200 883.050 ;
        RECT 162.000 880.500 163.800 880.950 ;
        RECT 158.700 880.050 160.200 880.200 ;
        RECT 158.100 877.950 160.200 880.050 ;
        RECT 159.300 876.000 160.200 877.950 ;
        RECT 161.100 877.500 165.000 879.300 ;
        RECT 161.100 877.200 163.200 877.500 ;
        RECT 159.300 874.950 160.800 876.000 ;
        RECT 154.800 873.600 156.900 874.500 ;
        RECT 111.000 872.400 114.600 873.600 ;
        RECT 77.100 861.000 78.900 867.000 ;
        RECT 80.100 861.600 81.900 867.600 ;
        RECT 83.100 861.000 84.900 867.600 ;
        RECT 95.100 861.600 96.900 867.600 ;
        RECT 98.100 861.000 99.900 867.600 ;
        RECT 111.000 861.600 112.800 872.400 ;
        RECT 116.100 861.000 117.900 873.600 ;
        RECT 131.100 872.700 138.900 873.600 ;
        RECT 131.100 861.600 132.900 872.700 ;
        RECT 134.100 861.000 135.900 871.800 ;
        RECT 137.100 861.600 138.900 872.700 ;
        RECT 140.100 861.600 141.900 873.600 ;
        RECT 152.100 872.400 156.900 873.600 ;
        RECT 159.600 873.600 160.800 874.950 ;
        RECT 164.400 873.600 166.500 875.700 ;
        RECT 182.400 873.600 183.300 880.950 ;
        RECT 187.950 879.150 189.750 880.950 ;
        RECT 206.400 873.600 207.300 880.950 ;
        RECT 211.950 879.150 213.750 880.950 ;
        RECT 230.100 873.600 231.300 880.950 ;
        RECT 236.100 879.150 237.900 880.950 ;
        RECT 248.100 873.600 249.300 880.950 ;
        RECT 251.100 876.300 252.000 887.700 ;
        RECT 270.000 887.700 271.800 888.600 ;
        RECT 253.500 880.950 255.600 883.050 ;
        RECT 253.800 879.150 255.600 880.950 ;
        RECT 266.400 880.950 268.500 883.050 ;
        RECT 266.400 879.150 268.200 880.950 ;
        RECT 250.200 875.400 252.000 876.300 ;
        RECT 270.000 876.300 270.900 887.700 ;
        RECT 272.700 883.050 273.900 890.400 ;
        RECT 287.100 883.050 288.900 884.850 ;
        RECT 293.700 883.050 294.900 890.400 ;
        RECT 314.100 889.950 321.900 891.300 ;
        RECT 323.100 890.400 324.900 896.400 ;
        RECT 335.100 890.400 336.900 896.400 ;
        RECT 295.950 888.450 298.050 889.050 ;
        RECT 301.950 888.450 304.050 889.050 ;
        RECT 295.950 887.550 304.050 888.450 ;
        RECT 323.100 888.300 324.300 890.400 ;
        RECT 295.950 886.950 298.050 887.550 ;
        RECT 301.950 886.950 304.050 887.550 ;
        RECT 320.700 887.400 324.300 888.300 ;
        RECT 335.700 888.300 336.900 890.400 ;
        RECT 338.100 891.300 339.900 896.400 ;
        RECT 341.100 892.200 342.900 897.000 ;
        RECT 344.100 891.300 345.900 896.400 ;
        RECT 356.100 893.400 357.900 897.000 ;
        RECT 359.100 893.400 360.900 896.400 ;
        RECT 338.100 889.950 345.900 891.300 ;
        RECT 346.950 891.450 349.050 892.050 ;
        RECT 355.950 891.450 358.050 892.050 ;
        RECT 346.950 890.550 358.050 891.450 ;
        RECT 346.950 889.950 349.050 890.550 ;
        RECT 355.950 889.950 358.050 890.550 ;
        RECT 335.700 887.400 339.300 888.300 ;
        RECT 298.950 883.050 300.750 884.850 ;
        RECT 317.100 883.050 318.900 884.850 ;
        RECT 320.700 883.050 321.900 887.400 ;
        RECT 323.100 883.050 324.900 884.850 ;
        RECT 335.100 883.050 336.900 884.850 ;
        RECT 338.100 883.050 339.300 887.400 ;
        RECT 341.100 883.050 342.900 884.850 ;
        RECT 359.100 883.050 360.300 893.400 ;
        RECT 374.100 890.400 375.900 896.400 ;
        RECT 374.700 888.300 375.900 890.400 ;
        RECT 377.100 891.300 378.900 896.400 ;
        RECT 380.100 892.200 381.900 897.000 ;
        RECT 383.100 891.300 384.900 896.400 ;
        RECT 377.100 889.950 384.900 891.300 ;
        RECT 398.100 890.400 399.900 896.400 ;
        RECT 401.100 890.400 402.900 897.000 ;
        RECT 404.100 893.400 405.900 896.400 ;
        RECT 374.700 887.400 378.300 888.300 ;
        RECT 374.100 883.050 375.900 884.850 ;
        RECT 377.100 883.050 378.300 887.400 ;
        RECT 380.100 883.050 381.900 884.850 ;
        RECT 398.100 883.050 399.300 890.400 ;
        RECT 404.700 889.500 405.900 893.400 ;
        RECT 416.100 891.300 417.900 896.400 ;
        RECT 419.100 892.200 420.900 897.000 ;
        RECT 422.100 891.300 423.900 896.400 ;
        RECT 416.100 889.950 423.900 891.300 ;
        RECT 425.100 890.400 426.900 896.400 ;
        RECT 440.700 895.200 441.900 897.000 ;
        RECT 400.200 888.600 405.900 889.500 ;
        RECT 400.200 887.700 402.000 888.600 ;
        RECT 425.100 888.300 426.300 890.400 ;
        RECT 440.100 889.200 441.900 895.200 ;
        RECT 444.600 890.700 446.400 895.200 ;
        RECT 449.700 894.600 450.900 897.000 ;
        RECT 444.300 889.800 446.400 890.700 ;
        RECT 449.100 889.800 450.900 894.600 ;
        RECT 452.100 892.200 453.900 895.200 ;
        RECT 467.100 893.400 468.900 896.400 ;
        RECT 470.100 893.400 471.900 897.000 ;
        RECT 271.800 880.950 273.900 883.050 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 382.950 880.950 385.050 883.050 ;
        RECT 398.100 880.950 400.200 883.050 ;
        RECT 270.000 875.400 271.800 876.300 ;
        RECT 250.200 874.500 255.900 875.400 ;
        RECT 152.100 861.600 153.900 872.400 ;
        RECT 155.100 861.000 156.900 871.500 ;
        RECT 159.600 861.600 161.400 873.600 ;
        RECT 164.400 872.700 168.900 873.600 ;
        RECT 164.100 861.000 165.900 871.500 ;
        RECT 167.100 861.600 168.900 872.700 ;
        RECT 182.100 861.600 183.900 873.600 ;
        RECT 185.100 872.700 192.900 873.600 ;
        RECT 185.100 861.600 186.900 872.700 ;
        RECT 188.100 861.000 189.900 871.800 ;
        RECT 191.100 861.600 192.900 872.700 ;
        RECT 206.100 861.600 207.900 873.600 ;
        RECT 209.100 872.700 216.900 873.600 ;
        RECT 209.100 861.600 210.900 872.700 ;
        RECT 212.100 861.000 213.900 871.800 ;
        RECT 215.100 861.600 216.900 872.700 ;
        RECT 230.100 872.100 232.500 873.600 ;
        RECT 228.000 869.100 229.800 870.900 ;
        RECT 227.700 861.000 229.500 867.600 ;
        RECT 230.700 861.600 232.500 872.100 ;
        RECT 235.800 861.000 237.600 873.600 ;
        RECT 248.100 861.600 249.900 873.600 ;
        RECT 251.100 861.000 252.900 871.800 ;
        RECT 254.700 867.600 255.900 874.500 ;
        RECT 254.100 861.600 255.900 867.600 ;
        RECT 266.100 874.500 271.800 875.400 ;
        RECT 266.100 867.600 267.300 874.500 ;
        RECT 272.700 873.600 273.900 880.950 ;
        RECT 290.100 879.150 291.900 880.950 ;
        RECT 294.000 875.400 294.900 880.950 ;
        RECT 295.950 879.150 297.750 880.950 ;
        RECT 314.100 879.150 315.900 880.950 ;
        RECT 290.100 874.500 294.900 875.400 ;
        RECT 266.100 861.600 267.900 867.600 ;
        RECT 269.100 861.000 270.900 871.800 ;
        RECT 272.100 861.600 273.900 873.600 ;
        RECT 287.100 862.500 288.900 873.600 ;
        RECT 290.100 863.400 291.900 874.500 ;
        RECT 320.700 873.600 321.900 880.950 ;
        RECT 322.950 876.450 325.050 877.050 ;
        RECT 328.950 876.450 331.050 877.050 ;
        RECT 322.950 875.550 331.050 876.450 ;
        RECT 322.950 874.950 325.050 875.550 ;
        RECT 328.950 874.950 331.050 875.550 ;
        RECT 293.100 872.400 300.900 873.300 ;
        RECT 293.100 862.500 294.900 872.400 ;
        RECT 287.100 861.600 294.900 862.500 ;
        RECT 296.100 861.000 297.900 871.500 ;
        RECT 299.100 861.600 300.900 872.400 ;
        RECT 314.400 861.000 316.200 873.600 ;
        RECT 319.500 872.100 321.900 873.600 ;
        RECT 338.100 873.600 339.300 880.950 ;
        RECT 344.100 879.150 345.900 880.950 ;
        RECT 356.100 879.150 357.900 880.950 ;
        RECT 338.100 872.100 340.500 873.600 ;
        RECT 319.500 861.600 321.300 872.100 ;
        RECT 322.200 869.100 324.000 870.900 ;
        RECT 336.000 869.100 337.800 870.900 ;
        RECT 322.500 861.000 324.300 867.600 ;
        RECT 335.700 861.000 337.500 867.600 ;
        RECT 338.700 861.600 340.500 872.100 ;
        RECT 343.800 861.000 345.600 873.600 ;
        RECT 359.100 867.600 360.300 880.950 ;
        RECT 377.100 873.600 378.300 880.950 ;
        RECT 383.100 879.150 384.900 880.950 ;
        RECT 398.100 873.600 399.300 880.950 ;
        RECT 401.100 876.300 402.000 887.700 ;
        RECT 422.700 887.400 426.300 888.300 ;
        RECT 419.100 883.050 420.900 884.850 ;
        RECT 422.700 883.050 423.900 887.400 ;
        RECT 425.100 883.050 426.900 884.850 ;
        RECT 444.300 883.050 445.200 889.800 ;
        RECT 453.000 888.900 453.900 892.200 ;
        RECT 403.500 880.950 405.600 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 421.950 880.950 424.050 883.050 ;
        RECT 424.950 880.950 427.050 883.050 ;
        RECT 440.100 880.950 442.200 883.050 ;
        RECT 443.100 880.950 445.200 883.050 ;
        RECT 446.700 888.000 453.900 888.900 ;
        RECT 446.700 880.950 447.900 888.000 ;
        RECT 452.100 883.050 453.900 884.850 ;
        RECT 467.700 883.050 468.900 893.400 ;
        RECT 482.100 890.400 483.900 896.400 ;
        RECT 485.100 891.300 486.900 897.000 ;
        RECT 489.600 890.400 491.400 896.400 ;
        RECT 494.100 891.300 495.900 897.000 ;
        RECT 497.100 890.400 498.900 896.400 ;
        RECT 509.700 893.400 511.500 897.000 ;
        RECT 512.700 891.600 514.500 896.400 ;
        RECT 509.400 890.400 514.500 891.600 ;
        RECT 517.200 890.400 519.000 897.000 ;
        RECT 533.100 890.400 534.900 896.400 ;
        RECT 482.100 889.500 486.900 890.400 ;
        RECT 484.800 888.300 486.900 889.500 ;
        RECT 489.900 888.900 491.100 890.400 ;
        RECT 488.100 886.800 491.100 888.900 ;
        RECT 497.100 888.600 498.300 890.400 ;
        RECT 486.900 883.800 489.000 885.900 ;
        RECT 448.800 880.950 450.900 883.050 ;
        RECT 451.800 880.950 453.900 883.050 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 482.100 880.950 484.200 883.050 ;
        RECT 486.900 882.000 488.700 883.800 ;
        RECT 489.900 881.100 491.100 886.800 ;
        RECT 492.000 887.700 498.300 888.600 ;
        RECT 492.000 885.600 494.100 887.700 ;
        RECT 492.000 883.800 493.800 885.600 ;
        RECT 496.800 883.050 498.600 884.850 ;
        RECT 509.400 883.050 510.300 890.400 ;
        RECT 533.700 888.300 534.900 890.400 ;
        RECT 536.100 891.300 537.900 896.400 ;
        RECT 539.100 892.200 540.900 897.000 ;
        RECT 542.100 891.300 543.900 896.400 ;
        RECT 536.100 889.950 543.900 891.300 ;
        RECT 557.400 890.400 559.200 897.000 ;
        RECT 562.500 889.200 564.300 896.400 ;
        RECT 578.100 891.300 579.900 896.400 ;
        RECT 581.100 892.200 582.900 897.000 ;
        RECT 584.100 891.300 585.900 896.400 ;
        RECT 578.100 889.950 585.900 891.300 ;
        RECT 587.100 890.400 588.900 896.400 ;
        RECT 560.100 888.300 564.300 889.200 ;
        RECT 587.100 888.300 588.300 890.400 ;
        RECT 533.700 887.400 537.300 888.300 ;
        RECT 529.950 885.450 532.050 886.050 ;
        RECT 511.950 883.050 513.750 884.850 ;
        RECT 518.100 883.050 519.900 884.850 ;
        RECT 524.550 884.550 532.050 885.450 ;
        RECT 496.800 882.300 498.900 883.050 ;
        RECT 403.800 879.150 405.600 880.950 ;
        RECT 416.100 879.150 417.900 880.950 ;
        RECT 400.200 875.400 402.000 876.300 ;
        RECT 400.200 874.500 405.900 875.400 ;
        RECT 377.100 872.100 379.500 873.600 ;
        RECT 375.000 869.100 376.800 870.900 ;
        RECT 356.100 861.000 357.900 867.600 ;
        RECT 359.100 861.600 360.900 867.600 ;
        RECT 374.700 861.000 376.500 867.600 ;
        RECT 377.700 861.600 379.500 872.100 ;
        RECT 382.800 861.000 384.600 873.600 ;
        RECT 398.100 861.600 399.900 873.600 ;
        RECT 401.100 861.000 402.900 871.800 ;
        RECT 404.700 867.600 405.900 874.500 ;
        RECT 422.700 873.600 423.900 880.950 ;
        RECT 440.400 879.150 442.200 880.950 ;
        RECT 404.100 861.600 405.900 867.600 ;
        RECT 416.400 861.000 418.200 873.600 ;
        RECT 421.500 872.100 423.900 873.600 ;
        RECT 421.500 861.600 423.300 872.100 ;
        RECT 424.200 869.100 426.000 870.900 ;
        RECT 424.500 861.000 426.300 867.600 ;
        RECT 440.100 861.000 441.900 873.600 ;
        RECT 444.300 873.000 445.200 880.950 ;
        RECT 446.100 879.150 447.900 880.950 ;
        RECT 449.100 879.150 450.900 880.950 ;
        RECT 446.100 874.800 447.300 879.150 ;
        RECT 446.100 873.900 453.900 874.800 ;
        RECT 444.300 872.100 446.400 873.000 ;
        RECT 444.600 861.600 446.400 872.100 ;
        RECT 449.100 861.000 450.900 873.000 ;
        RECT 453.000 868.800 453.900 873.900 ;
        RECT 452.100 862.800 453.900 868.800 ;
        RECT 467.700 867.600 468.900 880.950 ;
        RECT 470.100 879.150 471.900 880.950 ;
        RECT 482.400 879.150 484.200 880.950 ;
        RECT 488.700 880.200 491.100 881.100 ;
        RECT 492.000 880.950 498.900 882.300 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 511.950 880.950 514.050 883.050 ;
        RECT 514.950 880.950 517.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 492.000 880.500 493.800 880.950 ;
        RECT 488.700 880.050 490.200 880.200 ;
        RECT 488.100 877.950 490.200 880.050 ;
        RECT 489.300 876.000 490.200 877.950 ;
        RECT 491.100 877.500 495.000 879.300 ;
        RECT 491.100 877.200 493.200 877.500 ;
        RECT 489.300 874.950 490.800 876.000 ;
        RECT 484.800 873.600 486.900 874.500 ;
        RECT 482.100 872.400 486.900 873.600 ;
        RECT 489.600 873.600 490.800 874.950 ;
        RECT 494.400 873.600 496.500 875.700 ;
        RECT 509.400 873.600 510.300 880.950 ;
        RECT 514.950 879.150 516.750 880.950 ;
        RECT 524.550 879.450 525.450 884.550 ;
        RECT 529.950 883.950 532.050 884.550 ;
        RECT 533.100 883.050 534.900 884.850 ;
        RECT 536.100 883.050 537.300 887.400 ;
        RECT 539.100 883.050 540.900 884.850 ;
        RECT 557.250 883.050 559.050 884.850 ;
        RECT 560.100 883.050 561.300 888.300 ;
        RECT 584.700 887.400 588.300 888.300 ;
        RECT 602.100 887.400 603.900 897.000 ;
        RECT 608.700 888.000 610.500 896.400 ;
        RECT 623.100 891.300 624.900 896.400 ;
        RECT 626.100 892.200 627.900 897.000 ;
        RECT 629.100 891.300 630.900 896.400 ;
        RECT 623.100 889.950 630.900 891.300 ;
        RECT 632.100 890.400 633.900 896.400 ;
        RECT 647.100 890.400 648.900 897.000 ;
        RECT 650.100 890.400 651.900 896.400 ;
        RECT 665.100 893.400 666.900 896.400 ;
        RECT 668.100 893.400 669.900 897.000 ;
        RECT 632.100 888.300 633.300 890.400 ;
        RECT 563.100 883.050 564.900 884.850 ;
        RECT 581.100 883.050 582.900 884.850 ;
        RECT 584.700 883.050 585.900 887.400 ;
        RECT 608.700 886.800 612.000 888.000 ;
        RECT 587.100 883.050 588.900 884.850 ;
        RECT 602.100 883.050 603.900 884.850 ;
        RECT 608.100 883.050 609.900 884.850 ;
        RECT 611.100 883.050 612.000 886.800 ;
        RECT 629.700 887.400 633.300 888.300 ;
        RECT 626.100 883.050 627.900 884.850 ;
        RECT 629.700 883.050 630.900 887.400 ;
        RECT 632.100 883.050 633.900 884.850 ;
        RECT 647.100 883.050 648.900 884.850 ;
        RECT 650.100 883.050 651.300 890.400 ;
        RECT 665.700 883.050 666.900 893.400 ;
        RECT 683.100 890.400 684.900 896.400 ;
        RECT 686.100 890.400 687.900 897.000 ;
        RECT 689.100 893.400 690.900 896.400 ;
        RECT 683.100 883.050 684.300 890.400 ;
        RECT 689.700 889.500 690.900 893.400 ;
        RECT 704.400 890.400 706.200 897.000 ;
        RECT 685.200 888.600 690.900 889.500 ;
        RECT 709.500 889.200 711.300 896.400 ;
        RECT 722.100 891.300 723.900 896.400 ;
        RECT 725.100 892.200 726.900 897.000 ;
        RECT 728.100 891.300 729.900 896.400 ;
        RECT 722.100 889.950 729.900 891.300 ;
        RECT 731.100 890.400 732.900 896.400 ;
        RECT 743.100 893.400 744.900 897.000 ;
        RECT 746.100 893.400 747.900 896.400 ;
        RECT 749.100 893.400 750.900 897.000 ;
        RECT 685.200 887.700 687.000 888.600 ;
        RECT 532.950 880.950 535.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 559.950 880.950 562.050 883.050 ;
        RECT 562.950 880.950 565.050 883.050 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 583.950 880.950 586.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 604.950 880.950 607.050 883.050 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 646.950 880.950 649.050 883.050 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 683.100 880.950 685.200 883.050 ;
        RECT 521.550 878.550 525.450 879.450 ;
        RECT 511.950 876.450 514.050 877.050 ;
        RECT 521.550 876.450 522.450 878.550 ;
        RECT 511.950 875.550 522.450 876.450 ;
        RECT 511.950 874.950 514.050 875.550 ;
        RECT 536.100 873.600 537.300 880.950 ;
        RECT 542.100 879.150 543.900 880.950 ;
        RECT 467.100 861.600 468.900 867.600 ;
        RECT 470.100 861.000 471.900 867.600 ;
        RECT 482.100 861.600 483.900 872.400 ;
        RECT 485.100 861.000 486.900 871.500 ;
        RECT 489.600 861.600 491.400 873.600 ;
        RECT 494.400 872.700 498.900 873.600 ;
        RECT 494.100 861.000 495.900 871.500 ;
        RECT 497.100 861.600 498.900 872.700 ;
        RECT 509.100 861.600 510.900 873.600 ;
        RECT 512.100 872.700 519.900 873.600 ;
        RECT 512.100 861.600 513.900 872.700 ;
        RECT 515.100 861.000 516.900 871.800 ;
        RECT 518.100 861.600 519.900 872.700 ;
        RECT 536.100 872.100 538.500 873.600 ;
        RECT 534.000 869.100 535.800 870.900 ;
        RECT 533.700 861.000 535.500 867.600 ;
        RECT 536.700 861.600 538.500 872.100 ;
        RECT 541.800 861.000 543.600 873.600 ;
        RECT 560.100 867.600 561.300 880.950 ;
        RECT 578.100 879.150 579.900 880.950 ;
        RECT 584.700 873.600 585.900 880.950 ;
        RECT 605.100 879.150 606.900 880.950 ;
        RECT 557.100 861.000 558.900 867.600 ;
        RECT 560.100 861.600 561.900 867.600 ;
        RECT 563.100 861.000 564.900 867.600 ;
        RECT 578.400 861.000 580.200 873.600 ;
        RECT 583.500 872.100 585.900 873.600 ;
        RECT 583.500 861.600 585.300 872.100 ;
        RECT 586.200 869.100 588.000 870.900 ;
        RECT 611.100 868.800 612.000 880.950 ;
        RECT 623.100 879.150 624.900 880.950 ;
        RECT 629.700 873.600 630.900 880.950 ;
        RECT 650.100 873.600 651.300 880.950 ;
        RECT 605.400 867.900 612.000 868.800 ;
        RECT 605.400 867.600 606.900 867.900 ;
        RECT 586.500 861.000 588.300 867.600 ;
        RECT 602.100 861.000 603.900 867.600 ;
        RECT 605.100 861.600 606.900 867.600 ;
        RECT 611.100 867.600 612.000 867.900 ;
        RECT 608.100 861.000 609.900 867.000 ;
        RECT 611.100 861.600 612.900 867.600 ;
        RECT 623.400 861.000 625.200 873.600 ;
        RECT 628.500 872.100 630.900 873.600 ;
        RECT 628.500 861.600 630.300 872.100 ;
        RECT 631.200 869.100 633.000 870.900 ;
        RECT 631.500 861.000 633.300 867.600 ;
        RECT 647.100 861.000 648.900 873.600 ;
        RECT 650.100 861.600 651.900 873.600 ;
        RECT 665.700 867.600 666.900 880.950 ;
        RECT 668.100 879.150 669.900 880.950 ;
        RECT 683.100 873.600 684.300 880.950 ;
        RECT 686.100 876.300 687.000 887.700 ;
        RECT 707.100 888.300 711.300 889.200 ;
        RECT 731.100 888.300 732.300 890.400 ;
        RECT 704.250 883.050 706.050 884.850 ;
        RECT 707.100 883.050 708.300 888.300 ;
        RECT 728.700 887.400 732.300 888.300 ;
        RECT 710.100 883.050 711.900 884.850 ;
        RECT 725.100 883.050 726.900 884.850 ;
        RECT 728.700 883.050 729.900 887.400 ;
        RECT 731.100 883.050 732.900 884.850 ;
        RECT 746.700 883.050 747.600 893.400 ;
        RECT 761.100 891.300 762.900 896.400 ;
        RECT 764.100 892.200 765.900 897.000 ;
        RECT 767.100 891.300 768.900 896.400 ;
        RECT 761.100 889.950 768.900 891.300 ;
        RECT 770.100 890.400 771.900 896.400 ;
        RECT 770.100 888.300 771.300 890.400 ;
        RECT 785.700 889.200 787.500 896.400 ;
        RECT 790.800 890.400 792.600 897.000 ;
        RECT 807.000 890.400 808.800 897.000 ;
        RECT 811.500 891.600 813.300 896.400 ;
        RECT 814.500 893.400 816.300 897.000 ;
        RECT 827.700 893.400 829.500 897.000 ;
        RECT 830.700 891.600 832.500 896.400 ;
        RECT 811.500 890.400 816.600 891.600 ;
        RECT 785.700 888.300 789.900 889.200 ;
        RECT 767.700 887.400 771.300 888.300 ;
        RECT 751.950 885.450 756.000 886.050 ;
        RECT 751.950 883.950 756.450 885.450 ;
        RECT 688.500 880.950 690.600 883.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 742.950 880.950 745.050 883.050 ;
        RECT 745.950 880.950 748.050 883.050 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 688.800 879.150 690.600 880.950 ;
        RECT 685.200 875.400 687.000 876.300 ;
        RECT 694.950 876.450 697.050 877.050 ;
        RECT 703.950 876.450 706.050 877.050 ;
        RECT 694.950 875.550 706.050 876.450 ;
        RECT 685.200 874.500 690.900 875.400 ;
        RECT 694.950 874.950 697.050 875.550 ;
        RECT 703.950 874.950 706.050 875.550 ;
        RECT 665.100 861.600 666.900 867.600 ;
        RECT 668.100 861.000 669.900 867.600 ;
        RECT 683.100 861.600 684.900 873.600 ;
        RECT 686.100 861.000 687.900 871.800 ;
        RECT 689.700 867.600 690.900 874.500 ;
        RECT 707.100 867.600 708.300 880.950 ;
        RECT 722.100 879.150 723.900 880.950 ;
        RECT 728.700 873.600 729.900 880.950 ;
        RECT 743.100 879.150 744.900 880.950 ;
        RECT 746.700 873.600 747.600 880.950 ;
        RECT 748.950 879.150 750.750 880.950 ;
        RECT 755.550 876.450 756.450 883.950 ;
        RECT 764.100 883.050 765.900 884.850 ;
        RECT 767.700 883.050 768.900 887.400 ;
        RECT 772.950 885.450 777.000 886.050 ;
        RECT 770.100 883.050 771.900 884.850 ;
        RECT 772.950 883.950 777.450 885.450 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 763.950 880.950 766.050 883.050 ;
        RECT 766.950 880.950 769.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 761.100 879.150 762.900 880.950 ;
        RECT 763.950 876.450 766.050 877.050 ;
        RECT 755.550 875.550 766.050 876.450 ;
        RECT 763.950 874.950 766.050 875.550 ;
        RECT 767.700 873.600 768.900 880.950 ;
        RECT 776.550 876.900 777.450 883.950 ;
        RECT 785.100 883.050 786.900 884.850 ;
        RECT 788.700 883.050 789.900 888.300 ;
        RECT 790.950 883.050 792.750 884.850 ;
        RECT 806.100 883.050 807.900 884.850 ;
        RECT 812.250 883.050 814.050 884.850 ;
        RECT 815.700 883.050 816.600 890.400 ;
        RECT 827.400 890.400 832.500 891.600 ;
        RECT 835.200 890.400 837.000 897.000 ;
        RECT 827.400 883.050 828.300 890.400 ;
        RECT 848.100 887.400 849.900 897.000 ;
        RECT 854.700 888.000 856.500 896.400 ;
        RECT 874.500 888.000 876.300 896.400 ;
        RECT 854.700 886.800 858.000 888.000 ;
        RECT 829.950 883.050 831.750 884.850 ;
        RECT 836.100 883.050 837.900 884.850 ;
        RECT 848.100 883.050 849.900 884.850 ;
        RECT 854.100 883.050 855.900 884.850 ;
        RECT 857.100 883.050 858.000 886.800 ;
        RECT 873.000 886.800 876.300 888.000 ;
        RECT 881.100 887.400 882.900 897.000 ;
        RECT 895.500 888.000 897.300 896.400 ;
        RECT 894.000 886.800 897.300 888.000 ;
        RECT 902.100 887.400 903.900 897.000 ;
        RECT 915.000 890.400 916.800 897.000 ;
        RECT 919.500 891.600 921.300 896.400 ;
        RECT 922.500 893.400 924.300 897.000 ;
        RECT 919.500 890.400 924.600 891.600 ;
        RECT 873.000 883.050 873.900 886.800 ;
        RECT 888.000 885.450 892.050 886.050 ;
        RECT 875.100 883.050 876.900 884.850 ;
        RECT 881.100 883.050 882.900 884.850 ;
        RECT 887.550 883.950 892.050 885.450 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 826.950 880.950 829.050 883.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 847.950 880.950 850.050 883.050 ;
        RECT 850.950 880.950 853.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 871.950 880.950 874.050 883.050 ;
        RECT 874.950 880.950 877.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 775.950 874.800 778.050 876.900 ;
        RECT 689.100 861.600 690.900 867.600 ;
        RECT 704.100 861.000 705.900 867.600 ;
        RECT 707.100 861.600 708.900 867.600 ;
        RECT 710.100 861.000 711.900 867.600 ;
        RECT 722.400 861.000 724.200 873.600 ;
        RECT 727.500 872.100 729.900 873.600 ;
        RECT 744.000 872.400 747.600 873.600 ;
        RECT 727.500 861.600 729.300 872.100 ;
        RECT 730.200 869.100 732.000 870.900 ;
        RECT 730.500 861.000 732.300 867.600 ;
        RECT 744.000 861.600 745.800 872.400 ;
        RECT 749.100 861.000 750.900 873.600 ;
        RECT 761.400 861.000 763.200 873.600 ;
        RECT 766.500 872.100 768.900 873.600 ;
        RECT 766.500 861.600 768.300 872.100 ;
        RECT 769.200 869.100 771.000 870.900 ;
        RECT 788.700 867.600 789.900 880.950 ;
        RECT 809.250 879.150 811.050 880.950 ;
        RECT 815.700 873.600 816.600 880.950 ;
        RECT 827.400 873.600 828.300 880.950 ;
        RECT 832.950 879.150 834.750 880.950 ;
        RECT 851.100 879.150 852.900 880.950 ;
        RECT 806.100 872.700 813.900 873.600 ;
        RECT 769.500 861.000 771.300 867.600 ;
        RECT 785.100 861.000 786.900 867.600 ;
        RECT 788.100 861.600 789.900 867.600 ;
        RECT 791.100 861.000 792.900 867.600 ;
        RECT 806.100 861.600 807.900 872.700 ;
        RECT 809.100 861.000 810.900 871.800 ;
        RECT 812.100 861.600 813.900 872.700 ;
        RECT 815.100 861.600 816.900 873.600 ;
        RECT 827.100 861.600 828.900 873.600 ;
        RECT 830.100 872.700 837.900 873.600 ;
        RECT 830.100 861.600 831.900 872.700 ;
        RECT 833.100 861.000 834.900 871.800 ;
        RECT 836.100 861.600 837.900 872.700 ;
        RECT 857.100 868.800 858.000 880.950 ;
        RECT 851.400 867.900 858.000 868.800 ;
        RECT 851.400 867.600 852.900 867.900 ;
        RECT 848.100 861.000 849.900 867.600 ;
        RECT 851.100 861.600 852.900 867.600 ;
        RECT 857.100 867.600 858.000 867.900 ;
        RECT 873.000 868.800 873.900 880.950 ;
        RECT 878.100 879.150 879.900 880.950 ;
        RECT 887.550 880.050 888.450 883.950 ;
        RECT 894.000 883.050 894.900 886.800 ;
        RECT 904.950 885.450 909.000 886.050 ;
        RECT 896.100 883.050 897.900 884.850 ;
        RECT 902.100 883.050 903.900 884.850 ;
        RECT 904.950 883.950 909.450 885.450 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 901.950 880.950 904.050 883.050 ;
        RECT 887.550 878.550 892.050 880.050 ;
        RECT 888.000 877.950 892.050 878.550 ;
        RECT 894.000 868.800 894.900 880.950 ;
        RECT 899.100 879.150 900.900 880.950 ;
        RECT 908.550 879.450 909.450 883.950 ;
        RECT 914.100 883.050 915.900 884.850 ;
        RECT 920.250 883.050 922.050 884.850 ;
        RECT 923.700 883.050 924.600 890.400 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 919.950 880.950 922.050 883.050 ;
        RECT 922.950 880.950 925.050 883.050 ;
        RECT 908.550 878.550 912.450 879.450 ;
        RECT 917.250 879.150 919.050 880.950 ;
        RECT 901.950 876.450 904.050 876.750 ;
        RECT 911.550 876.450 912.450 878.550 ;
        RECT 919.950 876.450 922.050 877.050 ;
        RECT 901.950 875.550 922.050 876.450 ;
        RECT 901.950 874.650 904.050 875.550 ;
        RECT 919.950 874.950 922.050 875.550 ;
        RECT 923.700 873.600 924.600 880.950 ;
        RECT 914.100 872.700 921.900 873.600 ;
        RECT 873.000 867.900 879.600 868.800 ;
        RECT 873.000 867.600 873.900 867.900 ;
        RECT 854.100 861.000 855.900 867.000 ;
        RECT 857.100 861.600 858.900 867.600 ;
        RECT 872.100 861.600 873.900 867.600 ;
        RECT 878.100 867.600 879.600 867.900 ;
        RECT 894.000 867.900 900.600 868.800 ;
        RECT 894.000 867.600 894.900 867.900 ;
        RECT 875.100 861.000 876.900 867.000 ;
        RECT 878.100 861.600 879.900 867.600 ;
        RECT 881.100 861.000 882.900 867.600 ;
        RECT 893.100 861.600 894.900 867.600 ;
        RECT 899.100 867.600 900.600 867.900 ;
        RECT 896.100 861.000 897.900 867.000 ;
        RECT 899.100 861.600 900.900 867.600 ;
        RECT 902.100 861.000 903.900 867.600 ;
        RECT 914.100 861.600 915.900 872.700 ;
        RECT 917.100 861.000 918.900 871.800 ;
        RECT 920.100 861.600 921.900 872.700 ;
        RECT 923.100 861.600 924.900 873.600 ;
        RECT 11.100 851.400 12.900 858.000 ;
        RECT 14.100 851.400 15.900 857.400 ;
        RECT 17.100 852.000 18.900 858.000 ;
        RECT 14.400 851.100 15.900 851.400 ;
        RECT 20.100 851.400 21.900 857.400 ;
        RECT 35.100 851.400 36.900 858.000 ;
        RECT 38.100 851.400 39.900 857.400 ;
        RECT 41.100 851.400 42.900 858.000 ;
        RECT 56.100 851.400 57.900 857.400 ;
        RECT 59.100 852.000 60.900 858.000 ;
        RECT 20.100 851.100 21.000 851.400 ;
        RECT 14.400 850.200 21.000 851.100 ;
        RECT 10.950 843.450 13.050 844.050 ;
        RECT 16.950 843.450 19.050 844.200 ;
        RECT 10.950 842.550 19.050 843.450 ;
        RECT 10.950 841.950 13.050 842.550 ;
        RECT 16.950 842.100 19.050 842.550 ;
        RECT 14.100 838.050 15.900 839.850 ;
        RECT 20.100 838.050 21.000 850.200 ;
        RECT 25.950 843.450 28.050 844.050 ;
        RECT 34.950 843.450 37.050 844.050 ;
        RECT 25.950 842.550 37.050 843.450 ;
        RECT 25.950 841.950 28.050 842.550 ;
        RECT 34.950 841.950 37.050 842.550 ;
        RECT 38.700 838.050 39.900 851.400 ;
        RECT 57.000 851.100 57.900 851.400 ;
        RECT 62.100 851.400 63.900 857.400 ;
        RECT 65.100 851.400 66.900 858.000 ;
        RECT 77.100 851.400 78.900 857.400 ;
        RECT 80.100 852.000 81.900 858.000 ;
        RECT 62.100 851.100 63.600 851.400 ;
        RECT 57.000 850.200 63.600 851.100 ;
        RECT 78.000 851.100 78.900 851.400 ;
        RECT 83.100 851.400 84.900 857.400 ;
        RECT 86.100 851.400 87.900 858.000 ;
        RECT 101.100 851.400 102.900 858.000 ;
        RECT 104.100 851.400 105.900 857.400 ;
        RECT 107.100 851.400 108.900 858.000 ;
        RECT 122.100 851.400 123.900 858.000 ;
        RECT 125.100 851.400 126.900 857.400 ;
        RECT 137.700 851.400 139.500 858.000 ;
        RECT 83.100 851.100 84.600 851.400 ;
        RECT 78.000 850.200 84.600 851.100 ;
        RECT 57.000 838.050 57.900 850.200 ;
        RECT 67.950 840.450 72.000 841.050 ;
        RECT 62.100 838.050 63.900 839.850 ;
        RECT 67.950 838.950 72.450 840.450 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 11.100 834.150 12.900 835.950 ;
        RECT 17.100 834.150 18.900 835.950 ;
        RECT 20.100 832.200 21.000 835.950 ;
        RECT 35.100 834.150 36.900 835.950 ;
        RECT 11.100 822.000 12.900 831.600 ;
        RECT 17.700 831.000 21.000 832.200 ;
        RECT 17.700 822.600 19.500 831.000 ;
        RECT 38.700 830.700 39.900 835.950 ;
        RECT 40.950 834.150 42.750 835.950 ;
        RECT 57.000 832.200 57.900 835.950 ;
        RECT 59.100 834.150 60.900 835.950 ;
        RECT 65.100 834.150 66.900 835.950 ;
        RECT 57.000 831.000 60.300 832.200 ;
        RECT 71.550 832.050 72.450 838.950 ;
        RECT 78.000 838.050 78.900 850.200 ;
        RECT 83.100 838.050 84.900 839.850 ;
        RECT 104.100 838.050 105.300 851.400 ;
        RECT 122.100 838.050 123.900 839.850 ;
        RECT 125.100 838.050 126.300 851.400 ;
        RECT 138.000 848.100 139.800 849.900 ;
        RECT 140.700 846.900 142.500 857.400 ;
        RECT 140.100 845.400 142.500 846.900 ;
        RECT 145.800 845.400 147.600 858.000 ;
        RECT 158.100 846.300 159.900 857.400 ;
        RECT 161.100 847.500 162.900 858.000 ;
        RECT 158.100 845.400 162.600 846.300 ;
        RECT 165.600 845.400 167.400 857.400 ;
        RECT 170.100 847.500 171.900 858.000 ;
        RECT 173.100 846.600 174.900 857.400 ;
        RECT 185.100 851.400 186.900 858.000 ;
        RECT 188.100 851.400 189.900 857.400 ;
        RECT 191.100 851.400 192.900 858.000 ;
        RECT 132.000 840.450 136.050 841.050 ;
        RECT 131.550 838.950 136.050 840.450 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 79.950 835.950 82.050 838.050 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 78.000 832.200 78.900 835.950 ;
        RECT 80.100 834.150 81.900 835.950 ;
        RECT 86.100 834.150 87.900 835.950 ;
        RECT 101.250 834.150 103.050 835.950 ;
        RECT 35.700 829.800 39.900 830.700 ;
        RECT 35.700 822.600 37.500 829.800 ;
        RECT 40.800 822.000 42.600 828.600 ;
        RECT 58.500 822.600 60.300 831.000 ;
        RECT 65.100 822.000 66.900 831.600 ;
        RECT 70.950 829.950 73.050 832.050 ;
        RECT 78.000 831.000 81.300 832.200 ;
        RECT 79.500 822.600 81.300 831.000 ;
        RECT 86.100 822.000 87.900 831.600 ;
        RECT 91.950 831.450 94.050 832.050 ;
        RECT 100.950 831.450 103.050 832.050 ;
        RECT 91.950 830.550 103.050 831.450 ;
        RECT 91.950 829.950 94.050 830.550 ;
        RECT 100.950 829.950 103.050 830.550 ;
        RECT 104.100 830.700 105.300 835.950 ;
        RECT 107.100 834.150 108.900 835.950 ;
        RECT 104.100 829.800 108.300 830.700 ;
        RECT 101.400 822.000 103.200 828.600 ;
        RECT 106.500 822.600 108.300 829.800 ;
        RECT 125.100 825.600 126.300 835.950 ;
        RECT 131.550 835.050 132.450 838.950 ;
        RECT 140.100 838.050 141.300 845.400 ;
        RECT 160.500 843.300 162.600 845.400 ;
        RECT 166.200 844.050 167.400 845.400 ;
        RECT 170.100 845.400 174.900 846.600 ;
        RECT 170.100 844.500 172.200 845.400 ;
        RECT 166.200 843.000 167.700 844.050 ;
        RECT 163.800 841.500 165.900 841.800 ;
        RECT 146.100 838.050 147.900 839.850 ;
        RECT 162.000 839.700 165.900 841.500 ;
        RECT 166.800 841.050 167.700 843.000 ;
        RECT 166.800 838.950 168.900 841.050 ;
        RECT 166.800 838.800 168.300 838.950 ;
        RECT 163.200 838.050 165.000 838.500 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 158.100 836.700 165.000 838.050 ;
        RECT 165.900 837.900 168.300 838.800 ;
        RECT 172.800 838.050 174.600 839.850 ;
        RECT 188.100 838.050 189.300 851.400 ;
        RECT 206.100 845.400 207.900 857.400 ;
        RECT 209.100 846.300 210.900 857.400 ;
        RECT 212.100 847.200 213.900 858.000 ;
        RECT 215.100 846.300 216.900 857.400 ;
        RECT 227.700 851.400 229.500 858.000 ;
        RECT 228.000 848.100 229.800 849.900 ;
        RECT 230.700 846.900 232.500 857.400 ;
        RECT 209.100 845.400 216.900 846.300 ;
        RECT 230.100 845.400 232.500 846.900 ;
        RECT 235.800 845.400 237.600 858.000 ;
        RECT 248.100 851.400 249.900 858.000 ;
        RECT 251.100 851.400 252.900 857.400 ;
        RECT 254.100 851.400 255.900 858.000 ;
        RECT 202.950 840.450 205.050 841.050 ;
        RECT 197.550 839.550 205.050 840.450 ;
        RECT 158.100 835.950 160.200 836.700 ;
        RECT 131.550 833.550 136.050 835.050 ;
        RECT 137.100 834.150 138.900 835.950 ;
        RECT 132.000 832.950 136.050 833.550 ;
        RECT 140.100 831.600 141.300 835.950 ;
        RECT 143.100 834.150 144.900 835.950 ;
        RECT 158.400 834.150 160.200 835.950 ;
        RECT 163.200 833.400 165.000 835.200 ;
        RECT 137.700 830.700 141.300 831.600 ;
        RECT 162.900 831.300 165.000 833.400 ;
        RECT 137.700 828.600 138.900 830.700 ;
        RECT 158.700 830.400 165.000 831.300 ;
        RECT 165.900 832.200 167.100 837.900 ;
        RECT 168.300 835.200 170.100 837.000 ;
        RECT 172.800 835.950 174.900 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 168.000 833.100 170.100 835.200 ;
        RECT 185.250 834.150 187.050 835.950 ;
        RECT 122.100 822.000 123.900 825.600 ;
        RECT 125.100 822.600 126.900 825.600 ;
        RECT 137.100 822.600 138.900 828.600 ;
        RECT 140.100 827.700 147.900 829.050 ;
        RECT 158.700 828.600 159.900 830.400 ;
        RECT 165.900 830.100 168.900 832.200 ;
        RECT 188.100 830.700 189.300 835.950 ;
        RECT 191.100 834.150 192.900 835.950 ;
        RECT 197.550 835.050 198.450 839.550 ;
        RECT 202.950 838.950 205.050 839.550 ;
        RECT 206.400 838.050 207.300 845.400 ;
        RECT 222.000 840.450 226.050 841.050 ;
        RECT 211.950 838.050 213.750 839.850 ;
        RECT 221.550 838.950 226.050 840.450 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 193.950 833.550 198.450 835.050 ;
        RECT 193.950 832.950 198.000 833.550 ;
        RECT 165.900 828.600 167.100 830.100 ;
        RECT 170.100 829.500 172.200 830.700 ;
        RECT 188.100 829.800 192.300 830.700 ;
        RECT 170.100 828.600 174.900 829.500 ;
        RECT 140.100 822.600 141.900 827.700 ;
        RECT 143.100 822.000 144.900 826.800 ;
        RECT 146.100 822.600 147.900 827.700 ;
        RECT 158.100 822.600 159.900 828.600 ;
        RECT 161.100 822.000 162.900 827.700 ;
        RECT 165.600 822.600 167.400 828.600 ;
        RECT 170.100 822.000 171.900 827.700 ;
        RECT 173.100 822.600 174.900 828.600 ;
        RECT 185.400 822.000 187.200 828.600 ;
        RECT 190.500 822.600 192.300 829.800 ;
        RECT 206.400 828.600 207.300 835.950 ;
        RECT 208.950 834.150 210.750 835.950 ;
        RECT 215.100 834.150 216.900 835.950 ;
        RECT 211.950 831.450 214.050 832.050 ;
        RECT 221.550 831.450 222.450 838.950 ;
        RECT 230.100 838.050 231.300 845.400 ;
        RECT 236.100 838.050 237.900 839.850 ;
        RECT 251.100 838.050 252.300 851.400 ;
        RECT 270.000 846.600 271.800 857.400 ;
        RECT 270.000 845.400 273.600 846.600 ;
        RECT 275.100 845.400 276.900 858.000 ;
        RECT 287.100 846.300 288.900 857.400 ;
        RECT 290.100 847.500 291.900 858.000 ;
        RECT 294.600 846.300 296.400 857.400 ;
        RECT 298.800 847.500 300.900 858.000 ;
        RECT 302.100 846.600 303.900 857.400 ;
        RECT 269.100 838.050 270.900 839.850 ;
        RECT 272.700 838.050 273.600 845.400 ;
        RECT 287.100 845.100 291.900 846.300 ;
        RECT 294.600 845.400 297.900 846.300 ;
        RECT 289.800 844.200 291.900 845.100 ;
        RECT 289.800 843.300 295.200 844.200 ;
        RECT 293.400 841.500 295.200 843.300 ;
        RECT 296.700 841.050 297.900 845.400 ;
        RECT 298.800 845.400 303.900 846.600 ;
        RECT 317.100 846.300 318.900 857.400 ;
        RECT 320.100 847.500 321.900 858.000 ;
        RECT 317.100 845.400 321.600 846.300 ;
        RECT 324.600 845.400 326.400 857.400 ;
        RECT 329.100 847.500 330.900 858.000 ;
        RECT 332.100 846.600 333.900 857.400 ;
        RECT 298.800 844.500 300.900 845.400 ;
        RECT 319.500 843.300 321.600 845.400 ;
        RECT 325.200 844.050 326.400 845.400 ;
        RECT 329.100 845.400 333.900 846.600 ;
        RECT 347.100 846.300 348.900 857.400 ;
        RECT 350.100 847.200 351.900 858.000 ;
        RECT 353.100 846.300 354.900 857.400 ;
        RECT 347.100 845.400 354.900 846.300 ;
        RECT 356.100 845.400 357.900 857.400 ;
        RECT 368.700 851.400 370.500 858.000 ;
        RECT 369.000 848.100 370.800 849.900 ;
        RECT 371.700 846.900 373.500 857.400 ;
        RECT 371.100 845.400 373.500 846.900 ;
        RECT 376.800 845.400 378.600 858.000 ;
        RECT 389.100 846.300 390.900 857.400 ;
        RECT 392.100 847.200 393.900 858.000 ;
        RECT 395.100 846.300 396.900 857.400 ;
        RECT 389.100 845.400 396.900 846.300 ;
        RECT 398.100 845.400 399.900 857.400 ;
        RECT 413.400 845.400 415.200 858.000 ;
        RECT 418.500 846.900 420.300 857.400 ;
        RECT 421.500 851.400 423.300 858.000 ;
        RECT 421.200 848.100 423.000 849.900 ;
        RECT 418.500 845.400 420.900 846.900 ;
        RECT 435.000 846.600 436.800 857.400 ;
        RECT 435.000 845.400 438.600 846.600 ;
        RECT 440.100 845.400 441.900 858.000 ;
        RECT 455.100 851.400 456.900 858.000 ;
        RECT 458.100 851.400 459.900 857.400 ;
        RECT 461.100 851.400 462.900 858.000 ;
        RECT 476.700 851.400 478.500 858.000 ;
        RECT 329.100 844.500 331.200 845.400 ;
        RECT 325.200 843.000 326.700 844.050 ;
        RECT 322.800 841.500 324.900 841.800 ;
        RECT 296.100 840.300 298.200 841.050 ;
        RECT 274.950 838.050 276.750 839.850 ;
        RECT 291.900 838.200 293.700 840.000 ;
        RECT 295.200 838.950 298.200 840.300 ;
        RECT 226.950 835.950 229.050 838.050 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 247.950 835.950 250.050 838.050 ;
        RECT 250.950 835.950 253.050 838.050 ;
        RECT 253.950 835.950 256.050 838.050 ;
        RECT 268.950 835.950 271.050 838.050 ;
        RECT 271.950 835.950 274.050 838.050 ;
        RECT 274.950 835.950 277.050 838.050 ;
        RECT 227.100 834.150 228.900 835.950 ;
        RECT 230.100 831.600 231.300 835.950 ;
        RECT 233.100 834.150 234.900 835.950 ;
        RECT 248.250 834.150 250.050 835.950 ;
        RECT 211.950 830.550 222.450 831.450 ;
        RECT 227.700 830.700 231.300 831.600 ;
        RECT 251.100 830.700 252.300 835.950 ;
        RECT 254.100 834.150 255.900 835.950 ;
        RECT 211.950 829.950 214.050 830.550 ;
        RECT 227.700 828.600 228.900 830.700 ;
        RECT 251.100 829.800 255.300 830.700 ;
        RECT 206.400 827.400 211.500 828.600 ;
        RECT 206.700 822.000 208.500 825.600 ;
        RECT 209.700 822.600 211.500 827.400 ;
        RECT 214.200 822.000 216.000 828.600 ;
        RECT 227.100 822.600 228.900 828.600 ;
        RECT 230.100 827.700 237.900 829.050 ;
        RECT 230.100 822.600 231.900 827.700 ;
        RECT 233.100 822.000 234.900 826.800 ;
        RECT 236.100 822.600 237.900 827.700 ;
        RECT 248.400 822.000 250.200 828.600 ;
        RECT 253.500 822.600 255.300 829.800 ;
        RECT 272.700 825.600 273.600 835.950 ;
        RECT 287.100 835.800 289.200 838.050 ;
        RECT 291.900 836.100 294.000 838.200 ;
        RECT 287.400 835.200 289.200 835.800 ;
        RECT 287.400 834.000 294.000 835.200 ;
        RECT 291.900 833.100 294.000 834.000 ;
        RECT 289.500 831.000 291.600 831.600 ;
        RECT 292.500 831.300 294.300 833.100 ;
        RECT 295.200 832.200 296.100 838.950 ;
        RECT 301.800 838.050 303.600 839.850 ;
        RECT 321.000 839.700 324.900 841.500 ;
        RECT 325.800 841.050 326.700 843.000 ;
        RECT 325.800 838.950 327.900 841.050 ;
        RECT 325.800 838.800 327.300 838.950 ;
        RECT 322.200 838.050 324.000 838.500 ;
        RECT 297.000 836.100 298.800 837.900 ;
        RECT 297.000 834.000 299.100 836.100 ;
        RECT 301.800 835.950 303.900 838.050 ;
        RECT 317.100 836.700 324.000 838.050 ;
        RECT 324.900 837.900 327.300 838.800 ;
        RECT 331.800 838.050 333.600 839.850 ;
        RECT 350.250 838.050 352.050 839.850 ;
        RECT 356.700 838.050 357.600 845.400 ;
        RECT 371.100 838.050 372.300 845.400 ;
        RECT 377.100 838.050 378.900 839.850 ;
        RECT 392.250 838.050 394.050 839.850 ;
        RECT 398.700 838.050 399.600 845.400 ;
        RECT 409.950 840.450 412.050 841.050 ;
        RECT 404.550 839.550 412.050 840.450 ;
        RECT 317.100 835.950 319.200 836.700 ;
        RECT 317.400 834.150 319.200 835.950 ;
        RECT 322.200 833.400 324.000 835.200 ;
        RECT 287.100 829.500 291.600 831.000 ;
        RECT 295.200 830.100 298.200 832.200 ;
        RECT 287.100 828.600 288.600 829.500 ;
        RECT 269.100 822.000 270.900 825.600 ;
        RECT 272.100 822.600 273.900 825.600 ;
        RECT 275.100 822.000 276.900 825.600 ;
        RECT 287.100 822.600 288.900 828.600 ;
        RECT 295.200 828.000 296.100 830.100 ;
        RECT 299.400 829.500 301.500 831.900 ;
        RECT 321.900 831.300 324.000 833.400 ;
        RECT 317.700 830.400 324.000 831.300 ;
        RECT 324.900 832.200 326.100 837.900 ;
        RECT 327.300 835.200 329.100 837.000 ;
        RECT 331.800 835.950 333.900 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 352.950 835.950 355.050 838.050 ;
        RECT 355.950 835.950 358.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 376.950 835.950 379.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 394.950 835.950 397.050 838.050 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 327.000 833.100 329.100 835.200 ;
        RECT 347.100 834.150 348.900 835.950 ;
        RECT 353.250 834.150 355.050 835.950 ;
        RECT 299.400 828.600 303.900 829.500 ;
        RECT 317.700 828.600 318.900 830.400 ;
        RECT 324.900 830.100 327.900 832.200 ;
        RECT 334.950 831.450 337.050 832.050 ;
        RECT 349.950 831.450 352.050 832.050 ;
        RECT 324.900 828.600 326.100 830.100 ;
        RECT 329.100 829.500 331.200 830.700 ;
        RECT 334.950 830.550 352.050 831.450 ;
        RECT 334.950 829.950 337.050 830.550 ;
        RECT 349.950 829.950 352.050 830.550 ;
        RECT 329.100 828.600 333.900 829.500 ;
        RECT 356.700 828.600 357.600 835.950 ;
        RECT 368.100 834.150 369.900 835.950 ;
        RECT 371.100 831.600 372.300 835.950 ;
        RECT 374.100 834.150 375.900 835.950 ;
        RECT 389.100 834.150 390.900 835.950 ;
        RECT 395.250 834.150 397.050 835.950 ;
        RECT 368.700 830.700 372.300 831.600 ;
        RECT 368.700 828.600 369.900 830.700 ;
        RECT 290.100 822.000 291.900 827.700 ;
        RECT 294.300 822.600 296.100 828.000 ;
        RECT 298.800 822.000 300.600 827.700 ;
        RECT 302.100 822.600 303.900 828.600 ;
        RECT 317.100 822.600 318.900 828.600 ;
        RECT 320.100 822.000 321.900 827.700 ;
        RECT 324.600 822.600 326.400 828.600 ;
        RECT 329.100 822.000 330.900 827.700 ;
        RECT 332.100 822.600 333.900 828.600 ;
        RECT 348.000 822.000 349.800 828.600 ;
        RECT 352.500 827.400 357.600 828.600 ;
        RECT 352.500 822.600 354.300 827.400 ;
        RECT 355.500 822.000 357.300 825.600 ;
        RECT 368.100 822.600 369.900 828.600 ;
        RECT 371.100 827.700 378.900 829.050 ;
        RECT 398.700 828.600 399.600 835.950 ;
        RECT 404.550 835.050 405.450 839.550 ;
        RECT 409.950 838.950 412.050 839.550 ;
        RECT 413.100 838.050 414.900 839.850 ;
        RECT 419.700 838.050 420.900 845.400 ;
        RECT 434.100 838.050 435.900 839.850 ;
        RECT 437.700 838.050 438.600 845.400 ;
        RECT 439.950 838.050 441.750 839.850 ;
        RECT 458.700 838.050 459.900 851.400 ;
        RECT 477.000 848.100 478.800 849.900 ;
        RECT 479.700 846.900 481.500 857.400 ;
        RECT 479.100 845.400 481.500 846.900 ;
        RECT 484.800 845.400 486.600 858.000 ;
        RECT 497.700 851.400 499.500 858.000 ;
        RECT 498.000 848.100 499.800 849.900 ;
        RECT 500.700 846.900 502.500 857.400 ;
        RECT 500.100 845.400 502.500 846.900 ;
        RECT 505.800 845.400 507.600 858.000 ;
        RECT 521.100 845.400 522.900 858.000 ;
        RECT 526.200 846.600 528.000 857.400 ;
        RECT 539.100 851.400 540.900 857.400 ;
        RECT 542.100 851.400 543.900 858.000 ;
        RECT 554.100 851.400 555.900 858.000 ;
        RECT 557.100 851.400 558.900 857.400 ;
        RECT 560.100 851.400 561.900 858.000 ;
        RECT 524.400 845.400 528.000 846.600 ;
        RECT 471.000 840.450 475.050 841.050 ;
        RECT 470.550 838.950 475.050 840.450 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 415.950 835.950 418.050 838.050 ;
        RECT 418.950 835.950 421.050 838.050 ;
        RECT 421.950 835.950 424.050 838.050 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 400.950 833.550 405.450 835.050 ;
        RECT 416.100 834.150 417.900 835.950 ;
        RECT 400.950 832.950 405.000 833.550 ;
        RECT 419.700 831.600 420.900 835.950 ;
        RECT 422.100 834.150 423.900 835.950 ;
        RECT 419.700 830.700 423.300 831.600 ;
        RECT 371.100 822.600 372.900 827.700 ;
        RECT 374.100 822.000 375.900 826.800 ;
        RECT 377.100 822.600 378.900 827.700 ;
        RECT 390.000 822.000 391.800 828.600 ;
        RECT 394.500 827.400 399.600 828.600 ;
        RECT 413.100 827.700 420.900 829.050 ;
        RECT 394.500 822.600 396.300 827.400 ;
        RECT 397.500 822.000 399.300 825.600 ;
        RECT 413.100 822.600 414.900 827.700 ;
        RECT 416.100 822.000 417.900 826.800 ;
        RECT 419.100 822.600 420.900 827.700 ;
        RECT 422.100 828.600 423.300 830.700 ;
        RECT 422.100 822.600 423.900 828.600 ;
        RECT 437.700 825.600 438.600 835.950 ;
        RECT 455.100 834.150 456.900 835.950 ;
        RECT 458.700 830.700 459.900 835.950 ;
        RECT 460.950 834.150 462.750 835.950 ;
        RECT 470.550 835.050 471.450 838.950 ;
        RECT 479.100 838.050 480.300 845.400 ;
        RECT 481.950 843.450 484.050 844.050 ;
        RECT 481.950 842.550 489.450 843.450 ;
        RECT 481.950 841.950 484.050 842.550 ;
        RECT 488.550 840.450 489.450 842.550 ;
        RECT 485.100 838.050 486.900 839.850 ;
        RECT 488.550 839.550 492.450 840.450 ;
        RECT 475.950 835.950 478.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 470.550 833.550 475.050 835.050 ;
        RECT 476.100 834.150 477.900 835.950 ;
        RECT 471.000 832.950 475.050 833.550 ;
        RECT 479.100 831.600 480.300 835.950 ;
        RECT 482.100 834.150 483.900 835.950 ;
        RECT 491.550 834.450 492.450 839.550 ;
        RECT 500.100 838.050 501.300 845.400 ;
        RECT 506.100 838.050 507.900 839.850 ;
        RECT 521.250 838.050 523.050 839.850 ;
        RECT 524.400 838.050 525.300 845.400 ;
        RECT 527.100 838.050 528.900 839.850 ;
        RECT 539.700 838.050 540.900 851.400 ;
        RECT 542.100 838.050 543.900 839.850 ;
        RECT 557.100 838.050 558.300 851.400 ;
        RECT 572.400 845.400 574.200 858.000 ;
        RECT 577.500 846.900 579.300 857.400 ;
        RECT 580.500 851.400 582.300 858.000 ;
        RECT 596.700 851.400 598.500 858.000 ;
        RECT 580.200 848.100 582.000 849.900 ;
        RECT 597.000 848.100 598.800 849.900 ;
        RECT 599.700 846.900 601.500 857.400 ;
        RECT 577.500 845.400 579.900 846.900 ;
        RECT 572.100 838.050 573.900 839.850 ;
        RECT 578.700 838.050 579.900 845.400 ;
        RECT 599.100 845.400 601.500 846.900 ;
        RECT 604.800 845.400 606.600 858.000 ;
        RECT 617.100 851.400 618.900 858.000 ;
        RECT 620.100 851.400 621.900 857.400 ;
        RECT 623.100 851.400 624.900 858.000 ;
        RECT 638.100 851.400 639.900 857.400 ;
        RECT 641.100 851.400 642.900 858.000 ;
        RECT 599.100 838.050 600.300 845.400 ;
        RECT 612.000 840.450 616.050 841.050 ;
        RECT 605.100 838.050 606.900 839.850 ;
        RECT 611.550 838.950 616.050 840.450 ;
        RECT 496.950 835.950 499.050 838.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 520.950 835.950 523.050 838.050 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 571.950 835.950 574.050 838.050 ;
        RECT 574.950 835.950 577.050 838.050 ;
        RECT 577.950 835.950 580.050 838.050 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 595.950 835.950 598.050 838.050 ;
        RECT 598.950 835.950 601.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 491.550 834.000 495.450 834.450 ;
        RECT 497.100 834.150 498.900 835.950 ;
        RECT 491.550 833.550 496.050 834.000 ;
        RECT 455.700 829.800 459.900 830.700 ;
        RECT 476.700 830.700 480.300 831.600 ;
        RECT 434.100 822.000 435.900 825.600 ;
        RECT 437.100 822.600 438.900 825.600 ;
        RECT 440.100 822.000 441.900 825.600 ;
        RECT 455.700 822.600 457.500 829.800 ;
        RECT 476.700 828.600 477.900 830.700 ;
        RECT 493.950 829.950 496.050 833.550 ;
        RECT 500.100 831.600 501.300 835.950 ;
        RECT 503.100 834.150 504.900 835.950 ;
        RECT 497.700 830.700 501.300 831.600 ;
        RECT 460.800 822.000 462.600 828.600 ;
        RECT 476.100 822.600 477.900 828.600 ;
        RECT 479.100 827.700 486.900 829.050 ;
        RECT 497.700 828.600 498.900 830.700 ;
        RECT 479.100 822.600 480.900 827.700 ;
        RECT 482.100 822.000 483.900 826.800 ;
        RECT 485.100 822.600 486.900 827.700 ;
        RECT 497.100 822.600 498.900 828.600 ;
        RECT 500.100 827.700 507.900 829.050 ;
        RECT 500.100 822.600 501.900 827.700 ;
        RECT 503.100 822.000 504.900 826.800 ;
        RECT 506.100 822.600 507.900 827.700 ;
        RECT 524.400 825.600 525.300 835.950 ;
        RECT 526.950 831.450 529.050 831.750 ;
        RECT 532.950 831.450 535.050 832.050 ;
        RECT 526.950 830.550 535.050 831.450 ;
        RECT 526.950 829.650 529.050 830.550 ;
        RECT 532.950 829.950 535.050 830.550 ;
        RECT 539.700 825.600 540.900 835.950 ;
        RECT 554.250 834.150 556.050 835.950 ;
        RECT 557.100 830.700 558.300 835.950 ;
        RECT 560.100 834.150 561.900 835.950 ;
        RECT 575.100 834.150 576.900 835.950 ;
        RECT 578.700 831.600 579.900 835.950 ;
        RECT 581.100 834.150 582.900 835.950 ;
        RECT 596.100 834.150 597.900 835.950 ;
        RECT 599.100 831.600 600.300 835.950 ;
        RECT 602.100 834.150 603.900 835.950 ;
        RECT 611.550 835.050 612.450 838.950 ;
        RECT 620.100 838.050 621.300 851.400 ;
        RECT 638.700 838.050 639.900 851.400 ;
        RECT 653.100 850.200 654.900 856.200 ;
        RECT 653.100 845.100 654.000 850.200 ;
        RECT 656.100 846.000 657.900 858.000 ;
        RECT 660.600 846.900 662.400 857.400 ;
        RECT 660.600 846.000 662.700 846.900 ;
        RECT 653.100 844.200 660.900 845.100 ;
        RECT 659.700 839.850 660.900 844.200 ;
        RECT 641.100 838.050 642.900 839.850 ;
        RECT 656.100 838.050 657.900 839.850 ;
        RECT 659.100 838.050 660.900 839.850 ;
        RECT 661.800 838.050 662.700 846.000 ;
        RECT 665.100 845.400 666.900 858.000 ;
        RECT 677.100 851.400 678.900 858.000 ;
        RECT 680.100 851.400 681.900 857.400 ;
        RECT 683.100 851.400 684.900 858.000 ;
        RECT 698.100 851.400 699.900 857.400 ;
        RECT 664.800 838.050 666.600 839.850 ;
        RECT 680.700 838.050 681.900 851.400 ;
        RECT 698.100 844.500 699.300 851.400 ;
        RECT 701.100 847.200 702.900 858.000 ;
        RECT 704.100 845.400 705.900 857.400 ;
        RECT 698.100 843.600 703.800 844.500 ;
        RECT 702.000 842.700 703.800 843.600 ;
        RECT 698.400 838.050 700.200 839.850 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 653.100 835.950 655.200 838.050 ;
        RECT 656.100 835.950 658.200 838.050 ;
        RECT 611.550 833.550 616.050 835.050 ;
        RECT 617.250 834.150 619.050 835.950 ;
        RECT 612.000 832.950 616.050 833.550 ;
        RECT 578.700 830.700 582.300 831.600 ;
        RECT 557.100 829.800 561.300 830.700 ;
        RECT 521.100 822.000 522.900 825.600 ;
        RECT 524.100 822.600 525.900 825.600 ;
        RECT 527.100 822.000 528.900 825.600 ;
        RECT 539.100 822.600 540.900 825.600 ;
        RECT 542.100 822.000 543.900 825.600 ;
        RECT 554.400 822.000 556.200 828.600 ;
        RECT 559.500 822.600 561.300 829.800 ;
        RECT 572.100 827.700 579.900 829.050 ;
        RECT 572.100 822.600 573.900 827.700 ;
        RECT 575.100 822.000 576.900 826.800 ;
        RECT 578.100 822.600 579.900 827.700 ;
        RECT 581.100 828.600 582.300 830.700 ;
        RECT 596.700 830.700 600.300 831.600 ;
        RECT 620.100 830.700 621.300 835.950 ;
        RECT 623.100 834.150 624.900 835.950 ;
        RECT 596.700 828.600 597.900 830.700 ;
        RECT 620.100 829.800 624.300 830.700 ;
        RECT 581.100 822.600 582.900 828.600 ;
        RECT 596.100 822.600 597.900 828.600 ;
        RECT 599.100 827.700 606.900 829.050 ;
        RECT 599.100 822.600 600.900 827.700 ;
        RECT 602.100 822.000 603.900 826.800 ;
        RECT 605.100 822.600 606.900 827.700 ;
        RECT 617.400 822.000 619.200 828.600 ;
        RECT 622.500 822.600 624.300 829.800 ;
        RECT 638.700 825.600 639.900 835.950 ;
        RECT 653.100 834.150 654.900 835.950 ;
        RECT 659.100 831.000 660.300 838.050 ;
        RECT 653.100 830.100 660.300 831.000 ;
        RECT 661.800 835.950 663.900 838.050 ;
        RECT 664.800 835.950 666.900 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 682.950 835.950 685.050 838.050 ;
        RECT 698.400 835.950 700.500 838.050 ;
        RECT 653.100 826.800 654.000 830.100 ;
        RECT 661.800 829.200 662.700 835.950 ;
        RECT 677.100 834.150 678.900 835.950 ;
        RECT 680.700 830.700 681.900 835.950 ;
        RECT 682.950 834.150 684.750 835.950 ;
        RECT 677.700 829.800 681.900 830.700 ;
        RECT 702.000 831.300 702.900 842.700 ;
        RECT 704.700 838.050 705.900 845.400 ;
        RECT 716.100 851.400 717.900 857.400 ;
        RECT 716.100 844.500 717.300 851.400 ;
        RECT 719.100 847.200 720.900 858.000 ;
        RECT 722.100 845.400 723.900 857.400 ;
        RECT 737.100 851.400 738.900 858.000 ;
        RECT 740.100 851.400 741.900 857.400 ;
        RECT 716.100 843.600 721.800 844.500 ;
        RECT 720.000 842.700 721.800 843.600 ;
        RECT 703.800 835.950 705.900 838.050 ;
        RECT 716.400 838.050 718.200 839.850 ;
        RECT 716.400 835.950 718.500 838.050 ;
        RECT 702.000 830.400 703.800 831.300 ;
        RECT 638.100 822.600 639.900 825.600 ;
        RECT 641.100 822.000 642.900 825.600 ;
        RECT 653.100 823.800 654.900 826.800 ;
        RECT 656.100 824.400 657.900 829.200 ;
        RECT 660.600 828.300 662.700 829.200 ;
        RECT 656.100 822.000 657.300 824.400 ;
        RECT 660.600 823.800 662.400 828.300 ;
        RECT 665.100 823.800 666.900 829.800 ;
        RECT 665.100 822.000 666.300 823.800 ;
        RECT 677.700 822.600 679.500 829.800 ;
        RECT 698.100 829.500 703.800 830.400 ;
        RECT 682.800 822.000 684.600 828.600 ;
        RECT 698.100 825.600 699.300 829.500 ;
        RECT 704.700 828.600 705.900 835.950 ;
        RECT 720.000 831.300 720.900 842.700 ;
        RECT 722.700 838.050 723.900 845.400 ;
        RECT 737.100 838.050 738.900 839.850 ;
        RECT 740.100 838.050 741.300 851.400 ;
        RECT 752.100 845.400 753.900 857.400 ;
        RECT 755.100 846.300 756.900 857.400 ;
        RECT 758.100 847.200 759.900 858.000 ;
        RECT 761.100 846.300 762.900 857.400 ;
        RECT 776.100 851.400 777.900 858.000 ;
        RECT 779.100 851.400 780.900 857.400 ;
        RECT 782.100 852.000 783.900 858.000 ;
        RECT 779.400 851.100 780.900 851.400 ;
        RECT 785.100 851.400 786.900 857.400 ;
        RECT 797.100 851.400 798.900 858.000 ;
        RECT 800.100 851.400 801.900 857.400 ;
        RECT 803.100 851.400 804.900 858.000 ;
        RECT 785.100 851.100 786.000 851.400 ;
        RECT 779.400 850.200 786.000 851.100 ;
        RECT 755.100 845.400 762.900 846.300 ;
        RECT 752.400 838.050 753.300 845.400 ;
        RECT 757.950 838.050 759.750 839.850 ;
        RECT 779.100 838.050 780.900 839.850 ;
        RECT 785.100 838.050 786.000 850.200 ;
        RECT 800.700 838.050 801.900 851.400 ;
        RECT 818.400 845.400 820.200 858.000 ;
        RECT 823.500 846.900 825.300 857.400 ;
        RECT 826.500 851.400 828.300 858.000 ;
        RECT 826.200 848.100 828.000 849.900 ;
        RECT 823.500 845.400 825.900 846.900 ;
        RECT 839.400 845.400 841.200 858.000 ;
        RECT 844.500 846.900 846.300 857.400 ;
        RECT 847.500 851.400 849.300 858.000 ;
        RECT 847.200 848.100 849.000 849.900 ;
        RECT 844.500 845.400 846.900 846.900 ;
        RECT 863.400 845.400 865.200 858.000 ;
        RECT 868.500 846.900 870.300 857.400 ;
        RECT 871.500 851.400 873.300 858.000 ;
        RECT 871.200 848.100 873.000 849.900 ;
        RECT 868.500 845.400 870.900 846.900 ;
        RECT 884.400 845.400 886.200 858.000 ;
        RECT 889.500 846.900 891.300 857.400 ;
        RECT 892.500 851.400 894.300 858.000 ;
        RECT 892.200 848.100 894.000 849.900 ;
        RECT 906.600 846.900 908.400 857.400 ;
        RECT 889.500 845.400 891.900 846.900 ;
        RECT 818.100 838.050 819.900 839.850 ;
        RECT 824.700 838.050 825.900 845.400 ;
        RECT 839.100 838.050 840.900 839.850 ;
        RECT 845.700 838.050 846.900 845.400 ;
        RECT 853.950 843.450 856.050 844.050 ;
        RECT 859.950 843.450 862.050 844.050 ;
        RECT 853.950 842.550 862.050 843.450 ;
        RECT 853.950 841.950 856.050 842.550 ;
        RECT 859.950 841.950 862.050 842.550 ;
        RECT 850.950 840.450 853.050 841.050 ;
        RECT 856.950 840.450 859.050 841.050 ;
        RECT 850.950 839.550 859.050 840.450 ;
        RECT 850.950 838.950 853.050 839.550 ;
        RECT 856.950 838.950 859.050 839.550 ;
        RECT 863.100 838.050 864.900 839.850 ;
        RECT 869.700 838.050 870.900 845.400 ;
        RECT 884.100 838.050 885.900 839.850 ;
        RECT 890.700 838.050 891.900 845.400 ;
        RECT 906.000 845.400 908.400 846.900 ;
        RECT 909.600 845.400 911.400 858.000 ;
        RECT 914.100 845.400 915.900 857.400 ;
        RECT 906.000 838.050 907.200 845.400 ;
        RECT 914.700 843.900 915.900 845.400 ;
        RECT 908.100 842.700 915.900 843.900 ;
        RECT 908.100 842.100 909.900 842.700 ;
        RECT 721.800 835.950 723.900 838.050 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 796.950 835.950 799.050 838.050 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 820.950 835.950 823.050 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 905.100 835.950 907.200 838.050 ;
        RECT 720.000 830.400 721.800 831.300 ;
        RECT 698.100 822.600 699.900 825.600 ;
        RECT 701.100 822.000 702.900 828.600 ;
        RECT 704.100 822.600 705.900 828.600 ;
        RECT 716.100 829.500 721.800 830.400 ;
        RECT 716.100 825.600 717.300 829.500 ;
        RECT 722.700 828.600 723.900 835.950 ;
        RECT 716.100 822.600 717.900 825.600 ;
        RECT 719.100 822.000 720.900 828.600 ;
        RECT 722.100 822.600 723.900 828.600 ;
        RECT 740.100 825.600 741.300 835.950 ;
        RECT 752.400 828.600 753.300 835.950 ;
        RECT 754.950 834.150 756.750 835.950 ;
        RECT 761.100 834.150 762.900 835.950 ;
        RECT 776.100 834.150 777.900 835.950 ;
        RECT 782.100 834.150 783.900 835.950 ;
        RECT 785.100 832.200 786.000 835.950 ;
        RECT 797.100 834.150 798.900 835.950 ;
        RECT 752.400 827.400 757.500 828.600 ;
        RECT 737.100 822.000 738.900 825.600 ;
        RECT 740.100 822.600 741.900 825.600 ;
        RECT 752.700 822.000 754.500 825.600 ;
        RECT 755.700 822.600 757.500 827.400 ;
        RECT 760.200 822.000 762.000 828.600 ;
        RECT 776.100 822.000 777.900 831.600 ;
        RECT 782.700 831.000 786.000 832.200 ;
        RECT 782.700 822.600 784.500 831.000 ;
        RECT 800.700 830.700 801.900 835.950 ;
        RECT 802.950 834.150 804.750 835.950 ;
        RECT 821.100 834.150 822.900 835.950 ;
        RECT 824.700 831.600 825.900 835.950 ;
        RECT 827.100 834.150 828.900 835.950 ;
        RECT 842.100 834.150 843.900 835.950 ;
        RECT 845.700 831.600 846.900 835.950 ;
        RECT 848.100 834.150 849.900 835.950 ;
        RECT 866.100 834.150 867.900 835.950 ;
        RECT 869.700 831.600 870.900 835.950 ;
        RECT 872.100 834.150 873.900 835.950 ;
        RECT 887.100 834.150 888.900 835.950 ;
        RECT 890.700 831.600 891.900 835.950 ;
        RECT 893.100 834.150 894.900 835.950 ;
        RECT 824.700 830.700 828.300 831.600 ;
        RECT 845.700 830.700 849.300 831.600 ;
        RECT 869.700 830.700 873.300 831.600 ;
        RECT 890.700 830.700 894.300 831.600 ;
        RECT 797.700 829.800 801.900 830.700 ;
        RECT 797.700 822.600 799.500 829.800 ;
        RECT 802.800 822.000 804.600 828.600 ;
        RECT 818.100 827.700 825.900 829.050 ;
        RECT 818.100 822.600 819.900 827.700 ;
        RECT 821.100 822.000 822.900 826.800 ;
        RECT 824.100 822.600 825.900 827.700 ;
        RECT 827.100 828.600 828.300 830.700 ;
        RECT 827.100 822.600 828.900 828.600 ;
        RECT 839.100 827.700 846.900 829.050 ;
        RECT 839.100 822.600 840.900 827.700 ;
        RECT 842.100 822.000 843.900 826.800 ;
        RECT 845.100 822.600 846.900 827.700 ;
        RECT 848.100 828.600 849.300 830.700 ;
        RECT 848.100 822.600 849.900 828.600 ;
        RECT 863.100 827.700 870.900 829.050 ;
        RECT 863.100 822.600 864.900 827.700 ;
        RECT 866.100 822.000 867.900 826.800 ;
        RECT 869.100 822.600 870.900 827.700 ;
        RECT 872.100 828.600 873.300 830.700 ;
        RECT 872.100 822.600 873.900 828.600 ;
        RECT 884.100 827.700 891.900 829.050 ;
        RECT 884.100 822.600 885.900 827.700 ;
        RECT 887.100 822.000 888.900 826.800 ;
        RECT 890.100 822.600 891.900 827.700 ;
        RECT 893.100 828.600 894.300 830.700 ;
        RECT 905.100 828.600 906.000 835.950 ;
        RECT 908.400 831.600 909.300 842.100 ;
        RECT 910.200 838.050 912.000 839.850 ;
        RECT 910.500 835.950 912.600 838.050 ;
        RECT 913.800 835.950 915.900 838.050 ;
        RECT 913.800 834.150 915.600 835.950 ;
        RECT 907.200 830.700 909.300 831.600 ;
        RECT 907.200 829.800 912.600 830.700 ;
        RECT 893.100 822.600 894.900 828.600 ;
        RECT 905.100 822.600 906.900 828.600 ;
        RECT 908.100 822.000 909.900 828.000 ;
        RECT 911.700 825.600 912.600 829.800 ;
        RECT 911.100 822.600 912.900 825.600 ;
        RECT 914.100 822.600 915.900 825.600 ;
        RECT 914.700 822.000 915.900 822.600 ;
        RECT 14.100 812.400 15.900 818.400 ;
        RECT 14.700 810.300 15.900 812.400 ;
        RECT 17.100 813.300 18.900 818.400 ;
        RECT 20.100 814.200 21.900 819.000 ;
        RECT 23.100 813.300 24.900 818.400 ;
        RECT 17.100 811.950 24.900 813.300 ;
        RECT 38.700 811.200 40.500 818.400 ;
        RECT 43.800 812.400 45.600 819.000 ;
        RECT 56.400 812.400 58.200 819.000 ;
        RECT 61.500 811.200 63.300 818.400 ;
        RECT 74.100 812.400 75.900 818.400 ;
        RECT 38.700 810.300 42.900 811.200 ;
        RECT 55.950 810.450 58.050 811.050 ;
        RECT 14.700 809.400 18.300 810.300 ;
        RECT 14.100 805.050 15.900 806.850 ;
        RECT 17.100 805.050 18.300 809.400 ;
        RECT 20.100 805.050 21.900 806.850 ;
        RECT 38.100 805.050 39.900 806.850 ;
        RECT 41.700 805.050 42.900 810.300 ;
        RECT 50.550 809.550 58.050 810.450 ;
        RECT 43.950 805.050 45.750 806.850 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 7.950 798.450 10.050 799.050 ;
        RECT 13.950 798.450 16.050 799.050 ;
        RECT 7.950 797.550 16.050 798.450 ;
        RECT 7.950 796.950 10.050 797.550 ;
        RECT 13.950 796.950 16.050 797.550 ;
        RECT 17.100 795.600 18.300 802.950 ;
        RECT 23.100 801.150 24.900 802.950 ;
        RECT 17.100 794.100 19.500 795.600 ;
        RECT 15.000 791.100 16.800 792.900 ;
        RECT 14.700 783.000 16.500 789.600 ;
        RECT 17.700 783.600 19.500 794.100 ;
        RECT 22.800 783.000 24.600 795.600 ;
        RECT 41.700 789.600 42.900 802.950 ;
        RECT 50.550 801.450 51.450 809.550 ;
        RECT 55.950 808.950 58.050 809.550 ;
        RECT 59.100 810.300 63.300 811.200 ;
        RECT 74.700 810.300 75.900 812.400 ;
        RECT 77.100 813.300 78.900 818.400 ;
        RECT 80.100 814.200 81.900 819.000 ;
        RECT 83.100 813.300 84.900 818.400 ;
        RECT 77.100 811.950 84.900 813.300 ;
        RECT 95.700 811.200 97.500 818.400 ;
        RECT 100.800 812.400 102.600 819.000 ;
        RECT 116.100 812.400 117.900 818.400 ;
        RECT 95.700 810.300 99.900 811.200 ;
        RECT 56.250 805.050 58.050 806.850 ;
        RECT 59.100 805.050 60.300 810.300 ;
        RECT 74.700 809.400 78.300 810.300 ;
        RECT 62.100 805.050 63.900 806.850 ;
        RECT 74.100 805.050 75.900 806.850 ;
        RECT 77.100 805.050 78.300 809.400 ;
        RECT 80.100 805.050 81.900 806.850 ;
        RECT 95.100 805.050 96.900 806.850 ;
        RECT 98.700 805.050 99.900 810.300 ;
        RECT 109.950 807.450 112.050 811.050 ;
        RECT 116.700 810.300 117.900 812.400 ;
        RECT 119.100 813.300 120.900 818.400 ;
        RECT 122.100 814.200 123.900 819.000 ;
        RECT 125.100 813.300 126.900 818.400 ;
        RECT 137.100 815.400 138.900 818.400 ;
        RECT 140.100 815.400 141.900 819.000 ;
        RECT 119.100 811.950 126.900 813.300 ;
        RECT 116.700 809.400 120.300 810.300 ;
        RECT 107.550 807.000 112.050 807.450 ;
        RECT 100.950 805.050 102.750 806.850 ;
        RECT 107.550 806.550 111.450 807.000 ;
        RECT 55.950 802.950 58.050 805.050 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 76.950 802.950 79.050 805.050 ;
        RECT 79.950 802.950 82.050 805.050 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 50.550 800.550 54.450 801.450 ;
        RECT 53.550 799.050 54.450 800.550 ;
        RECT 53.550 797.550 58.050 799.050 ;
        RECT 54.000 796.950 58.050 797.550 ;
        RECT 59.100 789.600 60.300 802.950 ;
        RECT 77.100 795.600 78.300 802.950 ;
        RECT 83.100 801.150 84.900 802.950 ;
        RECT 77.100 794.100 79.500 795.600 ;
        RECT 75.000 791.100 76.800 792.900 ;
        RECT 38.100 783.000 39.900 789.600 ;
        RECT 41.100 783.600 42.900 789.600 ;
        RECT 44.100 783.000 45.900 789.600 ;
        RECT 56.100 783.000 57.900 789.600 ;
        RECT 59.100 783.600 60.900 789.600 ;
        RECT 62.100 783.000 63.900 789.600 ;
        RECT 74.700 783.000 76.500 789.600 ;
        RECT 77.700 783.600 79.500 794.100 ;
        RECT 82.800 783.000 84.600 795.600 ;
        RECT 98.700 789.600 99.900 802.950 ;
        RECT 107.550 802.050 108.450 806.550 ;
        RECT 116.100 805.050 117.900 806.850 ;
        RECT 119.100 805.050 120.300 809.400 ;
        RECT 122.100 805.050 123.900 806.850 ;
        RECT 137.700 805.050 138.900 815.400 ;
        RECT 155.100 812.400 156.900 818.400 ;
        RECT 155.700 810.300 156.900 812.400 ;
        RECT 158.100 813.300 159.900 818.400 ;
        RECT 161.100 814.200 162.900 819.000 ;
        RECT 164.100 813.300 165.900 818.400 ;
        RECT 179.100 815.400 180.900 819.000 ;
        RECT 182.100 815.400 183.900 818.400 ;
        RECT 194.100 815.400 195.900 818.400 ;
        RECT 197.100 815.400 198.900 819.000 ;
        RECT 158.100 811.950 165.900 813.300 ;
        RECT 155.700 809.400 159.300 810.300 ;
        RECT 155.100 805.050 156.900 806.850 ;
        RECT 158.100 805.050 159.300 809.400 ;
        RECT 161.100 805.050 162.900 806.850 ;
        RECT 182.100 805.050 183.300 815.400 ;
        RECT 194.700 805.050 195.900 815.400 ;
        RECT 210.000 812.400 211.800 819.000 ;
        RECT 214.500 813.600 216.300 818.400 ;
        RECT 217.500 815.400 219.300 819.000 ;
        RECT 233.700 815.400 235.500 819.000 ;
        RECT 236.700 813.600 238.500 818.400 ;
        RECT 214.500 812.400 219.600 813.600 ;
        RECT 211.950 810.450 214.050 811.200 ;
        RECT 206.550 809.550 214.050 810.450 ;
        RECT 206.550 807.450 207.450 809.550 ;
        RECT 211.950 809.100 214.050 809.550 ;
        RECT 203.550 806.550 207.450 807.450 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 181.950 802.950 184.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 103.950 800.550 108.450 802.050 ;
        RECT 103.950 799.950 108.000 800.550 ;
        RECT 119.100 795.600 120.300 802.950 ;
        RECT 125.100 801.150 126.900 802.950 ;
        RECT 119.100 794.100 121.500 795.600 ;
        RECT 117.000 791.100 118.800 792.900 ;
        RECT 95.100 783.000 96.900 789.600 ;
        RECT 98.100 783.600 99.900 789.600 ;
        RECT 101.100 783.000 102.900 789.600 ;
        RECT 116.700 783.000 118.500 789.600 ;
        RECT 119.700 783.600 121.500 794.100 ;
        RECT 124.800 783.000 126.600 795.600 ;
        RECT 137.700 789.600 138.900 802.950 ;
        RECT 140.100 801.150 141.900 802.950 ;
        RECT 158.100 795.600 159.300 802.950 ;
        RECT 164.100 801.150 165.900 802.950 ;
        RECT 179.100 801.150 180.900 802.950 ;
        RECT 158.100 794.100 160.500 795.600 ;
        RECT 156.000 791.100 157.800 792.900 ;
        RECT 137.100 783.600 138.900 789.600 ;
        RECT 140.100 783.000 141.900 789.600 ;
        RECT 155.700 783.000 157.500 789.600 ;
        RECT 158.700 783.600 160.500 794.100 ;
        RECT 163.800 783.000 165.600 795.600 ;
        RECT 182.100 789.600 183.300 802.950 ;
        RECT 194.700 789.600 195.900 802.950 ;
        RECT 197.100 801.150 198.900 802.950 ;
        RECT 203.550 802.050 204.450 806.550 ;
        RECT 209.100 805.050 210.900 806.850 ;
        RECT 215.250 805.050 217.050 806.850 ;
        RECT 218.700 805.050 219.600 812.400 ;
        RECT 233.400 812.400 238.500 813.600 ;
        RECT 241.200 812.400 243.000 819.000 ;
        RECT 257.100 813.000 258.900 818.400 ;
        RECT 260.100 813.900 261.900 819.000 ;
        RECT 263.100 817.500 270.900 818.400 ;
        RECT 263.100 813.000 264.900 817.500 ;
        RECT 233.400 805.050 234.300 812.400 ;
        RECT 257.100 812.100 264.900 813.000 ;
        RECT 266.100 812.400 267.900 816.600 ;
        RECT 269.100 812.400 270.900 817.500 ;
        RECT 281.100 812.400 282.900 818.400 ;
        RECT 241.950 810.450 244.050 811.050 ;
        RECT 247.950 810.450 250.050 811.050 ;
        RECT 266.400 810.900 267.300 812.400 ;
        RECT 241.950 809.550 250.050 810.450 ;
        RECT 241.950 808.950 244.050 809.550 ;
        RECT 247.950 808.950 250.050 809.550 ;
        RECT 262.950 809.700 267.300 810.900 ;
        RECT 281.700 810.300 282.900 812.400 ;
        RECT 284.100 813.300 285.900 818.400 ;
        RECT 287.100 814.200 288.900 819.000 ;
        RECT 290.100 813.300 291.900 818.400 ;
        RECT 284.100 811.950 291.900 813.300 ;
        RECT 305.100 813.300 306.900 818.400 ;
        RECT 308.100 814.200 309.900 819.000 ;
        RECT 311.100 813.300 312.900 818.400 ;
        RECT 305.100 811.950 312.900 813.300 ;
        RECT 314.100 812.400 315.900 818.400 ;
        RECT 314.100 810.300 315.300 812.400 ;
        RECT 326.700 811.200 328.500 818.400 ;
        RECT 331.800 812.400 333.600 819.000 ;
        RECT 349.500 812.400 351.300 819.000 ;
        RECT 354.000 812.400 355.800 818.400 ;
        RECT 358.500 812.400 360.300 819.000 ;
        RECT 371.100 812.400 372.900 818.400 ;
        RECT 326.700 810.300 330.900 811.200 ;
        RECT 235.950 805.050 237.750 806.850 ;
        RECT 242.100 805.050 243.900 806.850 ;
        RECT 260.250 805.050 262.050 806.850 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 217.950 802.950 220.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 262.950 805.050 264.000 809.700 ;
        RECT 281.700 809.400 285.300 810.300 ;
        RECT 265.950 805.050 267.750 806.850 ;
        RECT 281.100 805.050 282.900 806.850 ;
        RECT 284.100 805.050 285.300 809.400 ;
        RECT 311.700 809.400 315.300 810.300 ;
        RECT 292.950 807.450 297.000 808.050 ;
        RECT 300.000 807.450 304.050 808.050 ;
        RECT 287.100 805.050 288.900 806.850 ;
        RECT 292.950 805.950 297.450 807.450 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 203.550 800.550 208.050 802.050 ;
        RECT 212.250 801.150 214.050 802.950 ;
        RECT 204.000 799.950 208.050 800.550 ;
        RECT 218.700 795.600 219.600 802.950 ;
        RECT 233.400 795.600 234.300 802.950 ;
        RECT 238.950 801.150 240.750 802.950 ;
        RECT 257.100 801.150 258.900 802.950 ;
        RECT 241.950 798.450 244.050 798.750 ;
        RECT 247.950 798.450 250.050 799.050 ;
        RECT 241.950 797.550 250.050 798.450 ;
        RECT 241.950 796.650 244.050 797.550 ;
        RECT 247.950 796.950 250.050 797.550 ;
        RECT 209.100 794.700 216.900 795.600 ;
        RECT 179.100 783.000 180.900 789.600 ;
        RECT 182.100 783.600 183.900 789.600 ;
        RECT 194.100 783.600 195.900 789.600 ;
        RECT 197.100 783.000 198.900 789.600 ;
        RECT 209.100 783.600 210.900 794.700 ;
        RECT 212.100 783.000 213.900 793.800 ;
        RECT 215.100 783.600 216.900 794.700 ;
        RECT 218.100 783.600 219.900 795.600 ;
        RECT 233.100 783.600 234.900 795.600 ;
        RECT 236.100 794.700 243.900 795.600 ;
        RECT 236.100 783.600 237.900 794.700 ;
        RECT 239.100 783.000 240.900 793.800 ;
        RECT 242.100 783.600 243.900 794.700 ;
        RECT 247.950 795.450 250.050 795.900 ;
        RECT 253.950 795.450 256.050 796.050 ;
        RECT 262.950 795.600 264.000 802.950 ;
        RECT 268.950 801.150 270.750 802.950 ;
        RECT 271.950 798.450 274.050 799.050 ;
        RECT 280.950 798.450 283.050 799.050 ;
        RECT 271.950 797.550 283.050 798.450 ;
        RECT 271.950 796.950 274.050 797.550 ;
        RECT 280.950 796.950 283.050 797.550 ;
        RECT 284.100 795.600 285.300 802.950 ;
        RECT 290.100 801.150 291.900 802.950 ;
        RECT 296.550 802.050 297.450 805.950 ;
        RECT 292.950 800.550 297.450 802.050 ;
        RECT 299.550 805.950 304.050 807.450 ;
        RECT 299.550 801.450 300.450 805.950 ;
        RECT 308.100 805.050 309.900 806.850 ;
        RECT 311.700 805.050 312.900 809.400 ;
        RECT 314.100 805.050 315.900 806.850 ;
        RECT 326.100 805.050 327.900 806.850 ;
        RECT 329.700 805.050 330.900 810.300 ;
        RECT 331.950 805.050 333.750 806.850 ;
        RECT 347.100 805.050 348.900 806.850 ;
        RECT 353.700 805.050 354.900 812.400 ;
        RECT 371.700 810.300 372.900 812.400 ;
        RECT 374.100 813.300 375.900 818.400 ;
        RECT 377.100 814.200 378.900 819.000 ;
        RECT 380.100 813.300 381.900 818.400 ;
        RECT 374.100 811.950 381.900 813.300 ;
        RECT 395.100 812.400 396.900 818.400 ;
        RECT 395.700 810.300 396.900 812.400 ;
        RECT 398.100 813.300 399.900 818.400 ;
        RECT 401.100 814.200 402.900 819.000 ;
        RECT 404.100 813.300 405.900 818.400 ;
        RECT 398.100 811.950 405.900 813.300 ;
        RECT 419.100 810.600 420.900 818.400 ;
        RECT 423.600 812.400 425.400 819.000 ;
        RECT 426.600 814.200 428.400 818.400 ;
        RECT 426.600 812.400 429.300 814.200 ;
        RECT 425.700 810.600 427.500 811.500 ;
        RECT 371.700 809.400 375.300 810.300 ;
        RECT 395.700 809.400 399.300 810.300 ;
        RECT 419.100 809.700 427.500 810.600 ;
        RECT 358.950 805.050 360.750 806.850 ;
        RECT 371.100 805.050 372.900 806.850 ;
        RECT 374.100 805.050 375.300 809.400 ;
        RECT 382.950 807.450 385.050 808.050 ;
        RECT 388.950 807.450 391.050 808.050 ;
        RECT 377.100 805.050 378.900 806.850 ;
        RECT 382.950 806.550 391.050 807.450 ;
        RECT 382.950 805.950 385.050 806.550 ;
        RECT 388.950 805.950 391.050 806.550 ;
        RECT 395.100 805.050 396.900 806.850 ;
        RECT 398.100 805.050 399.300 809.400 ;
        RECT 401.100 805.050 402.900 806.850 ;
        RECT 419.250 805.050 421.050 806.850 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 313.950 802.950 316.050 805.050 ;
        RECT 325.950 802.950 328.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 419.100 802.950 421.200 805.050 ;
        RECT 299.550 800.550 303.450 801.450 ;
        RECT 305.100 801.150 306.900 802.950 ;
        RECT 292.950 799.950 297.000 800.550 ;
        RECT 302.550 798.450 303.450 800.550 ;
        RECT 307.950 798.450 310.050 799.050 ;
        RECT 302.550 797.550 310.050 798.450 ;
        RECT 307.950 796.950 310.050 797.550 ;
        RECT 311.700 795.600 312.900 802.950 ;
        RECT 247.950 794.550 256.050 795.450 ;
        RECT 247.950 793.800 250.050 794.550 ;
        RECT 253.950 793.950 256.050 794.550 ;
        RECT 257.100 783.000 258.900 795.600 ;
        RECT 261.600 783.600 264.900 795.600 ;
        RECT 267.600 783.000 269.400 795.600 ;
        RECT 284.100 794.100 286.500 795.600 ;
        RECT 282.000 791.100 283.800 792.900 ;
        RECT 281.700 783.000 283.500 789.600 ;
        RECT 284.700 783.600 286.500 794.100 ;
        RECT 289.800 783.000 291.600 795.600 ;
        RECT 305.400 783.000 307.200 795.600 ;
        RECT 310.500 794.100 312.900 795.600 ;
        RECT 310.500 783.600 312.300 794.100 ;
        RECT 313.200 791.100 315.000 792.900 ;
        RECT 329.700 789.600 330.900 802.950 ;
        RECT 350.100 801.150 351.900 802.950 ;
        RECT 354.000 797.400 354.900 802.950 ;
        RECT 355.950 801.150 357.750 802.950 ;
        RECT 350.100 796.500 354.900 797.400 ;
        RECT 313.500 783.000 315.300 789.600 ;
        RECT 326.100 783.000 327.900 789.600 ;
        RECT 329.100 783.600 330.900 789.600 ;
        RECT 332.100 783.000 333.900 789.600 ;
        RECT 347.100 784.500 348.900 795.600 ;
        RECT 350.100 785.400 351.900 796.500 ;
        RECT 374.100 795.600 375.300 802.950 ;
        RECT 380.100 801.150 381.900 802.950 ;
        RECT 398.100 795.600 399.300 802.950 ;
        RECT 404.100 801.150 405.900 802.950 ;
        RECT 353.100 794.400 360.900 795.300 ;
        RECT 353.100 784.500 354.900 794.400 ;
        RECT 347.100 783.600 354.900 784.500 ;
        RECT 356.100 783.000 357.900 793.500 ;
        RECT 359.100 783.600 360.900 794.400 ;
        RECT 374.100 794.100 376.500 795.600 ;
        RECT 372.000 791.100 373.800 792.900 ;
        RECT 371.700 783.000 373.500 789.600 ;
        RECT 374.700 783.600 376.500 794.100 ;
        RECT 379.800 783.000 381.600 795.600 ;
        RECT 398.100 794.100 400.500 795.600 ;
        RECT 396.000 791.100 397.800 792.900 ;
        RECT 395.700 783.000 397.500 789.600 ;
        RECT 398.700 783.600 400.500 794.100 ;
        RECT 403.800 783.000 405.600 795.600 ;
        RECT 422.100 789.600 423.000 809.700 ;
        RECT 428.400 805.050 429.300 812.400 ;
        RECT 440.100 813.300 441.900 818.400 ;
        RECT 443.100 814.200 444.900 819.000 ;
        RECT 446.100 813.300 447.900 818.400 ;
        RECT 440.100 811.950 447.900 813.300 ;
        RECT 449.100 812.400 450.900 818.400 ;
        RECT 449.100 810.300 450.300 812.400 ;
        RECT 461.700 811.200 463.500 818.400 ;
        RECT 466.800 812.400 468.600 819.000 ;
        RECT 482.700 812.400 484.500 819.000 ;
        RECT 487.200 812.400 489.000 818.400 ;
        RECT 491.700 812.400 493.500 819.000 ;
        RECT 509.100 813.300 510.900 818.400 ;
        RECT 512.100 814.200 513.900 819.000 ;
        RECT 515.100 813.300 516.900 818.400 ;
        RECT 461.700 810.300 465.900 811.200 ;
        RECT 484.950 810.450 487.050 811.050 ;
        RECT 446.700 809.400 450.300 810.300 ;
        RECT 443.100 805.050 444.900 806.850 ;
        RECT 446.700 805.050 447.900 809.400 ;
        RECT 449.100 805.050 450.900 806.850 ;
        RECT 461.100 805.050 462.900 806.850 ;
        RECT 464.700 805.050 465.900 810.300 ;
        RECT 473.550 809.550 487.050 810.450 ;
        RECT 466.950 805.050 468.750 806.850 ;
        RECT 424.500 802.950 426.600 805.050 ;
        RECT 427.800 802.950 429.900 805.050 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 445.950 802.950 448.050 805.050 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 424.200 801.150 426.000 802.950 ;
        RECT 428.400 795.600 429.300 802.950 ;
        RECT 440.100 801.150 441.900 802.950 ;
        RECT 446.700 795.600 447.900 802.950 ;
        RECT 419.100 783.000 420.900 789.600 ;
        RECT 422.100 783.600 423.900 789.600 ;
        RECT 425.100 783.000 426.900 795.000 ;
        RECT 428.100 783.600 429.900 795.600 ;
        RECT 440.400 783.000 442.200 795.600 ;
        RECT 445.500 794.100 447.900 795.600 ;
        RECT 445.500 783.600 447.300 794.100 ;
        RECT 448.200 791.100 450.000 792.900 ;
        RECT 464.700 789.600 465.900 802.950 ;
        RECT 473.550 802.050 474.450 809.550 ;
        RECT 484.950 808.950 487.050 809.550 ;
        RECT 482.250 805.050 484.050 806.850 ;
        RECT 488.100 805.050 489.300 812.400 ;
        RECT 509.100 811.950 516.900 813.300 ;
        RECT 518.100 812.400 519.900 818.400 ;
        RECT 535.500 812.400 537.300 819.000 ;
        RECT 540.000 812.400 541.800 818.400 ;
        RECT 544.500 812.400 546.300 819.000 ;
        RECT 518.100 810.300 519.300 812.400 ;
        RECT 515.700 809.400 519.300 810.300 ;
        RECT 520.950 810.450 523.050 811.050 ;
        RECT 532.950 810.450 535.050 811.200 ;
        RECT 520.950 809.550 535.050 810.450 ;
        RECT 504.000 807.450 508.050 808.050 ;
        RECT 494.100 805.050 495.900 806.850 ;
        RECT 503.550 805.950 508.050 807.450 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 469.950 800.550 474.450 802.050 ;
        RECT 485.250 801.150 487.050 802.950 ;
        RECT 469.950 799.950 474.000 800.550 ;
        RECT 488.100 797.400 489.000 802.950 ;
        RECT 491.100 801.150 492.900 802.950 ;
        RECT 503.550 802.050 504.450 805.950 ;
        RECT 512.100 805.050 513.900 806.850 ;
        RECT 515.700 805.050 516.900 809.400 ;
        RECT 520.950 808.950 523.050 809.550 ;
        RECT 532.950 809.100 535.050 809.550 ;
        RECT 529.950 807.450 532.050 808.050 ;
        RECT 518.100 805.050 519.900 806.850 ;
        RECT 524.550 806.550 532.050 807.450 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 503.550 800.550 508.050 802.050 ;
        RECT 509.100 801.150 510.900 802.950 ;
        RECT 504.000 799.950 508.050 800.550 ;
        RECT 488.100 796.500 492.900 797.400 ;
        RECT 508.950 796.950 514.050 799.050 ;
        RECT 482.100 794.400 489.900 795.300 ;
        RECT 448.500 783.000 450.300 789.600 ;
        RECT 461.100 783.000 462.900 789.600 ;
        RECT 464.100 783.600 465.900 789.600 ;
        RECT 467.100 783.000 468.900 789.600 ;
        RECT 482.100 783.600 483.900 794.400 ;
        RECT 485.100 783.000 486.900 793.500 ;
        RECT 488.100 784.500 489.900 794.400 ;
        RECT 491.100 785.400 492.900 796.500 ;
        RECT 515.700 795.600 516.900 802.950 ;
        RECT 524.550 802.050 525.450 806.550 ;
        RECT 529.950 805.950 532.050 806.550 ;
        RECT 533.100 805.050 534.900 806.850 ;
        RECT 539.700 805.050 540.900 812.400 ;
        RECT 557.700 811.200 559.500 818.400 ;
        RECT 562.800 812.400 564.600 819.000 ;
        RECT 575.100 815.400 576.900 818.400 ;
        RECT 578.100 815.400 579.900 819.000 ;
        RECT 557.700 810.300 561.900 811.200 ;
        RECT 544.950 805.050 546.750 806.850 ;
        RECT 557.100 805.050 558.900 806.850 ;
        RECT 560.700 805.050 561.900 810.300 ;
        RECT 562.950 805.050 564.750 806.850 ;
        RECT 575.700 805.050 576.900 815.400 ;
        RECT 594.000 812.400 595.800 819.000 ;
        RECT 598.500 813.600 600.300 818.400 ;
        RECT 601.500 815.400 603.300 819.000 ;
        RECT 598.500 812.400 603.600 813.600 ;
        RECT 593.100 805.050 594.900 806.850 ;
        RECT 599.250 805.050 601.050 806.850 ;
        RECT 602.700 805.050 603.600 812.400 ;
        RECT 617.700 811.200 619.500 818.400 ;
        RECT 622.800 812.400 624.600 819.000 ;
        RECT 640.500 812.400 642.300 819.000 ;
        RECT 645.000 812.400 646.800 818.400 ;
        RECT 649.500 812.400 651.300 819.000 ;
        RECT 662.100 815.400 663.900 819.000 ;
        RECT 665.100 815.400 666.900 818.400 ;
        RECT 610.950 808.950 613.050 811.050 ;
        RECT 617.700 810.300 621.900 811.200 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 592.950 802.950 595.050 805.050 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 520.950 800.550 525.450 802.050 ;
        RECT 536.100 801.150 537.900 802.950 ;
        RECT 520.950 799.950 525.000 800.550 ;
        RECT 520.950 798.450 523.050 798.900 ;
        RECT 532.950 798.450 535.050 799.050 ;
        RECT 520.950 797.550 535.050 798.450 ;
        RECT 520.950 796.800 523.050 797.550 ;
        RECT 532.950 796.950 535.050 797.550 ;
        RECT 540.000 797.400 540.900 802.950 ;
        RECT 541.950 801.150 543.750 802.950 ;
        RECT 536.100 796.500 540.900 797.400 ;
        RECT 544.950 798.450 547.050 799.050 ;
        RECT 553.950 798.450 556.050 799.050 ;
        RECT 544.950 797.550 556.050 798.450 ;
        RECT 544.950 796.950 547.050 797.550 ;
        RECT 553.950 796.950 556.050 797.550 ;
        RECT 494.100 784.500 495.900 795.600 ;
        RECT 488.100 783.600 495.900 784.500 ;
        RECT 509.400 783.000 511.200 795.600 ;
        RECT 514.500 794.100 516.900 795.600 ;
        RECT 514.500 783.600 516.300 794.100 ;
        RECT 517.200 791.100 519.000 792.900 ;
        RECT 517.500 783.000 519.300 789.600 ;
        RECT 520.950 789.450 523.050 789.900 ;
        RECT 529.950 789.450 532.050 790.050 ;
        RECT 520.950 788.550 532.050 789.450 ;
        RECT 520.950 787.800 523.050 788.550 ;
        RECT 529.950 787.950 532.050 788.550 ;
        RECT 533.100 784.500 534.900 795.600 ;
        RECT 536.100 785.400 537.900 796.500 ;
        RECT 539.100 794.400 546.900 795.300 ;
        RECT 539.100 784.500 540.900 794.400 ;
        RECT 533.100 783.600 540.900 784.500 ;
        RECT 542.100 783.000 543.900 793.500 ;
        RECT 545.100 783.600 546.900 794.400 ;
        RECT 560.700 789.600 561.900 802.950 ;
        RECT 575.700 789.600 576.900 802.950 ;
        RECT 578.100 801.150 579.900 802.950 ;
        RECT 596.250 801.150 598.050 802.950 ;
        RECT 602.700 795.600 603.600 802.950 ;
        RECT 611.550 802.050 612.450 808.950 ;
        RECT 617.100 805.050 618.900 806.850 ;
        RECT 620.700 805.050 621.900 810.300 ;
        RECT 625.950 807.450 630.000 808.050 ;
        RECT 622.950 805.050 624.750 806.850 ;
        RECT 625.950 805.950 630.450 807.450 ;
        RECT 616.950 802.950 619.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 611.550 800.550 616.050 802.050 ;
        RECT 612.000 799.950 616.050 800.550 ;
        RECT 593.100 794.700 600.900 795.600 ;
        RECT 557.100 783.000 558.900 789.600 ;
        RECT 560.100 783.600 561.900 789.600 ;
        RECT 563.100 783.000 564.900 789.600 ;
        RECT 575.100 783.600 576.900 789.600 ;
        RECT 578.100 783.000 579.900 789.600 ;
        RECT 593.100 783.600 594.900 794.700 ;
        RECT 596.100 783.000 597.900 793.800 ;
        RECT 599.100 783.600 600.900 794.700 ;
        RECT 602.100 783.600 603.900 795.600 ;
        RECT 620.700 789.600 621.900 802.950 ;
        RECT 629.550 801.450 630.450 805.950 ;
        RECT 638.100 805.050 639.900 806.850 ;
        RECT 644.700 805.050 645.900 812.400 ;
        RECT 649.950 805.050 651.750 806.850 ;
        RECT 665.100 805.050 666.300 815.400 ;
        RECT 677.400 812.400 679.200 819.000 ;
        RECT 682.500 811.200 684.300 818.400 ;
        RECT 698.400 812.400 700.200 819.000 ;
        RECT 703.500 811.200 705.300 818.400 ;
        RECT 716.700 812.400 718.500 819.000 ;
        RECT 721.200 812.400 723.000 818.400 ;
        RECT 725.700 812.400 727.500 819.000 ;
        RECT 740.100 815.400 741.900 818.400 ;
        RECT 743.100 815.400 744.900 819.000 ;
        RECT 680.100 810.300 684.300 811.200 ;
        RECT 701.100 810.300 705.300 811.200 ;
        RECT 672.000 807.450 676.050 808.050 ;
        RECT 671.550 805.950 676.050 807.450 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 640.950 802.950 643.050 805.050 ;
        RECT 643.950 802.950 646.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 634.950 801.450 637.050 802.050 ;
        RECT 629.550 800.550 637.050 801.450 ;
        RECT 641.100 801.150 642.900 802.950 ;
        RECT 634.950 799.950 637.050 800.550 ;
        RECT 628.950 798.450 631.050 798.900 ;
        RECT 637.950 798.450 640.050 799.050 ;
        RECT 628.950 797.550 640.050 798.450 ;
        RECT 628.950 796.800 631.050 797.550 ;
        RECT 637.950 796.950 640.050 797.550 ;
        RECT 645.000 797.400 645.900 802.950 ;
        RECT 646.950 801.150 648.750 802.950 ;
        RECT 662.100 801.150 663.900 802.950 ;
        RECT 641.100 796.500 645.900 797.400 ;
        RECT 617.100 783.000 618.900 789.600 ;
        RECT 620.100 783.600 621.900 789.600 ;
        RECT 623.100 783.000 624.900 789.600 ;
        RECT 638.100 784.500 639.900 795.600 ;
        RECT 641.100 785.400 642.900 796.500 ;
        RECT 644.100 794.400 651.900 795.300 ;
        RECT 644.100 784.500 645.900 794.400 ;
        RECT 638.100 783.600 645.900 784.500 ;
        RECT 647.100 783.000 648.900 793.500 ;
        RECT 650.100 783.600 651.900 794.400 ;
        RECT 665.100 789.600 666.300 802.950 ;
        RECT 671.550 802.050 672.450 805.950 ;
        RECT 677.250 805.050 679.050 806.850 ;
        RECT 680.100 805.050 681.300 810.300 ;
        RECT 683.100 805.050 684.900 806.850 ;
        RECT 698.250 805.050 700.050 806.850 ;
        RECT 701.100 805.050 702.300 810.300 ;
        RECT 704.100 805.050 705.900 806.850 ;
        RECT 716.250 805.050 718.050 806.850 ;
        RECT 722.100 805.050 723.300 812.400 ;
        RECT 728.100 805.050 729.900 806.850 ;
        RECT 740.700 805.050 741.900 815.400 ;
        RECT 755.400 812.400 757.200 819.000 ;
        RECT 760.500 811.200 762.300 818.400 ;
        RECT 776.100 812.400 777.900 818.400 ;
        RECT 742.950 810.450 745.050 811.050 ;
        RECT 751.950 810.450 754.050 811.050 ;
        RECT 742.950 809.550 754.050 810.450 ;
        RECT 742.950 808.950 745.050 809.550 ;
        RECT 751.950 808.950 754.050 809.550 ;
        RECT 758.100 810.300 762.300 811.200 ;
        RECT 776.700 810.300 777.900 812.400 ;
        RECT 779.100 813.300 780.900 818.400 ;
        RECT 782.100 814.200 783.900 819.000 ;
        RECT 785.100 813.300 786.900 818.400 ;
        RECT 779.100 811.950 786.900 813.300 ;
        RECT 800.100 813.300 801.900 818.400 ;
        RECT 803.100 814.200 804.900 819.000 ;
        RECT 806.100 813.300 807.900 818.400 ;
        RECT 800.100 811.950 807.900 813.300 ;
        RECT 809.100 812.400 810.900 818.400 ;
        RECT 821.100 815.400 822.900 819.000 ;
        RECT 824.100 815.400 825.900 818.400 ;
        RECT 809.100 810.300 810.300 812.400 ;
        RECT 755.250 805.050 757.050 806.850 ;
        RECT 758.100 805.050 759.300 810.300 ;
        RECT 776.700 809.400 780.300 810.300 ;
        RECT 761.100 805.050 762.900 806.850 ;
        RECT 776.100 805.050 777.900 806.850 ;
        RECT 779.100 805.050 780.300 809.400 ;
        RECT 806.700 809.400 810.300 810.300 ;
        RECT 795.000 807.450 799.050 808.050 ;
        RECT 782.100 805.050 783.900 806.850 ;
        RECT 794.550 805.950 799.050 807.450 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 667.950 800.550 672.450 802.050 ;
        RECT 667.950 799.950 672.000 800.550 ;
        RECT 680.100 789.600 681.300 802.950 ;
        RECT 685.950 795.450 688.050 796.050 ;
        RECT 694.950 795.450 697.050 796.050 ;
        RECT 685.950 794.550 697.050 795.450 ;
        RECT 685.950 793.950 688.050 794.550 ;
        RECT 694.950 793.950 697.050 794.550 ;
        RECT 701.100 789.600 702.300 802.950 ;
        RECT 719.250 801.150 721.050 802.950 ;
        RECT 722.100 797.400 723.000 802.950 ;
        RECT 725.100 801.150 726.900 802.950 ;
        RECT 722.100 796.500 726.900 797.400 ;
        RECT 716.100 794.400 723.900 795.300 ;
        RECT 662.100 783.000 663.900 789.600 ;
        RECT 665.100 783.600 666.900 789.600 ;
        RECT 677.100 783.000 678.900 789.600 ;
        RECT 680.100 783.600 681.900 789.600 ;
        RECT 683.100 783.000 684.900 789.600 ;
        RECT 698.100 783.000 699.900 789.600 ;
        RECT 701.100 783.600 702.900 789.600 ;
        RECT 704.100 783.000 705.900 789.600 ;
        RECT 716.100 783.600 717.900 794.400 ;
        RECT 719.100 783.000 720.900 793.500 ;
        RECT 722.100 784.500 723.900 794.400 ;
        RECT 725.100 785.400 726.900 796.500 ;
        RECT 728.100 784.500 729.900 795.600 ;
        RECT 740.700 789.600 741.900 802.950 ;
        RECT 743.100 801.150 744.900 802.950 ;
        RECT 758.100 789.600 759.300 802.950 ;
        RECT 779.100 795.600 780.300 802.950 ;
        RECT 785.100 801.150 786.900 802.950 ;
        RECT 790.950 802.050 793.050 805.050 ;
        RECT 787.950 801.000 793.050 802.050 ;
        RECT 794.550 802.050 795.450 805.950 ;
        RECT 803.100 805.050 804.900 806.850 ;
        RECT 806.700 805.050 807.900 809.400 ;
        RECT 816.000 807.450 820.050 808.050 ;
        RECT 809.100 805.050 810.900 806.850 ;
        RECT 815.550 805.950 820.050 807.450 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 787.950 800.550 792.450 801.000 ;
        RECT 794.550 800.550 799.050 802.050 ;
        RECT 800.100 801.150 801.900 802.950 ;
        RECT 787.950 799.950 792.000 800.550 ;
        RECT 795.000 799.950 799.050 800.550 ;
        RECT 806.700 795.600 807.900 802.950 ;
        RECT 815.550 802.050 816.450 805.950 ;
        RECT 824.100 805.050 825.300 815.400 ;
        RECT 839.100 809.400 840.900 819.000 ;
        RECT 845.700 810.000 847.500 818.400 ;
        RECT 865.500 810.000 867.300 818.400 ;
        RECT 845.700 808.800 849.000 810.000 ;
        RECT 839.100 805.050 840.900 806.850 ;
        RECT 845.100 805.050 846.900 806.850 ;
        RECT 848.100 805.050 849.000 808.800 ;
        RECT 864.000 808.800 867.300 810.000 ;
        RECT 872.100 809.400 873.900 819.000 ;
        RECT 888.000 812.400 889.800 819.000 ;
        RECT 892.500 813.600 894.300 818.400 ;
        RECT 895.500 815.400 897.300 819.000 ;
        RECT 911.100 815.400 912.900 819.000 ;
        RECT 914.100 815.400 915.900 818.400 ;
        RECT 917.100 815.400 918.900 819.000 ;
        RECT 892.500 812.400 897.600 813.600 ;
        RECT 864.000 805.050 864.900 808.800 ;
        RECT 874.950 807.450 879.000 808.050 ;
        RECT 874.950 807.000 879.450 807.450 ;
        RECT 866.100 805.050 867.900 806.850 ;
        RECT 872.100 805.050 873.900 806.850 ;
        RECT 874.950 805.950 880.050 807.000 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 841.950 802.950 844.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 865.950 802.950 868.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 811.950 800.550 816.450 802.050 ;
        RECT 821.100 801.150 822.900 802.950 ;
        RECT 811.950 799.950 816.000 800.550 ;
        RECT 779.100 794.100 781.500 795.600 ;
        RECT 777.000 791.100 778.800 792.900 ;
        RECT 722.100 783.600 729.900 784.500 ;
        RECT 740.100 783.600 741.900 789.600 ;
        RECT 743.100 783.000 744.900 789.600 ;
        RECT 755.100 783.000 756.900 789.600 ;
        RECT 758.100 783.600 759.900 789.600 ;
        RECT 761.100 783.000 762.900 789.600 ;
        RECT 776.700 783.000 778.500 789.600 ;
        RECT 779.700 783.600 781.500 794.100 ;
        RECT 784.800 783.000 786.600 795.600 ;
        RECT 800.400 783.000 802.200 795.600 ;
        RECT 805.500 794.100 807.900 795.600 ;
        RECT 805.500 783.600 807.300 794.100 ;
        RECT 808.200 791.100 810.000 792.900 ;
        RECT 824.100 789.600 825.300 802.950 ;
        RECT 842.100 801.150 843.900 802.950 ;
        RECT 848.100 790.800 849.000 802.950 ;
        RECT 842.400 789.900 849.000 790.800 ;
        RECT 842.400 789.600 843.900 789.900 ;
        RECT 808.500 783.000 810.300 789.600 ;
        RECT 821.100 783.000 822.900 789.600 ;
        RECT 824.100 783.600 825.900 789.600 ;
        RECT 839.100 783.000 840.900 789.600 ;
        RECT 842.100 783.600 843.900 789.600 ;
        RECT 848.100 789.600 849.000 789.900 ;
        RECT 864.000 790.800 864.900 802.950 ;
        RECT 869.100 801.150 870.900 802.950 ;
        RECT 877.950 802.800 880.050 805.950 ;
        RECT 887.100 805.050 888.900 806.850 ;
        RECT 893.250 805.050 895.050 806.850 ;
        RECT 896.700 805.050 897.600 812.400 ;
        RECT 914.700 805.050 915.600 815.400 ;
        RECT 916.950 810.450 919.050 811.050 ;
        RECT 928.950 810.450 931.050 811.050 ;
        RECT 916.950 809.550 931.050 810.450 ;
        RECT 916.950 808.950 919.050 809.550 ;
        RECT 928.950 808.950 931.050 809.550 ;
        RECT 886.950 802.950 889.050 805.050 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 895.950 802.950 898.050 805.050 ;
        RECT 910.950 802.950 913.050 805.050 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 890.250 801.150 892.050 802.950 ;
        RECT 896.700 795.600 897.600 802.950 ;
        RECT 911.100 801.150 912.900 802.950 ;
        RECT 914.700 795.600 915.600 802.950 ;
        RECT 916.950 801.150 918.750 802.950 ;
        RECT 887.100 794.700 894.900 795.600 ;
        RECT 864.000 789.900 870.600 790.800 ;
        RECT 864.000 789.600 864.900 789.900 ;
        RECT 845.100 783.000 846.900 789.000 ;
        RECT 848.100 783.600 849.900 789.600 ;
        RECT 863.100 783.600 864.900 789.600 ;
        RECT 869.100 789.600 870.600 789.900 ;
        RECT 866.100 783.000 867.900 789.000 ;
        RECT 869.100 783.600 870.900 789.600 ;
        RECT 872.100 783.000 873.900 789.600 ;
        RECT 887.100 783.600 888.900 794.700 ;
        RECT 890.100 783.000 891.900 793.800 ;
        RECT 893.100 783.600 894.900 794.700 ;
        RECT 896.100 783.600 897.900 795.600 ;
        RECT 912.000 794.400 915.600 795.600 ;
        RECT 912.000 783.600 913.800 794.400 ;
        RECT 917.100 783.000 918.900 795.600 ;
        RECT 14.100 773.400 15.900 780.000 ;
        RECT 17.100 773.400 18.900 779.400 ;
        RECT 20.100 773.400 21.900 780.000 ;
        RECT 32.100 773.400 33.900 779.400 ;
        RECT 35.100 774.000 36.900 780.000 ;
        RECT 17.100 760.050 18.300 773.400 ;
        RECT 33.000 773.100 33.900 773.400 ;
        RECT 38.100 773.400 39.900 779.400 ;
        RECT 41.100 773.400 42.900 780.000 ;
        RECT 38.100 773.100 39.600 773.400 ;
        RECT 33.000 772.200 39.600 773.100 ;
        RECT 33.000 760.050 33.900 772.200 ;
        RECT 53.100 768.300 54.900 779.400 ;
        RECT 56.100 769.500 57.900 780.000 ;
        RECT 53.100 767.400 57.600 768.300 ;
        RECT 60.600 767.400 62.400 779.400 ;
        RECT 65.100 769.500 66.900 780.000 ;
        RECT 68.100 768.600 69.900 779.400 ;
        RECT 55.500 765.300 57.600 767.400 ;
        RECT 61.200 766.050 62.400 767.400 ;
        RECT 65.100 767.400 69.900 768.600 ;
        RECT 80.100 778.500 87.900 779.400 ;
        RECT 80.100 767.400 81.900 778.500 ;
        RECT 65.100 766.500 67.200 767.400 ;
        RECT 83.100 766.500 84.900 777.600 ;
        RECT 86.100 768.600 87.900 778.500 ;
        RECT 89.100 769.500 90.900 780.000 ;
        RECT 92.100 768.600 93.900 779.400 ;
        RECT 108.600 768.900 110.400 779.400 ;
        RECT 86.100 767.700 93.900 768.600 ;
        RECT 108.000 767.400 110.400 768.900 ;
        RECT 111.600 767.400 113.400 780.000 ;
        RECT 116.100 767.400 117.900 779.400 ;
        RECT 131.700 773.400 133.500 780.000 ;
        RECT 132.000 770.100 133.800 771.900 ;
        RECT 134.700 768.900 136.500 779.400 ;
        RECT 61.200 765.000 62.700 766.050 ;
        RECT 83.100 765.600 87.900 766.500 ;
        RECT 58.800 763.500 60.900 763.800 ;
        RECT 38.100 760.050 39.900 761.850 ;
        RECT 57.000 761.700 60.900 763.500 ;
        RECT 61.800 763.050 62.700 765.000 ;
        RECT 61.800 760.950 63.900 763.050 ;
        RECT 61.800 760.800 63.300 760.950 ;
        RECT 58.200 760.050 60.000 760.500 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 53.100 758.700 60.000 760.050 ;
        RECT 60.900 759.900 63.300 760.800 ;
        RECT 67.800 760.050 69.600 761.850 ;
        RECT 83.100 760.050 84.900 761.850 ;
        RECT 87.000 760.050 87.900 765.600 ;
        RECT 88.950 760.050 90.750 761.850 ;
        RECT 108.000 760.050 109.200 767.400 ;
        RECT 116.700 765.900 117.900 767.400 ;
        RECT 110.100 764.700 117.900 765.900 ;
        RECT 134.100 767.400 136.500 768.900 ;
        RECT 139.800 767.400 141.600 780.000 ;
        RECT 142.950 768.450 145.050 772.050 ;
        RECT 148.950 768.450 151.050 769.050 ;
        RECT 142.950 768.000 151.050 768.450 ;
        RECT 143.550 767.550 151.050 768.000 ;
        RECT 110.100 764.100 111.900 764.700 ;
        RECT 53.100 757.950 55.200 758.700 ;
        RECT 14.250 756.150 16.050 757.950 ;
        RECT 17.100 752.700 18.300 757.950 ;
        RECT 20.100 756.150 21.900 757.950 ;
        RECT 33.000 754.200 33.900 757.950 ;
        RECT 35.100 756.150 36.900 757.950 ;
        RECT 41.100 756.150 42.900 757.950 ;
        RECT 46.950 754.950 49.050 757.050 ;
        RECT 53.400 756.150 55.200 757.950 ;
        RECT 58.200 755.400 60.000 757.200 ;
        RECT 33.000 753.000 36.300 754.200 ;
        RECT 17.100 751.800 21.300 752.700 ;
        RECT 14.400 744.000 16.200 750.600 ;
        RECT 19.500 744.600 21.300 751.800 ;
        RECT 34.500 744.600 36.300 753.000 ;
        RECT 41.100 744.000 42.900 753.600 ;
        RECT 47.550 751.050 48.450 754.950 ;
        RECT 57.900 753.300 60.000 755.400 ;
        RECT 53.700 752.400 60.000 753.300 ;
        RECT 60.900 754.200 62.100 759.900 ;
        RECT 63.300 757.200 65.100 759.000 ;
        RECT 67.800 757.950 69.900 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 91.950 757.950 94.050 760.050 ;
        RECT 107.100 757.950 109.200 760.050 ;
        RECT 63.000 755.100 65.100 757.200 ;
        RECT 80.100 756.150 81.900 757.950 ;
        RECT 47.550 749.550 52.050 751.050 ;
        RECT 53.700 750.600 54.900 752.400 ;
        RECT 60.900 752.100 63.900 754.200 ;
        RECT 60.900 750.600 62.100 752.100 ;
        RECT 65.100 751.500 67.200 752.700 ;
        RECT 65.100 750.600 69.900 751.500 ;
        RECT 86.700 750.600 87.900 757.950 ;
        RECT 91.950 756.150 93.750 757.950 ;
        RECT 88.950 753.450 91.050 754.050 ;
        RECT 100.950 753.450 103.050 754.050 ;
        RECT 88.950 752.550 103.050 753.450 ;
        RECT 88.950 751.950 91.050 752.550 ;
        RECT 100.950 751.950 103.050 752.550 ;
        RECT 107.100 750.600 108.000 757.950 ;
        RECT 110.400 753.600 111.300 764.100 ;
        RECT 112.200 760.050 114.000 761.850 ;
        RECT 134.100 760.050 135.300 767.400 ;
        RECT 148.950 766.950 151.050 767.550 ;
        RECT 152.100 767.400 153.900 779.400 ;
        RECT 155.100 768.300 156.900 779.400 ;
        RECT 158.100 769.200 159.900 780.000 ;
        RECT 161.100 768.300 162.900 779.400 ;
        RECT 176.100 773.400 177.900 779.400 ;
        RECT 179.100 773.400 180.900 780.000 ;
        RECT 194.100 773.400 195.900 779.400 ;
        RECT 197.100 773.400 198.900 780.000 ;
        RECT 209.700 773.400 211.500 780.000 ;
        RECT 155.100 767.400 162.900 768.300 ;
        RECT 140.100 760.050 141.900 761.850 ;
        RECT 152.400 760.050 153.300 767.400 ;
        RECT 160.950 765.450 163.050 766.050 ;
        RECT 166.950 765.450 169.050 766.050 ;
        RECT 160.950 764.550 169.050 765.450 ;
        RECT 160.950 763.950 163.050 764.550 ;
        RECT 166.950 763.950 169.050 764.550 ;
        RECT 157.950 760.050 159.750 761.850 ;
        RECT 176.700 760.050 177.900 773.400 ;
        RECT 179.100 760.050 180.900 761.850 ;
        RECT 194.700 760.050 195.900 773.400 ;
        RECT 210.000 770.100 211.800 771.900 ;
        RECT 212.700 768.900 214.500 779.400 ;
        RECT 212.100 767.400 214.500 768.900 ;
        RECT 217.800 767.400 219.600 780.000 ;
        RECT 230.700 773.400 232.500 780.000 ;
        RECT 231.000 770.100 232.800 771.900 ;
        RECT 233.700 768.900 235.500 779.400 ;
        RECT 233.100 767.400 235.500 768.900 ;
        RECT 238.800 767.400 240.600 780.000 ;
        RECT 254.400 767.400 256.200 780.000 ;
        RECT 259.500 768.900 261.300 779.400 ;
        RECT 262.500 773.400 264.300 780.000 ;
        RECT 262.200 770.100 264.000 771.900 ;
        RECT 259.500 767.400 261.900 768.900 ;
        RECT 275.100 767.400 276.900 779.400 ;
        RECT 278.100 768.300 279.900 779.400 ;
        RECT 281.100 769.200 282.900 780.000 ;
        RECT 284.100 768.300 285.900 779.400 ;
        RECT 299.100 773.400 300.900 780.000 ;
        RECT 302.100 773.400 303.900 779.400 ;
        RECT 278.100 767.400 285.900 768.300 ;
        RECT 199.950 762.450 202.050 766.050 ;
        RECT 199.950 762.000 204.450 762.450 ;
        RECT 197.100 760.050 198.900 761.850 ;
        RECT 200.550 761.550 204.450 762.000 ;
        RECT 112.500 757.950 114.600 760.050 ;
        RECT 115.800 757.950 117.900 760.050 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 133.950 757.950 136.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 154.950 757.950 157.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 115.800 756.150 117.600 757.950 ;
        RECT 131.100 756.150 132.900 757.950 ;
        RECT 109.200 752.700 111.300 753.600 ;
        RECT 109.200 751.800 114.600 752.700 ;
        RECT 48.000 748.950 52.050 749.550 ;
        RECT 53.100 744.600 54.900 750.600 ;
        RECT 56.100 744.000 57.900 749.700 ;
        RECT 60.600 744.600 62.400 750.600 ;
        RECT 65.100 744.000 66.900 749.700 ;
        RECT 68.100 744.600 69.900 750.600 ;
        RECT 82.500 744.000 84.300 750.600 ;
        RECT 87.000 744.600 88.800 750.600 ;
        RECT 91.500 744.000 93.300 750.600 ;
        RECT 107.100 744.600 108.900 750.600 ;
        RECT 110.100 744.000 111.900 750.000 ;
        RECT 113.700 747.600 114.600 751.800 ;
        RECT 115.950 750.450 118.050 754.050 ;
        RECT 134.100 753.600 135.300 757.950 ;
        RECT 137.100 756.150 138.900 757.950 ;
        RECT 131.700 752.700 135.300 753.600 ;
        RECT 124.950 750.450 127.050 751.050 ;
        RECT 131.700 750.600 132.900 752.700 ;
        RECT 115.950 750.000 127.050 750.450 ;
        RECT 116.550 749.550 127.050 750.000 ;
        RECT 124.950 748.950 127.050 749.550 ;
        RECT 113.100 744.600 114.900 747.600 ;
        RECT 116.100 744.600 117.900 747.600 ;
        RECT 131.100 744.600 132.900 750.600 ;
        RECT 134.100 749.700 141.900 751.050 ;
        RECT 134.100 744.600 135.900 749.700 ;
        RECT 116.700 744.000 117.900 744.600 ;
        RECT 137.100 744.000 138.900 748.800 ;
        RECT 140.100 744.600 141.900 749.700 ;
        RECT 152.400 750.600 153.300 757.950 ;
        RECT 154.950 756.150 156.750 757.950 ;
        RECT 161.100 756.150 162.900 757.950 ;
        RECT 152.400 749.400 157.500 750.600 ;
        RECT 152.700 744.000 154.500 747.600 ;
        RECT 155.700 744.600 157.500 749.400 ;
        RECT 160.200 744.000 162.000 750.600 ;
        RECT 176.700 747.600 177.900 757.950 ;
        RECT 194.700 747.600 195.900 757.950 ;
        RECT 203.550 757.050 204.450 761.550 ;
        RECT 212.100 760.050 213.300 767.400 ;
        RECT 218.100 760.050 219.900 761.850 ;
        RECT 233.100 760.050 234.300 767.400 ;
        RECT 235.950 765.450 238.050 766.050 ;
        RECT 256.950 765.450 259.050 766.050 ;
        RECT 235.950 764.550 259.050 765.450 ;
        RECT 235.950 763.950 238.050 764.550 ;
        RECT 256.950 763.950 259.050 764.550 ;
        RECT 239.100 760.050 240.900 761.850 ;
        RECT 254.100 760.050 255.900 761.850 ;
        RECT 260.700 760.050 261.900 767.400 ;
        RECT 271.950 762.450 274.050 766.050 ;
        RECT 269.550 762.000 274.050 762.450 ;
        RECT 269.550 761.550 273.450 762.000 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 253.950 757.950 256.050 760.050 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 203.550 755.550 208.050 757.050 ;
        RECT 209.100 756.150 210.900 757.950 ;
        RECT 204.000 754.950 208.050 755.550 ;
        RECT 212.100 753.600 213.300 757.950 ;
        RECT 215.100 756.150 216.900 757.950 ;
        RECT 230.100 756.150 231.900 757.950 ;
        RECT 233.100 753.600 234.300 757.950 ;
        RECT 236.100 756.150 237.900 757.950 ;
        RECT 257.100 756.150 258.900 757.950 ;
        RECT 209.700 752.700 213.300 753.600 ;
        RECT 230.700 752.700 234.300 753.600 ;
        RECT 260.700 753.600 261.900 757.950 ;
        RECT 263.100 756.150 264.900 757.950 ;
        RECT 269.550 757.050 270.450 761.550 ;
        RECT 275.400 760.050 276.300 767.400 ;
        RECT 298.950 765.450 301.050 766.050 ;
        RECT 293.550 764.550 301.050 765.450 ;
        RECT 280.950 760.050 282.750 761.850 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 269.550 755.550 274.050 757.050 ;
        RECT 270.000 754.950 274.050 755.550 ;
        RECT 260.700 752.700 264.300 753.600 ;
        RECT 209.700 750.600 210.900 752.700 ;
        RECT 176.100 744.600 177.900 747.600 ;
        RECT 179.100 744.000 180.900 747.600 ;
        RECT 194.100 744.600 195.900 747.600 ;
        RECT 197.100 744.000 198.900 747.600 ;
        RECT 209.100 744.600 210.900 750.600 ;
        RECT 212.100 749.700 219.900 751.050 ;
        RECT 230.700 750.600 231.900 752.700 ;
        RECT 212.100 744.600 213.900 749.700 ;
        RECT 215.100 744.000 216.900 748.800 ;
        RECT 218.100 744.600 219.900 749.700 ;
        RECT 230.100 744.600 231.900 750.600 ;
        RECT 233.100 749.700 240.900 751.050 ;
        RECT 233.100 744.600 234.900 749.700 ;
        RECT 236.100 744.000 237.900 748.800 ;
        RECT 239.100 744.600 240.900 749.700 ;
        RECT 254.100 749.700 261.900 751.050 ;
        RECT 254.100 744.600 255.900 749.700 ;
        RECT 257.100 744.000 258.900 748.800 ;
        RECT 260.100 744.600 261.900 749.700 ;
        RECT 263.100 750.600 264.300 752.700 ;
        RECT 275.400 750.600 276.300 757.950 ;
        RECT 277.950 756.150 279.750 757.950 ;
        RECT 284.100 756.150 285.900 757.950 ;
        RECT 288.000 756.450 292.050 757.050 ;
        RECT 287.550 754.950 292.050 756.450 ;
        RECT 277.950 753.450 280.050 754.050 ;
        RECT 287.550 753.450 288.450 754.950 ;
        RECT 293.550 754.050 294.450 764.550 ;
        RECT 298.950 763.950 301.050 764.550 ;
        RECT 299.100 757.950 301.200 760.050 ;
        RECT 299.250 756.150 301.050 757.950 ;
        RECT 291.000 753.900 294.450 754.050 ;
        RECT 277.950 752.550 288.450 753.450 ;
        RECT 289.950 752.550 294.450 753.900 ;
        RECT 302.100 753.300 303.000 773.400 ;
        RECT 305.100 768.000 306.900 780.000 ;
        RECT 308.100 767.400 309.900 779.400 ;
        RECT 320.400 767.400 322.200 780.000 ;
        RECT 325.500 768.900 327.300 779.400 ;
        RECT 328.500 773.400 330.300 780.000 ;
        RECT 344.100 778.500 351.900 779.400 ;
        RECT 328.200 770.100 330.000 771.900 ;
        RECT 325.500 767.400 327.900 768.900 ;
        RECT 344.100 767.400 345.900 778.500 ;
        RECT 304.200 760.050 306.000 761.850 ;
        RECT 308.400 760.050 309.300 767.400 ;
        RECT 310.950 763.950 313.050 766.050 ;
        RECT 304.500 757.950 306.600 760.050 ;
        RECT 307.800 757.950 309.900 760.050 ;
        RECT 277.950 751.950 280.050 752.550 ;
        RECT 289.950 751.950 294.000 752.550 ;
        RECT 299.100 752.400 307.500 753.300 ;
        RECT 289.950 751.800 292.050 751.950 ;
        RECT 263.100 744.600 264.900 750.600 ;
        RECT 275.400 749.400 280.500 750.600 ;
        RECT 275.700 744.000 277.500 747.600 ;
        RECT 278.700 744.600 280.500 749.400 ;
        RECT 283.200 744.000 285.000 750.600 ;
        RECT 286.950 747.450 289.050 748.050 ;
        RECT 292.950 747.450 295.050 748.050 ;
        RECT 286.950 746.550 295.050 747.450 ;
        RECT 286.950 745.950 289.050 746.550 ;
        RECT 292.950 745.950 295.050 746.550 ;
        RECT 299.100 744.600 300.900 752.400 ;
        RECT 305.700 751.500 307.500 752.400 ;
        RECT 308.400 750.600 309.300 757.950 ;
        RECT 311.550 756.450 312.450 763.950 ;
        RECT 320.100 760.050 321.900 761.850 ;
        RECT 326.700 760.050 327.900 767.400 ;
        RECT 347.100 766.500 348.900 777.600 ;
        RECT 350.100 768.600 351.900 778.500 ;
        RECT 353.100 769.500 354.900 780.000 ;
        RECT 356.100 768.600 357.900 779.400 ;
        RECT 350.100 767.700 357.900 768.600 ;
        RECT 368.100 768.600 369.900 779.400 ;
        RECT 371.100 769.500 372.900 780.000 ;
        RECT 374.100 778.500 381.900 779.400 ;
        RECT 374.100 768.600 375.900 778.500 ;
        RECT 368.100 767.700 375.900 768.600 ;
        RECT 377.100 766.500 378.900 777.600 ;
        RECT 380.100 767.400 381.900 778.500 ;
        RECT 392.700 773.400 394.500 780.000 ;
        RECT 393.000 770.100 394.800 771.900 ;
        RECT 395.700 768.900 397.500 779.400 ;
        RECT 395.100 767.400 397.500 768.900 ;
        RECT 400.800 767.400 402.600 780.000 ;
        RECT 416.700 773.400 418.500 780.000 ;
        RECT 417.000 770.100 418.800 771.900 ;
        RECT 419.700 768.900 421.500 779.400 ;
        RECT 419.100 767.400 421.500 768.900 ;
        RECT 424.800 767.400 426.600 780.000 ;
        RECT 440.100 773.400 441.900 780.000 ;
        RECT 443.100 773.400 444.900 779.400 ;
        RECT 446.100 773.400 447.900 780.000 ;
        RECT 347.100 765.600 351.900 766.500 ;
        RECT 339.000 762.450 343.050 763.050 ;
        RECT 338.550 760.950 343.050 762.450 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 316.950 756.450 319.050 757.050 ;
        RECT 311.550 755.550 319.050 756.450 ;
        RECT 323.100 756.150 324.900 757.950 ;
        RECT 316.950 754.950 319.050 755.550 ;
        RECT 326.700 753.600 327.900 757.950 ;
        RECT 329.100 756.150 330.900 757.950 ;
        RECT 338.550 756.900 339.450 760.950 ;
        RECT 347.100 760.050 348.900 761.850 ;
        RECT 351.000 760.050 351.900 765.600 ;
        RECT 374.100 765.600 378.900 766.500 ;
        RECT 352.950 760.050 354.750 761.850 ;
        RECT 371.250 760.050 373.050 761.850 ;
        RECT 374.100 760.050 375.000 765.600 ;
        RECT 390.000 765.450 394.050 766.050 ;
        RECT 389.550 763.950 394.050 765.450 ;
        RECT 389.550 762.450 390.450 763.950 ;
        RECT 377.100 760.050 378.900 761.850 ;
        RECT 386.550 761.550 390.450 762.450 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 346.950 757.950 349.050 760.050 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 337.950 754.800 340.050 756.900 ;
        RECT 344.100 756.150 345.900 757.950 ;
        RECT 326.700 752.700 330.300 753.600 ;
        RECT 303.600 744.000 305.400 750.600 ;
        RECT 306.600 748.800 309.300 750.600 ;
        RECT 320.100 749.700 327.900 751.050 ;
        RECT 306.600 744.600 308.400 748.800 ;
        RECT 320.100 744.600 321.900 749.700 ;
        RECT 323.100 744.000 324.900 748.800 ;
        RECT 326.100 744.600 327.900 749.700 ;
        RECT 329.100 750.600 330.300 752.700 ;
        RECT 331.950 753.450 334.050 754.050 ;
        RECT 346.950 753.450 349.050 753.750 ;
        RECT 331.950 752.550 349.050 753.450 ;
        RECT 331.950 751.950 334.050 752.550 ;
        RECT 346.950 751.650 349.050 752.550 ;
        RECT 350.700 750.600 351.900 757.950 ;
        RECT 355.950 756.150 357.750 757.950 ;
        RECT 368.250 756.150 370.050 757.950 ;
        RECT 374.100 750.600 375.300 757.950 ;
        RECT 380.100 756.150 381.900 757.950 ;
        RECT 386.550 757.050 387.450 761.550 ;
        RECT 395.100 760.050 396.300 767.400 ;
        RECT 401.100 760.050 402.900 761.850 ;
        RECT 419.100 760.050 420.300 767.400 ;
        RECT 435.000 762.450 439.050 763.050 ;
        RECT 425.100 760.050 426.900 761.850 ;
        RECT 434.550 760.950 439.050 762.450 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 418.950 757.950 421.050 760.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 386.550 755.550 391.050 757.050 ;
        RECT 392.100 756.150 393.900 757.950 ;
        RECT 387.000 754.950 391.050 755.550 ;
        RECT 395.100 753.600 396.300 757.950 ;
        RECT 398.100 756.150 399.900 757.950 ;
        RECT 416.100 756.150 417.900 757.950 ;
        RECT 419.100 753.600 420.300 757.950 ;
        RECT 422.100 756.150 423.900 757.950 ;
        RECT 434.550 757.050 435.450 760.950 ;
        RECT 443.100 760.050 444.300 773.400 ;
        RECT 458.100 767.400 459.900 779.400 ;
        RECT 461.100 768.000 462.900 780.000 ;
        RECT 464.100 773.400 465.900 779.400 ;
        RECT 467.100 773.400 468.900 780.000 ;
        RECT 479.100 773.400 480.900 780.000 ;
        RECT 482.100 773.400 483.900 779.400 ;
        RECT 485.100 774.000 486.900 780.000 ;
        RECT 458.700 760.050 459.600 767.400 ;
        RECT 462.000 760.050 463.800 761.850 ;
        RECT 439.950 757.950 442.050 760.050 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 458.100 757.950 460.200 760.050 ;
        RECT 461.400 757.950 463.500 760.050 ;
        RECT 434.550 755.550 439.050 757.050 ;
        RECT 440.250 756.150 442.050 757.950 ;
        RECT 435.000 754.950 439.050 755.550 ;
        RECT 392.700 752.700 396.300 753.600 ;
        RECT 416.700 752.700 420.300 753.600 ;
        RECT 443.100 752.700 444.300 757.950 ;
        RECT 446.100 756.150 447.900 757.950 ;
        RECT 392.700 750.600 393.900 752.700 ;
        RECT 329.100 744.600 330.900 750.600 ;
        RECT 346.500 744.000 348.300 750.600 ;
        RECT 351.000 744.600 352.800 750.600 ;
        RECT 355.500 744.000 357.300 750.600 ;
        RECT 368.700 744.000 370.500 750.600 ;
        RECT 373.200 744.600 375.000 750.600 ;
        RECT 377.700 744.000 379.500 750.600 ;
        RECT 392.100 744.600 393.900 750.600 ;
        RECT 395.100 749.700 402.900 751.050 ;
        RECT 416.700 750.600 417.900 752.700 ;
        RECT 443.100 751.800 447.300 752.700 ;
        RECT 395.100 744.600 396.900 749.700 ;
        RECT 398.100 744.000 399.900 748.800 ;
        RECT 401.100 744.600 402.900 749.700 ;
        RECT 416.100 744.600 417.900 750.600 ;
        RECT 419.100 749.700 426.900 751.050 ;
        RECT 419.100 744.600 420.900 749.700 ;
        RECT 422.100 744.000 423.900 748.800 ;
        RECT 425.100 744.600 426.900 749.700 ;
        RECT 440.400 744.000 442.200 750.600 ;
        RECT 445.500 744.600 447.300 751.800 ;
        RECT 458.700 750.600 459.600 757.950 ;
        RECT 465.000 753.300 465.900 773.400 ;
        RECT 482.400 773.100 483.900 773.400 ;
        RECT 488.100 773.400 489.900 779.400 ;
        RECT 488.100 773.100 489.000 773.400 ;
        RECT 482.400 772.200 489.000 773.100 ;
        RECT 482.100 760.050 483.900 761.850 ;
        RECT 488.100 760.050 489.000 772.200 ;
        RECT 500.100 767.400 501.900 780.000 ;
        RECT 503.100 767.400 504.900 779.400 ;
        RECT 515.400 767.400 517.200 780.000 ;
        RECT 520.500 768.900 522.300 779.400 ;
        RECT 523.500 773.400 525.300 780.000 ;
        RECT 539.100 773.400 540.900 780.000 ;
        RECT 542.100 773.400 543.900 779.400 ;
        RECT 545.100 773.400 546.900 780.000 ;
        RECT 560.700 773.400 562.500 780.000 ;
        RECT 523.200 770.100 525.000 771.900 ;
        RECT 520.500 767.400 522.900 768.900 ;
        RECT 493.950 763.950 496.050 766.050 ;
        RECT 466.800 757.950 468.900 760.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 484.950 757.950 487.050 760.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 466.950 756.150 468.750 757.950 ;
        RECT 479.100 756.150 480.900 757.950 ;
        RECT 485.100 756.150 486.900 757.950 ;
        RECT 488.100 754.200 489.000 757.950 ;
        RECT 494.550 757.050 495.450 763.950 ;
        RECT 503.100 760.050 504.300 767.400 ;
        RECT 515.100 760.050 516.900 761.850 ;
        RECT 521.700 760.050 522.900 767.400 ;
        RECT 542.100 760.050 543.300 773.400 ;
        RECT 561.000 770.100 562.800 771.900 ;
        RECT 563.700 768.900 565.500 779.400 ;
        RECT 563.100 767.400 565.500 768.900 ;
        RECT 568.800 767.400 570.600 780.000 ;
        RECT 581.100 767.400 582.900 780.000 ;
        RECT 586.200 768.600 588.000 779.400 ;
        RECT 602.100 773.400 603.900 779.400 ;
        RECT 605.100 773.400 606.900 780.000 ;
        RECT 584.400 767.400 588.000 768.600 ;
        RECT 555.000 762.450 559.050 763.050 ;
        RECT 554.550 760.950 559.050 762.450 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 490.950 755.550 495.450 757.050 ;
        RECT 500.100 756.150 501.900 757.950 ;
        RECT 490.950 754.950 495.000 755.550 ;
        RECT 460.500 752.400 468.900 753.300 ;
        RECT 460.500 751.500 462.300 752.400 ;
        RECT 458.700 748.800 461.400 750.600 ;
        RECT 459.600 744.600 461.400 748.800 ;
        RECT 462.600 744.000 464.400 750.600 ;
        RECT 467.100 744.600 468.900 752.400 ;
        RECT 479.100 744.000 480.900 753.600 ;
        RECT 485.700 753.000 489.000 754.200 ;
        RECT 485.700 744.600 487.500 753.000 ;
        RECT 503.100 750.600 504.300 757.950 ;
        RECT 518.100 756.150 519.900 757.950 ;
        RECT 521.700 753.600 522.900 757.950 ;
        RECT 524.100 756.150 525.900 757.950 ;
        RECT 539.250 756.150 541.050 757.950 ;
        RECT 521.700 752.700 525.300 753.600 ;
        RECT 500.100 744.000 501.900 750.600 ;
        RECT 503.100 744.600 504.900 750.600 ;
        RECT 515.100 749.700 522.900 751.050 ;
        RECT 515.100 744.600 516.900 749.700 ;
        RECT 518.100 744.000 519.900 748.800 ;
        RECT 521.100 744.600 522.900 749.700 ;
        RECT 524.100 750.600 525.300 752.700 ;
        RECT 542.100 752.700 543.300 757.950 ;
        RECT 545.100 756.150 546.900 757.950 ;
        RECT 547.950 756.450 550.050 757.050 ;
        RECT 554.550 756.450 555.450 760.950 ;
        RECT 563.100 760.050 564.300 767.400 ;
        RECT 571.950 762.450 576.000 763.050 ;
        RECT 569.100 760.050 570.900 761.850 ;
        RECT 571.950 760.950 576.450 762.450 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 562.950 757.950 565.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 547.950 755.550 555.450 756.450 ;
        RECT 560.100 756.150 561.900 757.950 ;
        RECT 547.950 754.950 550.050 755.550 ;
        RECT 563.100 753.600 564.300 757.950 ;
        RECT 566.100 756.150 567.900 757.950 ;
        RECT 575.550 757.050 576.450 760.950 ;
        RECT 581.250 760.050 583.050 761.850 ;
        RECT 584.400 760.050 585.300 767.400 ;
        RECT 598.950 762.450 601.050 763.050 ;
        RECT 587.100 760.050 588.900 761.850 ;
        RECT 593.550 761.550 601.050 762.450 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 586.950 757.950 589.050 760.050 ;
        RECT 571.950 755.550 576.450 757.050 ;
        RECT 571.950 754.950 576.000 755.550 ;
        RECT 560.700 752.700 564.300 753.600 ;
        RECT 542.100 751.800 546.300 752.700 ;
        RECT 524.100 744.600 525.900 750.600 ;
        RECT 539.400 744.000 541.200 750.600 ;
        RECT 544.500 744.600 546.300 751.800 ;
        RECT 560.700 750.600 561.900 752.700 ;
        RECT 560.100 744.600 561.900 750.600 ;
        RECT 563.100 749.700 570.900 751.050 ;
        RECT 563.100 744.600 564.900 749.700 ;
        RECT 566.100 744.000 567.900 748.800 ;
        RECT 569.100 744.600 570.900 749.700 ;
        RECT 584.400 747.600 585.300 757.950 ;
        RECT 593.550 757.050 594.450 761.550 ;
        RECT 598.950 760.950 601.050 761.550 ;
        RECT 602.700 760.050 603.900 773.400 ;
        RECT 617.100 767.400 618.900 779.400 ;
        RECT 620.100 767.400 621.900 780.000 ;
        RECT 632.100 767.400 633.900 779.400 ;
        RECT 636.600 767.400 638.400 780.000 ;
        RECT 639.600 768.900 641.400 779.400 ;
        RECT 656.100 773.400 657.900 780.000 ;
        RECT 659.100 773.400 660.900 779.400 ;
        RECT 662.100 773.400 663.900 780.000 ;
        RECT 639.600 767.400 642.000 768.900 ;
        RECT 605.100 760.050 606.900 761.850 ;
        RECT 617.700 760.050 618.900 767.400 ;
        RECT 632.100 765.900 633.300 767.400 ;
        RECT 632.100 764.700 639.900 765.900 ;
        RECT 638.100 764.100 639.900 764.700 ;
        RECT 625.950 760.950 628.050 763.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 589.950 755.550 594.450 757.050 ;
        RECT 589.950 754.950 594.000 755.550 ;
        RECT 602.700 747.600 603.900 757.950 ;
        RECT 617.700 750.600 618.900 757.950 ;
        RECT 620.100 756.150 621.900 757.950 ;
        RECT 626.550 757.050 627.450 760.950 ;
        RECT 636.000 760.050 637.800 761.850 ;
        RECT 632.100 757.950 634.200 760.050 ;
        RECT 635.400 757.950 637.500 760.050 ;
        RECT 622.950 755.550 627.450 757.050 ;
        RECT 632.400 756.150 634.200 757.950 ;
        RECT 622.950 754.950 627.000 755.550 ;
        RECT 638.700 753.600 639.600 764.100 ;
        RECT 640.800 760.050 642.000 767.400 ;
        RECT 646.950 768.450 649.050 769.050 ;
        RECT 652.950 768.450 655.050 769.050 ;
        RECT 646.950 767.550 655.050 768.450 ;
        RECT 646.950 766.950 649.050 767.550 ;
        RECT 652.950 766.950 655.050 767.550 ;
        RECT 659.700 760.050 660.900 773.400 ;
        RECT 677.400 767.400 679.200 780.000 ;
        RECT 682.500 768.900 684.300 779.400 ;
        RECT 685.500 773.400 687.300 780.000 ;
        RECT 701.100 773.400 702.900 779.400 ;
        RECT 704.100 774.000 705.900 780.000 ;
        RECT 702.000 773.100 702.900 773.400 ;
        RECT 707.100 773.400 708.900 779.400 ;
        RECT 710.100 773.400 711.900 780.000 ;
        RECT 707.100 773.100 708.600 773.400 ;
        RECT 702.000 772.200 708.600 773.100 ;
        RECT 685.200 770.100 687.000 771.900 ;
        RECT 682.500 767.400 684.900 768.900 ;
        RECT 677.100 760.050 678.900 761.850 ;
        RECT 683.700 760.050 684.900 767.400 ;
        RECT 702.000 760.050 702.900 772.200 ;
        RECT 703.950 768.450 706.050 769.050 ;
        RECT 709.950 768.450 712.050 769.050 ;
        RECT 703.950 767.550 712.050 768.450 ;
        RECT 703.950 766.950 706.050 767.550 ;
        RECT 709.950 766.950 712.050 767.550 ;
        RECT 725.400 767.400 727.200 780.000 ;
        RECT 730.500 768.900 732.300 779.400 ;
        RECT 733.500 773.400 735.300 780.000 ;
        RECT 749.100 773.400 750.900 780.000 ;
        RECT 752.100 773.400 753.900 779.400 ;
        RECT 733.200 770.100 735.000 771.900 ;
        RECT 730.500 767.400 732.900 768.900 ;
        RECT 715.950 765.450 718.050 766.050 ;
        RECT 724.950 765.450 727.050 766.050 ;
        RECT 715.950 764.550 727.050 765.450 ;
        RECT 715.950 763.950 718.050 764.550 ;
        RECT 724.950 763.950 727.050 764.550 ;
        RECT 707.100 760.050 708.900 761.850 ;
        RECT 725.100 760.050 726.900 761.850 ;
        RECT 731.700 760.050 732.900 767.400 ;
        RECT 640.800 757.950 642.900 760.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 749.100 757.950 751.200 760.050 ;
        RECT 638.700 752.700 640.800 753.600 ;
        RECT 635.400 751.800 640.800 752.700 ;
        RECT 581.100 744.000 582.900 747.600 ;
        RECT 584.100 744.600 585.900 747.600 ;
        RECT 587.100 744.000 588.900 747.600 ;
        RECT 602.100 744.600 603.900 747.600 ;
        RECT 605.100 744.000 606.900 747.600 ;
        RECT 617.100 744.600 618.900 750.600 ;
        RECT 620.100 744.000 621.900 750.600 ;
        RECT 635.400 747.600 636.300 751.800 ;
        RECT 642.000 750.600 642.900 757.950 ;
        RECT 656.100 756.150 657.900 757.950 ;
        RECT 659.700 752.700 660.900 757.950 ;
        RECT 661.950 756.150 663.750 757.950 ;
        RECT 680.100 756.150 681.900 757.950 ;
        RECT 683.700 753.600 684.900 757.950 ;
        RECT 686.100 756.150 687.900 757.950 ;
        RECT 702.000 754.200 702.900 757.950 ;
        RECT 704.100 756.150 705.900 757.950 ;
        RECT 710.100 756.150 711.900 757.950 ;
        RECT 728.100 756.150 729.900 757.950 ;
        RECT 683.700 752.700 687.300 753.600 ;
        RECT 702.000 753.000 705.300 754.200 ;
        RECT 731.700 753.600 732.900 757.950 ;
        RECT 734.100 756.150 735.900 757.950 ;
        RECT 749.250 756.150 751.050 757.950 ;
        RECT 632.100 744.600 633.900 747.600 ;
        RECT 635.100 744.600 636.900 747.600 ;
        RECT 632.100 744.000 633.300 744.600 ;
        RECT 638.100 744.000 639.900 750.000 ;
        RECT 641.100 744.600 642.900 750.600 ;
        RECT 656.700 751.800 660.900 752.700 ;
        RECT 656.700 744.600 658.500 751.800 ;
        RECT 661.800 744.000 663.600 750.600 ;
        RECT 677.100 749.700 684.900 751.050 ;
        RECT 677.100 744.600 678.900 749.700 ;
        RECT 680.100 744.000 681.900 748.800 ;
        RECT 683.100 744.600 684.900 749.700 ;
        RECT 686.100 750.600 687.300 752.700 ;
        RECT 686.100 744.600 687.900 750.600 ;
        RECT 703.500 744.600 705.300 753.000 ;
        RECT 710.100 744.000 711.900 753.600 ;
        RECT 731.700 752.700 735.300 753.600 ;
        RECT 752.100 753.300 753.000 773.400 ;
        RECT 755.100 768.000 756.900 780.000 ;
        RECT 758.100 767.400 759.900 779.400 ;
        RECT 773.100 767.400 774.900 779.400 ;
        RECT 776.100 768.300 777.900 779.400 ;
        RECT 779.100 769.200 780.900 780.000 ;
        RECT 782.100 768.300 783.900 779.400 ;
        RECT 776.100 767.400 783.900 768.300 ;
        RECT 797.100 768.600 798.900 779.400 ;
        RECT 800.100 769.500 801.900 780.000 ;
        RECT 803.100 778.500 810.900 779.400 ;
        RECT 803.100 768.600 804.900 778.500 ;
        RECT 797.100 767.700 804.900 768.600 ;
        RECT 754.200 760.050 756.000 761.850 ;
        RECT 758.400 760.050 759.300 767.400 ;
        RECT 773.400 760.050 774.300 767.400 ;
        RECT 806.100 766.500 807.900 777.600 ;
        RECT 809.100 767.400 810.900 778.500 ;
        RECT 821.100 773.400 822.900 779.400 ;
        RECT 824.100 774.000 825.900 780.000 ;
        RECT 822.000 773.100 822.900 773.400 ;
        RECT 827.100 773.400 828.900 779.400 ;
        RECT 830.100 773.400 831.900 780.000 ;
        RECT 842.700 773.400 844.500 780.000 ;
        RECT 827.100 773.100 828.600 773.400 ;
        RECT 822.000 772.200 828.600 773.100 ;
        RECT 803.100 765.600 807.900 766.500 ;
        RECT 793.950 762.450 796.050 763.050 ;
        RECT 778.950 760.050 780.750 761.850 ;
        RECT 788.550 761.550 796.050 762.450 ;
        RECT 754.500 757.950 756.600 760.050 ;
        RECT 757.800 757.950 759.900 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 725.100 749.700 732.900 751.050 ;
        RECT 725.100 744.600 726.900 749.700 ;
        RECT 728.100 744.000 729.900 748.800 ;
        RECT 731.100 744.600 732.900 749.700 ;
        RECT 734.100 750.600 735.300 752.700 ;
        RECT 749.100 752.400 757.500 753.300 ;
        RECT 734.100 744.600 735.900 750.600 ;
        RECT 749.100 744.600 750.900 752.400 ;
        RECT 755.700 751.500 757.500 752.400 ;
        RECT 758.400 750.600 759.300 757.950 ;
        RECT 753.600 744.000 755.400 750.600 ;
        RECT 756.600 748.800 759.300 750.600 ;
        RECT 773.400 750.600 774.300 757.950 ;
        RECT 775.950 756.150 777.750 757.950 ;
        RECT 782.100 756.150 783.900 757.950 ;
        RECT 788.550 757.050 789.450 761.550 ;
        RECT 793.950 760.950 796.050 761.550 ;
        RECT 800.250 760.050 802.050 761.850 ;
        RECT 803.100 760.050 804.000 765.600 ;
        RECT 806.100 760.050 807.900 761.850 ;
        RECT 822.000 760.050 822.900 772.200 ;
        RECT 843.000 770.100 844.800 771.900 ;
        RECT 823.950 768.450 826.050 769.050 ;
        RECT 841.950 768.450 844.050 769.050 ;
        RECT 845.700 768.900 847.500 779.400 ;
        RECT 823.950 767.550 844.050 768.450 ;
        RECT 823.950 766.950 826.050 767.550 ;
        RECT 841.950 766.950 844.050 767.550 ;
        RECT 845.100 767.400 847.500 768.900 ;
        RECT 850.800 767.400 852.600 780.000 ;
        RECT 866.100 773.400 867.900 779.400 ;
        RECT 869.100 774.000 870.900 780.000 ;
        RECT 867.000 773.100 867.900 773.400 ;
        RECT 872.100 773.400 873.900 779.400 ;
        RECT 875.100 773.400 876.900 780.000 ;
        RECT 872.100 773.100 873.600 773.400 ;
        RECT 867.000 772.200 873.600 773.100 ;
        RECT 829.950 765.450 832.050 765.900 ;
        RECT 841.950 765.450 844.050 766.050 ;
        RECT 829.950 764.550 844.050 765.450 ;
        RECT 829.950 763.800 832.050 764.550 ;
        RECT 841.950 763.950 844.050 764.550 ;
        RECT 827.100 760.050 828.900 761.850 ;
        RECT 845.100 760.050 846.300 767.400 ;
        RECT 851.100 760.050 852.900 761.850 ;
        RECT 867.000 760.050 867.900 772.200 ;
        RECT 887.100 767.400 888.900 779.400 ;
        RECT 890.100 768.300 891.900 779.400 ;
        RECT 893.100 769.200 894.900 780.000 ;
        RECT 896.100 768.300 897.900 779.400 ;
        RECT 911.100 773.400 912.900 779.400 ;
        RECT 914.100 774.000 915.900 780.000 ;
        RECT 890.100 767.400 897.900 768.300 ;
        RECT 912.000 773.100 912.900 773.400 ;
        RECT 917.100 773.400 918.900 779.400 ;
        RECT 920.100 773.400 921.900 780.000 ;
        RECT 917.100 773.100 918.600 773.400 ;
        RECT 912.000 772.200 918.600 773.100 ;
        RECT 872.100 760.050 873.900 761.850 ;
        RECT 887.400 760.050 888.300 767.400 ;
        RECT 892.950 760.050 894.750 761.850 ;
        RECT 912.000 760.050 912.900 772.200 ;
        RECT 916.950 765.450 919.050 766.050 ;
        RECT 916.950 764.550 924.450 765.450 ;
        RECT 916.950 763.950 919.050 764.550 ;
        RECT 923.550 762.450 924.450 764.550 ;
        RECT 917.100 760.050 918.900 761.850 ;
        RECT 923.550 761.550 927.450 762.450 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 865.950 757.950 868.050 760.050 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 871.950 757.950 874.050 760.050 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 889.950 757.950 892.050 760.050 ;
        RECT 892.950 757.950 895.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 913.950 757.950 916.050 760.050 ;
        RECT 916.950 757.950 919.050 760.050 ;
        RECT 919.950 757.950 922.050 760.050 ;
        RECT 784.950 755.550 789.450 757.050 ;
        RECT 797.250 756.150 799.050 757.950 ;
        RECT 784.950 754.950 789.000 755.550 ;
        RECT 803.100 750.600 804.300 757.950 ;
        RECT 809.100 756.150 810.900 757.950 ;
        RECT 822.000 754.200 822.900 757.950 ;
        RECT 824.100 756.150 825.900 757.950 ;
        RECT 830.100 756.150 831.900 757.950 ;
        RECT 842.100 756.150 843.900 757.950 ;
        RECT 805.950 753.450 808.050 754.050 ;
        RECT 814.950 753.450 817.050 754.050 ;
        RECT 805.950 752.550 817.050 753.450 ;
        RECT 822.000 753.000 825.300 754.200 ;
        RECT 845.100 753.600 846.300 757.950 ;
        RECT 848.100 756.150 849.900 757.950 ;
        RECT 805.950 751.950 808.050 752.550 ;
        RECT 814.950 751.950 817.050 752.550 ;
        RECT 773.400 749.400 778.500 750.600 ;
        RECT 756.600 744.600 758.400 748.800 ;
        RECT 773.700 744.000 775.500 747.600 ;
        RECT 776.700 744.600 778.500 749.400 ;
        RECT 781.200 744.000 783.000 750.600 ;
        RECT 797.700 744.000 799.500 750.600 ;
        RECT 802.200 744.600 804.000 750.600 ;
        RECT 806.700 744.000 808.500 750.600 ;
        RECT 823.500 744.600 825.300 753.000 ;
        RECT 830.100 744.000 831.900 753.600 ;
        RECT 842.700 752.700 846.300 753.600 ;
        RECT 867.000 754.200 867.900 757.950 ;
        RECT 869.100 756.150 870.900 757.950 ;
        RECT 875.100 756.150 876.900 757.950 ;
        RECT 867.000 753.000 870.300 754.200 ;
        RECT 842.700 750.600 843.900 752.700 ;
        RECT 842.100 744.600 843.900 750.600 ;
        RECT 845.100 749.700 852.900 751.050 ;
        RECT 845.100 744.600 846.900 749.700 ;
        RECT 848.100 744.000 849.900 748.800 ;
        RECT 851.100 744.600 852.900 749.700 ;
        RECT 868.500 744.600 870.300 753.000 ;
        RECT 875.100 744.000 876.900 753.600 ;
        RECT 887.400 750.600 888.300 757.950 ;
        RECT 889.950 756.150 891.750 757.950 ;
        RECT 896.100 756.150 897.900 757.950 ;
        RECT 912.000 754.200 912.900 757.950 ;
        RECT 914.100 756.150 915.900 757.950 ;
        RECT 920.100 756.150 921.900 757.950 ;
        RECT 926.550 757.050 927.450 761.550 ;
        RECT 922.950 755.550 927.450 757.050 ;
        RECT 922.950 754.950 927.000 755.550 ;
        RECT 912.000 753.000 915.300 754.200 ;
        RECT 887.400 749.400 892.500 750.600 ;
        RECT 887.700 744.000 889.500 747.600 ;
        RECT 890.700 744.600 892.500 749.400 ;
        RECT 895.200 744.000 897.000 750.600 ;
        RECT 913.500 744.600 915.300 753.000 ;
        RECT 920.100 744.000 921.900 753.600 ;
        RECT 11.100 737.400 12.900 741.000 ;
        RECT 14.100 737.400 15.900 740.400 ;
        RECT 17.100 737.400 18.900 741.000 ;
        RECT 29.100 737.400 30.900 740.400 ;
        RECT 32.100 737.400 33.900 741.000 ;
        RECT 47.100 737.400 48.900 741.000 ;
        RECT 50.100 737.400 51.900 740.400 ;
        RECT 53.100 737.400 54.900 741.000 ;
        RECT 68.100 737.400 69.900 740.400 ;
        RECT 71.100 737.400 72.900 741.000 ;
        RECT 83.100 737.400 84.900 740.400 ;
        RECT 86.100 737.400 87.900 741.000 ;
        RECT 14.400 727.050 15.300 737.400 ;
        RECT 29.700 727.050 30.900 737.400 ;
        RECT 31.950 735.450 34.050 736.050 ;
        RECT 46.950 735.450 49.050 736.050 ;
        RECT 31.950 734.550 49.050 735.450 ;
        RECT 31.950 733.950 34.050 734.550 ;
        RECT 46.950 733.950 49.050 734.550 ;
        RECT 50.400 727.050 51.300 737.400 ;
        RECT 68.700 727.050 69.900 737.400 ;
        RECT 83.700 727.050 84.900 737.400 ;
        RECT 101.100 734.400 102.900 740.400 ;
        RECT 101.700 732.300 102.900 734.400 ;
        RECT 104.100 735.300 105.900 740.400 ;
        RECT 107.100 736.200 108.900 741.000 ;
        RECT 110.100 735.300 111.900 740.400 ;
        RECT 104.100 733.950 111.900 735.300 ;
        RECT 122.100 734.400 123.900 740.400 ;
        RECT 122.700 732.300 123.900 734.400 ;
        RECT 125.100 735.300 126.900 740.400 ;
        RECT 128.100 736.200 129.900 741.000 ;
        RECT 131.100 735.300 132.900 740.400 ;
        RECT 125.100 733.950 132.900 735.300 ;
        RECT 143.100 734.400 144.900 740.400 ;
        RECT 146.100 735.300 147.900 741.000 ;
        RECT 150.600 734.400 152.400 740.400 ;
        RECT 155.100 735.300 156.900 741.000 ;
        RECT 158.100 734.400 159.900 740.400 ;
        RECT 170.100 737.400 171.900 741.000 ;
        RECT 173.100 737.400 174.900 740.400 ;
        RECT 176.100 737.400 177.900 741.000 ;
        RECT 191.100 737.400 192.900 740.400 ;
        RECT 194.100 737.400 195.900 741.000 ;
        RECT 206.700 737.400 208.500 741.000 ;
        RECT 143.100 733.500 147.900 734.400 ;
        RECT 145.800 732.300 147.900 733.500 ;
        RECT 150.900 732.900 152.100 734.400 ;
        RECT 101.700 731.400 105.300 732.300 ;
        RECT 122.700 731.400 126.300 732.300 ;
        RECT 96.000 729.450 100.050 730.050 ;
        RECT 95.550 727.950 100.050 729.450 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 46.950 724.950 49.050 727.050 ;
        RECT 49.950 724.950 52.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 67.950 724.950 70.050 727.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 11.250 723.150 13.050 724.950 ;
        RECT 14.400 717.600 15.300 724.950 ;
        RECT 17.100 723.150 18.900 724.950 ;
        RECT 11.100 705.000 12.900 717.600 ;
        RECT 14.400 716.400 18.000 717.600 ;
        RECT 16.200 705.600 18.000 716.400 ;
        RECT 29.700 711.600 30.900 724.950 ;
        RECT 32.100 723.150 33.900 724.950 ;
        RECT 47.250 723.150 49.050 724.950 ;
        RECT 50.400 717.600 51.300 724.950 ;
        RECT 53.100 723.150 54.900 724.950 ;
        RECT 29.100 705.600 30.900 711.600 ;
        RECT 32.100 705.000 33.900 711.600 ;
        RECT 47.100 705.000 48.900 717.600 ;
        RECT 50.400 716.400 54.000 717.600 ;
        RECT 52.200 705.600 54.000 716.400 ;
        RECT 68.700 711.600 69.900 724.950 ;
        RECT 71.100 723.150 72.900 724.950 ;
        RECT 83.700 711.600 84.900 724.950 ;
        RECT 86.100 723.150 87.900 724.950 ;
        RECT 95.550 724.050 96.450 727.950 ;
        RECT 101.100 727.050 102.900 728.850 ;
        RECT 104.100 727.050 105.300 731.400 ;
        RECT 107.100 727.050 108.900 728.850 ;
        RECT 122.100 727.050 123.900 728.850 ;
        RECT 125.100 727.050 126.300 731.400 ;
        RECT 149.100 730.800 152.100 732.900 ;
        RECT 158.100 732.600 159.300 734.400 ;
        RECT 128.100 727.050 129.900 728.850 ;
        RECT 147.900 727.800 150.000 729.900 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 143.100 724.950 145.200 727.050 ;
        RECT 147.900 726.000 149.700 727.800 ;
        RECT 150.900 725.100 152.100 730.800 ;
        RECT 153.000 731.700 159.300 732.600 ;
        RECT 153.000 729.600 155.100 731.700 ;
        RECT 153.000 727.800 154.800 729.600 ;
        RECT 157.800 727.050 159.600 728.850 ;
        RECT 173.400 727.050 174.300 737.400 ;
        RECT 191.700 727.050 192.900 737.400 ;
        RECT 209.700 735.600 211.500 740.400 ;
        RECT 206.400 734.400 211.500 735.600 ;
        RECT 214.200 734.400 216.000 741.000 ;
        RECT 230.100 734.400 231.900 740.400 ;
        RECT 206.400 727.050 207.300 734.400 ;
        RECT 230.700 732.300 231.900 734.400 ;
        RECT 233.100 735.300 234.900 740.400 ;
        RECT 236.100 736.200 237.900 741.000 ;
        RECT 239.100 735.300 240.900 740.400 ;
        RECT 251.100 737.400 252.900 740.400 ;
        RECT 254.100 737.400 255.900 741.000 ;
        RECT 233.100 733.950 240.900 735.300 ;
        RECT 230.700 731.400 234.300 732.300 ;
        RECT 208.950 727.050 210.750 728.850 ;
        RECT 215.100 727.050 216.900 728.850 ;
        RECT 230.100 727.050 231.900 728.850 ;
        RECT 233.100 727.050 234.300 731.400 ;
        RECT 241.950 729.450 246.000 730.050 ;
        RECT 236.100 727.050 237.900 728.850 ;
        RECT 241.950 727.950 246.450 729.450 ;
        RECT 157.800 726.300 159.900 727.050 ;
        RECT 95.550 722.550 100.050 724.050 ;
        RECT 96.000 721.950 100.050 722.550 ;
        RECT 104.100 717.600 105.300 724.950 ;
        RECT 110.100 723.150 111.900 724.950 ;
        RECT 112.950 720.450 115.050 721.050 ;
        RECT 121.950 720.450 124.050 721.050 ;
        RECT 112.950 719.550 124.050 720.450 ;
        RECT 112.950 718.950 115.050 719.550 ;
        RECT 121.950 718.950 124.050 719.550 ;
        RECT 125.100 717.600 126.300 724.950 ;
        RECT 131.100 723.150 132.900 724.950 ;
        RECT 143.400 723.150 145.200 724.950 ;
        RECT 149.700 724.200 152.100 725.100 ;
        RECT 153.000 724.950 159.900 726.300 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 205.950 724.950 208.050 727.050 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 153.000 724.500 154.800 724.950 ;
        RECT 149.700 724.050 151.200 724.200 ;
        RECT 149.100 721.950 151.200 724.050 ;
        RECT 127.950 720.450 130.050 721.050 ;
        RECT 139.950 720.450 142.050 721.050 ;
        RECT 127.950 719.550 142.050 720.450 ;
        RECT 127.950 718.950 130.050 719.550 ;
        RECT 139.950 718.950 142.050 719.550 ;
        RECT 150.300 720.000 151.200 721.950 ;
        RECT 152.100 721.500 156.000 723.300 ;
        RECT 170.250 723.150 172.050 724.950 ;
        RECT 152.100 721.200 154.200 721.500 ;
        RECT 150.300 718.950 151.800 720.000 ;
        RECT 145.800 717.600 147.900 718.500 ;
        RECT 104.100 716.100 106.500 717.600 ;
        RECT 102.000 713.100 103.800 714.900 ;
        RECT 68.100 705.600 69.900 711.600 ;
        RECT 71.100 705.000 72.900 711.600 ;
        RECT 83.100 705.600 84.900 711.600 ;
        RECT 86.100 705.000 87.900 711.600 ;
        RECT 101.700 705.000 103.500 711.600 ;
        RECT 104.700 705.600 106.500 716.100 ;
        RECT 109.800 705.000 111.600 717.600 ;
        RECT 125.100 716.100 127.500 717.600 ;
        RECT 123.000 713.100 124.800 714.900 ;
        RECT 122.700 705.000 124.500 711.600 ;
        RECT 125.700 705.600 127.500 716.100 ;
        RECT 130.800 705.000 132.600 717.600 ;
        RECT 143.100 716.400 147.900 717.600 ;
        RECT 150.600 717.600 151.800 718.950 ;
        RECT 155.400 717.600 157.500 719.700 ;
        RECT 173.400 717.600 174.300 724.950 ;
        RECT 176.100 723.150 177.900 724.950 ;
        RECT 143.100 705.600 144.900 716.400 ;
        RECT 146.100 705.000 147.900 715.500 ;
        RECT 150.600 705.600 152.400 717.600 ;
        RECT 155.400 716.700 159.900 717.600 ;
        RECT 155.100 705.000 156.900 715.500 ;
        RECT 158.100 705.600 159.900 716.700 ;
        RECT 170.100 705.000 171.900 717.600 ;
        RECT 173.400 716.400 177.000 717.600 ;
        RECT 175.200 705.600 177.000 716.400 ;
        RECT 191.700 711.600 192.900 724.950 ;
        RECT 194.100 723.150 195.900 724.950 ;
        RECT 206.400 717.600 207.300 724.950 ;
        RECT 211.950 723.150 213.750 724.950 ;
        RECT 208.950 720.450 211.050 720.750 ;
        RECT 223.950 720.450 226.050 721.050 ;
        RECT 208.950 719.550 226.050 720.450 ;
        RECT 208.950 718.650 211.050 719.550 ;
        RECT 223.950 718.950 226.050 719.550 ;
        RECT 233.100 717.600 234.300 724.950 ;
        RECT 239.100 723.150 240.900 724.950 ;
        RECT 245.550 724.050 246.450 727.950 ;
        RECT 251.700 727.050 252.900 737.400 ;
        RECT 269.100 734.400 270.900 740.400 ;
        RECT 269.700 732.300 270.900 734.400 ;
        RECT 272.100 735.300 273.900 740.400 ;
        RECT 275.100 736.200 276.900 741.000 ;
        RECT 278.100 735.300 279.900 740.400 ;
        RECT 272.100 733.950 279.900 735.300 ;
        RECT 293.100 732.600 294.900 740.400 ;
        RECT 297.600 734.400 299.400 741.000 ;
        RECT 300.600 736.200 302.400 740.400 ;
        RECT 300.600 734.400 303.300 736.200 ;
        RECT 299.700 732.600 301.500 733.500 ;
        RECT 269.700 731.400 273.300 732.300 ;
        RECT 293.100 731.700 301.500 732.600 ;
        RECT 269.100 727.050 270.900 728.850 ;
        RECT 272.100 727.050 273.300 731.400 ;
        RECT 275.100 727.050 276.900 728.850 ;
        RECT 293.250 727.050 295.050 728.850 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 293.100 724.950 295.200 727.050 ;
        RECT 241.950 722.550 246.450 724.050 ;
        RECT 241.950 721.950 246.000 722.550 ;
        RECT 191.100 705.600 192.900 711.600 ;
        RECT 194.100 705.000 195.900 711.600 ;
        RECT 206.100 705.600 207.900 717.600 ;
        RECT 209.100 716.700 216.900 717.600 ;
        RECT 209.100 705.600 210.900 716.700 ;
        RECT 212.100 705.000 213.900 715.800 ;
        RECT 215.100 705.600 216.900 716.700 ;
        RECT 233.100 716.100 235.500 717.600 ;
        RECT 231.000 713.100 232.800 714.900 ;
        RECT 230.700 705.000 232.500 711.600 ;
        RECT 233.700 705.600 235.500 716.100 ;
        RECT 238.800 705.000 240.600 717.600 ;
        RECT 251.700 711.600 252.900 724.950 ;
        RECT 254.100 723.150 255.900 724.950 ;
        RECT 272.100 717.600 273.300 724.950 ;
        RECT 278.100 723.150 279.900 724.950 ;
        RECT 272.100 716.100 274.500 717.600 ;
        RECT 270.000 713.100 271.800 714.900 ;
        RECT 251.100 705.600 252.900 711.600 ;
        RECT 254.100 705.000 255.900 711.600 ;
        RECT 269.700 705.000 271.500 711.600 ;
        RECT 272.700 705.600 274.500 716.100 ;
        RECT 277.800 705.000 279.600 717.600 ;
        RECT 296.100 711.600 297.000 731.700 ;
        RECT 302.400 727.050 303.300 734.400 ;
        RECT 314.100 735.300 315.900 740.400 ;
        RECT 317.100 736.200 318.900 741.000 ;
        RECT 320.100 735.300 321.900 740.400 ;
        RECT 314.100 733.950 321.900 735.300 ;
        RECT 323.100 734.400 324.900 740.400 ;
        RECT 323.100 732.300 324.300 734.400 ;
        RECT 335.700 733.200 337.500 740.400 ;
        RECT 340.800 734.400 342.600 741.000 ;
        RECT 353.100 734.400 354.900 740.400 ;
        RECT 335.700 732.300 339.900 733.200 ;
        RECT 320.700 731.400 324.300 732.300 ;
        RECT 317.100 727.050 318.900 728.850 ;
        RECT 320.700 727.050 321.900 731.400 ;
        RECT 323.100 727.050 324.900 728.850 ;
        RECT 335.100 727.050 336.900 728.850 ;
        RECT 338.700 727.050 339.900 732.300 ;
        RECT 353.700 732.300 354.900 734.400 ;
        RECT 356.100 735.300 357.900 740.400 ;
        RECT 359.100 736.200 360.900 741.000 ;
        RECT 362.100 735.300 363.900 740.400 ;
        RECT 356.100 733.950 363.900 735.300 ;
        RECT 374.700 734.400 376.500 741.000 ;
        RECT 379.200 734.400 381.000 740.400 ;
        RECT 383.700 734.400 385.500 741.000 ;
        RECT 398.400 734.400 400.200 741.000 ;
        RECT 353.700 731.400 357.300 732.300 ;
        RECT 340.950 727.050 342.750 728.850 ;
        RECT 353.100 727.050 354.900 728.850 ;
        RECT 356.100 727.050 357.300 731.400 ;
        RECT 359.100 727.050 360.900 728.850 ;
        RECT 374.250 727.050 376.050 728.850 ;
        RECT 380.100 727.050 381.300 734.400 ;
        RECT 403.500 733.200 405.300 740.400 ;
        RECT 419.400 734.400 421.200 741.000 ;
        RECT 424.500 733.200 426.300 740.400 ;
        RECT 440.100 734.400 441.900 740.400 ;
        RECT 401.100 732.300 405.300 733.200 ;
        RECT 422.100 732.300 426.300 733.200 ;
        RECT 440.700 732.300 441.900 734.400 ;
        RECT 443.100 735.300 444.900 740.400 ;
        RECT 446.100 736.200 447.900 741.000 ;
        RECT 449.100 735.300 450.900 740.400 ;
        RECT 462.600 736.200 464.400 740.400 ;
        RECT 443.100 733.950 450.900 735.300 ;
        RECT 461.700 734.400 464.400 736.200 ;
        RECT 465.600 734.400 467.400 741.000 ;
        RECT 386.100 727.050 387.900 728.850 ;
        RECT 398.250 727.050 400.050 728.850 ;
        RECT 401.100 727.050 402.300 732.300 ;
        RECT 404.100 727.050 405.900 728.850 ;
        RECT 419.250 727.050 421.050 728.850 ;
        RECT 422.100 727.050 423.300 732.300 ;
        RECT 440.700 731.400 444.300 732.300 ;
        RECT 425.100 727.050 426.900 728.850 ;
        RECT 440.100 727.050 441.900 728.850 ;
        RECT 443.100 727.050 444.300 731.400 ;
        RECT 446.100 727.050 447.900 728.850 ;
        RECT 461.700 727.050 462.600 734.400 ;
        RECT 463.500 732.600 465.300 733.500 ;
        RECT 470.100 732.600 471.900 740.400 ;
        RECT 463.500 731.700 471.900 732.600 ;
        RECT 485.700 733.200 487.500 740.400 ;
        RECT 490.800 734.400 492.600 741.000 ;
        RECT 505.500 734.400 507.300 741.000 ;
        RECT 510.000 734.400 511.800 740.400 ;
        RECT 514.500 734.400 516.300 741.000 ;
        RECT 485.700 732.300 489.900 733.200 ;
        RECT 298.500 724.950 300.600 727.050 ;
        RECT 301.800 724.950 303.900 727.050 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 334.950 724.950 337.050 727.050 ;
        RECT 337.950 724.950 340.050 727.050 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 385.950 724.950 388.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 461.100 724.950 463.200 727.050 ;
        RECT 464.400 724.950 466.500 727.050 ;
        RECT 298.200 723.150 300.000 724.950 ;
        RECT 302.400 717.600 303.300 724.950 ;
        RECT 314.100 723.150 315.900 724.950 ;
        RECT 320.700 717.600 321.900 724.950 ;
        RECT 325.950 720.450 328.050 721.050 ;
        RECT 334.950 720.450 337.050 721.050 ;
        RECT 325.950 719.550 337.050 720.450 ;
        RECT 325.950 718.950 328.050 719.550 ;
        RECT 334.950 718.950 337.050 719.550 ;
        RECT 293.100 705.000 294.900 711.600 ;
        RECT 296.100 705.600 297.900 711.600 ;
        RECT 299.100 705.000 300.900 717.000 ;
        RECT 302.100 705.600 303.900 717.600 ;
        RECT 314.400 705.000 316.200 717.600 ;
        RECT 319.500 716.100 321.900 717.600 ;
        RECT 319.500 705.600 321.300 716.100 ;
        RECT 322.200 713.100 324.000 714.900 ;
        RECT 338.700 711.600 339.900 724.950 ;
        RECT 356.100 717.600 357.300 724.950 ;
        RECT 362.100 723.150 363.900 724.950 ;
        RECT 377.250 723.150 379.050 724.950 ;
        RECT 358.950 720.450 361.050 721.050 ;
        RECT 376.950 720.450 379.050 721.050 ;
        RECT 358.950 719.550 379.050 720.450 ;
        RECT 358.950 718.950 361.050 719.550 ;
        RECT 376.950 718.950 379.050 719.550 ;
        RECT 380.100 719.400 381.000 724.950 ;
        RECT 383.100 723.150 384.900 724.950 ;
        RECT 385.950 720.450 388.050 721.050 ;
        RECT 391.950 720.450 394.050 721.050 ;
        RECT 385.950 719.550 394.050 720.450 ;
        RECT 380.100 718.500 384.900 719.400 ;
        RECT 385.950 718.950 388.050 719.550 ;
        RECT 391.950 718.950 394.050 719.550 ;
        RECT 356.100 716.100 358.500 717.600 ;
        RECT 354.000 713.100 355.800 714.900 ;
        RECT 322.500 705.000 324.300 711.600 ;
        RECT 335.100 705.000 336.900 711.600 ;
        RECT 338.100 705.600 339.900 711.600 ;
        RECT 341.100 705.000 342.900 711.600 ;
        RECT 353.700 705.000 355.500 711.600 ;
        RECT 356.700 705.600 358.500 716.100 ;
        RECT 361.800 705.000 363.600 717.600 ;
        RECT 374.100 716.400 381.900 717.300 ;
        RECT 374.100 705.600 375.900 716.400 ;
        RECT 377.100 705.000 378.900 715.500 ;
        RECT 380.100 706.500 381.900 716.400 ;
        RECT 383.100 707.400 384.900 718.500 ;
        RECT 386.100 706.500 387.900 717.600 ;
        RECT 401.100 711.600 402.300 724.950 ;
        RECT 422.100 711.600 423.300 724.950 ;
        RECT 443.100 717.600 444.300 724.950 ;
        RECT 449.100 723.150 450.900 724.950 ;
        RECT 448.950 720.450 451.050 721.050 ;
        RECT 454.950 720.450 457.050 721.050 ;
        RECT 448.950 719.550 457.050 720.450 ;
        RECT 448.950 718.950 451.050 719.550 ;
        RECT 454.950 718.950 457.050 719.550 ;
        RECT 461.700 717.600 462.600 724.950 ;
        RECT 465.000 723.150 466.800 724.950 ;
        RECT 443.100 716.100 445.500 717.600 ;
        RECT 441.000 713.100 442.800 714.900 ;
        RECT 380.100 705.600 387.900 706.500 ;
        RECT 398.100 705.000 399.900 711.600 ;
        RECT 401.100 705.600 402.900 711.600 ;
        RECT 404.100 705.000 405.900 711.600 ;
        RECT 419.100 705.000 420.900 711.600 ;
        RECT 422.100 705.600 423.900 711.600 ;
        RECT 425.100 705.000 426.900 711.600 ;
        RECT 440.700 705.000 442.500 711.600 ;
        RECT 443.700 705.600 445.500 716.100 ;
        RECT 448.800 705.000 450.600 717.600 ;
        RECT 461.100 705.600 462.900 717.600 ;
        RECT 464.100 705.000 465.900 717.000 ;
        RECT 468.000 711.600 468.900 731.700 ;
        RECT 469.950 727.050 471.750 728.850 ;
        RECT 485.100 727.050 486.900 728.850 ;
        RECT 488.700 727.050 489.900 732.300 ;
        RECT 498.000 729.450 502.050 730.050 ;
        RECT 490.950 727.050 492.750 728.850 ;
        RECT 497.550 727.950 502.050 729.450 ;
        RECT 469.800 724.950 471.900 727.050 ;
        RECT 484.950 724.950 487.050 727.050 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 488.700 711.600 489.900 724.950 ;
        RECT 497.550 724.050 498.450 727.950 ;
        RECT 503.100 727.050 504.900 728.850 ;
        RECT 509.700 727.050 510.900 734.400 ;
        RECT 529.500 732.000 531.300 740.400 ;
        RECT 528.000 730.800 531.300 732.000 ;
        RECT 536.100 731.400 537.900 741.000 ;
        RECT 548.100 734.400 549.900 740.400 ;
        RECT 551.100 734.400 552.900 741.000 ;
        RECT 563.100 737.400 564.900 740.400 ;
        RECT 566.100 737.400 567.900 741.000 ;
        RECT 514.950 727.050 516.750 728.850 ;
        RECT 528.000 727.050 528.900 730.800 ;
        RECT 530.100 727.050 531.900 728.850 ;
        RECT 536.100 727.050 537.900 728.850 ;
        RECT 548.700 727.050 549.900 734.400 ;
        RECT 551.100 727.050 552.900 728.850 ;
        RECT 563.700 727.050 564.900 737.400 ;
        RECT 581.100 734.400 582.900 740.400 ;
        RECT 584.100 735.000 585.900 741.000 ;
        RECT 590.700 740.400 591.900 741.000 ;
        RECT 587.100 737.400 588.900 740.400 ;
        RECT 590.100 737.400 591.900 740.400 ;
        RECT 602.100 737.400 603.900 740.400 ;
        RECT 568.950 729.450 573.000 730.050 ;
        RECT 568.950 727.950 573.450 729.450 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 497.550 722.550 502.050 724.050 ;
        RECT 506.100 723.150 507.900 724.950 ;
        RECT 498.000 721.950 502.050 722.550 ;
        RECT 510.000 719.400 510.900 724.950 ;
        RECT 511.950 723.150 513.750 724.950 ;
        RECT 506.100 718.500 510.900 719.400 ;
        RECT 467.100 705.600 468.900 711.600 ;
        RECT 470.100 705.000 471.900 711.600 ;
        RECT 485.100 705.000 486.900 711.600 ;
        RECT 488.100 705.600 489.900 711.600 ;
        RECT 491.100 705.000 492.900 711.600 ;
        RECT 503.100 706.500 504.900 717.600 ;
        RECT 506.100 707.400 507.900 718.500 ;
        RECT 509.100 716.400 516.900 717.300 ;
        RECT 509.100 706.500 510.900 716.400 ;
        RECT 503.100 705.600 510.900 706.500 ;
        RECT 512.100 705.000 513.900 715.500 ;
        RECT 515.100 705.600 516.900 716.400 ;
        RECT 528.000 712.800 528.900 724.950 ;
        RECT 533.100 723.150 534.900 724.950 ;
        RECT 548.700 717.600 549.900 724.950 ;
        RECT 528.000 711.900 534.600 712.800 ;
        RECT 528.000 711.600 528.900 711.900 ;
        RECT 527.100 705.600 528.900 711.600 ;
        RECT 533.100 711.600 534.600 711.900 ;
        RECT 530.100 705.000 531.900 711.000 ;
        RECT 533.100 705.600 534.900 711.600 ;
        RECT 536.100 705.000 537.900 711.600 ;
        RECT 548.100 705.600 549.900 717.600 ;
        RECT 551.100 705.000 552.900 717.600 ;
        RECT 563.700 711.600 564.900 724.950 ;
        RECT 566.100 723.150 567.900 724.950 ;
        RECT 572.550 724.050 573.450 727.950 ;
        RECT 581.100 727.050 582.000 734.400 ;
        RECT 587.700 733.200 588.600 737.400 ;
        RECT 583.200 732.300 588.600 733.200 ;
        RECT 602.100 733.500 603.300 737.400 ;
        RECT 605.100 734.400 606.900 741.000 ;
        RECT 608.100 734.400 609.900 740.400 ;
        RECT 602.100 732.600 607.800 733.500 ;
        RECT 583.200 731.400 585.300 732.300 ;
        RECT 581.100 724.950 583.200 727.050 ;
        RECT 568.950 722.550 573.450 724.050 ;
        RECT 568.950 721.950 573.000 722.550 ;
        RECT 582.000 717.600 583.200 724.950 ;
        RECT 584.400 720.900 585.300 731.400 ;
        RECT 606.000 731.700 607.800 732.600 ;
        RECT 589.800 727.050 591.600 728.850 ;
        RECT 586.500 724.950 588.600 727.050 ;
        RECT 589.800 724.950 591.900 727.050 ;
        RECT 602.400 724.950 604.500 727.050 ;
        RECT 586.200 723.150 588.000 724.950 ;
        RECT 602.400 723.150 604.200 724.950 ;
        RECT 584.100 720.300 585.900 720.900 ;
        RECT 606.000 720.300 606.900 731.700 ;
        RECT 608.700 727.050 609.900 734.400 ;
        RECT 620.100 735.300 621.900 740.400 ;
        RECT 623.100 736.200 624.900 741.000 ;
        RECT 626.100 735.300 627.900 740.400 ;
        RECT 620.100 733.950 627.900 735.300 ;
        RECT 629.100 734.400 630.900 740.400 ;
        RECT 641.100 737.400 642.900 740.400 ;
        RECT 644.100 737.400 645.900 741.000 ;
        RECT 629.100 732.300 630.300 734.400 ;
        RECT 626.700 731.400 630.300 732.300 ;
        RECT 623.100 727.050 624.900 728.850 ;
        RECT 626.700 727.050 627.900 731.400 ;
        RECT 629.100 727.050 630.900 728.850 ;
        RECT 634.950 727.950 637.050 730.050 ;
        RECT 607.800 724.950 609.900 727.050 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 622.950 724.950 625.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 584.100 719.100 591.900 720.300 ;
        RECT 606.000 719.400 607.800 720.300 ;
        RECT 590.700 717.600 591.900 719.100 ;
        RECT 582.000 716.100 584.400 717.600 ;
        RECT 563.100 705.600 564.900 711.600 ;
        RECT 566.100 705.000 567.900 711.600 ;
        RECT 582.600 705.600 584.400 716.100 ;
        RECT 585.600 705.000 587.400 717.600 ;
        RECT 590.100 705.600 591.900 717.600 ;
        RECT 602.100 718.500 607.800 719.400 ;
        RECT 602.100 711.600 603.300 718.500 ;
        RECT 608.700 717.600 609.900 724.950 ;
        RECT 613.950 720.450 616.050 724.050 ;
        RECT 620.100 723.150 621.900 724.950 ;
        RECT 619.950 720.450 622.050 721.050 ;
        RECT 613.950 720.000 622.050 720.450 ;
        RECT 614.550 719.550 622.050 720.000 ;
        RECT 619.950 718.950 622.050 719.550 ;
        RECT 626.700 717.600 627.900 724.950 ;
        RECT 635.550 724.050 636.450 727.950 ;
        RECT 641.700 727.050 642.900 737.400 ;
        RECT 656.400 734.400 658.200 741.000 ;
        RECT 661.500 733.200 663.300 740.400 ;
        RECT 659.100 732.300 663.300 733.200 ;
        RECT 646.950 729.450 651.000 730.050 ;
        RECT 646.950 727.950 651.450 729.450 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 634.950 721.950 637.050 724.050 ;
        RECT 628.950 720.450 631.050 721.050 ;
        RECT 637.950 720.450 640.050 721.050 ;
        RECT 628.950 719.550 640.050 720.450 ;
        RECT 628.950 718.950 631.050 719.550 ;
        RECT 637.950 718.950 640.050 719.550 ;
        RECT 602.100 705.600 603.900 711.600 ;
        RECT 605.100 705.000 606.900 715.800 ;
        RECT 608.100 705.600 609.900 717.600 ;
        RECT 620.400 705.000 622.200 717.600 ;
        RECT 625.500 716.100 627.900 717.600 ;
        RECT 625.500 705.600 627.300 716.100 ;
        RECT 628.200 713.100 630.000 714.900 ;
        RECT 641.700 711.600 642.900 724.950 ;
        RECT 644.100 723.150 645.900 724.950 ;
        RECT 650.550 724.050 651.450 727.950 ;
        RECT 656.250 727.050 658.050 728.850 ;
        RECT 659.100 727.050 660.300 732.300 ;
        RECT 674.100 731.400 675.900 741.000 ;
        RECT 680.700 732.000 682.500 740.400 ;
        RECT 695.100 734.400 696.900 740.400 ;
        RECT 695.700 732.300 696.900 734.400 ;
        RECT 698.100 735.300 699.900 740.400 ;
        RECT 701.100 736.200 702.900 741.000 ;
        RECT 704.100 735.300 705.900 740.400 ;
        RECT 716.100 737.400 717.900 741.000 ;
        RECT 719.100 737.400 720.900 740.400 ;
        RECT 731.100 737.400 732.900 740.400 ;
        RECT 734.100 737.400 735.900 741.000 ;
        RECT 698.100 733.950 705.900 735.300 ;
        RECT 680.700 730.800 684.000 732.000 ;
        RECT 695.700 731.400 699.300 732.300 ;
        RECT 662.100 727.050 663.900 728.850 ;
        RECT 674.100 727.050 675.900 728.850 ;
        RECT 680.100 727.050 681.900 728.850 ;
        RECT 683.100 727.050 684.000 730.800 ;
        RECT 690.000 729.450 694.050 730.050 ;
        RECT 689.550 727.950 694.050 729.450 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 646.950 722.550 651.450 724.050 ;
        RECT 646.950 721.950 651.000 722.550 ;
        RECT 659.100 711.600 660.300 724.950 ;
        RECT 677.100 723.150 678.900 724.950 ;
        RECT 683.100 712.800 684.000 724.950 ;
        RECT 689.550 724.050 690.450 727.950 ;
        RECT 695.100 727.050 696.900 728.850 ;
        RECT 698.100 727.050 699.300 731.400 ;
        RECT 701.100 727.050 702.900 728.850 ;
        RECT 719.100 727.050 720.300 737.400 ;
        RECT 721.950 729.450 726.000 730.050 ;
        RECT 721.950 729.000 726.450 729.450 ;
        RECT 721.950 727.950 727.050 729.000 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 685.950 722.550 690.450 724.050 ;
        RECT 685.950 721.950 690.000 722.550 ;
        RECT 698.100 717.600 699.300 724.950 ;
        RECT 704.100 723.150 705.900 724.950 ;
        RECT 716.100 723.150 717.900 724.950 ;
        RECT 698.100 716.100 700.500 717.600 ;
        RECT 696.000 713.100 697.800 714.900 ;
        RECT 677.400 711.900 684.000 712.800 ;
        RECT 677.400 711.600 678.900 711.900 ;
        RECT 628.500 705.000 630.300 711.600 ;
        RECT 641.100 705.600 642.900 711.600 ;
        RECT 644.100 705.000 645.900 711.600 ;
        RECT 656.100 705.000 657.900 711.600 ;
        RECT 659.100 705.600 660.900 711.600 ;
        RECT 662.100 705.000 663.900 711.600 ;
        RECT 674.100 705.000 675.900 711.600 ;
        RECT 677.100 705.600 678.900 711.600 ;
        RECT 683.100 711.600 684.000 711.900 ;
        RECT 680.100 705.000 681.900 711.000 ;
        RECT 683.100 705.600 684.900 711.600 ;
        RECT 695.700 705.000 697.500 711.600 ;
        RECT 698.700 705.600 700.500 716.100 ;
        RECT 703.800 705.000 705.600 717.600 ;
        RECT 719.100 711.600 720.300 724.950 ;
        RECT 724.950 724.800 727.050 727.950 ;
        RECT 731.700 727.050 732.900 737.400 ;
        RECT 751.500 732.000 753.300 740.400 ;
        RECT 750.000 730.800 753.300 732.000 ;
        RECT 758.100 731.400 759.900 741.000 ;
        RECT 770.100 731.400 771.900 741.000 ;
        RECT 776.700 732.000 778.500 740.400 ;
        RECT 784.950 738.450 787.050 738.900 ;
        RECT 790.950 738.450 793.050 739.050 ;
        RECT 784.950 737.550 793.050 738.450 ;
        RECT 784.950 736.800 787.050 737.550 ;
        RECT 790.950 736.950 793.050 737.550 ;
        RECT 794.100 734.400 795.900 740.400 ;
        RECT 794.700 732.300 795.900 734.400 ;
        RECT 797.100 735.300 798.900 740.400 ;
        RECT 800.100 736.200 801.900 741.000 ;
        RECT 803.100 735.300 804.900 740.400 ;
        RECT 815.700 737.400 817.500 741.000 ;
        RECT 818.700 735.600 820.500 740.400 ;
        RECT 797.100 733.950 804.900 735.300 ;
        RECT 815.400 734.400 820.500 735.600 ;
        RECT 823.200 734.400 825.000 741.000 ;
        RECT 776.700 730.800 780.000 732.000 ;
        RECT 794.700 731.400 798.300 732.300 ;
        RECT 750.000 727.050 750.900 730.800 ;
        RECT 765.000 729.450 769.050 730.050 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 758.100 727.050 759.900 728.850 ;
        RECT 764.550 727.950 769.050 729.450 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 754.950 724.950 757.050 727.050 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 731.700 711.600 732.900 724.950 ;
        RECT 734.100 723.150 735.900 724.950 ;
        RECT 750.000 712.800 750.900 724.950 ;
        RECT 755.100 723.150 756.900 724.950 ;
        RECT 764.550 723.450 765.450 727.950 ;
        RECT 770.100 727.050 771.900 728.850 ;
        RECT 776.100 727.050 777.900 728.850 ;
        RECT 779.100 727.050 780.000 730.800 ;
        RECT 794.100 727.050 795.900 728.850 ;
        RECT 797.100 727.050 798.300 731.400 ;
        RECT 805.950 729.450 810.000 730.050 ;
        RECT 800.100 727.050 801.900 728.850 ;
        RECT 805.950 727.950 810.450 729.450 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 761.550 722.550 765.450 723.450 ;
        RECT 773.100 723.150 774.900 724.950 ;
        RECT 751.950 720.450 754.050 721.050 ;
        RECT 761.550 720.450 762.450 722.550 ;
        RECT 751.950 719.550 762.450 720.450 ;
        RECT 751.950 718.950 754.050 719.550 ;
        RECT 779.100 712.800 780.000 724.950 ;
        RECT 797.100 717.600 798.300 724.950 ;
        RECT 803.100 723.150 804.900 724.950 ;
        RECT 809.550 724.050 810.450 727.950 ;
        RECT 815.400 727.050 816.300 734.400 ;
        RECT 839.100 731.400 840.900 741.000 ;
        RECT 845.700 732.000 847.500 740.400 ;
        RECT 850.950 732.450 853.050 733.050 ;
        RECT 856.950 732.450 859.050 732.900 ;
        RECT 845.700 730.800 849.000 732.000 ;
        RECT 850.950 731.550 859.050 732.450 ;
        RECT 862.500 732.000 864.300 740.400 ;
        RECT 850.950 730.950 853.050 731.550 ;
        RECT 856.950 730.800 859.050 731.550 ;
        RECT 861.000 730.800 864.300 732.000 ;
        RECT 869.100 731.400 870.900 741.000 ;
        RECT 881.100 734.400 882.900 740.400 ;
        RECT 881.700 732.300 882.900 734.400 ;
        RECT 884.100 735.300 885.900 740.400 ;
        RECT 887.100 736.200 888.900 741.000 ;
        RECT 890.100 735.300 891.900 740.400 ;
        RECT 884.100 733.950 891.900 735.300 ;
        RECT 881.700 731.400 885.300 732.300 ;
        RECT 905.100 731.400 906.900 741.000 ;
        RECT 911.700 732.000 913.500 740.400 ;
        RECT 826.950 729.450 831.000 730.050 ;
        RECT 817.950 727.050 819.750 728.850 ;
        RECT 824.100 727.050 825.900 728.850 ;
        RECT 826.950 727.950 831.450 729.450 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 805.950 722.550 810.450 724.050 ;
        RECT 805.950 721.950 810.000 722.550 ;
        RECT 815.400 717.600 816.300 724.950 ;
        RECT 820.950 723.150 822.750 724.950 ;
        RECT 830.550 723.450 831.450 727.950 ;
        RECT 839.100 727.050 840.900 728.850 ;
        RECT 845.100 727.050 846.900 728.850 ;
        RECT 848.100 727.050 849.000 730.800 ;
        RECT 861.000 727.050 861.900 730.800 ;
        RECT 871.950 729.450 876.000 730.050 ;
        RECT 863.100 727.050 864.900 728.850 ;
        RECT 869.100 727.050 870.900 728.850 ;
        RECT 871.950 727.950 876.450 729.450 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 859.950 724.950 862.050 727.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 835.950 723.450 838.050 724.050 ;
        RECT 830.550 722.550 838.050 723.450 ;
        RECT 842.100 723.150 843.900 724.950 ;
        RECT 835.950 721.950 838.050 722.550 ;
        RECT 817.950 720.450 820.050 721.050 ;
        RECT 832.950 720.450 835.050 721.050 ;
        RECT 844.950 720.450 847.050 721.050 ;
        RECT 817.950 719.550 847.050 720.450 ;
        RECT 817.950 718.950 820.050 719.550 ;
        RECT 832.950 718.950 835.050 719.550 ;
        RECT 844.950 718.950 847.050 719.550 ;
        RECT 797.100 716.100 799.500 717.600 ;
        RECT 795.000 713.100 796.800 714.900 ;
        RECT 750.000 711.900 756.600 712.800 ;
        RECT 750.000 711.600 750.900 711.900 ;
        RECT 716.100 705.000 717.900 711.600 ;
        RECT 719.100 705.600 720.900 711.600 ;
        RECT 731.100 705.600 732.900 711.600 ;
        RECT 734.100 705.000 735.900 711.600 ;
        RECT 749.100 705.600 750.900 711.600 ;
        RECT 755.100 711.600 756.600 711.900 ;
        RECT 773.400 711.900 780.000 712.800 ;
        RECT 773.400 711.600 774.900 711.900 ;
        RECT 752.100 705.000 753.900 711.000 ;
        RECT 755.100 705.600 756.900 711.600 ;
        RECT 758.100 705.000 759.900 711.600 ;
        RECT 770.100 705.000 771.900 711.600 ;
        RECT 773.100 705.600 774.900 711.600 ;
        RECT 779.100 711.600 780.000 711.900 ;
        RECT 776.100 705.000 777.900 711.000 ;
        RECT 779.100 705.600 780.900 711.600 ;
        RECT 794.700 705.000 796.500 711.600 ;
        RECT 797.700 705.600 799.500 716.100 ;
        RECT 802.800 705.000 804.600 717.600 ;
        RECT 815.100 705.600 816.900 717.600 ;
        RECT 818.100 716.700 825.900 717.600 ;
        RECT 818.100 705.600 819.900 716.700 ;
        RECT 821.100 705.000 822.900 715.800 ;
        RECT 824.100 705.600 825.900 716.700 ;
        RECT 848.100 712.800 849.000 724.950 ;
        RECT 842.400 711.900 849.000 712.800 ;
        RECT 842.400 711.600 843.900 711.900 ;
        RECT 839.100 705.000 840.900 711.600 ;
        RECT 842.100 705.600 843.900 711.600 ;
        RECT 848.100 711.600 849.000 711.900 ;
        RECT 861.000 712.800 861.900 724.950 ;
        RECT 866.100 723.150 867.900 724.950 ;
        RECT 875.550 724.050 876.450 727.950 ;
        RECT 881.100 727.050 882.900 728.850 ;
        RECT 884.100 727.050 885.300 731.400 ;
        RECT 911.700 730.800 915.000 732.000 ;
        RECT 887.100 727.050 888.900 728.850 ;
        RECT 905.100 727.050 906.900 728.850 ;
        RECT 911.100 727.050 912.900 728.850 ;
        RECT 914.100 727.050 915.000 730.800 ;
        RECT 880.950 724.950 883.050 727.050 ;
        RECT 883.950 724.950 886.050 727.050 ;
        RECT 886.950 724.950 889.050 727.050 ;
        RECT 889.950 724.950 892.050 727.050 ;
        RECT 904.950 724.950 907.050 727.050 ;
        RECT 907.950 724.950 910.050 727.050 ;
        RECT 910.950 724.950 913.050 727.050 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 871.950 722.550 876.450 724.050 ;
        RECT 871.950 721.950 876.000 722.550 ;
        RECT 865.950 720.450 868.050 721.050 ;
        RECT 880.950 720.450 883.050 721.050 ;
        RECT 865.950 719.550 883.050 720.450 ;
        RECT 865.950 718.950 868.050 719.550 ;
        RECT 880.950 718.950 883.050 719.550 ;
        RECT 884.100 717.600 885.300 724.950 ;
        RECT 890.100 723.150 891.900 724.950 ;
        RECT 908.100 723.150 909.900 724.950 ;
        RECT 884.100 716.100 886.500 717.600 ;
        RECT 882.000 713.100 883.800 714.900 ;
        RECT 861.000 711.900 867.600 712.800 ;
        RECT 861.000 711.600 861.900 711.900 ;
        RECT 845.100 705.000 846.900 711.000 ;
        RECT 848.100 705.600 849.900 711.600 ;
        RECT 860.100 705.600 861.900 711.600 ;
        RECT 866.100 711.600 867.600 711.900 ;
        RECT 863.100 705.000 864.900 711.000 ;
        RECT 866.100 705.600 867.900 711.600 ;
        RECT 869.100 705.000 870.900 711.600 ;
        RECT 881.700 705.000 883.500 711.600 ;
        RECT 884.700 705.600 886.500 716.100 ;
        RECT 889.800 705.000 891.600 717.600 ;
        RECT 914.100 712.800 915.000 724.950 ;
        RECT 908.400 711.900 915.000 712.800 ;
        RECT 908.400 711.600 909.900 711.900 ;
        RECT 905.100 705.000 906.900 711.600 ;
        RECT 908.100 705.600 909.900 711.600 ;
        RECT 914.100 711.600 915.000 711.900 ;
        RECT 911.100 705.000 912.900 711.000 ;
        RECT 914.100 705.600 915.900 711.600 ;
        RECT 14.100 689.400 15.900 701.400 ;
        RECT 18.600 689.400 20.400 702.000 ;
        RECT 21.600 690.900 23.400 701.400 ;
        RECT 21.600 689.400 24.000 690.900 ;
        RECT 38.400 689.400 40.200 702.000 ;
        RECT 43.500 690.900 45.300 701.400 ;
        RECT 46.500 695.400 48.300 702.000 ;
        RECT 46.200 692.100 48.000 693.900 ;
        RECT 43.500 689.400 45.900 690.900 ;
        RECT 59.100 689.400 60.900 702.000 ;
        RECT 64.200 690.600 66.000 701.400 ;
        RECT 77.100 695.400 78.900 702.000 ;
        RECT 80.100 695.400 81.900 701.400 ;
        RECT 62.400 689.400 66.000 690.600 ;
        RECT 14.100 687.900 15.300 689.400 ;
        RECT 14.100 686.700 21.900 687.900 ;
        RECT 20.100 686.100 21.900 686.700 ;
        RECT 18.000 682.050 19.800 683.850 ;
        RECT 14.100 679.950 16.200 682.050 ;
        RECT 17.400 679.950 19.500 682.050 ;
        RECT 14.400 678.150 16.200 679.950 ;
        RECT 20.700 675.600 21.600 686.100 ;
        RECT 22.800 682.050 24.000 689.400 ;
        RECT 38.100 682.050 39.900 683.850 ;
        RECT 44.700 682.050 45.900 689.400 ;
        RECT 54.000 684.450 58.050 685.050 ;
        RECT 53.550 682.950 58.050 684.450 ;
        RECT 22.800 679.950 24.900 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 20.700 674.700 22.800 675.600 ;
        RECT 17.400 673.800 22.800 674.700 ;
        RECT 17.400 669.600 18.300 673.800 ;
        RECT 24.000 672.600 24.900 679.950 ;
        RECT 41.100 678.150 42.900 679.950 ;
        RECT 44.700 675.600 45.900 679.950 ;
        RECT 47.100 678.150 48.900 679.950 ;
        RECT 53.550 679.050 54.450 682.950 ;
        RECT 59.250 682.050 61.050 683.850 ;
        RECT 62.400 682.050 63.300 689.400 ;
        RECT 73.950 685.950 76.050 688.050 ;
        RECT 65.100 682.050 66.900 683.850 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 53.550 677.550 58.050 679.050 ;
        RECT 54.000 676.950 58.050 677.550 ;
        RECT 44.700 674.700 48.300 675.600 ;
        RECT 14.100 666.600 15.900 669.600 ;
        RECT 17.100 666.600 18.900 669.600 ;
        RECT 14.100 666.000 15.300 666.600 ;
        RECT 20.100 666.000 21.900 672.000 ;
        RECT 23.100 666.600 24.900 672.600 ;
        RECT 38.100 671.700 45.900 673.050 ;
        RECT 38.100 666.600 39.900 671.700 ;
        RECT 41.100 666.000 42.900 670.800 ;
        RECT 44.100 666.600 45.900 671.700 ;
        RECT 47.100 672.600 48.300 674.700 ;
        RECT 47.100 666.600 48.900 672.600 ;
        RECT 62.400 669.600 63.300 679.950 ;
        RECT 67.950 678.450 70.050 679.050 ;
        RECT 74.550 678.450 75.450 685.950 ;
        RECT 77.100 679.950 79.200 682.050 ;
        RECT 67.950 677.550 75.450 678.450 ;
        RECT 77.250 678.150 79.050 679.950 ;
        RECT 67.950 676.950 70.050 677.550 ;
        RECT 80.100 675.300 81.000 695.400 ;
        RECT 83.100 690.000 84.900 702.000 ;
        RECT 86.100 689.400 87.900 701.400 ;
        RECT 101.100 689.400 102.900 702.000 ;
        RECT 106.200 690.600 108.000 701.400 ;
        RECT 119.100 695.400 120.900 702.000 ;
        RECT 122.100 695.400 123.900 701.400 ;
        RECT 125.100 695.400 126.900 702.000 ;
        RECT 140.700 695.400 142.500 702.000 ;
        RECT 104.400 689.400 108.000 690.600 ;
        RECT 82.200 682.050 84.000 683.850 ;
        RECT 86.400 682.050 87.300 689.400 ;
        RECT 101.250 682.050 103.050 683.850 ;
        RECT 104.400 682.050 105.300 689.400 ;
        RECT 109.950 684.450 114.000 685.050 ;
        RECT 107.100 682.050 108.900 683.850 ;
        RECT 109.950 682.950 114.450 684.450 ;
        RECT 82.500 679.950 84.600 682.050 ;
        RECT 85.800 679.950 87.900 682.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 77.100 674.400 85.500 675.300 ;
        RECT 59.100 666.000 60.900 669.600 ;
        RECT 62.100 666.600 63.900 669.600 ;
        RECT 65.100 666.000 66.900 669.600 ;
        RECT 77.100 666.600 78.900 674.400 ;
        RECT 83.700 673.500 85.500 674.400 ;
        RECT 86.400 672.600 87.300 679.950 ;
        RECT 81.600 666.000 83.400 672.600 ;
        RECT 84.600 670.800 87.300 672.600 ;
        RECT 84.600 666.600 86.400 670.800 ;
        RECT 104.400 669.600 105.300 679.950 ;
        RECT 113.550 675.900 114.450 682.950 ;
        RECT 122.100 682.050 123.300 695.400 ;
        RECT 141.000 692.100 142.800 693.900 ;
        RECT 143.700 690.900 145.500 701.400 ;
        RECT 143.100 689.400 145.500 690.900 ;
        RECT 148.800 689.400 150.600 702.000 ;
        RECT 161.100 689.400 162.900 702.000 ;
        RECT 166.200 690.600 168.000 701.400 ;
        RECT 164.400 689.400 168.000 690.600 ;
        RECT 179.400 689.400 181.200 702.000 ;
        RECT 184.500 690.900 186.300 701.400 ;
        RECT 187.500 695.400 189.300 702.000 ;
        RECT 203.100 695.400 204.900 702.000 ;
        RECT 206.100 695.400 207.900 701.400 ;
        RECT 209.100 695.400 210.900 702.000 ;
        RECT 212.700 695.400 214.500 702.000 ;
        RECT 215.700 696.300 217.500 701.400 ;
        RECT 215.400 695.400 217.500 696.300 ;
        RECT 218.700 695.400 220.500 702.000 ;
        RECT 187.200 692.100 189.000 693.900 ;
        RECT 184.500 689.400 186.900 690.900 ;
        RECT 143.100 682.050 144.300 689.400 ;
        RECT 149.100 682.050 150.900 683.850 ;
        RECT 161.250 682.050 163.050 683.850 ;
        RECT 164.400 682.050 165.300 689.400 ;
        RECT 167.100 682.050 168.900 683.850 ;
        RECT 179.100 682.050 180.900 683.850 ;
        RECT 185.700 682.050 186.900 689.400 ;
        RECT 187.950 687.450 190.050 688.050 ;
        RECT 193.950 687.450 196.050 688.050 ;
        RECT 187.950 686.550 196.050 687.450 ;
        RECT 187.950 685.950 190.050 686.550 ;
        RECT 193.950 685.950 196.050 686.550 ;
        RECT 206.700 682.050 207.900 695.400 ;
        RECT 215.400 694.500 216.300 695.400 ;
        RECT 212.700 693.600 216.300 694.500 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 121.950 679.950 124.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 145.950 679.950 148.050 682.050 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 679.950 169.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 119.250 678.150 121.050 679.950 ;
        RECT 112.950 673.800 115.050 675.900 ;
        RECT 122.100 674.700 123.300 679.950 ;
        RECT 125.100 678.150 126.900 679.950 ;
        RECT 140.100 678.150 141.900 679.950 ;
        RECT 143.100 675.600 144.300 679.950 ;
        RECT 146.100 678.150 147.900 679.950 ;
        RECT 140.700 674.700 144.300 675.600 ;
        RECT 122.100 673.800 126.300 674.700 ;
        RECT 101.100 666.000 102.900 669.600 ;
        RECT 104.100 666.600 105.900 669.600 ;
        RECT 107.100 666.000 108.900 669.600 ;
        RECT 119.400 666.000 121.200 672.600 ;
        RECT 124.500 666.600 126.300 673.800 ;
        RECT 140.700 672.600 141.900 674.700 ;
        RECT 140.100 666.600 141.900 672.600 ;
        RECT 143.100 671.700 150.900 673.050 ;
        RECT 143.100 666.600 144.900 671.700 ;
        RECT 146.100 666.000 147.900 670.800 ;
        RECT 149.100 666.600 150.900 671.700 ;
        RECT 164.400 669.600 165.300 679.950 ;
        RECT 182.100 678.150 183.900 679.950 ;
        RECT 185.700 675.600 186.900 679.950 ;
        RECT 188.100 678.150 189.900 679.950 ;
        RECT 203.100 678.150 204.900 679.950 ;
        RECT 185.700 674.700 189.300 675.600 ;
        RECT 206.700 674.700 207.900 679.950 ;
        RECT 208.950 678.150 210.750 679.950 ;
        RECT 179.100 671.700 186.900 673.050 ;
        RECT 161.100 666.000 162.900 669.600 ;
        RECT 164.100 666.600 165.900 669.600 ;
        RECT 167.100 666.000 168.900 669.600 ;
        RECT 179.100 666.600 180.900 671.700 ;
        RECT 182.100 666.000 183.900 670.800 ;
        RECT 185.100 666.600 186.900 671.700 ;
        RECT 188.100 672.600 189.300 674.700 ;
        RECT 203.700 673.800 207.900 674.700 ;
        RECT 212.700 677.400 213.900 693.600 ;
        RECT 217.200 692.400 219.000 692.700 ;
        RECT 221.700 692.400 223.500 701.400 ;
        RECT 224.700 695.400 226.500 702.000 ;
        RECT 228.300 698.400 230.100 701.400 ;
        RECT 231.300 698.400 233.100 701.400 ;
        RECT 228.300 696.300 230.400 698.400 ;
        RECT 231.300 696.300 233.400 698.400 ;
        RECT 234.300 695.400 236.100 701.400 ;
        RECT 237.300 695.400 239.100 702.000 ;
        RECT 233.700 693.300 235.800 695.400 ;
        RECT 241.200 693.900 243.000 701.400 ;
        RECT 244.200 695.400 246.000 702.000 ;
        RECT 247.200 695.400 249.000 701.400 ;
        RECT 250.200 698.400 252.000 701.400 ;
        RECT 253.200 698.400 255.000 701.400 ;
        RECT 256.200 698.400 258.000 701.400 ;
        RECT 250.200 696.300 252.300 698.400 ;
        RECT 253.200 696.300 255.300 698.400 ;
        RECT 256.200 696.300 258.300 698.400 ;
        RECT 259.200 695.400 261.000 702.000 ;
        RECT 262.200 695.400 264.000 701.400 ;
        RECT 265.200 695.400 267.000 702.000 ;
        RECT 268.200 695.400 270.000 701.400 ;
        RECT 271.200 695.400 273.000 702.000 ;
        RECT 274.500 695.400 276.300 701.400 ;
        RECT 277.500 695.400 279.300 702.000 ;
        RECT 290.100 695.400 291.900 702.000 ;
        RECT 293.100 695.400 294.900 701.400 ;
        RECT 296.100 695.400 297.900 702.000 ;
        RECT 308.700 695.400 310.500 702.000 ;
        RECT 217.200 691.200 236.400 692.400 ;
        RECT 241.200 691.800 244.500 693.900 ;
        RECT 247.200 691.500 249.900 695.400 ;
        RECT 253.200 694.500 255.300 695.400 ;
        RECT 253.200 693.300 261.300 694.500 ;
        RECT 259.500 692.700 261.300 693.300 ;
        RECT 262.200 692.400 263.400 695.400 ;
        RECT 268.800 694.500 270.000 695.400 ;
        RECT 268.800 693.600 272.700 694.500 ;
        RECT 266.100 692.400 267.900 693.000 ;
        RECT 217.200 690.900 219.000 691.200 ;
        RECT 235.200 690.600 236.400 691.200 ;
        RECT 250.800 690.600 252.900 691.500 ;
        RECT 220.500 689.700 222.300 690.300 ;
        RECT 230.400 689.700 232.500 690.300 ;
        RECT 220.500 688.500 232.500 689.700 ;
        RECT 235.200 689.400 252.900 690.600 ;
        RECT 256.200 690.300 258.300 691.500 ;
        RECT 262.200 691.200 267.900 692.400 ;
        RECT 271.800 690.300 272.700 693.600 ;
        RECT 256.200 689.400 272.700 690.300 ;
        RECT 230.400 688.200 232.500 688.500 ;
        RECT 235.200 687.300 270.900 688.500 ;
        RECT 235.200 686.700 236.400 687.300 ;
        RECT 269.100 686.700 270.900 687.300 ;
        RECT 222.900 685.800 236.400 686.700 ;
        RECT 247.800 685.800 249.900 686.100 ;
        RECT 222.900 685.050 224.700 685.800 ;
        RECT 214.800 682.950 216.900 685.050 ;
        RECT 220.800 683.250 224.700 685.050 ;
        RECT 242.400 684.300 244.500 685.200 ;
        RECT 220.800 682.950 222.900 683.250 ;
        RECT 233.400 683.100 244.500 684.300 ;
        RECT 246.000 684.000 249.900 685.800 ;
        RECT 254.100 684.300 255.900 686.100 ;
        RECT 255.000 683.100 255.900 684.300 ;
        RECT 215.100 681.300 216.900 682.950 ;
        RECT 233.400 682.500 235.200 683.100 ;
        RECT 242.400 682.200 255.900 683.100 ;
        RECT 258.600 682.800 263.700 684.600 ;
        RECT 265.800 682.950 267.900 685.050 ;
        RECT 258.600 681.300 259.500 682.800 ;
        RECT 215.100 680.100 259.500 681.300 ;
        RECT 265.800 680.100 267.300 682.950 ;
        RECT 230.400 677.400 232.200 679.200 ;
        RECT 238.800 678.000 240.900 679.050 ;
        RECT 260.700 678.600 267.300 680.100 ;
        RECT 212.700 676.200 229.500 677.400 ;
        RECT 188.100 666.600 189.900 672.600 ;
        RECT 203.700 666.600 205.500 673.800 ;
        RECT 212.700 672.600 213.900 676.200 ;
        RECT 227.400 675.300 229.500 676.200 ;
        RECT 216.900 674.700 218.700 675.300 ;
        RECT 216.900 673.500 225.300 674.700 ;
        RECT 223.800 672.600 225.300 673.500 ;
        RECT 230.400 674.400 231.300 677.400 ;
        RECT 235.800 677.100 240.900 678.000 ;
        RECT 235.800 676.200 237.600 677.100 ;
        RECT 238.800 676.950 240.900 677.100 ;
        RECT 245.100 677.100 262.200 678.600 ;
        RECT 245.100 676.500 247.200 677.100 ;
        RECT 245.100 674.700 246.900 676.500 ;
        RECT 263.100 675.900 270.900 677.700 ;
        RECT 230.400 673.200 237.600 674.400 ;
        RECT 232.800 672.600 234.600 673.200 ;
        RECT 236.700 672.600 237.600 673.200 ;
        RECT 252.300 672.600 258.900 674.400 ;
        RECT 263.100 672.600 264.600 675.900 ;
        RECT 271.800 672.600 272.700 689.400 ;
        RECT 208.800 666.000 210.600 672.600 ;
        RECT 212.700 666.600 214.500 672.600 ;
        RECT 218.100 666.000 219.900 672.600 ;
        RECT 223.500 666.600 225.300 672.600 ;
        RECT 227.700 669.600 229.800 671.700 ;
        RECT 230.700 669.600 232.800 671.700 ;
        RECT 233.700 669.600 235.800 671.700 ;
        RECT 236.700 671.400 239.400 672.600 ;
        RECT 237.600 670.500 239.400 671.400 ;
        RECT 241.200 670.500 243.900 672.600 ;
        RECT 227.700 666.600 229.500 669.600 ;
        RECT 230.700 666.600 232.500 669.600 ;
        RECT 233.700 666.600 235.500 669.600 ;
        RECT 236.700 666.000 238.500 669.600 ;
        RECT 241.200 666.600 243.000 670.500 ;
        RECT 247.200 669.600 249.300 671.700 ;
        RECT 250.200 669.600 252.300 671.700 ;
        RECT 253.200 669.600 255.300 671.700 ;
        RECT 256.200 669.600 258.300 671.700 ;
        RECT 260.400 671.400 264.600 672.600 ;
        RECT 244.200 666.000 246.000 669.600 ;
        RECT 247.200 666.600 249.000 669.600 ;
        RECT 250.200 666.600 252.000 669.600 ;
        RECT 253.200 666.600 255.000 669.600 ;
        RECT 256.200 666.600 258.000 669.600 ;
        RECT 260.400 666.600 262.200 671.400 ;
        RECT 265.500 666.000 267.300 672.600 ;
        RECT 270.900 666.600 272.700 672.600 ;
        RECT 274.500 685.050 276.000 695.400 ;
        RECT 274.500 682.950 276.900 685.050 ;
        RECT 274.500 669.600 276.000 682.950 ;
        RECT 293.100 682.050 294.300 695.400 ;
        RECT 309.000 692.100 310.800 693.900 ;
        RECT 311.700 690.900 313.500 701.400 ;
        RECT 311.100 689.400 313.500 690.900 ;
        RECT 316.800 689.400 318.600 702.000 ;
        RECT 320.700 695.400 322.500 702.000 ;
        RECT 323.700 696.300 325.500 701.400 ;
        RECT 323.400 695.400 325.500 696.300 ;
        RECT 326.700 695.400 328.500 702.000 ;
        RECT 323.400 694.500 324.300 695.400 ;
        RECT 320.700 693.600 324.300 694.500 ;
        RECT 311.100 682.050 312.300 689.400 ;
        RECT 317.100 682.050 318.900 683.850 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 290.250 678.150 292.050 679.950 ;
        RECT 293.100 674.700 294.300 679.950 ;
        RECT 296.100 678.150 297.900 679.950 ;
        RECT 308.100 678.150 309.900 679.950 ;
        RECT 311.100 675.600 312.300 679.950 ;
        RECT 314.100 678.150 315.900 679.950 ;
        RECT 308.700 674.700 312.300 675.600 ;
        RECT 320.700 677.400 321.900 693.600 ;
        RECT 325.200 692.400 327.000 692.700 ;
        RECT 329.700 692.400 331.500 701.400 ;
        RECT 332.700 695.400 334.500 702.000 ;
        RECT 336.300 698.400 338.100 701.400 ;
        RECT 339.300 698.400 341.100 701.400 ;
        RECT 336.300 696.300 338.400 698.400 ;
        RECT 339.300 696.300 341.400 698.400 ;
        RECT 342.300 695.400 344.100 701.400 ;
        RECT 345.300 695.400 347.100 702.000 ;
        RECT 341.700 693.300 343.800 695.400 ;
        RECT 349.200 693.900 351.000 701.400 ;
        RECT 352.200 695.400 354.000 702.000 ;
        RECT 355.200 695.400 357.000 701.400 ;
        RECT 358.200 698.400 360.000 701.400 ;
        RECT 361.200 698.400 363.000 701.400 ;
        RECT 364.200 698.400 366.000 701.400 ;
        RECT 358.200 696.300 360.300 698.400 ;
        RECT 361.200 696.300 363.300 698.400 ;
        RECT 364.200 696.300 366.300 698.400 ;
        RECT 367.200 695.400 369.000 702.000 ;
        RECT 370.200 695.400 372.000 701.400 ;
        RECT 373.200 695.400 375.000 702.000 ;
        RECT 376.200 695.400 378.000 701.400 ;
        RECT 379.200 695.400 381.000 702.000 ;
        RECT 382.500 695.400 384.300 701.400 ;
        RECT 385.500 695.400 387.300 702.000 ;
        RECT 398.100 695.400 399.900 702.000 ;
        RECT 401.100 695.400 402.900 701.400 ;
        RECT 404.100 695.400 405.900 702.000 ;
        RECT 419.700 695.400 421.500 702.000 ;
        RECT 325.200 691.200 344.400 692.400 ;
        RECT 349.200 691.800 352.500 693.900 ;
        RECT 355.200 691.500 357.900 695.400 ;
        RECT 361.200 694.500 363.300 695.400 ;
        RECT 361.200 693.300 369.300 694.500 ;
        RECT 367.500 692.700 369.300 693.300 ;
        RECT 370.200 692.400 371.400 695.400 ;
        RECT 376.800 694.500 378.000 695.400 ;
        RECT 376.800 693.600 380.700 694.500 ;
        RECT 374.100 692.400 375.900 693.000 ;
        RECT 325.200 690.900 327.000 691.200 ;
        RECT 343.200 690.600 344.400 691.200 ;
        RECT 358.800 690.600 360.900 691.500 ;
        RECT 328.500 689.700 330.300 690.300 ;
        RECT 338.400 689.700 340.500 690.300 ;
        RECT 328.500 688.500 340.500 689.700 ;
        RECT 343.200 689.400 360.900 690.600 ;
        RECT 364.200 690.300 366.300 691.500 ;
        RECT 370.200 691.200 375.900 692.400 ;
        RECT 379.800 690.300 380.700 693.600 ;
        RECT 364.200 689.400 380.700 690.300 ;
        RECT 338.400 688.200 340.500 688.500 ;
        RECT 343.200 687.300 378.900 688.500 ;
        RECT 343.200 686.700 344.400 687.300 ;
        RECT 377.100 686.700 378.900 687.300 ;
        RECT 330.900 685.800 344.400 686.700 ;
        RECT 355.800 685.800 357.900 686.100 ;
        RECT 330.900 685.050 332.700 685.800 ;
        RECT 322.800 682.950 324.900 685.050 ;
        RECT 328.800 683.250 332.700 685.050 ;
        RECT 350.400 684.300 352.500 685.200 ;
        RECT 328.800 682.950 330.900 683.250 ;
        RECT 341.400 683.100 352.500 684.300 ;
        RECT 354.000 684.000 357.900 685.800 ;
        RECT 362.100 684.300 363.900 686.100 ;
        RECT 363.000 683.100 363.900 684.300 ;
        RECT 323.100 681.300 324.900 682.950 ;
        RECT 341.400 682.500 343.200 683.100 ;
        RECT 350.400 682.200 363.900 683.100 ;
        RECT 366.600 682.800 371.700 684.600 ;
        RECT 373.800 682.950 375.900 685.050 ;
        RECT 366.600 681.300 367.500 682.800 ;
        RECT 323.100 680.100 367.500 681.300 ;
        RECT 373.800 680.100 375.300 682.950 ;
        RECT 338.400 677.400 340.200 679.200 ;
        RECT 346.800 678.000 348.900 679.050 ;
        RECT 368.700 678.600 375.300 680.100 ;
        RECT 320.700 676.200 337.500 677.400 ;
        RECT 293.100 673.800 297.300 674.700 ;
        RECT 274.500 666.600 276.300 669.600 ;
        RECT 277.500 666.000 279.300 669.600 ;
        RECT 290.400 666.000 292.200 672.600 ;
        RECT 295.500 666.600 297.300 673.800 ;
        RECT 308.700 672.600 309.900 674.700 ;
        RECT 308.100 666.600 309.900 672.600 ;
        RECT 311.100 671.700 318.900 673.050 ;
        RECT 311.100 666.600 312.900 671.700 ;
        RECT 314.100 666.000 315.900 670.800 ;
        RECT 317.100 666.600 318.900 671.700 ;
        RECT 320.700 672.600 321.900 676.200 ;
        RECT 335.400 675.300 337.500 676.200 ;
        RECT 324.900 674.700 326.700 675.300 ;
        RECT 324.900 673.500 333.300 674.700 ;
        RECT 331.800 672.600 333.300 673.500 ;
        RECT 338.400 674.400 339.300 677.400 ;
        RECT 343.800 677.100 348.900 678.000 ;
        RECT 343.800 676.200 345.600 677.100 ;
        RECT 346.800 676.950 348.900 677.100 ;
        RECT 353.100 677.100 370.200 678.600 ;
        RECT 353.100 676.500 355.200 677.100 ;
        RECT 353.100 674.700 354.900 676.500 ;
        RECT 371.100 675.900 378.900 677.700 ;
        RECT 338.400 673.200 345.600 674.400 ;
        RECT 340.800 672.600 342.600 673.200 ;
        RECT 344.700 672.600 345.600 673.200 ;
        RECT 360.300 672.600 366.900 674.400 ;
        RECT 371.100 672.600 372.600 675.900 ;
        RECT 379.800 672.600 380.700 689.400 ;
        RECT 320.700 666.600 322.500 672.600 ;
        RECT 326.100 666.000 327.900 672.600 ;
        RECT 331.500 666.600 333.300 672.600 ;
        RECT 335.700 669.600 337.800 671.700 ;
        RECT 338.700 669.600 340.800 671.700 ;
        RECT 341.700 669.600 343.800 671.700 ;
        RECT 344.700 671.400 347.400 672.600 ;
        RECT 345.600 670.500 347.400 671.400 ;
        RECT 349.200 670.500 351.900 672.600 ;
        RECT 335.700 666.600 337.500 669.600 ;
        RECT 338.700 666.600 340.500 669.600 ;
        RECT 341.700 666.600 343.500 669.600 ;
        RECT 344.700 666.000 346.500 669.600 ;
        RECT 349.200 666.600 351.000 670.500 ;
        RECT 355.200 669.600 357.300 671.700 ;
        RECT 358.200 669.600 360.300 671.700 ;
        RECT 361.200 669.600 363.300 671.700 ;
        RECT 364.200 669.600 366.300 671.700 ;
        RECT 368.400 671.400 372.600 672.600 ;
        RECT 352.200 666.000 354.000 669.600 ;
        RECT 355.200 666.600 357.000 669.600 ;
        RECT 358.200 666.600 360.000 669.600 ;
        RECT 361.200 666.600 363.000 669.600 ;
        RECT 364.200 666.600 366.000 669.600 ;
        RECT 368.400 666.600 370.200 671.400 ;
        RECT 373.500 666.000 375.300 672.600 ;
        RECT 378.900 666.600 380.700 672.600 ;
        RECT 382.500 685.050 384.000 695.400 ;
        RECT 382.500 682.950 384.900 685.050 ;
        RECT 382.500 669.600 384.000 682.950 ;
        RECT 401.700 682.050 402.900 695.400 ;
        RECT 420.000 692.100 421.800 693.900 ;
        RECT 422.700 690.900 424.500 701.400 ;
        RECT 422.100 689.400 424.500 690.900 ;
        RECT 427.800 689.400 429.600 702.000 ;
        RECT 443.100 689.400 444.900 701.400 ;
        RECT 446.100 690.000 447.900 702.000 ;
        RECT 449.100 695.400 450.900 701.400 ;
        RECT 452.100 695.400 453.900 702.000 ;
        RECT 464.100 695.400 465.900 702.000 ;
        RECT 467.100 695.400 468.900 701.400 ;
        RECT 470.100 695.400 471.900 702.000 ;
        RECT 482.100 695.400 483.900 702.000 ;
        RECT 485.100 695.400 486.900 701.400 ;
        RECT 422.100 682.050 423.300 689.400 ;
        RECT 424.950 687.450 427.050 688.050 ;
        RECT 433.950 687.450 436.050 688.050 ;
        RECT 424.950 686.550 436.050 687.450 ;
        RECT 424.950 685.950 427.050 686.550 ;
        RECT 433.950 685.950 436.050 686.550 ;
        RECT 428.100 682.050 429.900 683.850 ;
        RECT 443.700 682.050 444.600 689.400 ;
        RECT 447.000 682.050 448.800 683.850 ;
        RECT 397.950 679.950 400.050 682.050 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 443.100 679.950 445.200 682.050 ;
        RECT 446.400 679.950 448.500 682.050 ;
        RECT 398.100 678.150 399.900 679.950 ;
        RECT 401.700 674.700 402.900 679.950 ;
        RECT 403.950 678.150 405.750 679.950 ;
        RECT 419.100 678.150 420.900 679.950 ;
        RECT 398.700 673.800 402.900 674.700 ;
        RECT 403.950 675.450 406.050 676.050 ;
        RECT 412.950 675.450 415.050 676.050 ;
        RECT 422.100 675.600 423.300 679.950 ;
        RECT 425.100 678.150 426.900 679.950 ;
        RECT 403.950 674.550 415.050 675.450 ;
        RECT 403.950 673.950 406.050 674.550 ;
        RECT 412.950 673.950 415.050 674.550 ;
        RECT 419.700 674.700 423.300 675.600 ;
        RECT 382.500 666.600 384.300 669.600 ;
        RECT 385.500 666.000 387.300 669.600 ;
        RECT 398.700 666.600 400.500 673.800 ;
        RECT 419.700 672.600 420.900 674.700 ;
        RECT 403.800 666.000 405.600 672.600 ;
        RECT 419.100 666.600 420.900 672.600 ;
        RECT 422.100 671.700 429.900 673.050 ;
        RECT 422.100 666.600 423.900 671.700 ;
        RECT 425.100 666.000 426.900 670.800 ;
        RECT 428.100 666.600 429.900 671.700 ;
        RECT 443.700 672.600 444.600 679.950 ;
        RECT 450.000 675.300 450.900 695.400 ;
        RECT 467.100 682.050 468.300 695.400 ;
        RECT 482.100 682.050 483.900 683.850 ;
        RECT 485.100 682.050 486.300 695.400 ;
        RECT 501.000 690.600 502.800 701.400 ;
        RECT 501.000 689.400 504.600 690.600 ;
        RECT 506.100 689.400 507.900 702.000 ;
        RECT 521.700 695.400 523.500 702.000 ;
        RECT 522.000 692.100 523.800 693.900 ;
        RECT 524.700 690.900 526.500 701.400 ;
        RECT 524.100 689.400 526.500 690.900 ;
        RECT 529.800 689.400 531.600 702.000 ;
        RECT 542.100 689.400 543.900 701.400 ;
        RECT 545.100 691.200 546.900 702.000 ;
        RECT 548.100 695.400 549.900 701.400 ;
        RECT 500.100 682.050 501.900 683.850 ;
        RECT 503.700 682.050 504.600 689.400 ;
        RECT 505.950 682.050 507.750 683.850 ;
        RECT 524.100 682.050 525.300 689.400 ;
        RECT 530.100 682.050 531.900 683.850 ;
        RECT 542.100 682.050 543.300 689.400 ;
        RECT 548.700 688.500 549.900 695.400 ;
        RECT 560.100 689.400 561.900 701.400 ;
        RECT 563.100 690.300 564.900 701.400 ;
        RECT 566.100 691.200 567.900 702.000 ;
        RECT 569.100 690.300 570.900 701.400 ;
        RECT 581.100 695.400 582.900 702.000 ;
        RECT 584.100 695.400 585.900 701.400 ;
        RECT 587.100 696.000 588.900 702.000 ;
        RECT 584.400 695.100 585.900 695.400 ;
        RECT 590.100 695.400 591.900 701.400 ;
        RECT 605.100 695.400 606.900 702.000 ;
        RECT 608.100 695.400 609.900 701.400 ;
        RECT 623.100 695.400 624.900 702.000 ;
        RECT 626.100 695.400 627.900 701.400 ;
        RECT 629.100 695.400 630.900 702.000 ;
        RECT 641.100 695.400 642.900 702.000 ;
        RECT 644.100 695.400 645.900 701.400 ;
        RECT 647.100 695.400 648.900 702.000 ;
        RECT 662.100 695.400 663.900 702.000 ;
        RECT 665.100 695.400 666.900 701.400 ;
        RECT 668.100 695.400 669.900 702.000 ;
        RECT 683.100 695.400 684.900 701.400 ;
        RECT 686.100 695.400 687.900 702.000 ;
        RECT 698.100 700.500 705.900 701.400 ;
        RECT 590.100 695.100 591.000 695.400 ;
        RECT 584.400 694.200 591.000 695.100 ;
        RECT 563.100 689.400 570.900 690.300 ;
        RECT 544.200 687.600 549.900 688.500 ;
        RECT 544.200 686.700 546.000 687.600 ;
        RECT 451.800 679.950 453.900 682.050 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 520.950 679.950 523.050 682.050 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 542.100 679.950 544.200 682.050 ;
        RECT 451.950 678.150 453.750 679.950 ;
        RECT 464.250 678.150 466.050 679.950 ;
        RECT 445.500 674.400 453.900 675.300 ;
        RECT 445.500 673.500 447.300 674.400 ;
        RECT 443.700 670.800 446.400 672.600 ;
        RECT 444.600 666.600 446.400 670.800 ;
        RECT 447.600 666.000 449.400 672.600 ;
        RECT 452.100 666.600 453.900 674.400 ;
        RECT 467.100 674.700 468.300 679.950 ;
        RECT 470.100 678.150 471.900 679.950 ;
        RECT 467.100 673.800 471.300 674.700 ;
        RECT 464.400 666.000 466.200 672.600 ;
        RECT 469.500 666.600 471.300 673.800 ;
        RECT 485.100 669.600 486.300 679.950 ;
        RECT 503.700 669.600 504.600 679.950 ;
        RECT 508.950 678.450 511.050 679.050 ;
        RECT 514.950 678.450 517.050 679.050 ;
        RECT 508.950 677.550 517.050 678.450 ;
        RECT 521.100 678.150 522.900 679.950 ;
        RECT 508.950 676.950 511.050 677.550 ;
        RECT 514.950 676.950 517.050 677.550 ;
        RECT 524.100 675.600 525.300 679.950 ;
        RECT 527.100 678.150 528.900 679.950 ;
        RECT 521.700 674.700 525.300 675.600 ;
        RECT 521.700 672.600 522.900 674.700 ;
        RECT 482.100 666.000 483.900 669.600 ;
        RECT 485.100 666.600 486.900 669.600 ;
        RECT 500.100 666.000 501.900 669.600 ;
        RECT 503.100 666.600 504.900 669.600 ;
        RECT 506.100 666.000 507.900 669.600 ;
        RECT 521.100 666.600 522.900 672.600 ;
        RECT 524.100 671.700 531.900 673.050 ;
        RECT 524.100 666.600 525.900 671.700 ;
        RECT 527.100 666.000 528.900 670.800 ;
        RECT 530.100 666.600 531.900 671.700 ;
        RECT 542.100 672.600 543.300 679.950 ;
        RECT 545.100 675.300 546.000 686.700 ;
        RECT 547.800 682.050 549.600 683.850 ;
        RECT 560.400 682.050 561.300 689.400 ;
        RECT 568.950 687.450 571.050 688.050 ;
        RECT 580.950 687.450 583.050 688.200 ;
        RECT 586.950 687.450 589.050 688.050 ;
        RECT 568.950 686.550 589.050 687.450 ;
        RECT 568.950 685.950 571.050 686.550 ;
        RECT 580.950 686.100 583.050 686.550 ;
        RECT 586.950 685.950 589.050 686.550 ;
        RECT 565.950 682.050 567.750 683.850 ;
        RECT 584.100 682.050 585.900 683.850 ;
        RECT 590.100 682.050 591.000 694.200 ;
        RECT 605.100 682.050 606.900 683.850 ;
        RECT 608.100 682.050 609.300 695.400 ;
        RECT 626.100 682.050 627.300 695.400 ;
        RECT 636.000 684.450 640.050 685.050 ;
        RECT 635.550 682.950 640.050 684.450 ;
        RECT 547.500 679.950 549.600 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 607.950 679.950 610.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 628.950 679.950 631.050 682.050 ;
        RECT 544.200 674.400 546.000 675.300 ;
        RECT 544.200 673.500 549.900 674.400 ;
        RECT 542.100 666.600 543.900 672.600 ;
        RECT 545.100 666.000 546.900 672.600 ;
        RECT 548.700 669.600 549.900 673.500 ;
        RECT 560.400 672.600 561.300 679.950 ;
        RECT 562.950 678.150 564.750 679.950 ;
        RECT 569.100 678.150 570.900 679.950 ;
        RECT 581.100 678.150 582.900 679.950 ;
        RECT 587.100 678.150 588.900 679.950 ;
        RECT 590.100 676.200 591.000 679.950 ;
        RECT 562.950 675.450 565.050 676.050 ;
        RECT 574.950 675.450 577.050 676.050 ;
        RECT 562.950 674.550 577.050 675.450 ;
        RECT 562.950 673.950 565.050 674.550 ;
        RECT 574.950 673.950 577.050 674.550 ;
        RECT 560.400 671.400 565.500 672.600 ;
        RECT 548.100 666.600 549.900 669.600 ;
        RECT 560.700 666.000 562.500 669.600 ;
        RECT 563.700 666.600 565.500 671.400 ;
        RECT 568.200 666.000 570.000 672.600 ;
        RECT 581.100 666.000 582.900 675.600 ;
        RECT 587.700 675.000 591.000 676.200 ;
        RECT 592.950 675.450 595.050 676.050 ;
        RECT 604.950 675.450 607.050 676.050 ;
        RECT 587.700 666.600 589.500 675.000 ;
        RECT 592.950 674.550 607.050 675.450 ;
        RECT 592.950 673.950 595.050 674.550 ;
        RECT 604.950 673.950 607.050 674.550 ;
        RECT 608.100 669.600 609.300 679.950 ;
        RECT 623.250 678.150 625.050 679.950 ;
        RECT 626.100 674.700 627.300 679.950 ;
        RECT 629.100 678.150 630.900 679.950 ;
        RECT 635.550 679.050 636.450 682.950 ;
        RECT 644.700 682.050 645.900 695.400 ;
        RECT 665.100 682.050 666.300 695.400 ;
        RECT 683.700 682.050 684.900 695.400 ;
        RECT 698.100 691.200 699.900 700.500 ;
        RECT 701.100 691.800 702.900 699.600 ;
        RECT 688.950 684.450 691.050 685.050 ;
        RECT 697.950 684.450 700.050 685.050 ;
        RECT 686.100 682.050 687.900 683.850 ;
        RECT 688.950 683.550 700.050 684.450 ;
        RECT 688.950 682.950 691.050 683.550 ;
        RECT 697.950 682.950 700.050 683.550 ;
        RECT 701.700 682.050 702.900 691.800 ;
        RECT 704.100 691.800 705.900 700.500 ;
        RECT 707.100 700.500 714.900 701.400 ;
        RECT 707.100 692.700 708.900 700.500 ;
        RECT 710.100 691.800 711.900 699.600 ;
        RECT 704.100 690.900 711.900 691.800 ;
        RECT 713.100 691.500 714.900 700.500 ;
        RECT 716.100 692.400 717.900 702.000 ;
        RECT 719.100 691.500 720.900 701.400 ;
        RECT 731.700 695.400 733.500 702.000 ;
        RECT 732.000 692.100 733.800 693.900 ;
        RECT 713.100 690.600 720.900 691.500 ;
        RECT 734.700 690.900 736.500 701.400 ;
        RECT 734.100 689.400 736.500 690.900 ;
        RECT 739.800 689.400 741.600 702.000 ;
        RECT 755.100 695.400 756.900 702.000 ;
        RECT 758.100 695.400 759.900 701.400 ;
        RECT 773.100 695.400 774.900 702.000 ;
        RECT 776.100 695.400 777.900 701.400 ;
        RECT 779.100 696.000 780.900 702.000 ;
        RECT 718.950 687.450 721.050 688.050 ;
        RECT 724.950 687.450 727.050 688.050 ;
        RECT 718.950 686.550 727.050 687.450 ;
        RECT 718.950 685.950 721.050 686.550 ;
        RECT 724.950 685.950 727.050 686.550 ;
        RECT 706.950 682.050 708.750 683.850 ;
        RECT 716.100 682.050 717.900 683.850 ;
        RECT 734.100 682.050 735.300 689.400 ;
        RECT 740.100 682.050 741.900 683.850 ;
        RECT 755.100 682.050 756.900 683.850 ;
        RECT 758.100 682.050 759.300 695.400 ;
        RECT 776.400 695.100 777.900 695.400 ;
        RECT 782.100 695.400 783.900 701.400 ;
        RECT 797.100 695.400 798.900 702.000 ;
        RECT 800.100 695.400 801.900 701.400 ;
        RECT 803.100 695.400 804.900 702.000 ;
        RECT 782.100 695.100 783.000 695.400 ;
        RECT 776.400 694.200 783.000 695.100 ;
        RECT 776.100 682.050 777.900 683.850 ;
        RECT 782.100 682.050 783.000 694.200 ;
        RECT 800.700 682.050 801.900 695.400 ;
        RECT 818.100 690.300 819.900 701.400 ;
        RECT 821.100 691.200 822.900 702.000 ;
        RECT 824.100 690.300 825.900 701.400 ;
        RECT 818.100 689.400 825.900 690.300 ;
        RECT 827.100 689.400 828.900 701.400 ;
        RECT 839.100 695.400 840.900 702.000 ;
        RECT 842.100 695.400 843.900 701.400 ;
        RECT 845.100 696.000 846.900 702.000 ;
        RECT 842.400 695.100 843.900 695.400 ;
        RECT 848.100 695.400 849.900 701.400 ;
        RECT 860.100 695.400 861.900 702.000 ;
        RECT 863.100 695.400 864.900 701.400 ;
        RECT 866.100 695.400 867.900 702.000 ;
        RECT 878.100 695.400 879.900 701.400 ;
        RECT 881.100 696.000 882.900 702.000 ;
        RECT 848.100 695.100 849.000 695.400 ;
        RECT 842.400 694.200 849.000 695.100 ;
        RECT 813.000 684.450 817.050 685.050 ;
        RECT 812.550 682.950 817.050 684.450 ;
        RECT 640.950 679.950 643.050 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 664.950 679.950 667.050 682.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 701.400 679.950 703.500 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 716.100 679.950 718.200 682.050 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 733.950 679.950 736.050 682.050 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 631.950 677.550 636.450 679.050 ;
        RECT 641.100 678.150 642.900 679.950 ;
        RECT 631.950 676.950 636.000 677.550 ;
        RECT 644.700 674.700 645.900 679.950 ;
        RECT 646.950 678.150 648.750 679.950 ;
        RECT 662.250 678.150 664.050 679.950 ;
        RECT 626.100 673.800 630.300 674.700 ;
        RECT 605.100 666.000 606.900 669.600 ;
        RECT 608.100 666.600 609.900 669.600 ;
        RECT 623.400 666.000 625.200 672.600 ;
        RECT 628.500 666.600 630.300 673.800 ;
        RECT 641.700 673.800 645.900 674.700 ;
        RECT 665.100 674.700 666.300 679.950 ;
        RECT 668.100 678.150 669.900 679.950 ;
        RECT 665.100 673.800 669.300 674.700 ;
        RECT 641.700 666.600 643.500 673.800 ;
        RECT 646.800 666.000 648.600 672.600 ;
        RECT 662.400 666.000 664.200 672.600 ;
        RECT 667.500 666.600 669.300 673.800 ;
        RECT 683.700 669.600 684.900 679.950 ;
        RECT 701.700 671.400 702.900 679.950 ;
        RECT 710.250 678.150 712.050 679.950 ;
        RECT 731.100 678.150 732.900 679.950 ;
        RECT 706.950 675.450 709.050 676.050 ;
        RECT 721.950 675.450 724.050 676.050 ;
        RECT 727.950 675.450 730.050 676.050 ;
        RECT 734.100 675.600 735.300 679.950 ;
        RECT 737.100 678.150 738.900 679.950 ;
        RECT 706.950 674.550 730.050 675.450 ;
        RECT 706.950 673.950 709.050 674.550 ;
        RECT 721.950 673.950 724.050 674.550 ;
        RECT 727.950 673.950 730.050 674.550 ;
        RECT 731.700 674.700 735.300 675.600 ;
        RECT 731.700 672.600 732.900 674.700 ;
        RECT 701.700 670.500 714.300 671.400 ;
        RECT 706.200 669.600 707.100 670.500 ;
        RECT 713.400 669.600 714.300 670.500 ;
        RECT 683.100 666.600 684.900 669.600 ;
        RECT 686.100 666.000 687.900 669.600 ;
        RECT 706.200 666.600 708.900 669.600 ;
        RECT 710.100 666.000 711.900 669.600 ;
        RECT 713.100 666.600 714.900 669.600 ;
        RECT 716.100 666.000 718.200 669.600 ;
        RECT 731.100 666.600 732.900 672.600 ;
        RECT 734.100 671.700 741.900 673.050 ;
        RECT 734.100 666.600 735.900 671.700 ;
        RECT 737.100 666.000 738.900 670.800 ;
        RECT 740.100 666.600 741.900 671.700 ;
        RECT 758.100 669.600 759.300 679.950 ;
        RECT 773.100 678.150 774.900 679.950 ;
        RECT 779.100 678.150 780.900 679.950 ;
        RECT 782.100 676.200 783.000 679.950 ;
        RECT 797.100 678.150 798.900 679.950 ;
        RECT 755.100 666.000 756.900 669.600 ;
        RECT 758.100 666.600 759.900 669.600 ;
        RECT 773.100 666.000 774.900 675.600 ;
        RECT 779.700 675.000 783.000 676.200 ;
        RECT 779.700 666.600 781.500 675.000 ;
        RECT 800.700 674.700 801.900 679.950 ;
        RECT 802.950 678.150 804.750 679.950 ;
        RECT 797.700 673.800 801.900 674.700 ;
        RECT 802.950 675.450 805.050 676.050 ;
        RECT 812.550 675.450 813.450 682.950 ;
        RECT 821.250 682.050 823.050 683.850 ;
        RECT 827.700 682.050 828.600 689.400 ;
        RECT 829.950 687.450 832.050 688.050 ;
        RECT 838.950 687.450 841.050 688.200 ;
        RECT 844.950 687.450 847.050 688.050 ;
        RECT 829.950 686.550 847.050 687.450 ;
        RECT 829.950 685.950 832.050 686.550 ;
        RECT 838.950 686.100 841.050 686.550 ;
        RECT 844.950 685.950 847.050 686.550 ;
        RECT 842.100 682.050 843.900 683.850 ;
        RECT 848.100 682.050 849.000 694.200 ;
        RECT 863.100 682.050 864.300 695.400 ;
        RECT 879.000 695.100 879.900 695.400 ;
        RECT 884.100 695.400 885.900 701.400 ;
        RECT 887.100 695.400 888.900 702.000 ;
        RECT 884.100 695.100 885.600 695.400 ;
        RECT 879.000 694.200 885.600 695.100 ;
        RECT 873.000 684.450 877.050 685.050 ;
        RECT 872.550 682.950 877.050 684.450 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 823.950 679.950 826.050 682.050 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 844.950 679.950 847.050 682.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 818.100 678.150 819.900 679.950 ;
        RECT 824.250 678.150 826.050 679.950 ;
        RECT 802.950 674.550 813.450 675.450 ;
        RECT 802.950 673.950 805.050 674.550 ;
        RECT 797.700 666.600 799.500 673.800 ;
        RECT 827.700 672.600 828.600 679.950 ;
        RECT 839.100 678.150 840.900 679.950 ;
        RECT 845.100 678.150 846.900 679.950 ;
        RECT 848.100 676.200 849.000 679.950 ;
        RECT 860.250 678.150 862.050 679.950 ;
        RECT 802.800 666.000 804.600 672.600 ;
        RECT 819.000 666.000 820.800 672.600 ;
        RECT 823.500 671.400 828.600 672.600 ;
        RECT 823.500 666.600 825.300 671.400 ;
        RECT 826.500 666.000 828.300 669.600 ;
        RECT 839.100 666.000 840.900 675.600 ;
        RECT 845.700 675.000 849.000 676.200 ;
        RECT 845.700 666.600 847.500 675.000 ;
        RECT 863.100 674.700 864.300 679.950 ;
        RECT 866.100 678.150 867.900 679.950 ;
        RECT 872.550 679.050 873.450 682.950 ;
        RECT 879.000 682.050 879.900 694.200 ;
        RECT 886.950 690.450 889.050 691.050 ;
        RECT 895.950 690.450 898.050 691.050 ;
        RECT 886.950 689.550 898.050 690.450 ;
        RECT 886.950 688.950 889.050 689.550 ;
        RECT 895.950 688.950 898.050 689.550 ;
        RECT 899.100 690.300 900.900 701.400 ;
        RECT 902.100 691.200 903.900 702.000 ;
        RECT 905.100 690.300 906.900 701.400 ;
        RECT 899.100 689.400 906.900 690.300 ;
        RECT 908.100 689.400 909.900 701.400 ;
        RECT 923.100 695.400 924.900 701.400 ;
        RECT 926.100 696.000 927.900 702.000 ;
        RECT 924.000 695.100 924.900 695.400 ;
        RECT 929.100 695.400 930.900 701.400 ;
        RECT 932.100 695.400 933.900 702.000 ;
        RECT 929.100 695.100 930.600 695.400 ;
        RECT 924.000 694.200 930.600 695.100 ;
        RECT 883.950 687.450 886.050 688.050 ;
        RECT 883.950 686.550 894.450 687.450 ;
        RECT 883.950 685.950 886.050 686.550 ;
        RECT 884.100 682.050 885.900 683.850 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 868.950 677.550 873.450 679.050 ;
        RECT 868.950 676.950 873.000 677.550 ;
        RECT 879.000 676.200 879.900 679.950 ;
        RECT 881.100 678.150 882.900 679.950 ;
        RECT 887.100 678.150 888.900 679.950 ;
        RECT 893.550 679.050 894.450 686.550 ;
        RECT 902.250 682.050 904.050 683.850 ;
        RECT 908.700 682.050 909.600 689.400 ;
        RECT 918.000 684.450 922.050 685.050 ;
        RECT 917.550 682.950 922.050 684.450 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 889.950 677.550 894.450 679.050 ;
        RECT 899.100 678.150 900.900 679.950 ;
        RECT 905.250 678.150 907.050 679.950 ;
        RECT 889.950 676.950 894.000 677.550 ;
        RECT 879.000 675.000 882.300 676.200 ;
        RECT 863.100 673.800 867.300 674.700 ;
        RECT 860.400 666.000 862.200 672.600 ;
        RECT 865.500 666.600 867.300 673.800 ;
        RECT 880.500 666.600 882.300 675.000 ;
        RECT 887.100 666.000 888.900 675.600 ;
        RECT 908.700 672.600 909.600 679.950 ;
        RECT 917.550 679.050 918.450 682.950 ;
        RECT 924.000 682.050 924.900 694.200 ;
        RECT 929.100 682.050 930.900 683.850 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 925.950 679.950 928.050 682.050 ;
        RECT 928.950 679.950 931.050 682.050 ;
        RECT 931.950 679.950 934.050 682.050 ;
        RECT 917.550 677.550 922.050 679.050 ;
        RECT 918.000 676.950 922.050 677.550 ;
        RECT 924.000 676.200 924.900 679.950 ;
        RECT 926.100 678.150 927.900 679.950 ;
        RECT 932.100 678.150 933.900 679.950 ;
        RECT 924.000 675.000 927.300 676.200 ;
        RECT 900.000 666.000 901.800 672.600 ;
        RECT 904.500 671.400 909.600 672.600 ;
        RECT 904.500 666.600 906.300 671.400 ;
        RECT 907.500 666.000 909.300 669.600 ;
        RECT 925.500 666.600 927.300 675.000 ;
        RECT 932.100 666.000 933.900 675.600 ;
        RECT 14.100 659.400 15.900 663.000 ;
        RECT 17.100 659.400 18.900 662.400 ;
        RECT 20.100 659.400 21.900 663.000 ;
        RECT 35.100 659.400 36.900 663.000 ;
        RECT 38.100 659.400 39.900 662.400 ;
        RECT 17.400 649.050 18.300 659.400 ;
        RECT 38.100 649.050 39.300 659.400 ;
        RECT 50.100 657.300 51.900 662.400 ;
        RECT 53.100 658.200 54.900 663.000 ;
        RECT 56.100 657.300 57.900 662.400 ;
        RECT 50.100 655.950 57.900 657.300 ;
        RECT 59.100 656.400 60.900 662.400 ;
        RECT 71.100 659.400 72.900 662.400 ;
        RECT 74.100 659.400 75.900 663.000 ;
        RECT 86.100 659.400 87.900 663.000 ;
        RECT 89.100 659.400 90.900 662.400 ;
        RECT 92.100 659.400 93.900 663.000 ;
        RECT 104.100 659.400 105.900 663.000 ;
        RECT 107.100 659.400 108.900 662.400 ;
        RECT 122.100 659.400 123.900 663.000 ;
        RECT 125.100 659.400 126.900 662.400 ;
        RECT 128.100 659.400 129.900 663.000 ;
        RECT 140.100 659.400 141.900 662.400 ;
        RECT 143.100 659.400 144.900 663.000 ;
        RECT 158.100 659.400 159.900 663.000 ;
        RECT 161.100 659.400 162.900 662.400 ;
        RECT 164.100 659.400 165.900 663.000 ;
        RECT 59.100 654.300 60.300 656.400 ;
        RECT 56.700 653.400 60.300 654.300 ;
        RECT 53.100 649.050 54.900 650.850 ;
        RECT 56.700 649.050 57.900 653.400 ;
        RECT 59.100 649.050 60.900 650.850 ;
        RECT 71.700 649.050 72.900 659.400 ;
        RECT 89.700 649.050 90.600 659.400 ;
        RECT 107.100 649.050 108.300 659.400 ;
        RECT 125.400 649.050 126.300 659.400 ;
        RECT 140.700 649.050 141.900 659.400 ;
        RECT 161.700 649.050 162.600 659.400 ;
        RECT 178.500 656.400 180.300 663.000 ;
        RECT 183.000 656.400 184.800 662.400 ;
        RECT 187.500 656.400 189.300 663.000 ;
        RECT 200.100 656.400 201.900 663.000 ;
        RECT 203.100 656.400 204.900 662.400 ;
        RECT 206.100 656.400 207.900 663.000 ;
        RECT 221.100 659.400 222.900 663.000 ;
        RECT 224.100 659.400 225.900 662.400 ;
        RECT 239.100 659.400 240.900 663.000 ;
        RECT 242.100 659.400 243.900 662.400 ;
        RECT 245.100 659.400 246.900 663.000 ;
        RECT 176.100 649.050 177.900 650.850 ;
        RECT 182.700 649.050 183.900 656.400 ;
        RECT 187.950 649.050 189.750 650.850 ;
        RECT 203.550 649.050 204.600 656.400 ;
        RECT 205.800 649.050 207.600 650.850 ;
        RECT 224.100 649.050 225.300 659.400 ;
        RECT 242.400 649.050 243.300 659.400 ;
        RECT 248.700 656.400 250.500 662.400 ;
        RECT 254.100 656.400 255.900 663.000 ;
        RECT 259.500 656.400 261.300 662.400 ;
        RECT 263.700 659.400 265.500 662.400 ;
        RECT 266.700 659.400 268.500 662.400 ;
        RECT 269.700 659.400 271.500 662.400 ;
        RECT 272.700 659.400 274.500 663.000 ;
        RECT 263.700 657.300 265.800 659.400 ;
        RECT 266.700 657.300 268.800 659.400 ;
        RECT 269.700 657.300 271.800 659.400 ;
        RECT 277.200 658.500 279.000 662.400 ;
        RECT 280.200 659.400 282.000 663.000 ;
        RECT 283.200 659.400 285.000 662.400 ;
        RECT 286.200 659.400 288.000 662.400 ;
        RECT 289.200 659.400 291.000 662.400 ;
        RECT 292.200 659.400 294.000 662.400 ;
        RECT 273.600 657.600 275.400 658.500 ;
        RECT 272.700 656.400 275.400 657.600 ;
        RECT 277.200 656.400 279.900 658.500 ;
        RECT 283.200 657.300 285.300 659.400 ;
        RECT 286.200 657.300 288.300 659.400 ;
        RECT 289.200 657.300 291.300 659.400 ;
        RECT 292.200 657.300 294.300 659.400 ;
        RECT 296.400 657.600 298.200 662.400 ;
        RECT 296.400 656.400 300.600 657.600 ;
        RECT 301.500 656.400 303.300 663.000 ;
        RECT 306.900 656.400 308.700 662.400 ;
        RECT 248.700 652.800 249.900 656.400 ;
        RECT 259.800 655.500 261.300 656.400 ;
        RECT 268.800 655.800 270.600 656.400 ;
        RECT 272.700 655.800 273.600 656.400 ;
        RECT 252.900 654.300 261.300 655.500 ;
        RECT 266.400 654.600 273.600 655.800 ;
        RECT 288.300 654.600 294.900 656.400 ;
        RECT 252.900 653.700 254.700 654.300 ;
        RECT 263.400 652.800 265.500 653.700 ;
        RECT 248.700 651.600 265.500 652.800 ;
        RECT 266.400 651.600 267.300 654.600 ;
        RECT 271.800 651.900 273.600 652.800 ;
        RECT 281.100 652.500 282.900 654.300 ;
        RECT 299.100 653.100 300.600 656.400 ;
        RECT 274.800 651.900 276.900 652.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 70.950 646.950 73.050 649.050 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 88.950 646.950 91.050 649.050 ;
        RECT 91.950 646.950 94.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 121.950 646.950 124.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 142.950 646.950 145.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 160.950 646.950 163.050 649.050 ;
        RECT 163.950 646.950 166.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 187.950 646.950 190.050 649.050 ;
        RECT 200.400 646.950 204.600 649.050 ;
        RECT 205.500 646.950 207.600 649.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 241.950 646.950 244.050 649.050 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 14.250 645.150 16.050 646.950 ;
        RECT 17.400 639.600 18.300 646.950 ;
        RECT 20.100 645.150 21.900 646.950 ;
        RECT 35.100 645.150 36.900 646.950 ;
        RECT 14.100 627.000 15.900 639.600 ;
        RECT 17.400 638.400 21.000 639.600 ;
        RECT 19.200 627.600 21.000 638.400 ;
        RECT 38.100 633.600 39.300 646.950 ;
        RECT 50.100 645.150 51.900 646.950 ;
        RECT 56.700 639.600 57.900 646.950 ;
        RECT 35.100 627.000 36.900 633.600 ;
        RECT 38.100 627.600 39.900 633.600 ;
        RECT 50.400 627.000 52.200 639.600 ;
        RECT 55.500 638.100 57.900 639.600 ;
        RECT 55.500 627.600 57.300 638.100 ;
        RECT 58.200 635.100 60.000 636.900 ;
        RECT 71.700 633.600 72.900 646.950 ;
        RECT 74.100 645.150 75.900 646.950 ;
        RECT 86.100 645.150 87.900 646.950 ;
        RECT 89.700 639.600 90.600 646.950 ;
        RECT 91.950 645.150 93.750 646.950 ;
        RECT 104.100 645.150 105.900 646.950 ;
        RECT 87.000 638.400 90.600 639.600 ;
        RECT 58.500 627.000 60.300 633.600 ;
        RECT 71.100 627.600 72.900 633.600 ;
        RECT 74.100 627.000 75.900 633.600 ;
        RECT 87.000 627.600 88.800 638.400 ;
        RECT 92.100 627.000 93.900 639.600 ;
        RECT 107.100 633.600 108.300 646.950 ;
        RECT 122.250 645.150 124.050 646.950 ;
        RECT 125.400 639.600 126.300 646.950 ;
        RECT 128.100 645.150 129.900 646.950 ;
        RECT 104.100 627.000 105.900 633.600 ;
        RECT 107.100 627.600 108.900 633.600 ;
        RECT 122.100 627.000 123.900 639.600 ;
        RECT 125.400 638.400 129.000 639.600 ;
        RECT 127.200 627.600 129.000 638.400 ;
        RECT 140.700 633.600 141.900 646.950 ;
        RECT 143.100 645.150 144.900 646.950 ;
        RECT 158.100 645.150 159.900 646.950 ;
        RECT 161.700 639.600 162.600 646.950 ;
        RECT 163.950 645.150 165.750 646.950 ;
        RECT 179.100 645.150 180.900 646.950 ;
        RECT 183.000 641.400 183.900 646.950 ;
        RECT 184.950 645.150 186.750 646.950 ;
        RECT 179.100 640.500 183.900 641.400 ;
        RECT 187.950 642.450 190.050 643.050 ;
        RECT 199.950 642.450 202.050 643.050 ;
        RECT 187.950 641.550 202.050 642.450 ;
        RECT 187.950 640.950 190.050 641.550 ;
        RECT 199.950 640.950 202.050 641.550 ;
        RECT 159.000 638.400 162.600 639.600 ;
        RECT 140.100 627.600 141.900 633.600 ;
        RECT 143.100 627.000 144.900 633.600 ;
        RECT 159.000 627.600 160.800 638.400 ;
        RECT 164.100 627.000 165.900 639.600 ;
        RECT 176.100 628.500 177.900 639.600 ;
        RECT 179.100 629.400 180.900 640.500 ;
        RECT 203.550 639.600 204.600 646.950 ;
        RECT 221.100 645.150 222.900 646.950 ;
        RECT 182.100 638.400 189.900 639.300 ;
        RECT 182.100 628.500 183.900 638.400 ;
        RECT 176.100 627.600 183.900 628.500 ;
        RECT 185.100 627.000 186.900 637.500 ;
        RECT 188.100 627.600 189.900 638.400 ;
        RECT 200.100 627.000 201.900 639.600 ;
        RECT 203.100 627.600 204.900 639.600 ;
        RECT 206.100 627.000 207.900 639.600 ;
        RECT 224.100 633.600 225.300 646.950 ;
        RECT 239.250 645.150 241.050 646.950 ;
        RECT 242.400 639.600 243.300 646.950 ;
        RECT 245.100 645.150 246.900 646.950 ;
        RECT 221.100 627.000 222.900 633.600 ;
        RECT 224.100 627.600 225.900 633.600 ;
        RECT 239.100 627.000 240.900 639.600 ;
        RECT 242.400 638.400 246.000 639.600 ;
        RECT 244.200 627.600 246.000 638.400 ;
        RECT 248.700 635.400 249.900 651.600 ;
        RECT 266.400 649.800 268.200 651.600 ;
        RECT 271.800 651.000 276.900 651.900 ;
        RECT 274.800 649.950 276.900 651.000 ;
        RECT 281.100 651.900 283.200 652.500 ;
        RECT 281.100 650.400 298.200 651.900 ;
        RECT 299.100 651.300 306.900 653.100 ;
        RECT 296.700 648.900 303.300 650.400 ;
        RECT 251.100 647.700 295.500 648.900 ;
        RECT 251.100 646.050 252.900 647.700 ;
        RECT 250.800 643.950 252.900 646.050 ;
        RECT 256.800 645.750 258.900 646.050 ;
        RECT 269.400 645.900 271.200 646.500 ;
        RECT 278.400 645.900 291.900 646.800 ;
        RECT 256.800 643.950 260.700 645.750 ;
        RECT 269.400 644.700 280.500 645.900 ;
        RECT 258.900 643.200 260.700 643.950 ;
        RECT 278.400 643.800 280.500 644.700 ;
        RECT 282.000 643.200 285.900 645.000 ;
        RECT 291.000 644.700 291.900 645.900 ;
        RECT 258.900 642.300 272.400 643.200 ;
        RECT 283.800 642.900 285.900 643.200 ;
        RECT 290.100 642.900 291.900 644.700 ;
        RECT 294.600 646.200 295.500 647.700 ;
        RECT 294.600 644.400 299.700 646.200 ;
        RECT 301.800 646.050 303.300 648.900 ;
        RECT 301.800 643.950 303.900 646.050 ;
        RECT 271.200 641.700 272.400 642.300 ;
        RECT 305.100 641.700 306.900 642.300 ;
        RECT 266.400 640.500 268.500 640.800 ;
        RECT 271.200 640.500 306.900 641.700 ;
        RECT 256.500 639.300 268.500 640.500 ;
        RECT 307.800 639.600 308.700 656.400 ;
        RECT 256.500 638.700 258.300 639.300 ;
        RECT 266.400 638.700 268.500 639.300 ;
        RECT 271.200 638.400 288.900 639.600 ;
        RECT 253.200 637.800 255.000 638.100 ;
        RECT 271.200 637.800 272.400 638.400 ;
        RECT 253.200 636.600 272.400 637.800 ;
        RECT 286.800 637.500 288.900 638.400 ;
        RECT 292.200 638.700 308.700 639.600 ;
        RECT 292.200 637.500 294.300 638.700 ;
        RECT 253.200 636.300 255.000 636.600 ;
        RECT 248.700 634.500 252.300 635.400 ;
        RECT 251.400 633.600 252.300 634.500 ;
        RECT 248.700 627.000 250.500 633.600 ;
        RECT 251.400 632.700 253.500 633.600 ;
        RECT 251.700 627.600 253.500 632.700 ;
        RECT 254.700 627.000 256.500 633.600 ;
        RECT 257.700 627.600 259.500 636.600 ;
        RECT 269.700 633.600 271.800 635.700 ;
        RECT 277.200 635.100 280.500 637.200 ;
        RECT 260.700 627.000 262.500 633.600 ;
        RECT 264.300 630.600 266.400 632.700 ;
        RECT 267.300 630.600 269.400 632.700 ;
        RECT 264.300 627.600 266.100 630.600 ;
        RECT 267.300 627.600 269.100 630.600 ;
        RECT 270.300 627.600 272.100 633.600 ;
        RECT 273.300 627.000 275.100 633.600 ;
        RECT 277.200 627.600 279.000 635.100 ;
        RECT 283.200 633.600 285.900 637.500 ;
        RECT 298.200 636.600 303.900 637.800 ;
        RECT 295.500 635.700 297.300 636.300 ;
        RECT 289.200 634.500 297.300 635.700 ;
        RECT 289.200 633.600 291.300 634.500 ;
        RECT 298.200 633.600 299.400 636.600 ;
        RECT 302.100 636.000 303.900 636.600 ;
        RECT 307.800 635.400 308.700 638.700 ;
        RECT 304.800 634.500 308.700 635.400 ;
        RECT 310.500 659.400 312.300 662.400 ;
        RECT 313.500 659.400 315.300 663.000 ;
        RECT 310.500 646.050 312.000 659.400 ;
        RECT 329.100 656.400 330.900 662.400 ;
        RECT 329.700 654.300 330.900 656.400 ;
        RECT 332.100 657.300 333.900 662.400 ;
        RECT 335.100 658.200 336.900 663.000 ;
        RECT 338.100 657.300 339.900 662.400 ;
        RECT 332.100 655.950 339.900 657.300 ;
        RECT 353.700 655.200 355.500 662.400 ;
        RECT 358.800 656.400 360.600 663.000 ;
        RECT 371.100 659.400 372.900 663.000 ;
        RECT 374.100 659.400 375.900 662.400 ;
        RECT 340.950 654.450 343.050 655.050 ;
        RECT 346.950 654.450 349.050 655.050 ;
        RECT 329.700 653.400 333.300 654.300 ;
        RECT 329.100 649.050 330.900 650.850 ;
        RECT 332.100 649.050 333.300 653.400 ;
        RECT 340.950 653.550 349.050 654.450 ;
        RECT 353.700 654.300 357.900 655.200 ;
        RECT 340.950 652.950 343.050 653.550 ;
        RECT 346.950 652.950 349.050 653.550 ;
        RECT 335.100 649.050 336.900 650.850 ;
        RECT 353.100 649.050 354.900 650.850 ;
        RECT 356.700 649.050 357.900 654.300 ;
        RECT 358.950 649.050 360.750 650.850 ;
        RECT 374.100 649.050 375.300 659.400 ;
        RECT 386.400 656.400 388.200 663.000 ;
        RECT 391.500 655.200 393.300 662.400 ;
        RECT 407.100 656.400 408.900 662.400 ;
        RECT 389.100 654.300 393.300 655.200 ;
        RECT 407.700 654.300 408.900 656.400 ;
        RECT 410.100 657.300 411.900 662.400 ;
        RECT 413.100 658.200 414.900 663.000 ;
        RECT 416.100 657.300 417.900 662.400 ;
        RECT 418.950 660.450 421.050 661.050 ;
        RECT 424.950 660.450 427.050 661.050 ;
        RECT 418.950 659.550 427.050 660.450 ;
        RECT 418.950 658.950 421.050 659.550 ;
        RECT 424.950 658.950 427.050 659.550 ;
        RECT 410.100 655.950 417.900 657.300 ;
        RECT 428.100 656.400 429.900 662.400 ;
        RECT 431.100 656.400 432.900 663.000 ;
        RECT 434.100 659.400 435.900 662.400 ;
        RECT 449.100 659.400 450.900 663.000 ;
        RECT 452.100 659.400 453.900 662.400 ;
        RECT 386.250 649.050 388.050 650.850 ;
        RECT 389.100 649.050 390.300 654.300 ;
        RECT 407.700 653.400 411.300 654.300 ;
        RECT 392.100 649.050 393.900 650.850 ;
        RECT 407.100 649.050 408.900 650.850 ;
        RECT 410.100 649.050 411.300 653.400 ;
        RECT 413.100 649.050 414.900 650.850 ;
        RECT 428.100 649.050 429.300 656.400 ;
        RECT 434.700 655.500 435.900 659.400 ;
        RECT 430.200 654.600 435.900 655.500 ;
        RECT 430.200 653.700 432.000 654.600 ;
        RECT 328.950 646.950 331.050 649.050 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 352.950 646.950 355.050 649.050 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 373.950 646.950 376.050 649.050 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 428.100 646.950 430.200 649.050 ;
        RECT 310.500 643.950 312.900 646.050 ;
        RECT 304.800 633.600 306.000 634.500 ;
        RECT 310.500 633.600 312.000 643.950 ;
        RECT 332.100 639.600 333.300 646.950 ;
        RECT 338.100 645.150 339.900 646.950 ;
        RECT 332.100 638.100 334.500 639.600 ;
        RECT 330.000 635.100 331.800 636.900 ;
        RECT 280.200 627.000 282.000 633.600 ;
        RECT 283.200 627.600 285.000 633.600 ;
        RECT 286.200 630.600 288.300 632.700 ;
        RECT 289.200 630.600 291.300 632.700 ;
        RECT 292.200 630.600 294.300 632.700 ;
        RECT 286.200 627.600 288.000 630.600 ;
        RECT 289.200 627.600 291.000 630.600 ;
        RECT 292.200 627.600 294.000 630.600 ;
        RECT 295.200 627.000 297.000 633.600 ;
        RECT 298.200 627.600 300.000 633.600 ;
        RECT 301.200 627.000 303.000 633.600 ;
        RECT 304.200 627.600 306.000 633.600 ;
        RECT 307.200 627.000 309.000 633.600 ;
        RECT 310.500 627.600 312.300 633.600 ;
        RECT 313.500 627.000 315.300 633.600 ;
        RECT 329.700 627.000 331.500 633.600 ;
        RECT 332.700 627.600 334.500 638.100 ;
        RECT 337.800 627.000 339.600 639.600 ;
        RECT 356.700 633.600 357.900 646.950 ;
        RECT 371.100 645.150 372.900 646.950 ;
        RECT 374.100 633.600 375.300 646.950 ;
        RECT 389.100 633.600 390.300 646.950 ;
        RECT 410.100 639.600 411.300 646.950 ;
        RECT 416.100 645.150 417.900 646.950 ;
        RECT 428.100 639.600 429.300 646.950 ;
        RECT 431.100 642.300 432.000 653.700 ;
        RECT 452.100 649.050 453.300 659.400 ;
        RECT 467.700 655.200 469.500 662.400 ;
        RECT 472.800 656.400 474.600 663.000 ;
        RECT 485.100 657.300 486.900 662.400 ;
        RECT 488.100 658.200 489.900 663.000 ;
        RECT 491.100 657.300 492.900 662.400 ;
        RECT 485.100 655.950 492.900 657.300 ;
        RECT 494.100 656.400 495.900 662.400 ;
        RECT 497.700 656.400 499.500 662.400 ;
        RECT 503.100 656.400 504.900 663.000 ;
        RECT 508.500 656.400 510.300 662.400 ;
        RECT 512.700 659.400 514.500 662.400 ;
        RECT 515.700 659.400 517.500 662.400 ;
        RECT 518.700 659.400 520.500 662.400 ;
        RECT 521.700 659.400 523.500 663.000 ;
        RECT 512.700 657.300 514.800 659.400 ;
        RECT 515.700 657.300 517.800 659.400 ;
        RECT 518.700 657.300 520.800 659.400 ;
        RECT 526.200 658.500 528.000 662.400 ;
        RECT 529.200 659.400 531.000 663.000 ;
        RECT 532.200 659.400 534.000 662.400 ;
        RECT 535.200 659.400 537.000 662.400 ;
        RECT 538.200 659.400 540.000 662.400 ;
        RECT 541.200 659.400 543.000 662.400 ;
        RECT 522.600 657.600 524.400 658.500 ;
        RECT 521.700 656.400 524.400 657.600 ;
        RECT 526.200 656.400 528.900 658.500 ;
        RECT 532.200 657.300 534.300 659.400 ;
        RECT 535.200 657.300 537.300 659.400 ;
        RECT 538.200 657.300 540.300 659.400 ;
        RECT 541.200 657.300 543.300 659.400 ;
        RECT 545.400 657.600 547.200 662.400 ;
        RECT 545.400 656.400 549.600 657.600 ;
        RECT 550.500 656.400 552.300 663.000 ;
        RECT 555.900 656.400 557.700 662.400 ;
        RECT 467.700 654.300 471.900 655.200 ;
        RECT 467.100 649.050 468.900 650.850 ;
        RECT 470.700 649.050 471.900 654.300 ;
        RECT 475.950 651.450 478.050 655.050 ;
        RECT 494.100 654.300 495.300 656.400 ;
        RECT 491.700 653.400 495.300 654.300 ;
        RECT 475.950 651.000 480.450 651.450 ;
        RECT 472.950 649.050 474.750 650.850 ;
        RECT 476.550 650.550 480.450 651.000 ;
        RECT 433.500 646.950 435.600 649.050 ;
        RECT 448.950 646.950 451.050 649.050 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 466.950 646.950 469.050 649.050 ;
        RECT 469.950 646.950 472.050 649.050 ;
        RECT 472.950 646.950 475.050 649.050 ;
        RECT 433.800 645.150 435.600 646.950 ;
        RECT 449.100 645.150 450.900 646.950 ;
        RECT 430.200 641.400 432.000 642.300 ;
        RECT 430.200 640.500 435.900 641.400 ;
        RECT 410.100 638.100 412.500 639.600 ;
        RECT 408.000 635.100 409.800 636.900 ;
        RECT 353.100 627.000 354.900 633.600 ;
        RECT 356.100 627.600 357.900 633.600 ;
        RECT 359.100 627.000 360.900 633.600 ;
        RECT 371.100 627.000 372.900 633.600 ;
        RECT 374.100 627.600 375.900 633.600 ;
        RECT 386.100 627.000 387.900 633.600 ;
        RECT 389.100 627.600 390.900 633.600 ;
        RECT 392.100 627.000 393.900 633.600 ;
        RECT 407.700 627.000 409.500 633.600 ;
        RECT 410.700 627.600 412.500 638.100 ;
        RECT 415.800 627.000 417.600 639.600 ;
        RECT 428.100 627.600 429.900 639.600 ;
        RECT 431.100 627.000 432.900 637.800 ;
        RECT 434.700 633.600 435.900 640.500 ;
        RECT 452.100 633.600 453.300 646.950 ;
        RECT 454.950 645.450 457.050 646.050 ;
        RECT 460.950 645.450 463.050 646.050 ;
        RECT 454.950 644.550 463.050 645.450 ;
        RECT 454.950 643.950 457.050 644.550 ;
        RECT 460.950 643.950 463.050 644.550 ;
        RECT 434.100 627.600 435.900 633.600 ;
        RECT 449.100 627.000 450.900 633.600 ;
        RECT 452.100 627.600 453.900 633.600 ;
        RECT 457.950 633.450 460.050 633.900 ;
        RECT 463.950 633.450 466.050 634.050 ;
        RECT 470.700 633.600 471.900 646.950 ;
        RECT 479.550 645.450 480.450 650.550 ;
        RECT 488.100 649.050 489.900 650.850 ;
        RECT 491.700 649.050 492.900 653.400 ;
        RECT 497.700 652.800 498.900 656.400 ;
        RECT 508.800 655.500 510.300 656.400 ;
        RECT 517.800 655.800 519.600 656.400 ;
        RECT 521.700 655.800 522.600 656.400 ;
        RECT 501.900 654.300 510.300 655.500 ;
        RECT 515.400 654.600 522.600 655.800 ;
        RECT 537.300 654.600 543.900 656.400 ;
        RECT 501.900 653.700 503.700 654.300 ;
        RECT 512.400 652.800 514.500 653.700 ;
        RECT 497.700 651.600 514.500 652.800 ;
        RECT 515.400 651.600 516.300 654.600 ;
        RECT 520.800 651.900 522.600 652.800 ;
        RECT 530.100 652.500 531.900 654.300 ;
        RECT 548.100 653.100 549.600 656.400 ;
        RECT 523.800 651.900 525.900 652.050 ;
        RECT 494.100 649.050 495.900 650.850 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 479.550 645.000 483.450 645.450 ;
        RECT 485.100 645.150 486.900 646.950 ;
        RECT 479.550 644.550 484.050 645.000 ;
        RECT 481.950 640.950 484.050 644.550 ;
        RECT 491.700 639.600 492.900 646.950 ;
        RECT 457.950 632.550 466.050 633.450 ;
        RECT 457.950 631.800 460.050 632.550 ;
        RECT 463.950 631.950 466.050 632.550 ;
        RECT 467.100 627.000 468.900 633.600 ;
        RECT 470.100 627.600 471.900 633.600 ;
        RECT 473.100 627.000 474.900 633.600 ;
        RECT 485.400 627.000 487.200 639.600 ;
        RECT 490.500 638.100 492.900 639.600 ;
        RECT 490.500 627.600 492.300 638.100 ;
        RECT 493.200 635.100 495.000 636.900 ;
        RECT 497.700 635.400 498.900 651.600 ;
        RECT 515.400 649.800 517.200 651.600 ;
        RECT 520.800 651.000 525.900 651.900 ;
        RECT 523.800 649.950 525.900 651.000 ;
        RECT 530.100 651.900 532.200 652.500 ;
        RECT 530.100 650.400 547.200 651.900 ;
        RECT 548.100 651.300 555.900 653.100 ;
        RECT 545.700 648.900 552.300 650.400 ;
        RECT 500.100 647.700 544.500 648.900 ;
        RECT 500.100 646.050 501.900 647.700 ;
        RECT 499.800 643.950 501.900 646.050 ;
        RECT 505.800 645.750 507.900 646.050 ;
        RECT 518.400 645.900 520.200 646.500 ;
        RECT 527.400 645.900 540.900 646.800 ;
        RECT 505.800 643.950 509.700 645.750 ;
        RECT 518.400 644.700 529.500 645.900 ;
        RECT 507.900 643.200 509.700 643.950 ;
        RECT 527.400 643.800 529.500 644.700 ;
        RECT 531.000 643.200 534.900 645.000 ;
        RECT 540.000 644.700 540.900 645.900 ;
        RECT 507.900 642.300 521.400 643.200 ;
        RECT 532.800 642.900 534.900 643.200 ;
        RECT 539.100 642.900 540.900 644.700 ;
        RECT 543.600 646.200 544.500 647.700 ;
        RECT 543.600 644.400 548.700 646.200 ;
        RECT 550.800 646.050 552.300 648.900 ;
        RECT 550.800 643.950 552.900 646.050 ;
        RECT 520.200 641.700 521.400 642.300 ;
        RECT 554.100 641.700 555.900 642.300 ;
        RECT 515.400 640.500 517.500 640.800 ;
        RECT 520.200 640.500 555.900 641.700 ;
        RECT 505.500 639.300 517.500 640.500 ;
        RECT 556.800 639.600 557.700 656.400 ;
        RECT 505.500 638.700 507.300 639.300 ;
        RECT 515.400 638.700 517.500 639.300 ;
        RECT 520.200 638.400 537.900 639.600 ;
        RECT 502.200 637.800 504.000 638.100 ;
        RECT 520.200 637.800 521.400 638.400 ;
        RECT 502.200 636.600 521.400 637.800 ;
        RECT 535.800 637.500 537.900 638.400 ;
        RECT 541.200 638.700 557.700 639.600 ;
        RECT 541.200 637.500 543.300 638.700 ;
        RECT 502.200 636.300 504.000 636.600 ;
        RECT 497.700 634.500 501.300 635.400 ;
        RECT 500.400 633.600 501.300 634.500 ;
        RECT 493.500 627.000 495.300 633.600 ;
        RECT 497.700 627.000 499.500 633.600 ;
        RECT 500.400 632.700 502.500 633.600 ;
        RECT 500.700 627.600 502.500 632.700 ;
        RECT 503.700 627.000 505.500 633.600 ;
        RECT 506.700 627.600 508.500 636.600 ;
        RECT 518.700 633.600 520.800 635.700 ;
        RECT 526.200 635.100 529.500 637.200 ;
        RECT 509.700 627.000 511.500 633.600 ;
        RECT 513.300 630.600 515.400 632.700 ;
        RECT 516.300 630.600 518.400 632.700 ;
        RECT 513.300 627.600 515.100 630.600 ;
        RECT 516.300 627.600 518.100 630.600 ;
        RECT 519.300 627.600 521.100 633.600 ;
        RECT 522.300 627.000 524.100 633.600 ;
        RECT 526.200 627.600 528.000 635.100 ;
        RECT 532.200 633.600 534.900 637.500 ;
        RECT 547.200 636.600 552.900 637.800 ;
        RECT 544.500 635.700 546.300 636.300 ;
        RECT 538.200 634.500 546.300 635.700 ;
        RECT 538.200 633.600 540.300 634.500 ;
        RECT 547.200 633.600 548.400 636.600 ;
        RECT 551.100 636.000 552.900 636.600 ;
        RECT 556.800 635.400 557.700 638.700 ;
        RECT 553.800 634.500 557.700 635.400 ;
        RECT 559.500 659.400 561.300 662.400 ;
        RECT 562.500 659.400 564.300 663.000 ;
        RECT 575.100 659.400 576.900 663.000 ;
        RECT 578.100 659.400 579.900 662.400 ;
        RECT 559.500 646.050 561.000 659.400 ;
        RECT 565.950 657.450 568.050 658.050 ;
        RECT 571.950 657.450 574.050 658.050 ;
        RECT 565.950 656.550 574.050 657.450 ;
        RECT 565.950 655.950 568.050 656.550 ;
        RECT 571.950 655.950 574.050 656.550 ;
        RECT 568.950 654.450 571.050 655.050 ;
        RECT 574.950 654.450 577.050 655.050 ;
        RECT 568.950 653.550 577.050 654.450 ;
        RECT 568.950 652.950 571.050 653.550 ;
        RECT 574.950 652.950 577.050 653.550 ;
        RECT 578.100 649.050 579.300 659.400 ;
        RECT 593.100 656.400 594.900 662.400 ;
        RECT 593.700 654.300 594.900 656.400 ;
        RECT 596.100 657.300 597.900 662.400 ;
        RECT 599.100 658.200 600.900 663.000 ;
        RECT 602.100 657.300 603.900 662.400 ;
        RECT 596.100 655.950 603.900 657.300 ;
        RECT 617.700 655.200 619.500 662.400 ;
        RECT 622.800 656.400 624.600 663.000 ;
        RECT 638.100 659.400 639.900 663.000 ;
        RECT 641.100 659.400 642.900 662.400 ;
        RECT 644.100 659.400 645.900 663.000 ;
        RECT 617.700 654.300 621.900 655.200 ;
        RECT 593.700 653.400 597.300 654.300 ;
        RECT 593.100 649.050 594.900 650.850 ;
        RECT 596.100 649.050 597.300 653.400 ;
        RECT 599.100 649.050 600.900 650.850 ;
        RECT 617.100 649.050 618.900 650.850 ;
        RECT 620.700 649.050 621.900 654.300 ;
        RECT 622.950 649.050 624.750 650.850 ;
        RECT 641.400 649.050 642.300 659.400 ;
        RECT 659.400 656.400 661.200 663.000 ;
        RECT 664.500 655.200 666.300 662.400 ;
        RECT 677.700 659.400 679.500 663.000 ;
        RECT 680.700 657.600 682.500 662.400 ;
        RECT 662.100 654.300 666.300 655.200 ;
        RECT 677.400 656.400 682.500 657.600 ;
        RECT 685.200 656.400 687.000 663.000 ;
        RECT 659.250 649.050 661.050 650.850 ;
        RECT 662.100 649.050 663.300 654.300 ;
        RECT 665.100 649.050 666.900 650.850 ;
        RECT 677.400 649.050 678.300 656.400 ;
        RECT 698.100 653.400 699.900 663.000 ;
        RECT 704.700 654.000 706.500 662.400 ;
        RECT 724.500 654.000 726.300 662.400 ;
        RECT 704.700 652.800 708.000 654.000 ;
        RECT 679.950 649.050 681.750 650.850 ;
        RECT 686.100 649.050 687.900 650.850 ;
        RECT 698.100 649.050 699.900 650.850 ;
        RECT 704.100 649.050 705.900 650.850 ;
        RECT 707.100 649.050 708.000 652.800 ;
        RECT 723.000 652.800 726.300 654.000 ;
        RECT 731.100 653.400 732.900 663.000 ;
        RECT 746.100 657.300 747.900 662.400 ;
        RECT 749.100 658.200 750.900 663.000 ;
        RECT 752.100 657.300 753.900 662.400 ;
        RECT 746.100 655.950 753.900 657.300 ;
        RECT 755.100 656.400 756.900 662.400 ;
        RECT 770.100 659.400 771.900 663.000 ;
        RECT 773.100 659.400 774.900 662.400 ;
        RECT 776.100 659.400 777.900 663.000 ;
        RECT 755.100 654.300 756.300 656.400 ;
        RECT 752.700 653.400 756.300 654.300 ;
        RECT 723.000 649.050 723.900 652.800 ;
        RECT 725.100 649.050 726.900 650.850 ;
        RECT 731.100 649.050 732.900 650.850 ;
        RECT 739.950 649.950 742.050 652.050 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 598.950 646.950 601.050 649.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 619.950 646.950 622.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 640.950 646.950 643.050 649.050 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 658.950 646.950 661.050 649.050 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 706.950 646.950 709.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 559.500 643.950 561.900 646.050 ;
        RECT 575.100 645.150 576.900 646.950 ;
        RECT 553.800 633.600 555.000 634.500 ;
        RECT 559.500 633.600 561.000 643.950 ;
        RECT 578.100 633.600 579.300 646.950 ;
        RECT 596.100 639.600 597.300 646.950 ;
        RECT 602.100 645.150 603.900 646.950 ;
        RECT 596.100 638.100 598.500 639.600 ;
        RECT 594.000 635.100 595.800 636.900 ;
        RECT 529.200 627.000 531.000 633.600 ;
        RECT 532.200 627.600 534.000 633.600 ;
        RECT 535.200 630.600 537.300 632.700 ;
        RECT 538.200 630.600 540.300 632.700 ;
        RECT 541.200 630.600 543.300 632.700 ;
        RECT 535.200 627.600 537.000 630.600 ;
        RECT 538.200 627.600 540.000 630.600 ;
        RECT 541.200 627.600 543.000 630.600 ;
        RECT 544.200 627.000 546.000 633.600 ;
        RECT 547.200 627.600 549.000 633.600 ;
        RECT 550.200 627.000 552.000 633.600 ;
        RECT 553.200 627.600 555.000 633.600 ;
        RECT 556.200 627.000 558.000 633.600 ;
        RECT 559.500 627.600 561.300 633.600 ;
        RECT 562.500 627.000 564.300 633.600 ;
        RECT 575.100 627.000 576.900 633.600 ;
        RECT 578.100 627.600 579.900 633.600 ;
        RECT 593.700 627.000 595.500 633.600 ;
        RECT 596.700 627.600 598.500 638.100 ;
        RECT 601.800 627.000 603.600 639.600 ;
        RECT 620.700 633.600 621.900 646.950 ;
        RECT 638.250 645.150 640.050 646.950 ;
        RECT 628.950 642.450 631.050 643.050 ;
        RECT 637.950 642.450 640.050 643.050 ;
        RECT 628.950 641.550 640.050 642.450 ;
        RECT 628.950 640.950 631.050 641.550 ;
        RECT 637.950 640.950 640.050 641.550 ;
        RECT 641.400 639.600 642.300 646.950 ;
        RECT 644.100 645.150 645.900 646.950 ;
        RECT 617.100 627.000 618.900 633.600 ;
        RECT 620.100 627.600 621.900 633.600 ;
        RECT 623.100 627.000 624.900 633.600 ;
        RECT 638.100 627.000 639.900 639.600 ;
        RECT 641.400 638.400 645.000 639.600 ;
        RECT 643.200 627.600 645.000 638.400 ;
        RECT 662.100 633.600 663.300 646.950 ;
        RECT 677.400 639.600 678.300 646.950 ;
        RECT 682.950 645.150 684.750 646.950 ;
        RECT 701.100 645.150 702.900 646.950 ;
        RECT 679.950 642.450 682.050 643.050 ;
        RECT 691.950 642.450 694.050 643.050 ;
        RECT 703.950 642.450 706.050 643.050 ;
        RECT 679.950 641.550 706.050 642.450 ;
        RECT 679.950 640.950 682.050 641.550 ;
        RECT 691.950 640.950 694.050 641.550 ;
        RECT 703.950 640.950 706.050 641.550 ;
        RECT 659.100 627.000 660.900 633.600 ;
        RECT 662.100 627.600 663.900 633.600 ;
        RECT 665.100 627.000 666.900 633.600 ;
        RECT 677.100 627.600 678.900 639.600 ;
        RECT 680.100 638.700 687.900 639.600 ;
        RECT 680.100 627.600 681.900 638.700 ;
        RECT 683.100 627.000 684.900 637.800 ;
        RECT 686.100 627.600 687.900 638.700 ;
        RECT 707.100 634.800 708.000 646.950 ;
        RECT 701.400 633.900 708.000 634.800 ;
        RECT 701.400 633.600 702.900 633.900 ;
        RECT 698.100 627.000 699.900 633.600 ;
        RECT 701.100 627.600 702.900 633.600 ;
        RECT 707.100 633.600 708.000 633.900 ;
        RECT 723.000 634.800 723.900 646.950 ;
        RECT 728.100 645.150 729.900 646.950 ;
        RECT 733.950 645.450 736.050 646.050 ;
        RECT 740.550 645.450 741.450 649.950 ;
        RECT 749.100 649.050 750.900 650.850 ;
        RECT 752.700 649.050 753.900 653.400 ;
        RECT 760.950 651.450 763.050 652.050 ;
        RECT 766.950 651.450 769.050 652.050 ;
        RECT 755.100 649.050 756.900 650.850 ;
        RECT 760.950 650.550 769.050 651.450 ;
        RECT 760.950 649.950 763.050 650.550 ;
        RECT 766.950 649.950 769.050 650.550 ;
        RECT 773.700 649.050 774.600 659.400 ;
        RECT 791.400 656.400 793.200 663.000 ;
        RECT 796.500 655.200 798.300 662.400 ;
        RECT 812.100 657.300 813.900 662.400 ;
        RECT 815.100 658.200 816.900 663.000 ;
        RECT 818.100 657.300 819.900 662.400 ;
        RECT 812.100 655.950 819.900 657.300 ;
        RECT 821.100 656.400 822.900 662.400 ;
        RECT 833.100 659.400 834.900 663.000 ;
        RECT 836.100 659.400 837.900 662.400 ;
        RECT 794.100 654.300 798.300 655.200 ;
        RECT 821.100 654.300 822.300 656.400 ;
        RECT 791.250 649.050 793.050 650.850 ;
        RECT 794.100 649.050 795.300 654.300 ;
        RECT 818.700 653.400 822.300 654.300 ;
        RECT 797.100 649.050 798.900 650.850 ;
        RECT 815.100 649.050 816.900 650.850 ;
        RECT 818.700 649.050 819.900 653.400 ;
        RECT 821.100 649.050 822.900 650.850 ;
        RECT 836.100 649.050 837.300 659.400 ;
        RECT 848.100 657.300 849.900 662.400 ;
        RECT 851.100 658.200 852.900 663.000 ;
        RECT 854.100 657.300 855.900 662.400 ;
        RECT 848.100 655.950 855.900 657.300 ;
        RECT 857.100 656.400 858.900 662.400 ;
        RECT 869.700 659.400 871.500 663.000 ;
        RECT 872.700 657.600 874.500 662.400 ;
        RECT 869.400 656.400 874.500 657.600 ;
        RECT 877.200 656.400 879.000 663.000 ;
        RECT 890.100 659.400 891.900 662.400 ;
        RECT 893.100 659.400 894.900 663.000 ;
        RECT 857.100 654.300 858.300 656.400 ;
        RECT 854.700 653.400 858.300 654.300 ;
        RECT 843.000 651.450 847.050 652.050 ;
        RECT 842.550 649.950 847.050 651.450 ;
        RECT 745.950 646.950 748.050 649.050 ;
        RECT 748.950 646.950 751.050 649.050 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 775.950 646.950 778.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 733.950 644.550 741.450 645.450 ;
        RECT 746.100 645.150 747.900 646.950 ;
        RECT 733.950 643.950 736.050 644.550 ;
        RECT 752.700 639.600 753.900 646.950 ;
        RECT 770.100 645.150 771.900 646.950 ;
        RECT 773.700 639.600 774.600 646.950 ;
        RECT 775.950 645.150 777.750 646.950 ;
        RECT 723.000 633.900 729.600 634.800 ;
        RECT 723.000 633.600 723.900 633.900 ;
        RECT 704.100 627.000 705.900 633.000 ;
        RECT 707.100 627.600 708.900 633.600 ;
        RECT 722.100 627.600 723.900 633.600 ;
        RECT 728.100 633.600 729.600 633.900 ;
        RECT 725.100 627.000 726.900 633.000 ;
        RECT 728.100 627.600 729.900 633.600 ;
        RECT 731.100 627.000 732.900 633.600 ;
        RECT 746.400 627.000 748.200 639.600 ;
        RECT 751.500 638.100 753.900 639.600 ;
        RECT 771.000 638.400 774.600 639.600 ;
        RECT 751.500 627.600 753.300 638.100 ;
        RECT 754.200 635.100 756.000 636.900 ;
        RECT 754.500 627.000 756.300 633.600 ;
        RECT 771.000 627.600 772.800 638.400 ;
        RECT 776.100 627.000 777.900 639.600 ;
        RECT 794.100 633.600 795.300 646.950 ;
        RECT 812.100 645.150 813.900 646.950 ;
        RECT 818.700 639.600 819.900 646.950 ;
        RECT 833.100 645.150 834.900 646.950 ;
        RECT 796.950 636.450 799.050 636.900 ;
        RECT 802.950 636.450 805.050 637.050 ;
        RECT 796.950 635.550 805.050 636.450 ;
        RECT 796.950 634.800 799.050 635.550 ;
        RECT 802.950 634.950 805.050 635.550 ;
        RECT 791.100 627.000 792.900 633.600 ;
        RECT 794.100 627.600 795.900 633.600 ;
        RECT 797.100 627.000 798.900 633.600 ;
        RECT 812.400 627.000 814.200 639.600 ;
        RECT 817.500 638.100 819.900 639.600 ;
        RECT 817.500 627.600 819.300 638.100 ;
        RECT 820.200 635.100 822.000 636.900 ;
        RECT 836.100 633.600 837.300 646.950 ;
        RECT 842.550 646.050 843.450 649.950 ;
        RECT 851.100 649.050 852.900 650.850 ;
        RECT 854.700 649.050 855.900 653.400 ;
        RECT 864.000 651.450 868.050 652.050 ;
        RECT 857.100 649.050 858.900 650.850 ;
        RECT 863.550 649.950 868.050 651.450 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 850.950 646.950 853.050 649.050 ;
        RECT 853.950 646.950 856.050 649.050 ;
        RECT 856.950 646.950 859.050 649.050 ;
        RECT 842.550 644.550 847.050 646.050 ;
        RECT 848.100 645.150 849.900 646.950 ;
        RECT 843.000 643.950 847.050 644.550 ;
        RECT 854.700 639.600 855.900 646.950 ;
        RECT 863.550 646.050 864.450 649.950 ;
        RECT 869.400 649.050 870.300 656.400 ;
        RECT 871.950 649.050 873.750 650.850 ;
        RECT 878.100 649.050 879.900 650.850 ;
        RECT 890.700 649.050 891.900 659.400 ;
        RECT 892.950 657.450 895.050 658.050 ;
        RECT 901.950 657.450 904.050 658.050 ;
        RECT 892.950 656.550 904.050 657.450 ;
        RECT 892.950 655.950 895.050 656.550 ;
        RECT 901.950 655.950 904.050 656.550 ;
        RECT 908.100 657.300 909.900 662.400 ;
        RECT 911.100 658.200 912.900 663.000 ;
        RECT 914.100 657.300 915.900 662.400 ;
        RECT 908.100 655.950 915.900 657.300 ;
        RECT 917.100 656.400 918.900 662.400 ;
        RECT 922.950 660.450 925.050 661.050 ;
        RECT 931.950 660.450 934.050 661.050 ;
        RECT 922.950 659.550 934.050 660.450 ;
        RECT 922.950 658.950 925.050 659.550 ;
        RECT 931.950 658.950 934.050 659.550 ;
        RECT 892.950 654.450 895.050 655.050 ;
        RECT 892.950 653.550 903.450 654.450 ;
        RECT 917.100 654.300 918.300 656.400 ;
        RECT 928.950 654.450 931.050 655.050 ;
        RECT 892.950 652.950 895.050 653.550 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 874.950 646.950 877.050 649.050 ;
        RECT 877.950 646.950 880.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 859.950 644.550 864.450 646.050 ;
        RECT 859.950 643.950 864.000 644.550 ;
        RECT 856.950 642.450 859.050 643.050 ;
        RECT 865.950 642.450 868.050 643.050 ;
        RECT 856.950 641.550 868.050 642.450 ;
        RECT 856.950 640.950 859.050 641.550 ;
        RECT 865.950 640.950 868.050 641.550 ;
        RECT 869.400 639.600 870.300 646.950 ;
        RECT 874.950 645.150 876.750 646.950 ;
        RECT 820.500 627.000 822.300 633.600 ;
        RECT 833.100 627.000 834.900 633.600 ;
        RECT 836.100 627.600 837.900 633.600 ;
        RECT 848.400 627.000 850.200 639.600 ;
        RECT 853.500 638.100 855.900 639.600 ;
        RECT 853.500 627.600 855.300 638.100 ;
        RECT 856.200 635.100 858.000 636.900 ;
        RECT 856.500 627.000 858.300 633.600 ;
        RECT 869.100 627.600 870.900 639.600 ;
        RECT 872.100 638.700 879.900 639.600 ;
        RECT 872.100 627.600 873.900 638.700 ;
        RECT 875.100 627.000 876.900 637.800 ;
        RECT 878.100 627.600 879.900 638.700 ;
        RECT 890.700 633.600 891.900 646.950 ;
        RECT 893.100 645.150 894.900 646.950 ;
        RECT 902.550 646.050 903.450 653.550 ;
        RECT 914.700 653.400 918.300 654.300 ;
        RECT 923.550 653.550 931.050 654.450 ;
        RECT 911.100 649.050 912.900 650.850 ;
        RECT 914.700 649.050 915.900 653.400 ;
        RECT 917.100 649.050 918.900 650.850 ;
        RECT 907.950 646.950 910.050 649.050 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 916.950 646.950 919.050 649.050 ;
        RECT 902.550 644.550 907.050 646.050 ;
        RECT 908.100 645.150 909.900 646.950 ;
        RECT 903.000 643.950 907.050 644.550 ;
        RECT 892.950 642.450 895.050 643.050 ;
        RECT 910.950 642.450 913.050 643.050 ;
        RECT 892.950 641.550 913.050 642.450 ;
        RECT 892.950 640.950 895.050 641.550 ;
        RECT 910.950 640.950 913.050 641.550 ;
        RECT 914.700 639.600 915.900 646.950 ;
        RECT 923.550 646.050 924.450 653.550 ;
        RECT 928.950 652.950 931.050 653.550 ;
        RECT 919.950 644.550 924.450 646.050 ;
        RECT 919.950 643.950 924.000 644.550 ;
        RECT 890.100 627.600 891.900 633.600 ;
        RECT 893.100 627.000 894.900 633.600 ;
        RECT 908.400 627.000 910.200 639.600 ;
        RECT 913.500 638.100 915.900 639.600 ;
        RECT 913.500 627.600 915.300 638.100 ;
        RECT 916.200 635.100 918.000 636.900 ;
        RECT 916.500 627.000 918.300 633.600 ;
        RECT 14.100 611.400 15.900 624.000 ;
        RECT 17.100 610.500 18.900 623.400 ;
        RECT 20.100 611.400 21.900 624.000 ;
        RECT 23.100 611.400 24.900 623.400 ;
        RECT 26.100 611.400 27.900 624.000 ;
        RECT 38.100 611.400 39.900 623.400 ;
        RECT 41.100 612.300 42.900 623.400 ;
        RECT 44.100 613.200 45.900 624.000 ;
        RECT 47.100 612.300 48.900 623.400 ;
        RECT 41.100 611.400 48.900 612.300 ;
        RECT 63.000 612.600 64.800 623.400 ;
        RECT 63.000 611.400 66.600 612.600 ;
        RECT 68.100 611.400 69.900 624.000 ;
        RECT 80.700 617.400 82.500 624.000 ;
        RECT 81.000 614.100 82.800 615.900 ;
        RECT 83.700 612.900 85.500 623.400 ;
        RECT 83.100 611.400 85.500 612.900 ;
        RECT 88.800 611.400 90.600 624.000 ;
        RECT 104.100 611.400 105.900 624.000 ;
        RECT 109.200 612.600 111.000 623.400 ;
        RECT 115.950 615.450 118.050 616.050 ;
        RECT 121.950 615.450 124.050 616.050 ;
        RECT 115.950 614.550 124.050 615.450 ;
        RECT 115.950 613.950 118.050 614.550 ;
        RECT 121.950 613.950 124.050 614.550 ;
        RECT 107.400 611.400 111.000 612.600 ;
        RECT 125.100 611.400 126.900 623.400 ;
        RECT 129.600 611.400 131.400 624.000 ;
        RECT 132.600 612.900 134.400 623.400 ;
        RECT 146.100 617.400 147.900 623.400 ;
        RECT 149.100 617.400 150.900 624.000 ;
        RECT 132.600 611.400 135.000 612.900 ;
        RECT 23.100 610.500 24.300 611.400 ;
        RECT 17.100 609.600 24.300 610.500 ;
        RECT 17.100 604.050 18.900 605.850 ;
        RECT 23.100 604.050 24.300 609.600 ;
        RECT 34.950 606.450 37.050 607.050 ;
        RECT 29.550 605.550 37.050 606.450 ;
        RECT 17.100 601.950 19.200 604.050 ;
        RECT 23.100 601.950 25.200 604.050 ;
        RECT 23.100 596.700 24.300 601.950 ;
        RECT 29.550 601.050 30.450 605.550 ;
        RECT 34.950 604.950 37.050 605.550 ;
        RECT 38.400 604.050 39.300 611.400 ;
        RECT 43.950 604.050 45.750 605.850 ;
        RECT 62.100 604.050 63.900 605.850 ;
        RECT 65.700 604.050 66.600 611.400 ;
        RECT 67.950 604.050 69.750 605.850 ;
        RECT 83.100 604.050 84.300 611.400 ;
        RECT 89.100 604.050 90.900 605.850 ;
        RECT 104.250 604.050 106.050 605.850 ;
        RECT 107.400 604.050 108.300 611.400 ;
        RECT 125.100 609.900 126.300 611.400 ;
        RECT 125.100 608.700 132.900 609.900 ;
        RECT 131.100 608.100 132.900 608.700 ;
        RECT 110.100 604.050 111.900 605.850 ;
        RECT 129.000 604.050 130.800 605.850 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 46.950 601.950 49.050 604.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 85.950 601.950 88.050 604.050 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 106.950 601.950 109.050 604.050 ;
        RECT 109.950 601.950 112.050 604.050 ;
        RECT 125.100 601.950 127.200 604.050 ;
        RECT 128.400 601.950 130.500 604.050 ;
        RECT 25.950 599.550 30.450 601.050 ;
        RECT 25.950 598.950 30.000 599.550 ;
        RECT 17.100 595.500 24.300 596.700 ;
        RECT 17.100 594.600 18.300 595.500 ;
        RECT 23.100 594.600 24.300 595.500 ;
        RECT 38.400 594.600 39.300 601.950 ;
        RECT 40.950 600.150 42.750 601.950 ;
        RECT 47.100 600.150 48.900 601.950 ;
        RECT 14.100 588.000 15.900 594.600 ;
        RECT 17.100 588.600 18.900 594.600 ;
        RECT 20.100 588.000 21.900 594.600 ;
        RECT 23.100 588.600 24.900 594.600 ;
        RECT 26.100 588.000 27.900 594.600 ;
        RECT 38.400 593.400 43.500 594.600 ;
        RECT 38.700 588.000 40.500 591.600 ;
        RECT 41.700 588.600 43.500 593.400 ;
        RECT 46.200 588.000 48.000 594.600 ;
        RECT 65.700 591.600 66.600 601.950 ;
        RECT 80.100 600.150 81.900 601.950 ;
        RECT 83.100 597.600 84.300 601.950 ;
        RECT 86.100 600.150 87.900 601.950 ;
        RECT 80.700 596.700 84.300 597.600 ;
        RECT 80.700 594.600 81.900 596.700 ;
        RECT 62.100 588.000 63.900 591.600 ;
        RECT 65.100 588.600 66.900 591.600 ;
        RECT 68.100 588.000 69.900 591.600 ;
        RECT 80.100 588.600 81.900 594.600 ;
        RECT 83.100 593.700 90.900 595.050 ;
        RECT 83.100 588.600 84.900 593.700 ;
        RECT 86.100 588.000 87.900 592.800 ;
        RECT 89.100 588.600 90.900 593.700 ;
        RECT 107.400 591.600 108.300 601.950 ;
        RECT 125.400 600.150 127.200 601.950 ;
        RECT 131.700 597.600 132.600 608.100 ;
        RECT 133.800 604.050 135.000 611.400 ;
        RECT 146.700 604.050 147.900 617.400 ;
        RECT 162.600 611.400 164.400 624.000 ;
        RECT 167.100 611.400 170.400 623.400 ;
        RECT 173.100 611.400 174.900 624.000 ;
        RECT 188.100 622.500 195.900 623.400 ;
        RECT 188.100 611.400 189.900 622.500 ;
        RECT 149.100 604.050 150.900 605.850 ;
        RECT 161.250 604.050 163.050 605.850 ;
        RECT 168.000 604.050 169.050 611.400 ;
        RECT 191.100 610.500 192.900 621.600 ;
        RECT 194.100 612.600 195.900 622.500 ;
        RECT 197.100 613.500 198.900 624.000 ;
        RECT 200.100 612.600 201.900 623.400 ;
        RECT 212.100 617.400 213.900 623.400 ;
        RECT 215.100 617.400 216.900 624.000 ;
        RECT 194.100 611.700 201.900 612.600 ;
        RECT 172.950 609.450 175.050 610.050 ;
        RECT 181.950 609.450 184.050 610.050 ;
        RECT 191.100 609.600 195.900 610.500 ;
        RECT 172.950 608.550 184.050 609.450 ;
        RECT 172.950 607.950 175.050 608.550 ;
        RECT 181.950 607.950 184.050 608.550 ;
        RECT 175.950 606.450 180.000 607.050 ;
        RECT 183.000 606.450 187.050 607.050 ;
        RECT 173.100 604.050 174.900 605.850 ;
        RECT 175.950 604.950 180.450 606.450 ;
        RECT 133.800 601.950 135.900 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 148.950 601.950 151.050 604.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 131.700 596.700 133.800 597.600 ;
        RECT 128.400 595.800 133.800 596.700 ;
        RECT 109.950 594.450 112.050 594.900 ;
        RECT 115.950 594.450 118.050 595.050 ;
        RECT 109.950 593.550 118.050 594.450 ;
        RECT 109.950 592.800 112.050 593.550 ;
        RECT 115.950 592.950 118.050 593.550 ;
        RECT 128.400 591.600 129.300 595.800 ;
        RECT 135.000 594.600 135.900 601.950 ;
        RECT 104.100 588.000 105.900 591.600 ;
        RECT 107.100 588.600 108.900 591.600 ;
        RECT 110.100 588.000 111.900 591.600 ;
        RECT 125.100 588.600 126.900 591.600 ;
        RECT 128.100 588.600 129.900 591.600 ;
        RECT 125.100 588.000 126.300 588.600 ;
        RECT 131.100 588.000 132.900 594.000 ;
        RECT 134.100 588.600 135.900 594.600 ;
        RECT 146.700 591.600 147.900 601.950 ;
        RECT 164.250 600.150 166.050 601.950 ;
        RECT 151.950 597.450 154.050 598.050 ;
        RECT 160.950 597.450 163.050 598.050 ;
        RECT 151.950 596.550 163.050 597.450 ;
        RECT 168.000 597.300 169.050 601.950 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 169.950 600.150 171.750 601.950 ;
        RECT 179.550 597.900 180.450 604.950 ;
        RECT 182.550 604.950 187.050 606.450 ;
        RECT 182.550 601.050 183.450 604.950 ;
        RECT 191.100 604.050 192.900 605.850 ;
        RECT 195.000 604.050 195.900 609.600 ;
        RECT 202.950 606.450 207.000 607.050 ;
        RECT 196.950 604.050 198.750 605.850 ;
        RECT 202.950 604.950 207.450 606.450 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 182.550 599.550 187.050 601.050 ;
        RECT 188.100 600.150 189.900 601.950 ;
        RECT 183.000 598.950 187.050 599.550 ;
        RECT 151.950 595.950 154.050 596.550 ;
        RECT 160.950 595.950 163.050 596.550 ;
        RECT 164.700 596.100 169.050 597.300 ;
        RECT 151.950 594.450 154.050 594.900 ;
        RECT 157.950 594.450 160.050 595.050 ;
        RECT 164.700 594.600 165.600 596.100 ;
        RECT 178.950 595.800 181.050 597.900 ;
        RECT 151.950 593.550 160.050 594.450 ;
        RECT 151.950 592.800 154.050 593.550 ;
        RECT 157.950 592.950 160.050 593.550 ;
        RECT 146.100 588.600 147.900 591.600 ;
        RECT 149.100 588.000 150.900 591.600 ;
        RECT 161.100 589.500 162.900 594.600 ;
        RECT 164.100 590.400 165.900 594.600 ;
        RECT 167.100 594.000 174.900 594.900 ;
        RECT 194.700 594.600 195.900 601.950 ;
        RECT 199.950 600.150 201.750 601.950 ;
        RECT 206.550 600.450 207.450 604.950 ;
        RECT 212.700 604.050 213.900 617.400 ;
        RECT 227.100 611.400 228.900 623.400 ;
        RECT 230.100 613.200 231.900 624.000 ;
        RECT 233.100 617.400 234.900 623.400 ;
        RECT 245.100 617.400 246.900 624.000 ;
        RECT 248.100 617.400 249.900 623.400 ;
        RECT 251.100 617.400 252.900 624.000 ;
        RECT 266.700 617.400 268.500 624.000 ;
        RECT 217.950 606.450 222.000 607.050 ;
        RECT 215.100 604.050 216.900 605.850 ;
        RECT 217.950 604.950 222.450 606.450 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 203.550 599.550 207.450 600.450 ;
        RECT 196.950 597.450 199.050 598.050 ;
        RECT 203.550 597.450 204.450 599.550 ;
        RECT 196.950 596.550 204.450 597.450 ;
        RECT 196.950 595.950 199.050 596.550 ;
        RECT 167.100 589.500 168.900 594.000 ;
        RECT 161.100 588.600 168.900 589.500 ;
        RECT 170.100 588.000 171.900 593.100 ;
        RECT 173.100 588.600 174.900 594.000 ;
        RECT 190.500 588.000 192.300 594.600 ;
        RECT 195.000 588.600 196.800 594.600 ;
        RECT 199.500 588.000 201.300 594.600 ;
        RECT 212.700 591.600 213.900 601.950 ;
        RECT 221.550 601.050 222.450 604.950 ;
        RECT 217.950 599.550 222.450 601.050 ;
        RECT 227.100 604.050 228.300 611.400 ;
        RECT 233.700 610.500 234.900 617.400 ;
        RECT 229.200 609.600 234.900 610.500 ;
        RECT 229.200 608.700 231.000 609.600 ;
        RECT 227.100 601.950 229.200 604.050 ;
        RECT 217.950 598.950 222.000 599.550 ;
        RECT 227.100 594.600 228.300 601.950 ;
        RECT 230.100 597.300 231.000 608.700 ;
        RECT 232.800 604.050 234.600 605.850 ;
        RECT 248.700 604.050 249.900 617.400 ;
        RECT 267.000 614.100 268.800 615.900 ;
        RECT 269.700 612.900 271.500 623.400 ;
        RECT 269.100 611.400 271.500 612.900 ;
        RECT 274.800 611.400 276.600 624.000 ;
        RECT 290.400 611.400 292.200 624.000 ;
        RECT 295.500 612.900 297.300 623.400 ;
        RECT 298.500 617.400 300.300 624.000 ;
        RECT 311.100 617.400 312.900 624.000 ;
        RECT 314.100 617.400 315.900 623.400 ;
        RECT 317.100 617.400 318.900 624.000 ;
        RECT 332.100 617.400 333.900 624.000 ;
        RECT 335.100 617.400 336.900 623.400 ;
        RECT 298.200 614.100 300.000 615.900 ;
        RECT 295.500 611.400 297.900 612.900 ;
        RECT 269.100 604.050 270.300 611.400 ;
        RECT 275.100 604.050 276.900 605.850 ;
        RECT 290.100 604.050 291.900 605.850 ;
        RECT 296.700 604.050 297.900 611.400 ;
        RECT 306.000 606.450 310.050 607.050 ;
        RECT 305.550 604.950 310.050 606.450 ;
        RECT 232.500 601.950 234.600 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 245.100 600.150 246.900 601.950 ;
        RECT 229.200 596.400 231.000 597.300 ;
        RECT 248.700 596.700 249.900 601.950 ;
        RECT 250.950 600.150 252.750 601.950 ;
        RECT 266.100 600.150 267.900 601.950 ;
        RECT 229.200 595.500 234.900 596.400 ;
        RECT 212.100 588.600 213.900 591.600 ;
        RECT 215.100 588.000 216.900 591.600 ;
        RECT 227.100 588.600 228.900 594.600 ;
        RECT 230.100 588.000 231.900 594.600 ;
        RECT 233.700 591.600 234.900 595.500 ;
        RECT 233.100 588.600 234.900 591.600 ;
        RECT 245.700 595.800 249.900 596.700 ;
        RECT 250.950 597.450 253.050 598.050 ;
        RECT 259.950 597.450 262.050 598.050 ;
        RECT 269.100 597.600 270.300 601.950 ;
        RECT 272.100 600.150 273.900 601.950 ;
        RECT 293.100 600.150 294.900 601.950 ;
        RECT 250.950 596.550 262.050 597.450 ;
        RECT 250.950 595.950 253.050 596.550 ;
        RECT 259.950 595.950 262.050 596.550 ;
        RECT 266.700 596.700 270.300 597.600 ;
        RECT 296.700 597.600 297.900 601.950 ;
        RECT 299.100 600.150 300.900 601.950 ;
        RECT 305.550 601.050 306.450 604.950 ;
        RECT 314.100 604.050 315.300 617.400 ;
        RECT 319.950 606.450 324.000 607.050 ;
        RECT 319.950 604.950 324.450 606.450 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 313.950 601.950 316.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 301.950 599.550 306.450 601.050 ;
        RECT 311.250 600.150 313.050 601.950 ;
        RECT 301.950 598.950 306.000 599.550 ;
        RECT 296.700 596.700 300.300 597.600 ;
        RECT 245.700 588.600 247.500 595.800 ;
        RECT 266.700 594.600 267.900 596.700 ;
        RECT 250.800 588.000 252.600 594.600 ;
        RECT 266.100 588.600 267.900 594.600 ;
        RECT 269.100 593.700 276.900 595.050 ;
        RECT 269.100 588.600 270.900 593.700 ;
        RECT 272.100 588.000 273.900 592.800 ;
        RECT 275.100 588.600 276.900 593.700 ;
        RECT 290.100 593.700 297.900 595.050 ;
        RECT 290.100 588.600 291.900 593.700 ;
        RECT 293.100 588.000 294.900 592.800 ;
        RECT 296.100 588.600 297.900 593.700 ;
        RECT 299.100 594.600 300.300 596.700 ;
        RECT 314.100 596.700 315.300 601.950 ;
        RECT 317.100 600.150 318.900 601.950 ;
        RECT 323.550 601.050 324.450 604.950 ;
        RECT 332.100 604.050 333.900 605.850 ;
        RECT 335.100 604.050 336.300 617.400 ;
        RECT 347.400 611.400 349.200 624.000 ;
        RECT 352.500 612.900 354.300 623.400 ;
        RECT 355.500 617.400 357.300 624.000 ;
        RECT 368.700 617.400 370.500 624.000 ;
        RECT 355.200 614.100 357.000 615.900 ;
        RECT 369.000 614.100 370.800 615.900 ;
        RECT 371.700 612.900 373.500 623.400 ;
        RECT 352.500 611.400 354.900 612.900 ;
        RECT 347.100 604.050 348.900 605.850 ;
        RECT 353.700 604.050 354.900 611.400 ;
        RECT 371.100 611.400 373.500 612.900 ;
        RECT 376.800 611.400 378.600 624.000 ;
        RECT 389.100 611.400 390.900 623.400 ;
        RECT 392.100 612.300 393.900 623.400 ;
        RECT 395.100 613.200 396.900 624.000 ;
        RECT 398.100 612.300 399.900 623.400 ;
        RECT 392.100 611.400 399.900 612.300 ;
        RECT 413.400 611.400 415.200 624.000 ;
        RECT 418.500 612.900 420.300 623.400 ;
        RECT 421.500 617.400 423.300 624.000 ;
        RECT 434.100 617.400 435.900 624.000 ;
        RECT 437.100 617.400 438.900 623.400 ;
        RECT 440.100 617.400 441.900 624.000 ;
        RECT 452.100 617.400 453.900 623.400 ;
        RECT 421.200 614.100 423.000 615.900 ;
        RECT 418.500 611.400 420.900 612.900 ;
        RECT 363.000 606.450 367.050 607.050 ;
        RECT 362.550 604.950 367.050 606.450 ;
        RECT 331.950 601.950 334.050 604.050 ;
        RECT 334.950 601.950 337.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 319.950 599.550 324.450 601.050 ;
        RECT 319.950 598.950 324.000 599.550 ;
        RECT 314.100 595.800 318.300 596.700 ;
        RECT 299.100 588.600 300.900 594.600 ;
        RECT 311.400 588.000 313.200 594.600 ;
        RECT 316.500 588.600 318.300 595.800 ;
        RECT 335.100 591.600 336.300 601.950 ;
        RECT 350.100 600.150 351.900 601.950 ;
        RECT 353.700 597.600 354.900 601.950 ;
        RECT 356.100 600.150 357.900 601.950 ;
        RECT 362.550 601.050 363.450 604.950 ;
        RECT 371.100 604.050 372.300 611.400 ;
        RECT 377.100 604.050 378.900 605.850 ;
        RECT 382.950 604.950 385.050 607.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 358.950 599.550 363.450 601.050 ;
        RECT 368.100 600.150 369.900 601.950 ;
        RECT 358.950 598.950 363.000 599.550 ;
        RECT 371.100 597.600 372.300 601.950 ;
        RECT 374.100 600.150 375.900 601.950 ;
        RECT 383.550 601.050 384.450 604.950 ;
        RECT 389.400 604.050 390.300 611.400 ;
        RECT 391.950 609.450 394.050 610.200 ;
        RECT 406.950 609.450 409.050 610.050 ;
        RECT 412.950 609.450 415.050 610.050 ;
        RECT 415.950 609.450 418.050 610.050 ;
        RECT 391.950 608.550 402.450 609.450 ;
        RECT 391.950 608.100 394.050 608.550 ;
        RECT 401.550 606.450 402.450 608.550 ;
        RECT 406.950 608.550 418.050 609.450 ;
        RECT 406.950 607.950 409.050 608.550 ;
        RECT 412.950 607.950 415.050 608.550 ;
        RECT 415.950 607.950 418.050 608.550 ;
        RECT 394.950 604.050 396.750 605.850 ;
        RECT 401.550 605.550 405.450 606.450 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 379.950 599.550 384.450 601.050 ;
        RECT 379.950 598.950 384.000 599.550 ;
        RECT 353.700 596.700 357.300 597.600 ;
        RECT 347.100 593.700 354.900 595.050 ;
        RECT 332.100 588.000 333.900 591.600 ;
        RECT 335.100 588.600 336.900 591.600 ;
        RECT 347.100 588.600 348.900 593.700 ;
        RECT 350.100 588.000 351.900 592.800 ;
        RECT 353.100 588.600 354.900 593.700 ;
        RECT 356.100 594.600 357.300 596.700 ;
        RECT 368.700 596.700 372.300 597.600 ;
        RECT 368.700 594.600 369.900 596.700 ;
        RECT 356.100 588.600 357.900 594.600 ;
        RECT 368.100 588.600 369.900 594.600 ;
        RECT 371.100 593.700 378.900 595.050 ;
        RECT 371.100 588.600 372.900 593.700 ;
        RECT 374.100 588.000 375.900 592.800 ;
        RECT 377.100 588.600 378.900 593.700 ;
        RECT 389.400 594.600 390.300 601.950 ;
        RECT 391.950 600.150 393.750 601.950 ;
        RECT 398.100 600.150 399.900 601.950 ;
        RECT 404.550 600.450 405.450 605.550 ;
        RECT 413.100 604.050 414.900 605.850 ;
        RECT 419.700 604.050 420.900 611.400 ;
        RECT 437.700 604.050 438.900 617.400 ;
        RECT 452.100 610.500 453.300 617.400 ;
        RECT 455.100 613.200 456.900 624.000 ;
        RECT 458.100 611.400 459.900 623.400 ;
        RECT 461.700 617.400 463.500 624.000 ;
        RECT 464.700 617.400 466.500 623.400 ;
        RECT 468.000 617.400 469.800 624.000 ;
        RECT 471.000 617.400 472.800 623.400 ;
        RECT 474.000 617.400 475.800 624.000 ;
        RECT 477.000 617.400 478.800 623.400 ;
        RECT 480.000 617.400 481.800 624.000 ;
        RECT 483.000 620.400 484.800 623.400 ;
        RECT 486.000 620.400 487.800 623.400 ;
        RECT 489.000 620.400 490.800 623.400 ;
        RECT 482.700 618.300 484.800 620.400 ;
        RECT 485.700 618.300 487.800 620.400 ;
        RECT 488.700 618.300 490.800 620.400 ;
        RECT 492.000 617.400 493.800 623.400 ;
        RECT 495.000 617.400 496.800 624.000 ;
        RECT 452.100 609.600 457.800 610.500 ;
        RECT 456.000 608.700 457.800 609.600 ;
        RECT 452.400 604.050 454.200 605.850 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 415.950 601.950 418.050 604.050 ;
        RECT 418.950 601.950 421.050 604.050 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 439.950 601.950 442.050 604.050 ;
        RECT 452.400 601.950 454.500 604.050 ;
        RECT 409.950 600.450 412.050 601.050 ;
        RECT 404.550 599.550 412.050 600.450 ;
        RECT 416.100 600.150 417.900 601.950 ;
        RECT 409.950 598.950 412.050 599.550 ;
        RECT 391.950 597.450 394.050 598.050 ;
        RECT 403.950 597.450 406.050 598.050 ;
        RECT 391.950 596.550 406.050 597.450 ;
        RECT 419.700 597.600 420.900 601.950 ;
        RECT 422.100 600.150 423.900 601.950 ;
        RECT 434.100 600.150 435.900 601.950 ;
        RECT 419.700 596.700 423.300 597.600 ;
        RECT 437.700 596.700 438.900 601.950 ;
        RECT 439.950 600.150 441.750 601.950 ;
        RECT 391.950 595.950 394.050 596.550 ;
        RECT 403.950 595.950 406.050 596.550 ;
        RECT 389.400 593.400 394.500 594.600 ;
        RECT 389.700 588.000 391.500 591.600 ;
        RECT 392.700 588.600 394.500 593.400 ;
        RECT 397.200 588.000 399.000 594.600 ;
        RECT 413.100 593.700 420.900 595.050 ;
        RECT 413.100 588.600 414.900 593.700 ;
        RECT 416.100 588.000 417.900 592.800 ;
        RECT 419.100 588.600 420.900 593.700 ;
        RECT 422.100 594.600 423.300 596.700 ;
        RECT 434.700 595.800 438.900 596.700 ;
        RECT 456.000 597.300 456.900 608.700 ;
        RECT 458.700 604.050 459.900 611.400 ;
        RECT 465.000 607.050 466.500 617.400 ;
        RECT 471.000 616.500 472.200 617.400 ;
        RECT 464.100 604.950 466.500 607.050 ;
        RECT 457.800 601.950 459.900 604.050 ;
        RECT 456.000 596.400 457.800 597.300 ;
        RECT 422.100 588.600 423.900 594.600 ;
        RECT 434.700 588.600 436.500 595.800 ;
        RECT 452.100 595.500 457.800 596.400 ;
        RECT 439.800 588.000 441.600 594.600 ;
        RECT 452.100 591.600 453.300 595.500 ;
        RECT 458.700 594.600 459.900 601.950 ;
        RECT 452.100 588.600 453.900 591.600 ;
        RECT 455.100 588.000 456.900 594.600 ;
        RECT 458.100 588.600 459.900 594.600 ;
        RECT 465.000 591.600 466.500 604.950 ;
        RECT 461.700 588.000 463.500 591.600 ;
        RECT 464.700 588.600 466.500 591.600 ;
        RECT 468.300 615.600 472.200 616.500 ;
        RECT 468.300 612.300 469.200 615.600 ;
        RECT 473.100 614.400 474.900 615.000 ;
        RECT 477.600 614.400 478.800 617.400 ;
        RECT 485.700 616.500 487.800 617.400 ;
        RECT 479.700 615.300 487.800 616.500 ;
        RECT 479.700 614.700 481.500 615.300 ;
        RECT 473.100 613.200 478.800 614.400 ;
        RECT 491.100 613.500 493.800 617.400 ;
        RECT 498.000 615.900 499.800 623.400 ;
        RECT 501.900 617.400 503.700 624.000 ;
        RECT 504.900 617.400 506.700 623.400 ;
        RECT 507.900 620.400 509.700 623.400 ;
        RECT 510.900 620.400 512.700 623.400 ;
        RECT 507.600 618.300 509.700 620.400 ;
        RECT 510.600 618.300 512.700 620.400 ;
        RECT 514.500 617.400 516.300 624.000 ;
        RECT 496.500 613.800 499.800 615.900 ;
        RECT 505.200 615.300 507.300 617.400 ;
        RECT 517.500 614.400 519.300 623.400 ;
        RECT 520.500 617.400 522.300 624.000 ;
        RECT 523.500 618.300 525.300 623.400 ;
        RECT 523.500 617.400 525.600 618.300 ;
        RECT 526.500 617.400 528.300 624.000 ;
        RECT 524.700 616.500 525.600 617.400 ;
        RECT 524.700 615.600 528.300 616.500 ;
        RECT 522.000 614.400 523.800 614.700 ;
        RECT 482.700 612.300 484.800 613.500 ;
        RECT 468.300 611.400 484.800 612.300 ;
        RECT 488.100 612.600 490.200 613.500 ;
        RECT 504.600 613.200 523.800 614.400 ;
        RECT 504.600 612.600 505.800 613.200 ;
        RECT 522.000 612.900 523.800 613.200 ;
        RECT 488.100 611.400 505.800 612.600 ;
        RECT 508.500 611.700 510.600 612.300 ;
        RECT 518.700 611.700 520.500 612.300 ;
        RECT 468.300 594.600 469.200 611.400 ;
        RECT 508.500 610.500 520.500 611.700 ;
        RECT 470.100 609.300 505.800 610.500 ;
        RECT 508.500 610.200 510.600 610.500 ;
        RECT 470.100 608.700 471.900 609.300 ;
        RECT 504.600 608.700 505.800 609.300 ;
        RECT 473.100 604.950 475.200 607.050 ;
        RECT 473.700 602.100 475.200 604.950 ;
        RECT 477.300 604.800 482.400 606.600 ;
        RECT 481.500 603.300 482.400 604.800 ;
        RECT 485.100 606.300 486.900 608.100 ;
        RECT 491.100 607.800 493.200 608.100 ;
        RECT 504.600 607.800 518.100 608.700 ;
        RECT 485.100 605.100 486.000 606.300 ;
        RECT 491.100 606.000 495.000 607.800 ;
        RECT 496.500 606.300 498.600 607.200 ;
        RECT 516.300 607.050 518.100 607.800 ;
        RECT 496.500 605.100 507.600 606.300 ;
        RECT 516.300 605.250 520.200 607.050 ;
        RECT 485.100 604.200 498.600 605.100 ;
        RECT 505.800 604.500 507.600 605.100 ;
        RECT 518.100 604.950 520.200 605.250 ;
        RECT 524.100 604.950 526.200 607.050 ;
        RECT 524.100 603.300 525.900 604.950 ;
        RECT 481.500 602.100 525.900 603.300 ;
        RECT 473.700 600.600 480.300 602.100 ;
        RECT 470.100 597.900 477.900 599.700 ;
        RECT 478.800 599.100 495.900 600.600 ;
        RECT 493.800 598.500 495.900 599.100 ;
        RECT 500.100 600.000 502.200 601.050 ;
        RECT 500.100 599.100 505.200 600.000 ;
        RECT 508.800 599.400 510.600 601.200 ;
        RECT 527.100 599.400 528.300 615.600 ;
        RECT 542.400 611.400 544.200 624.000 ;
        RECT 547.500 612.900 549.300 623.400 ;
        RECT 550.500 617.400 552.300 624.000 ;
        RECT 563.100 617.400 564.900 624.000 ;
        RECT 566.100 617.400 567.900 623.400 ;
        RECT 569.100 617.400 570.900 624.000 ;
        RECT 572.700 617.400 574.500 624.000 ;
        RECT 575.700 618.300 577.500 623.400 ;
        RECT 575.400 617.400 577.500 618.300 ;
        RECT 578.700 617.400 580.500 624.000 ;
        RECT 550.200 614.100 552.000 615.900 ;
        RECT 547.500 611.400 549.900 612.900 ;
        RECT 537.000 606.450 541.050 607.050 ;
        RECT 536.550 604.950 541.050 606.450 ;
        RECT 500.100 598.950 502.200 599.100 ;
        RECT 476.400 594.600 477.900 597.900 ;
        RECT 494.100 596.700 495.900 598.500 ;
        RECT 503.400 598.200 505.200 599.100 ;
        RECT 509.700 596.400 510.600 599.400 ;
        RECT 511.500 598.200 528.300 599.400 ;
        RECT 529.950 600.450 532.050 600.900 ;
        RECT 536.550 600.450 537.450 604.950 ;
        RECT 542.100 604.050 543.900 605.850 ;
        RECT 548.700 604.050 549.900 611.400 ;
        RECT 566.700 604.050 567.900 617.400 ;
        RECT 575.400 616.500 576.300 617.400 ;
        RECT 572.700 615.600 576.300 616.500 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 529.950 599.550 537.450 600.450 ;
        RECT 545.100 600.150 546.900 601.950 ;
        RECT 529.950 598.800 532.050 599.550 ;
        RECT 511.500 597.300 513.600 598.200 ;
        RECT 522.300 596.700 524.100 597.300 ;
        RECT 482.100 594.600 488.700 596.400 ;
        RECT 503.400 595.200 510.600 596.400 ;
        RECT 515.700 595.500 524.100 596.700 ;
        RECT 503.400 594.600 504.300 595.200 ;
        RECT 506.400 594.600 508.200 595.200 ;
        RECT 515.700 594.600 517.200 595.500 ;
        RECT 527.100 594.600 528.300 598.200 ;
        RECT 548.700 597.600 549.900 601.950 ;
        RECT 551.100 600.150 552.900 601.950 ;
        RECT 563.100 600.150 564.900 601.950 ;
        RECT 548.700 596.700 552.300 597.600 ;
        RECT 566.700 596.700 567.900 601.950 ;
        RECT 568.950 600.150 570.750 601.950 ;
        RECT 468.300 588.600 470.100 594.600 ;
        RECT 473.700 588.000 475.500 594.600 ;
        RECT 476.400 593.400 480.600 594.600 ;
        RECT 478.800 588.600 480.600 593.400 ;
        RECT 482.700 591.600 484.800 593.700 ;
        RECT 485.700 591.600 487.800 593.700 ;
        RECT 488.700 591.600 490.800 593.700 ;
        RECT 491.700 591.600 493.800 593.700 ;
        RECT 497.100 592.500 499.800 594.600 ;
        RECT 501.600 593.400 504.300 594.600 ;
        RECT 501.600 592.500 503.400 593.400 ;
        RECT 483.000 588.600 484.800 591.600 ;
        RECT 486.000 588.600 487.800 591.600 ;
        RECT 489.000 588.600 490.800 591.600 ;
        RECT 492.000 588.600 493.800 591.600 ;
        RECT 495.000 588.000 496.800 591.600 ;
        RECT 498.000 588.600 499.800 592.500 ;
        RECT 505.200 591.600 507.300 593.700 ;
        RECT 508.200 591.600 510.300 593.700 ;
        RECT 511.200 591.600 513.300 593.700 ;
        RECT 502.500 588.000 504.300 591.600 ;
        RECT 505.500 588.600 507.300 591.600 ;
        RECT 508.500 588.600 510.300 591.600 ;
        RECT 511.500 588.600 513.300 591.600 ;
        RECT 515.700 588.600 517.500 594.600 ;
        RECT 521.100 588.000 522.900 594.600 ;
        RECT 526.500 588.600 528.300 594.600 ;
        RECT 542.100 593.700 549.900 595.050 ;
        RECT 542.100 588.600 543.900 593.700 ;
        RECT 545.100 588.000 546.900 592.800 ;
        RECT 548.100 588.600 549.900 593.700 ;
        RECT 551.100 594.600 552.300 596.700 ;
        RECT 563.700 595.800 567.900 596.700 ;
        RECT 572.700 599.400 573.900 615.600 ;
        RECT 577.200 614.400 579.000 614.700 ;
        RECT 581.700 614.400 583.500 623.400 ;
        RECT 584.700 617.400 586.500 624.000 ;
        RECT 588.300 620.400 590.100 623.400 ;
        RECT 591.300 620.400 593.100 623.400 ;
        RECT 588.300 618.300 590.400 620.400 ;
        RECT 591.300 618.300 593.400 620.400 ;
        RECT 594.300 617.400 596.100 623.400 ;
        RECT 597.300 617.400 599.100 624.000 ;
        RECT 593.700 615.300 595.800 617.400 ;
        RECT 601.200 615.900 603.000 623.400 ;
        RECT 604.200 617.400 606.000 624.000 ;
        RECT 607.200 617.400 609.000 623.400 ;
        RECT 610.200 620.400 612.000 623.400 ;
        RECT 613.200 620.400 615.000 623.400 ;
        RECT 616.200 620.400 618.000 623.400 ;
        RECT 610.200 618.300 612.300 620.400 ;
        RECT 613.200 618.300 615.300 620.400 ;
        RECT 616.200 618.300 618.300 620.400 ;
        RECT 619.200 617.400 621.000 624.000 ;
        RECT 622.200 617.400 624.000 623.400 ;
        RECT 625.200 617.400 627.000 624.000 ;
        RECT 628.200 617.400 630.000 623.400 ;
        RECT 631.200 617.400 633.000 624.000 ;
        RECT 634.500 617.400 636.300 623.400 ;
        RECT 637.500 617.400 639.300 624.000 ;
        RECT 650.100 617.400 651.900 624.000 ;
        RECT 653.100 617.400 654.900 623.400 ;
        RECT 668.100 617.400 669.900 624.000 ;
        RECT 671.100 617.400 672.900 623.400 ;
        RECT 674.100 617.400 675.900 624.000 ;
        RECT 577.200 613.200 596.400 614.400 ;
        RECT 601.200 613.800 604.500 615.900 ;
        RECT 607.200 613.500 609.900 617.400 ;
        RECT 613.200 616.500 615.300 617.400 ;
        RECT 613.200 615.300 621.300 616.500 ;
        RECT 619.500 614.700 621.300 615.300 ;
        RECT 622.200 614.400 623.400 617.400 ;
        RECT 628.800 616.500 630.000 617.400 ;
        RECT 628.800 615.600 632.700 616.500 ;
        RECT 626.100 614.400 627.900 615.000 ;
        RECT 577.200 612.900 579.000 613.200 ;
        RECT 595.200 612.600 596.400 613.200 ;
        RECT 610.800 612.600 612.900 613.500 ;
        RECT 580.500 611.700 582.300 612.300 ;
        RECT 590.400 611.700 592.500 612.300 ;
        RECT 580.500 610.500 592.500 611.700 ;
        RECT 595.200 611.400 612.900 612.600 ;
        RECT 616.200 612.300 618.300 613.500 ;
        RECT 622.200 613.200 627.900 614.400 ;
        RECT 631.800 612.300 632.700 615.600 ;
        RECT 616.200 611.400 632.700 612.300 ;
        RECT 590.400 610.200 592.500 610.500 ;
        RECT 595.200 609.300 630.900 610.500 ;
        RECT 595.200 608.700 596.400 609.300 ;
        RECT 629.100 608.700 630.900 609.300 ;
        RECT 582.900 607.800 596.400 608.700 ;
        RECT 607.800 607.800 609.900 608.100 ;
        RECT 582.900 607.050 584.700 607.800 ;
        RECT 574.800 604.950 576.900 607.050 ;
        RECT 580.800 605.250 584.700 607.050 ;
        RECT 602.400 606.300 604.500 607.200 ;
        RECT 580.800 604.950 582.900 605.250 ;
        RECT 593.400 605.100 604.500 606.300 ;
        RECT 606.000 606.000 609.900 607.800 ;
        RECT 614.100 606.300 615.900 608.100 ;
        RECT 615.000 605.100 615.900 606.300 ;
        RECT 575.100 603.300 576.900 604.950 ;
        RECT 593.400 604.500 595.200 605.100 ;
        RECT 602.400 604.200 615.900 605.100 ;
        RECT 618.600 604.800 623.700 606.600 ;
        RECT 625.800 604.950 627.900 607.050 ;
        RECT 618.600 603.300 619.500 604.800 ;
        RECT 575.100 602.100 619.500 603.300 ;
        RECT 625.800 602.100 627.300 604.950 ;
        RECT 590.400 599.400 592.200 601.200 ;
        RECT 598.800 600.000 600.900 601.050 ;
        RECT 620.700 600.600 627.300 602.100 ;
        RECT 572.700 598.200 589.500 599.400 ;
        RECT 551.100 588.600 552.900 594.600 ;
        RECT 563.700 588.600 565.500 595.800 ;
        RECT 572.700 594.600 573.900 598.200 ;
        RECT 587.400 597.300 589.500 598.200 ;
        RECT 576.900 596.700 578.700 597.300 ;
        RECT 576.900 595.500 585.300 596.700 ;
        RECT 583.800 594.600 585.300 595.500 ;
        RECT 590.400 596.400 591.300 599.400 ;
        RECT 595.800 599.100 600.900 600.000 ;
        RECT 595.800 598.200 597.600 599.100 ;
        RECT 598.800 598.950 600.900 599.100 ;
        RECT 605.100 599.100 622.200 600.600 ;
        RECT 605.100 598.500 607.200 599.100 ;
        RECT 605.100 596.700 606.900 598.500 ;
        RECT 623.100 597.900 630.900 599.700 ;
        RECT 590.400 595.200 597.600 596.400 ;
        RECT 592.800 594.600 594.600 595.200 ;
        RECT 596.700 594.600 597.600 595.200 ;
        RECT 612.300 594.600 618.900 596.400 ;
        RECT 623.100 594.600 624.600 597.900 ;
        RECT 631.800 594.600 632.700 611.400 ;
        RECT 568.800 588.000 570.600 594.600 ;
        RECT 572.700 588.600 574.500 594.600 ;
        RECT 578.100 588.000 579.900 594.600 ;
        RECT 583.500 588.600 585.300 594.600 ;
        RECT 587.700 591.600 589.800 593.700 ;
        RECT 590.700 591.600 592.800 593.700 ;
        RECT 593.700 591.600 595.800 593.700 ;
        RECT 596.700 593.400 599.400 594.600 ;
        RECT 597.600 592.500 599.400 593.400 ;
        RECT 601.200 592.500 603.900 594.600 ;
        RECT 587.700 588.600 589.500 591.600 ;
        RECT 590.700 588.600 592.500 591.600 ;
        RECT 593.700 588.600 595.500 591.600 ;
        RECT 596.700 588.000 598.500 591.600 ;
        RECT 601.200 588.600 603.000 592.500 ;
        RECT 607.200 591.600 609.300 593.700 ;
        RECT 610.200 591.600 612.300 593.700 ;
        RECT 613.200 591.600 615.300 593.700 ;
        RECT 616.200 591.600 618.300 593.700 ;
        RECT 620.400 593.400 624.600 594.600 ;
        RECT 604.200 588.000 606.000 591.600 ;
        RECT 607.200 588.600 609.000 591.600 ;
        RECT 610.200 588.600 612.000 591.600 ;
        RECT 613.200 588.600 615.000 591.600 ;
        RECT 616.200 588.600 618.000 591.600 ;
        RECT 620.400 588.600 622.200 593.400 ;
        RECT 625.500 588.000 627.300 594.600 ;
        RECT 630.900 588.600 632.700 594.600 ;
        RECT 634.500 607.050 636.000 617.400 ;
        RECT 634.500 604.950 636.900 607.050 ;
        RECT 634.500 591.600 636.000 604.950 ;
        RECT 650.100 604.050 651.900 605.850 ;
        RECT 653.100 604.050 654.300 617.400 ;
        RECT 658.950 607.950 661.050 610.050 ;
        RECT 649.950 601.950 652.050 604.050 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 653.100 591.600 654.300 601.950 ;
        RECT 659.550 598.050 660.450 607.950 ;
        RECT 671.700 604.050 672.900 617.400 ;
        RECT 673.950 612.450 676.050 613.050 ;
        RECT 685.950 612.450 688.050 613.050 ;
        RECT 673.950 611.550 688.050 612.450 ;
        RECT 673.950 610.950 676.050 611.550 ;
        RECT 685.950 610.950 688.050 611.550 ;
        RECT 689.100 611.400 690.900 623.400 ;
        RECT 692.100 613.200 693.900 624.000 ;
        RECT 695.100 617.400 696.900 623.400 ;
        RECT 710.700 617.400 712.500 624.000 ;
        RECT 689.100 604.050 690.300 611.400 ;
        RECT 695.700 610.500 696.900 617.400 ;
        RECT 711.000 614.100 712.800 615.900 ;
        RECT 713.700 612.900 715.500 623.400 ;
        RECT 691.200 609.600 696.900 610.500 ;
        RECT 713.100 611.400 715.500 612.900 ;
        RECT 718.800 611.400 720.600 624.000 ;
        RECT 731.100 611.400 732.900 623.400 ;
        RECT 734.100 612.300 735.900 623.400 ;
        RECT 737.100 613.200 738.900 624.000 ;
        RECT 740.100 612.300 741.900 623.400 ;
        RECT 734.100 611.400 741.900 612.300 ;
        RECT 755.100 611.400 756.900 624.000 ;
        RECT 760.200 612.600 762.000 623.400 ;
        RECT 773.100 617.400 774.900 624.000 ;
        RECT 776.100 617.400 777.900 623.400 ;
        RECT 779.100 617.400 780.900 624.000 ;
        RECT 791.100 617.400 792.900 623.400 ;
        RECT 794.100 617.400 795.900 624.000 ;
        RECT 758.400 611.400 762.000 612.600 ;
        RECT 691.200 608.700 693.000 609.600 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 689.100 601.950 691.200 604.050 ;
        RECT 668.100 600.150 669.900 601.950 ;
        RECT 659.550 597.900 663.000 598.050 ;
        RECT 659.550 596.550 664.050 597.900 ;
        RECT 671.700 596.700 672.900 601.950 ;
        RECT 673.950 600.150 675.750 601.950 ;
        RECT 660.000 595.950 664.050 596.550 ;
        RECT 661.950 595.800 664.050 595.950 ;
        RECT 668.700 595.800 672.900 596.700 ;
        RECT 634.500 588.600 636.300 591.600 ;
        RECT 637.500 588.000 639.300 591.600 ;
        RECT 650.100 588.000 651.900 591.600 ;
        RECT 653.100 588.600 654.900 591.600 ;
        RECT 668.700 588.600 670.500 595.800 ;
        RECT 689.100 594.600 690.300 601.950 ;
        RECT 692.100 597.300 693.000 608.700 ;
        RECT 694.800 604.050 696.600 605.850 ;
        RECT 713.100 604.050 714.300 611.400 ;
        RECT 727.950 606.450 730.050 610.050 ;
        RECT 725.550 606.000 730.050 606.450 ;
        RECT 719.100 604.050 720.900 605.850 ;
        RECT 725.550 605.550 729.450 606.000 ;
        RECT 694.500 601.950 696.600 604.050 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 715.950 601.950 718.050 604.050 ;
        RECT 718.950 601.950 721.050 604.050 ;
        RECT 710.100 600.150 711.900 601.950 ;
        RECT 713.100 597.600 714.300 601.950 ;
        RECT 716.100 600.150 717.900 601.950 ;
        RECT 725.550 601.050 726.450 605.550 ;
        RECT 731.400 604.050 732.300 611.400 ;
        RECT 742.950 606.450 745.050 607.050 ;
        RECT 748.950 606.450 751.050 607.050 ;
        RECT 736.950 604.050 738.750 605.850 ;
        RECT 742.950 605.550 751.050 606.450 ;
        RECT 742.950 604.950 745.050 605.550 ;
        RECT 748.950 604.950 751.050 605.550 ;
        RECT 755.250 604.050 757.050 605.850 ;
        RECT 758.400 604.050 759.300 611.400 ;
        RECT 763.950 609.450 766.050 610.050 ;
        RECT 772.950 609.450 775.050 610.050 ;
        RECT 763.950 608.550 775.050 609.450 ;
        RECT 763.950 607.950 766.050 608.550 ;
        RECT 772.950 607.950 775.050 608.550 ;
        RECT 768.000 606.450 772.050 607.050 ;
        RECT 761.100 604.050 762.900 605.850 ;
        RECT 767.550 604.950 772.050 606.450 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 721.950 599.550 726.450 601.050 ;
        RECT 721.950 598.950 726.000 599.550 ;
        RECT 691.200 596.400 693.000 597.300 ;
        RECT 710.700 596.700 714.300 597.600 ;
        RECT 691.200 595.500 696.900 596.400 ;
        RECT 673.800 588.000 675.600 594.600 ;
        RECT 689.100 588.600 690.900 594.600 ;
        RECT 692.100 588.000 693.900 594.600 ;
        RECT 695.700 591.600 696.900 595.500 ;
        RECT 710.700 594.600 711.900 596.700 ;
        RECT 695.100 588.600 696.900 591.600 ;
        RECT 710.100 588.600 711.900 594.600 ;
        RECT 713.100 593.700 720.900 595.050 ;
        RECT 713.100 588.600 714.900 593.700 ;
        RECT 716.100 588.000 717.900 592.800 ;
        RECT 719.100 588.600 720.900 593.700 ;
        RECT 731.400 594.600 732.300 601.950 ;
        RECT 733.950 600.150 735.750 601.950 ;
        RECT 740.100 600.150 741.900 601.950 ;
        RECT 731.400 593.400 736.500 594.600 ;
        RECT 731.700 588.000 733.500 591.600 ;
        RECT 734.700 588.600 736.500 593.400 ;
        RECT 739.200 588.000 741.000 594.600 ;
        RECT 758.400 591.600 759.300 601.950 ;
        RECT 767.550 601.050 768.450 604.950 ;
        RECT 776.700 604.050 777.900 617.400 ;
        RECT 791.700 604.050 792.900 617.400 ;
        RECT 809.100 612.600 810.900 623.400 ;
        RECT 812.100 613.500 813.900 624.000 ;
        RECT 815.100 622.500 822.900 623.400 ;
        RECT 815.100 612.600 816.900 622.500 ;
        RECT 809.100 611.700 816.900 612.600 ;
        RECT 818.100 610.500 819.900 621.600 ;
        RECT 821.100 611.400 822.900 622.500 ;
        RECT 833.100 617.400 834.900 623.400 ;
        RECT 836.100 618.000 837.900 624.000 ;
        RECT 834.000 617.100 834.900 617.400 ;
        RECT 839.100 617.400 840.900 623.400 ;
        RECT 842.100 617.400 843.900 624.000 ;
        RECT 854.100 622.500 861.900 623.400 ;
        RECT 839.100 617.100 840.600 617.400 ;
        RECT 834.000 616.200 840.600 617.100 ;
        RECT 815.100 609.600 819.900 610.500 ;
        RECT 796.950 606.450 801.000 607.050 ;
        RECT 794.100 604.050 795.900 605.850 ;
        RECT 796.950 604.950 801.450 606.450 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 763.950 599.550 768.450 601.050 ;
        RECT 773.100 600.150 774.900 601.950 ;
        RECT 763.950 598.950 768.000 599.550 ;
        RECT 776.700 596.700 777.900 601.950 ;
        RECT 778.950 600.150 780.750 601.950 ;
        RECT 773.700 595.800 777.900 596.700 ;
        RECT 755.100 588.000 756.900 591.600 ;
        RECT 758.100 588.600 759.900 591.600 ;
        RECT 761.100 588.000 762.900 591.600 ;
        RECT 773.700 588.600 775.500 595.800 ;
        RECT 778.800 588.000 780.600 594.600 ;
        RECT 791.700 591.600 792.900 601.950 ;
        RECT 800.550 600.900 801.450 604.950 ;
        RECT 812.250 604.050 814.050 605.850 ;
        RECT 815.100 604.050 816.000 609.600 ;
        RECT 818.100 604.050 819.900 605.850 ;
        RECT 834.000 604.050 834.900 616.200 ;
        RECT 854.100 611.400 855.900 622.500 ;
        RECT 857.100 610.500 858.900 621.600 ;
        RECT 860.100 612.600 861.900 622.500 ;
        RECT 863.100 613.500 864.900 624.000 ;
        RECT 866.100 612.600 867.900 623.400 ;
        RECT 860.100 611.700 867.900 612.600 ;
        RECT 881.100 611.400 882.900 623.400 ;
        RECT 884.100 612.000 885.900 624.000 ;
        RECT 887.100 617.400 888.900 623.400 ;
        RECT 890.100 617.400 891.900 624.000 ;
        RECT 857.100 609.600 861.900 610.500 ;
        RECT 839.100 604.050 840.900 605.850 ;
        RECT 857.100 604.050 858.900 605.850 ;
        RECT 861.000 604.050 861.900 609.600 ;
        RECT 862.950 609.450 865.050 610.050 ;
        RECT 877.950 609.450 880.050 610.050 ;
        RECT 862.950 608.550 880.050 609.450 ;
        RECT 862.950 607.950 865.050 608.550 ;
        RECT 877.950 607.950 880.050 608.550 ;
        RECT 862.950 604.050 864.750 605.850 ;
        RECT 881.700 604.050 882.600 611.400 ;
        RECT 885.000 604.050 886.800 605.850 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 881.100 601.950 883.200 604.050 ;
        RECT 884.400 601.950 886.500 604.050 ;
        RECT 799.950 598.800 802.050 600.900 ;
        RECT 809.250 600.150 811.050 601.950 ;
        RECT 815.100 594.600 816.300 601.950 ;
        RECT 821.100 600.150 822.900 601.950 ;
        RECT 834.000 598.200 834.900 601.950 ;
        RECT 836.100 600.150 837.900 601.950 ;
        RECT 842.100 600.150 843.900 601.950 ;
        RECT 854.100 600.150 855.900 601.950 ;
        RECT 834.000 597.000 837.300 598.200 ;
        RECT 791.100 588.600 792.900 591.600 ;
        RECT 794.100 588.000 795.900 591.600 ;
        RECT 809.700 588.000 811.500 594.600 ;
        RECT 814.200 588.600 816.000 594.600 ;
        RECT 818.700 588.000 820.500 594.600 ;
        RECT 835.500 588.600 837.300 597.000 ;
        RECT 842.100 588.000 843.900 597.600 ;
        RECT 860.700 594.600 861.900 601.950 ;
        RECT 865.950 600.150 867.750 601.950 ;
        RECT 881.700 594.600 882.600 601.950 ;
        RECT 888.000 597.300 888.900 617.400 ;
        RECT 902.400 611.400 904.200 624.000 ;
        RECT 907.500 612.900 909.300 623.400 ;
        RECT 910.500 617.400 912.300 624.000 ;
        RECT 926.100 617.400 927.900 624.000 ;
        RECT 929.100 617.400 930.900 623.400 ;
        RECT 932.100 617.400 933.900 624.000 ;
        RECT 910.200 614.100 912.000 615.900 ;
        RECT 925.950 615.450 928.050 616.050 ;
        RECT 917.550 615.000 928.050 615.450 ;
        RECT 916.950 614.550 928.050 615.000 ;
        RECT 907.500 611.400 909.900 612.900 ;
        RECT 902.100 604.050 903.900 605.850 ;
        RECT 908.700 604.050 909.900 611.400 ;
        RECT 916.950 610.950 919.050 614.550 ;
        RECT 925.950 613.950 928.050 614.550 ;
        RECT 921.000 606.450 925.050 607.050 ;
        RECT 920.550 604.950 925.050 606.450 ;
        RECT 889.800 601.950 891.900 604.050 ;
        RECT 901.950 601.950 904.050 604.050 ;
        RECT 904.950 601.950 907.050 604.050 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 889.950 600.150 891.750 601.950 ;
        RECT 905.100 600.150 906.900 601.950 ;
        RECT 908.700 597.600 909.900 601.950 ;
        RECT 911.100 600.150 912.900 601.950 ;
        RECT 913.950 600.450 916.050 601.050 ;
        RECT 920.550 600.450 921.450 604.950 ;
        RECT 929.100 604.050 930.300 617.400 ;
        RECT 925.950 601.950 928.050 604.050 ;
        RECT 928.950 601.950 931.050 604.050 ;
        RECT 931.950 601.950 934.050 604.050 ;
        RECT 913.950 599.550 921.450 600.450 ;
        RECT 926.250 600.150 928.050 601.950 ;
        RECT 913.950 598.950 916.050 599.550 ;
        RECT 883.500 596.400 891.900 597.300 ;
        RECT 908.700 596.700 912.300 597.600 ;
        RECT 883.500 595.500 885.300 596.400 ;
        RECT 856.500 588.000 858.300 594.600 ;
        RECT 861.000 588.600 862.800 594.600 ;
        RECT 865.500 588.000 867.300 594.600 ;
        RECT 881.700 592.800 884.400 594.600 ;
        RECT 882.600 588.600 884.400 592.800 ;
        RECT 885.600 588.000 887.400 594.600 ;
        RECT 890.100 588.600 891.900 596.400 ;
        RECT 902.100 593.700 909.900 595.050 ;
        RECT 902.100 588.600 903.900 593.700 ;
        RECT 905.100 588.000 906.900 592.800 ;
        RECT 908.100 588.600 909.900 593.700 ;
        RECT 911.100 594.600 912.300 596.700 ;
        RECT 929.100 596.700 930.300 601.950 ;
        RECT 932.100 600.150 933.900 601.950 ;
        RECT 929.100 595.800 933.300 596.700 ;
        RECT 911.100 588.600 912.900 594.600 ;
        RECT 926.400 588.000 928.200 594.600 ;
        RECT 931.500 588.600 933.300 595.800 ;
        RECT 11.100 578.400 12.900 584.400 ;
        RECT 14.100 578.400 15.900 585.000 ;
        RECT 17.100 581.400 18.900 584.400 ;
        RECT 11.100 571.050 12.300 578.400 ;
        RECT 17.700 577.500 18.900 581.400 ;
        RECT 29.100 579.300 30.900 584.400 ;
        RECT 32.100 580.200 33.900 585.000 ;
        RECT 35.100 579.300 36.900 584.400 ;
        RECT 29.100 577.950 36.900 579.300 ;
        RECT 38.100 578.400 39.900 584.400 ;
        RECT 13.200 576.600 18.900 577.500 ;
        RECT 13.200 575.700 15.000 576.600 ;
        RECT 38.100 576.300 39.300 578.400 ;
        RECT 50.700 577.200 52.500 584.400 ;
        RECT 55.800 578.400 57.600 585.000 ;
        RECT 71.700 578.400 73.500 585.000 ;
        RECT 76.200 578.400 78.000 584.400 ;
        RECT 80.700 578.400 82.500 585.000 ;
        RECT 95.100 581.400 96.900 584.400 ;
        RECT 98.100 581.400 99.900 585.000 ;
        RECT 50.700 576.300 54.900 577.200 ;
        RECT 11.100 568.950 13.200 571.050 ;
        RECT 11.100 561.600 12.300 568.950 ;
        RECT 14.100 564.300 15.000 575.700 ;
        RECT 35.700 575.400 39.300 576.300 ;
        RECT 32.100 571.050 33.900 572.850 ;
        RECT 35.700 571.050 36.900 575.400 ;
        RECT 40.950 573.450 45.000 574.050 ;
        RECT 38.100 571.050 39.900 572.850 ;
        RECT 40.950 571.950 45.450 573.450 ;
        RECT 16.500 568.950 18.600 571.050 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 16.800 567.150 18.600 568.950 ;
        RECT 29.100 567.150 30.900 568.950 ;
        RECT 13.200 563.400 15.000 564.300 ;
        RECT 13.200 562.500 18.900 563.400 ;
        RECT 11.100 549.600 12.900 561.600 ;
        RECT 14.100 549.000 15.900 559.800 ;
        RECT 17.700 555.600 18.900 562.500 ;
        RECT 35.700 561.600 36.900 568.950 ;
        RECT 44.550 568.050 45.450 571.950 ;
        RECT 50.100 571.050 51.900 572.850 ;
        RECT 53.700 571.050 54.900 576.300 ;
        RECT 64.950 576.450 67.050 577.050 ;
        RECT 73.950 576.450 76.050 577.050 ;
        RECT 64.950 575.550 76.050 576.450 ;
        RECT 64.950 574.950 67.050 575.550 ;
        RECT 73.950 574.950 76.050 575.550 ;
        RECT 55.950 571.050 57.750 572.850 ;
        RECT 71.250 571.050 73.050 572.850 ;
        RECT 77.100 571.050 78.300 578.400 ;
        RECT 83.100 571.050 84.900 572.850 ;
        RECT 95.700 571.050 96.900 581.400 ;
        RECT 110.100 579.300 111.900 584.400 ;
        RECT 113.100 580.200 114.900 585.000 ;
        RECT 116.100 579.300 117.900 584.400 ;
        RECT 110.100 577.950 117.900 579.300 ;
        RECT 119.100 578.400 120.900 584.400 ;
        RECT 119.100 576.300 120.300 578.400 ;
        RECT 124.950 577.950 127.050 580.050 ;
        RECT 116.700 575.400 120.300 576.300 ;
        RECT 105.000 573.450 109.050 574.050 ;
        RECT 104.550 571.950 109.050 573.450 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 44.550 566.550 49.050 568.050 ;
        RECT 45.000 565.950 49.050 566.550 ;
        RECT 17.100 549.600 18.900 555.600 ;
        RECT 29.400 549.000 31.200 561.600 ;
        RECT 34.500 560.100 36.900 561.600 ;
        RECT 34.500 549.600 36.300 560.100 ;
        RECT 37.200 557.100 39.000 558.900 ;
        RECT 53.700 555.600 54.900 568.950 ;
        RECT 74.250 567.150 76.050 568.950 ;
        RECT 55.950 564.450 58.050 565.050 ;
        RECT 73.950 564.450 76.050 565.050 ;
        RECT 55.950 563.550 76.050 564.450 ;
        RECT 55.950 562.950 58.050 563.550 ;
        RECT 73.950 562.950 76.050 563.550 ;
        RECT 77.100 563.400 78.000 568.950 ;
        RECT 80.100 567.150 81.900 568.950 ;
        RECT 77.100 562.500 81.900 563.400 ;
        RECT 71.100 560.400 78.900 561.300 ;
        RECT 37.500 549.000 39.300 555.600 ;
        RECT 50.100 549.000 51.900 555.600 ;
        RECT 53.100 549.600 54.900 555.600 ;
        RECT 56.100 549.000 57.900 555.600 ;
        RECT 71.100 549.600 72.900 560.400 ;
        RECT 74.100 549.000 75.900 559.500 ;
        RECT 77.100 550.500 78.900 560.400 ;
        RECT 80.100 551.400 81.900 562.500 ;
        RECT 83.100 550.500 84.900 561.600 ;
        RECT 95.700 555.600 96.900 568.950 ;
        RECT 98.100 567.150 99.900 568.950 ;
        RECT 104.550 568.050 105.450 571.950 ;
        RECT 113.100 571.050 114.900 572.850 ;
        RECT 116.700 571.050 117.900 575.400 ;
        RECT 119.100 571.050 120.900 572.850 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 100.950 566.550 105.450 568.050 ;
        RECT 110.100 567.150 111.900 568.950 ;
        RECT 100.950 565.950 105.000 566.550 ;
        RECT 116.700 561.600 117.900 568.950 ;
        RECT 125.550 568.050 126.450 577.950 ;
        RECT 131.100 575.400 132.900 585.000 ;
        RECT 137.700 576.000 139.500 584.400 ;
        RECT 152.100 579.300 153.900 584.400 ;
        RECT 155.100 580.200 156.900 585.000 ;
        RECT 158.100 579.300 159.900 584.400 ;
        RECT 152.100 577.950 159.900 579.300 ;
        RECT 161.100 578.400 162.900 584.400 ;
        RECT 177.600 580.200 179.400 584.400 ;
        RECT 176.700 578.400 179.400 580.200 ;
        RECT 180.600 578.400 182.400 585.000 ;
        RECT 161.100 576.300 162.300 578.400 ;
        RECT 137.700 574.800 141.000 576.000 ;
        RECT 131.100 571.050 132.900 572.850 ;
        RECT 137.100 571.050 138.900 572.850 ;
        RECT 140.100 571.050 141.000 574.800 ;
        RECT 158.700 575.400 162.300 576.300 ;
        RECT 142.950 573.450 147.000 574.050 ;
        RECT 142.950 571.950 147.450 573.450 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 125.550 566.550 130.050 568.050 ;
        RECT 134.100 567.150 135.900 568.950 ;
        RECT 126.000 565.950 130.050 566.550 ;
        RECT 77.100 549.600 84.900 550.500 ;
        RECT 95.100 549.600 96.900 555.600 ;
        RECT 98.100 549.000 99.900 555.600 ;
        RECT 110.400 549.000 112.200 561.600 ;
        RECT 115.500 560.100 117.900 561.600 ;
        RECT 115.500 549.600 117.300 560.100 ;
        RECT 118.200 557.100 120.000 558.900 ;
        RECT 140.100 556.800 141.000 568.950 ;
        RECT 146.550 567.450 147.450 571.950 ;
        RECT 155.100 571.050 156.900 572.850 ;
        RECT 158.700 571.050 159.900 575.400 ;
        RECT 161.100 571.050 162.900 572.850 ;
        RECT 176.700 571.050 177.600 578.400 ;
        RECT 178.500 576.600 180.300 577.500 ;
        RECT 185.100 576.600 186.900 584.400 ;
        RECT 200.700 581.400 202.500 585.000 ;
        RECT 203.700 579.600 205.500 584.400 ;
        RECT 178.500 575.700 186.900 576.600 ;
        RECT 200.400 578.400 205.500 579.600 ;
        RECT 208.200 578.400 210.000 585.000 ;
        RECT 221.100 581.400 222.900 584.400 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 176.100 568.950 178.200 571.050 ;
        RECT 179.400 568.950 181.500 571.050 ;
        RECT 146.550 566.550 150.450 567.450 ;
        RECT 152.100 567.150 153.900 568.950 ;
        RECT 149.550 565.050 150.450 566.550 ;
        RECT 149.550 563.550 154.050 565.050 ;
        RECT 150.000 562.950 154.050 563.550 ;
        RECT 158.700 561.600 159.900 568.950 ;
        RECT 160.950 564.450 163.050 565.050 ;
        RECT 172.950 564.450 175.050 564.900 ;
        RECT 160.950 563.550 175.050 564.450 ;
        RECT 160.950 562.950 163.050 563.550 ;
        RECT 172.950 562.800 175.050 563.550 ;
        RECT 176.700 561.600 177.600 568.950 ;
        RECT 180.000 567.150 181.800 568.950 ;
        RECT 134.400 555.900 141.000 556.800 ;
        RECT 134.400 555.600 135.900 555.900 ;
        RECT 118.500 549.000 120.300 555.600 ;
        RECT 131.100 549.000 132.900 555.600 ;
        RECT 134.100 549.600 135.900 555.600 ;
        RECT 140.100 555.600 141.000 555.900 ;
        RECT 137.100 549.000 138.900 555.000 ;
        RECT 140.100 549.600 141.900 555.600 ;
        RECT 152.400 549.000 154.200 561.600 ;
        RECT 157.500 560.100 159.900 561.600 ;
        RECT 157.500 549.600 159.300 560.100 ;
        RECT 160.200 557.100 162.000 558.900 ;
        RECT 160.500 549.000 162.300 555.600 ;
        RECT 176.100 549.600 177.900 561.600 ;
        RECT 179.100 549.000 180.900 561.000 ;
        RECT 183.000 555.600 183.900 575.700 ;
        RECT 184.950 571.050 186.750 572.850 ;
        RECT 200.400 571.050 201.300 578.400 ;
        RECT 221.100 577.500 222.300 581.400 ;
        RECT 224.100 578.400 225.900 585.000 ;
        RECT 227.100 578.400 228.900 584.400 ;
        RECT 221.100 576.600 226.800 577.500 ;
        RECT 225.000 575.700 226.800 576.600 ;
        RECT 211.950 573.450 216.000 574.050 ;
        RECT 202.950 571.050 204.750 572.850 ;
        RECT 209.100 571.050 210.900 572.850 ;
        RECT 211.950 571.950 216.450 573.450 ;
        RECT 184.800 568.950 186.900 571.050 ;
        RECT 199.950 568.950 202.050 571.050 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 200.400 561.600 201.300 568.950 ;
        RECT 205.950 567.150 207.750 568.950 ;
        RECT 215.550 568.050 216.450 571.950 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 221.400 568.950 223.500 571.050 ;
        RECT 211.950 566.550 216.450 568.050 ;
        RECT 211.950 565.950 216.000 566.550 ;
        RECT 208.950 564.450 211.050 564.750 ;
        RECT 218.550 564.450 219.450 568.950 ;
        RECT 221.400 567.150 223.200 568.950 ;
        RECT 208.950 563.550 219.450 564.450 ;
        RECT 225.000 564.300 225.900 575.700 ;
        RECT 227.700 571.050 228.900 578.400 ;
        RECT 226.800 568.950 228.900 571.050 ;
        RECT 208.950 562.650 211.050 563.550 ;
        RECT 225.000 563.400 226.800 564.300 ;
        RECT 221.100 562.500 226.800 563.400 ;
        RECT 182.100 549.600 183.900 555.600 ;
        RECT 185.100 549.000 186.900 555.600 ;
        RECT 200.100 549.600 201.900 561.600 ;
        RECT 203.100 560.700 210.900 561.600 ;
        RECT 203.100 549.600 204.900 560.700 ;
        RECT 206.100 549.000 207.900 559.800 ;
        RECT 209.100 549.600 210.900 560.700 ;
        RECT 221.100 555.600 222.300 562.500 ;
        RECT 227.700 561.600 228.900 568.950 ;
        RECT 221.100 549.600 222.900 555.600 ;
        RECT 224.100 549.000 225.900 559.800 ;
        RECT 227.100 549.600 228.900 561.600 ;
        RECT 230.700 578.400 232.500 584.400 ;
        RECT 236.100 578.400 237.900 585.000 ;
        RECT 241.500 578.400 243.300 584.400 ;
        RECT 245.700 581.400 247.500 584.400 ;
        RECT 248.700 581.400 250.500 584.400 ;
        RECT 251.700 581.400 253.500 584.400 ;
        RECT 254.700 581.400 256.500 585.000 ;
        RECT 245.700 579.300 247.800 581.400 ;
        RECT 248.700 579.300 250.800 581.400 ;
        RECT 251.700 579.300 253.800 581.400 ;
        RECT 259.200 580.500 261.000 584.400 ;
        RECT 262.200 581.400 264.000 585.000 ;
        RECT 265.200 581.400 267.000 584.400 ;
        RECT 268.200 581.400 270.000 584.400 ;
        RECT 271.200 581.400 273.000 584.400 ;
        RECT 274.200 581.400 276.000 584.400 ;
        RECT 255.600 579.600 257.400 580.500 ;
        RECT 254.700 578.400 257.400 579.600 ;
        RECT 259.200 578.400 261.900 580.500 ;
        RECT 265.200 579.300 267.300 581.400 ;
        RECT 268.200 579.300 270.300 581.400 ;
        RECT 271.200 579.300 273.300 581.400 ;
        RECT 274.200 579.300 276.300 581.400 ;
        RECT 278.400 579.600 280.200 584.400 ;
        RECT 278.400 578.400 282.600 579.600 ;
        RECT 283.500 578.400 285.300 585.000 ;
        RECT 288.900 578.400 290.700 584.400 ;
        RECT 230.700 574.800 231.900 578.400 ;
        RECT 241.800 577.500 243.300 578.400 ;
        RECT 250.800 577.800 252.600 578.400 ;
        RECT 254.700 577.800 255.600 578.400 ;
        RECT 234.900 576.300 243.300 577.500 ;
        RECT 248.400 576.600 255.600 577.800 ;
        RECT 270.300 576.600 276.900 578.400 ;
        RECT 234.900 575.700 236.700 576.300 ;
        RECT 245.400 574.800 247.500 575.700 ;
        RECT 230.700 573.600 247.500 574.800 ;
        RECT 248.400 573.600 249.300 576.600 ;
        RECT 253.800 573.900 255.600 574.800 ;
        RECT 263.100 574.500 264.900 576.300 ;
        RECT 281.100 575.100 282.600 578.400 ;
        RECT 256.800 573.900 258.900 574.050 ;
        RECT 230.700 557.400 231.900 573.600 ;
        RECT 248.400 571.800 250.200 573.600 ;
        RECT 253.800 573.000 258.900 573.900 ;
        RECT 256.800 571.950 258.900 573.000 ;
        RECT 263.100 573.900 265.200 574.500 ;
        RECT 263.100 572.400 280.200 573.900 ;
        RECT 281.100 573.300 288.900 575.100 ;
        RECT 278.700 570.900 285.300 572.400 ;
        RECT 233.100 569.700 277.500 570.900 ;
        RECT 233.100 568.050 234.900 569.700 ;
        RECT 232.800 565.950 234.900 568.050 ;
        RECT 238.800 567.750 240.900 568.050 ;
        RECT 251.400 567.900 253.200 568.500 ;
        RECT 260.400 567.900 273.900 568.800 ;
        RECT 238.800 565.950 242.700 567.750 ;
        RECT 251.400 566.700 262.500 567.900 ;
        RECT 240.900 565.200 242.700 565.950 ;
        RECT 260.400 565.800 262.500 566.700 ;
        RECT 264.000 565.200 267.900 567.000 ;
        RECT 273.000 566.700 273.900 567.900 ;
        RECT 240.900 564.300 254.400 565.200 ;
        RECT 265.800 564.900 267.900 565.200 ;
        RECT 272.100 564.900 273.900 566.700 ;
        RECT 276.600 568.200 277.500 569.700 ;
        RECT 276.600 566.400 281.700 568.200 ;
        RECT 283.800 568.050 285.300 570.900 ;
        RECT 283.800 565.950 285.900 568.050 ;
        RECT 253.200 563.700 254.400 564.300 ;
        RECT 287.100 563.700 288.900 564.300 ;
        RECT 248.400 562.500 250.500 562.800 ;
        RECT 253.200 562.500 288.900 563.700 ;
        RECT 238.500 561.300 250.500 562.500 ;
        RECT 289.800 561.600 290.700 578.400 ;
        RECT 238.500 560.700 240.300 561.300 ;
        RECT 248.400 560.700 250.500 561.300 ;
        RECT 253.200 560.400 270.900 561.600 ;
        RECT 235.200 559.800 237.000 560.100 ;
        RECT 253.200 559.800 254.400 560.400 ;
        RECT 235.200 558.600 254.400 559.800 ;
        RECT 268.800 559.500 270.900 560.400 ;
        RECT 274.200 560.700 290.700 561.600 ;
        RECT 274.200 559.500 276.300 560.700 ;
        RECT 235.200 558.300 237.000 558.600 ;
        RECT 230.700 556.500 234.300 557.400 ;
        RECT 233.400 555.600 234.300 556.500 ;
        RECT 230.700 549.000 232.500 555.600 ;
        RECT 233.400 554.700 235.500 555.600 ;
        RECT 233.700 549.600 235.500 554.700 ;
        RECT 236.700 549.000 238.500 555.600 ;
        RECT 239.700 549.600 241.500 558.600 ;
        RECT 251.700 555.600 253.800 557.700 ;
        RECT 259.200 557.100 262.500 559.200 ;
        RECT 242.700 549.000 244.500 555.600 ;
        RECT 246.300 552.600 248.400 554.700 ;
        RECT 249.300 552.600 251.400 554.700 ;
        RECT 246.300 549.600 248.100 552.600 ;
        RECT 249.300 549.600 251.100 552.600 ;
        RECT 252.300 549.600 254.100 555.600 ;
        RECT 255.300 549.000 257.100 555.600 ;
        RECT 259.200 549.600 261.000 557.100 ;
        RECT 265.200 555.600 267.900 559.500 ;
        RECT 280.200 558.600 285.900 559.800 ;
        RECT 277.500 557.700 279.300 558.300 ;
        RECT 271.200 556.500 279.300 557.700 ;
        RECT 271.200 555.600 273.300 556.500 ;
        RECT 280.200 555.600 281.400 558.600 ;
        RECT 284.100 558.000 285.900 558.600 ;
        RECT 289.800 557.400 290.700 560.700 ;
        RECT 286.800 556.500 290.700 557.400 ;
        RECT 292.500 581.400 294.300 584.400 ;
        RECT 295.500 581.400 297.300 585.000 ;
        RECT 292.500 568.050 294.000 581.400 ;
        RECT 308.400 578.400 310.200 585.000 ;
        RECT 313.500 577.200 315.300 584.400 ;
        RECT 329.100 578.400 330.900 584.400 ;
        RECT 311.100 576.300 315.300 577.200 ;
        RECT 329.700 576.300 330.900 578.400 ;
        RECT 332.100 579.300 333.900 584.400 ;
        RECT 335.100 580.200 336.900 585.000 ;
        RECT 338.100 579.300 339.900 584.400 ;
        RECT 332.100 577.950 339.900 579.300 ;
        RECT 353.100 579.300 354.900 584.400 ;
        RECT 356.100 580.200 357.900 585.000 ;
        RECT 359.100 579.300 360.900 584.400 ;
        RECT 353.100 577.950 360.900 579.300 ;
        RECT 362.100 578.400 363.900 584.400 ;
        RECT 362.100 576.300 363.300 578.400 ;
        RECT 374.700 577.200 376.500 584.400 ;
        RECT 379.800 578.400 381.600 585.000 ;
        RECT 395.700 577.200 397.500 584.400 ;
        RECT 400.800 578.400 402.600 585.000 ;
        RECT 413.100 579.300 414.900 584.400 ;
        RECT 416.100 580.200 417.900 585.000 ;
        RECT 419.100 579.300 420.900 584.400 ;
        RECT 413.100 577.950 420.900 579.300 ;
        RECT 422.100 578.400 423.900 584.400 ;
        RECT 425.700 578.400 427.500 584.400 ;
        RECT 431.100 578.400 432.900 585.000 ;
        RECT 436.500 578.400 438.300 584.400 ;
        RECT 440.700 581.400 442.500 584.400 ;
        RECT 443.700 581.400 445.500 584.400 ;
        RECT 446.700 581.400 448.500 584.400 ;
        RECT 449.700 581.400 451.500 585.000 ;
        RECT 440.700 579.300 442.800 581.400 ;
        RECT 443.700 579.300 445.800 581.400 ;
        RECT 446.700 579.300 448.800 581.400 ;
        RECT 454.200 580.500 456.000 584.400 ;
        RECT 457.200 581.400 459.000 585.000 ;
        RECT 460.200 581.400 462.000 584.400 ;
        RECT 463.200 581.400 465.000 584.400 ;
        RECT 466.200 581.400 468.000 584.400 ;
        RECT 469.200 581.400 471.000 584.400 ;
        RECT 450.600 579.600 452.400 580.500 ;
        RECT 449.700 578.400 452.400 579.600 ;
        RECT 454.200 578.400 456.900 580.500 ;
        RECT 460.200 579.300 462.300 581.400 ;
        RECT 463.200 579.300 465.300 581.400 ;
        RECT 466.200 579.300 468.300 581.400 ;
        RECT 469.200 579.300 471.300 581.400 ;
        RECT 473.400 579.600 475.200 584.400 ;
        RECT 473.400 578.400 477.600 579.600 ;
        RECT 478.500 578.400 480.300 585.000 ;
        RECT 483.900 578.400 485.700 584.400 ;
        RECT 374.700 576.300 378.900 577.200 ;
        RECT 395.700 576.300 399.900 577.200 ;
        RECT 422.100 576.300 423.300 578.400 ;
        RECT 295.950 571.950 298.050 574.050 ;
        RECT 292.500 565.950 294.900 568.050 ;
        RECT 296.550 567.450 297.450 571.950 ;
        RECT 308.250 571.050 310.050 572.850 ;
        RECT 311.100 571.050 312.300 576.300 ;
        RECT 329.700 575.400 333.300 576.300 ;
        RECT 324.000 573.450 328.050 574.050 ;
        RECT 314.100 571.050 315.900 572.850 ;
        RECT 323.550 571.950 328.050 573.450 ;
        RECT 307.950 568.950 310.050 571.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 304.950 567.450 307.050 568.050 ;
        RECT 296.550 566.550 307.050 567.450 ;
        RECT 304.950 565.950 307.050 566.550 ;
        RECT 286.800 555.600 288.000 556.500 ;
        RECT 292.500 555.600 294.000 565.950 ;
        RECT 311.100 555.600 312.300 568.950 ;
        RECT 323.550 568.050 324.450 571.950 ;
        RECT 329.100 571.050 330.900 572.850 ;
        RECT 332.100 571.050 333.300 575.400 ;
        RECT 359.700 575.400 363.300 576.300 ;
        RECT 349.950 573.450 352.050 574.050 ;
        RECT 335.100 571.050 336.900 572.850 ;
        RECT 344.550 572.550 352.050 573.450 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 323.550 566.550 328.050 568.050 ;
        RECT 324.000 565.950 328.050 566.550 ;
        RECT 332.100 561.600 333.300 568.950 ;
        RECT 338.100 567.150 339.900 568.950 ;
        RECT 344.550 568.050 345.450 572.550 ;
        RECT 349.950 571.950 352.050 572.550 ;
        RECT 356.100 571.050 357.900 572.850 ;
        RECT 359.700 571.050 360.900 575.400 ;
        RECT 364.950 573.450 369.000 574.050 ;
        RECT 362.100 571.050 363.900 572.850 ;
        RECT 364.950 571.950 369.450 573.450 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 355.950 568.950 358.050 571.050 ;
        RECT 358.950 568.950 361.050 571.050 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 340.950 566.550 345.450 568.050 ;
        RECT 353.100 567.150 354.900 568.950 ;
        RECT 340.950 565.950 345.000 566.550 ;
        RECT 359.700 561.600 360.900 568.950 ;
        RECT 368.550 568.050 369.450 571.950 ;
        RECT 374.100 571.050 375.900 572.850 ;
        RECT 377.700 571.050 378.900 576.300 ;
        RECT 390.000 573.450 394.050 574.050 ;
        RECT 379.950 571.050 381.750 572.850 ;
        RECT 389.550 571.950 394.050 573.450 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 376.950 568.950 379.050 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 364.950 566.550 369.450 568.050 ;
        RECT 364.950 565.950 369.000 566.550 ;
        RECT 361.950 564.450 364.050 564.750 ;
        RECT 373.950 564.450 376.050 565.050 ;
        RECT 361.950 563.550 376.050 564.450 ;
        RECT 361.950 562.650 364.050 563.550 ;
        RECT 373.950 562.950 376.050 563.550 ;
        RECT 332.100 560.100 334.500 561.600 ;
        RECT 330.000 557.100 331.800 558.900 ;
        RECT 262.200 549.000 264.000 555.600 ;
        RECT 265.200 549.600 267.000 555.600 ;
        RECT 268.200 552.600 270.300 554.700 ;
        RECT 271.200 552.600 273.300 554.700 ;
        RECT 274.200 552.600 276.300 554.700 ;
        RECT 268.200 549.600 270.000 552.600 ;
        RECT 271.200 549.600 273.000 552.600 ;
        RECT 274.200 549.600 276.000 552.600 ;
        RECT 277.200 549.000 279.000 555.600 ;
        RECT 280.200 549.600 282.000 555.600 ;
        RECT 283.200 549.000 285.000 555.600 ;
        RECT 286.200 549.600 288.000 555.600 ;
        RECT 289.200 549.000 291.000 555.600 ;
        RECT 292.500 549.600 294.300 555.600 ;
        RECT 295.500 549.000 297.300 555.600 ;
        RECT 308.100 549.000 309.900 555.600 ;
        RECT 311.100 549.600 312.900 555.600 ;
        RECT 314.100 549.000 315.900 555.600 ;
        RECT 329.700 549.000 331.500 555.600 ;
        RECT 332.700 549.600 334.500 560.100 ;
        RECT 337.800 549.000 339.600 561.600 ;
        RECT 353.400 549.000 355.200 561.600 ;
        RECT 358.500 560.100 360.900 561.600 ;
        RECT 358.500 549.600 360.300 560.100 ;
        RECT 361.200 557.100 363.000 558.900 ;
        RECT 377.700 555.600 378.900 568.950 ;
        RECT 379.950 564.450 382.050 565.050 ;
        RECT 389.550 564.450 390.450 571.950 ;
        RECT 395.100 571.050 396.900 572.850 ;
        RECT 398.700 571.050 399.900 576.300 ;
        RECT 419.700 575.400 423.300 576.300 ;
        RECT 400.950 571.050 402.750 572.850 ;
        RECT 416.100 571.050 417.900 572.850 ;
        RECT 419.700 571.050 420.900 575.400 ;
        RECT 425.700 574.800 426.900 578.400 ;
        RECT 436.800 577.500 438.300 578.400 ;
        RECT 445.800 577.800 447.600 578.400 ;
        RECT 449.700 577.800 450.600 578.400 ;
        RECT 429.900 576.300 438.300 577.500 ;
        RECT 443.400 576.600 450.600 577.800 ;
        RECT 465.300 576.600 471.900 578.400 ;
        RECT 429.900 575.700 431.700 576.300 ;
        RECT 440.400 574.800 442.500 575.700 ;
        RECT 425.700 573.600 442.500 574.800 ;
        RECT 443.400 573.600 444.300 576.600 ;
        RECT 448.800 573.900 450.600 574.800 ;
        RECT 458.100 574.500 459.900 576.300 ;
        RECT 476.100 575.100 477.600 578.400 ;
        RECT 451.800 573.900 453.900 574.050 ;
        RECT 422.100 571.050 423.900 572.850 ;
        RECT 394.950 568.950 397.050 571.050 ;
        RECT 397.950 568.950 400.050 571.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 418.950 568.950 421.050 571.050 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 379.950 563.550 390.450 564.450 ;
        RECT 379.950 562.950 382.050 563.550 ;
        RECT 398.700 555.600 399.900 568.950 ;
        RECT 413.100 567.150 414.900 568.950 ;
        RECT 419.700 561.600 420.900 568.950 ;
        RECT 361.500 549.000 363.300 555.600 ;
        RECT 374.100 549.000 375.900 555.600 ;
        RECT 377.100 549.600 378.900 555.600 ;
        RECT 380.100 549.000 381.900 555.600 ;
        RECT 395.100 549.000 396.900 555.600 ;
        RECT 398.100 549.600 399.900 555.600 ;
        RECT 401.100 549.000 402.900 555.600 ;
        RECT 413.400 549.000 415.200 561.600 ;
        RECT 418.500 560.100 420.900 561.600 ;
        RECT 418.500 549.600 420.300 560.100 ;
        RECT 421.200 557.100 423.000 558.900 ;
        RECT 425.700 557.400 426.900 573.600 ;
        RECT 443.400 571.800 445.200 573.600 ;
        RECT 448.800 573.000 453.900 573.900 ;
        RECT 451.800 571.950 453.900 573.000 ;
        RECT 458.100 573.900 460.200 574.500 ;
        RECT 458.100 572.400 475.200 573.900 ;
        RECT 476.100 573.300 483.900 575.100 ;
        RECT 473.700 570.900 480.300 572.400 ;
        RECT 428.100 569.700 472.500 570.900 ;
        RECT 428.100 568.050 429.900 569.700 ;
        RECT 427.800 565.950 429.900 568.050 ;
        RECT 433.800 567.750 435.900 568.050 ;
        RECT 446.400 567.900 448.200 568.500 ;
        RECT 455.400 567.900 468.900 568.800 ;
        RECT 433.800 565.950 437.700 567.750 ;
        RECT 446.400 566.700 457.500 567.900 ;
        RECT 435.900 565.200 437.700 565.950 ;
        RECT 455.400 565.800 457.500 566.700 ;
        RECT 459.000 565.200 462.900 567.000 ;
        RECT 468.000 566.700 468.900 567.900 ;
        RECT 435.900 564.300 449.400 565.200 ;
        RECT 460.800 564.900 462.900 565.200 ;
        RECT 467.100 564.900 468.900 566.700 ;
        RECT 471.600 568.200 472.500 569.700 ;
        RECT 471.600 566.400 476.700 568.200 ;
        RECT 478.800 568.050 480.300 570.900 ;
        RECT 478.800 565.950 480.900 568.050 ;
        RECT 448.200 563.700 449.400 564.300 ;
        RECT 482.100 563.700 483.900 564.300 ;
        RECT 443.400 562.500 445.500 562.800 ;
        RECT 448.200 562.500 483.900 563.700 ;
        RECT 433.500 561.300 445.500 562.500 ;
        RECT 484.800 561.600 485.700 578.400 ;
        RECT 433.500 560.700 435.300 561.300 ;
        RECT 443.400 560.700 445.500 561.300 ;
        RECT 448.200 560.400 465.900 561.600 ;
        RECT 430.200 559.800 432.000 560.100 ;
        RECT 448.200 559.800 449.400 560.400 ;
        RECT 430.200 558.600 449.400 559.800 ;
        RECT 463.800 559.500 465.900 560.400 ;
        RECT 469.200 560.700 485.700 561.600 ;
        RECT 469.200 559.500 471.300 560.700 ;
        RECT 430.200 558.300 432.000 558.600 ;
        RECT 425.700 556.500 429.300 557.400 ;
        RECT 428.400 555.600 429.300 556.500 ;
        RECT 421.500 549.000 423.300 555.600 ;
        RECT 425.700 549.000 427.500 555.600 ;
        RECT 428.400 554.700 430.500 555.600 ;
        RECT 428.700 549.600 430.500 554.700 ;
        RECT 431.700 549.000 433.500 555.600 ;
        RECT 434.700 549.600 436.500 558.600 ;
        RECT 446.700 555.600 448.800 557.700 ;
        RECT 454.200 557.100 457.500 559.200 ;
        RECT 437.700 549.000 439.500 555.600 ;
        RECT 441.300 552.600 443.400 554.700 ;
        RECT 444.300 552.600 446.400 554.700 ;
        RECT 441.300 549.600 443.100 552.600 ;
        RECT 444.300 549.600 446.100 552.600 ;
        RECT 447.300 549.600 449.100 555.600 ;
        RECT 450.300 549.000 452.100 555.600 ;
        RECT 454.200 549.600 456.000 557.100 ;
        RECT 460.200 555.600 462.900 559.500 ;
        RECT 475.200 558.600 480.900 559.800 ;
        RECT 472.500 557.700 474.300 558.300 ;
        RECT 466.200 556.500 474.300 557.700 ;
        RECT 466.200 555.600 468.300 556.500 ;
        RECT 475.200 555.600 476.400 558.600 ;
        RECT 479.100 558.000 480.900 558.600 ;
        RECT 484.800 557.400 485.700 560.700 ;
        RECT 481.800 556.500 485.700 557.400 ;
        RECT 487.500 581.400 489.300 584.400 ;
        RECT 490.500 581.400 492.300 585.000 ;
        RECT 506.100 581.400 507.900 584.400 ;
        RECT 487.500 568.050 489.000 581.400 ;
        RECT 506.100 577.500 507.300 581.400 ;
        RECT 509.100 578.400 510.900 585.000 ;
        RECT 512.100 578.400 513.900 584.400 ;
        RECT 506.100 576.600 511.800 577.500 ;
        RECT 510.000 575.700 511.800 576.600 ;
        RECT 506.400 568.950 508.500 571.050 ;
        RECT 487.500 565.950 489.900 568.050 ;
        RECT 506.400 567.150 508.200 568.950 ;
        RECT 481.800 555.600 483.000 556.500 ;
        RECT 487.500 555.600 489.000 565.950 ;
        RECT 510.000 564.300 510.900 575.700 ;
        RECT 512.700 571.050 513.900 578.400 ;
        RECT 527.100 579.300 528.900 584.400 ;
        RECT 530.100 580.200 531.900 585.000 ;
        RECT 533.100 579.300 534.900 584.400 ;
        RECT 527.100 577.950 534.900 579.300 ;
        RECT 536.100 578.400 537.900 584.400 ;
        RECT 548.400 578.400 550.200 585.000 ;
        RECT 536.100 576.300 537.300 578.400 ;
        RECT 553.500 577.200 555.300 584.400 ;
        RECT 566.100 579.300 567.900 584.400 ;
        RECT 569.100 580.200 570.900 585.000 ;
        RECT 572.100 579.300 573.900 584.400 ;
        RECT 566.100 577.950 573.900 579.300 ;
        RECT 575.100 578.400 576.900 584.400 ;
        RECT 533.700 575.400 537.300 576.300 ;
        RECT 551.100 576.300 555.300 577.200 ;
        RECT 575.100 576.300 576.300 578.400 ;
        RECT 590.700 577.200 592.500 584.400 ;
        RECT 595.800 578.400 597.600 585.000 ;
        RECT 611.400 578.400 613.200 585.000 ;
        RECT 616.500 577.200 618.300 584.400 ;
        RECT 629.100 581.400 630.900 584.400 ;
        RECT 632.100 581.400 633.900 585.000 ;
        RECT 590.700 576.300 594.900 577.200 ;
        RECT 530.100 571.050 531.900 572.850 ;
        RECT 533.700 571.050 534.900 575.400 ;
        RECT 543.000 573.450 547.050 574.050 ;
        RECT 536.100 571.050 537.900 572.850 ;
        RECT 542.550 571.950 547.050 573.450 ;
        RECT 511.800 568.950 513.900 571.050 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 510.000 563.400 511.800 564.300 ;
        RECT 506.100 562.500 511.800 563.400 ;
        RECT 506.100 555.600 507.300 562.500 ;
        RECT 512.700 561.600 513.900 568.950 ;
        RECT 527.100 567.150 528.900 568.950 ;
        RECT 533.700 561.600 534.900 568.950 ;
        RECT 542.550 568.050 543.450 571.950 ;
        RECT 548.250 571.050 550.050 572.850 ;
        RECT 551.100 571.050 552.300 576.300 ;
        RECT 572.700 575.400 576.300 576.300 ;
        RECT 554.100 571.050 555.900 572.850 ;
        RECT 569.100 571.050 570.900 572.850 ;
        RECT 572.700 571.050 573.900 575.400 ;
        RECT 575.100 571.050 576.900 572.850 ;
        RECT 580.950 571.950 583.050 574.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 538.950 566.550 543.450 568.050 ;
        RECT 538.950 565.950 543.000 566.550 ;
        RECT 457.200 549.000 459.000 555.600 ;
        RECT 460.200 549.600 462.000 555.600 ;
        RECT 463.200 552.600 465.300 554.700 ;
        RECT 466.200 552.600 468.300 554.700 ;
        RECT 469.200 552.600 471.300 554.700 ;
        RECT 463.200 549.600 465.000 552.600 ;
        RECT 466.200 549.600 468.000 552.600 ;
        RECT 469.200 549.600 471.000 552.600 ;
        RECT 472.200 549.000 474.000 555.600 ;
        RECT 475.200 549.600 477.000 555.600 ;
        RECT 478.200 549.000 480.000 555.600 ;
        RECT 481.200 549.600 483.000 555.600 ;
        RECT 484.200 549.000 486.000 555.600 ;
        RECT 487.500 549.600 489.300 555.600 ;
        RECT 490.500 549.000 492.300 555.600 ;
        RECT 506.100 549.600 507.900 555.600 ;
        RECT 509.100 549.000 510.900 559.800 ;
        RECT 512.100 549.600 513.900 561.600 ;
        RECT 527.400 549.000 529.200 561.600 ;
        RECT 532.500 560.100 534.900 561.600 ;
        RECT 532.500 549.600 534.300 560.100 ;
        RECT 535.200 557.100 537.000 558.900 ;
        RECT 551.100 555.600 552.300 568.950 ;
        RECT 566.100 567.150 567.900 568.950 ;
        RECT 572.700 561.600 573.900 568.950 ;
        RECT 581.550 568.050 582.450 571.950 ;
        RECT 590.100 571.050 591.900 572.850 ;
        RECT 593.700 571.050 594.900 576.300 ;
        RECT 614.100 576.300 618.300 577.200 ;
        RECT 595.950 571.050 597.750 572.850 ;
        RECT 611.250 571.050 613.050 572.850 ;
        RECT 614.100 571.050 615.300 576.300 ;
        RECT 617.100 571.050 618.900 572.850 ;
        RECT 629.700 571.050 630.900 581.400 ;
        RECT 644.100 575.400 645.900 585.000 ;
        RECT 650.700 576.000 652.500 584.400 ;
        RECT 668.100 578.400 669.900 584.400 ;
        RECT 668.700 576.300 669.900 578.400 ;
        RECT 671.100 579.300 672.900 584.400 ;
        RECT 674.100 580.200 675.900 585.000 ;
        RECT 677.100 579.300 678.900 584.400 ;
        RECT 671.100 577.950 678.900 579.300 ;
        RECT 689.100 581.400 690.900 584.400 ;
        RECT 689.100 577.500 690.300 581.400 ;
        RECT 692.100 578.400 693.900 585.000 ;
        RECT 695.100 578.400 696.900 584.400 ;
        RECT 710.100 581.400 711.900 585.000 ;
        RECT 713.100 581.400 714.900 584.400 ;
        RECT 689.100 576.600 694.800 577.500 ;
        RECT 650.700 574.800 654.000 576.000 ;
        RECT 668.700 575.400 672.300 576.300 ;
        RECT 644.100 571.050 645.900 572.850 ;
        RECT 650.100 571.050 651.900 572.850 ;
        RECT 653.100 571.050 654.000 574.800 ;
        RECT 668.100 571.050 669.900 572.850 ;
        RECT 671.100 571.050 672.300 575.400 ;
        RECT 693.000 575.700 694.800 576.600 ;
        RECT 674.100 571.050 675.900 572.850 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 595.950 568.950 598.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 689.400 568.950 691.500 571.050 ;
        RECT 577.950 566.550 582.450 568.050 ;
        RECT 577.950 565.950 582.000 566.550 ;
        RECT 535.500 549.000 537.300 555.600 ;
        RECT 548.100 549.000 549.900 555.600 ;
        RECT 551.100 549.600 552.900 555.600 ;
        RECT 554.100 549.000 555.900 555.600 ;
        RECT 566.400 549.000 568.200 561.600 ;
        RECT 571.500 560.100 573.900 561.600 ;
        RECT 571.500 549.600 573.300 560.100 ;
        RECT 574.200 557.100 576.000 558.900 ;
        RECT 593.700 555.600 594.900 568.950 ;
        RECT 595.950 564.450 598.050 565.050 ;
        RECT 601.950 564.450 604.050 565.050 ;
        RECT 595.950 563.550 604.050 564.450 ;
        RECT 595.950 562.950 598.050 563.550 ;
        RECT 601.950 562.950 604.050 563.550 ;
        RECT 614.100 555.600 615.300 568.950 ;
        RECT 629.700 555.600 630.900 568.950 ;
        RECT 632.100 567.150 633.900 568.950 ;
        RECT 647.100 567.150 648.900 568.950 ;
        RECT 643.950 564.450 646.050 564.750 ;
        RECT 649.950 564.450 652.050 565.050 ;
        RECT 643.950 563.550 652.050 564.450 ;
        RECT 643.950 562.650 646.050 563.550 ;
        RECT 649.950 562.950 652.050 563.550 ;
        RECT 653.100 556.800 654.000 568.950 ;
        RECT 671.100 561.600 672.300 568.950 ;
        RECT 677.100 567.150 678.900 568.950 ;
        RECT 689.400 567.150 691.200 568.950 ;
        RECT 673.950 564.450 676.050 565.050 ;
        RECT 679.950 564.450 682.050 565.050 ;
        RECT 673.950 563.550 682.050 564.450 ;
        RECT 673.950 562.950 676.050 563.550 ;
        RECT 679.950 562.950 682.050 563.550 ;
        RECT 693.000 564.300 693.900 575.700 ;
        RECT 695.700 571.050 696.900 578.400 ;
        RECT 713.100 571.050 714.300 581.400 ;
        RECT 728.100 579.300 729.900 584.400 ;
        RECT 731.100 580.200 732.900 585.000 ;
        RECT 734.100 579.300 735.900 584.400 ;
        RECT 728.100 577.950 735.900 579.300 ;
        RECT 737.100 578.400 738.900 584.400 ;
        RECT 737.100 576.300 738.300 578.400 ;
        RECT 734.700 575.400 738.300 576.300 ;
        RECT 739.950 576.450 742.050 580.050 ;
        RECT 750.000 578.400 751.800 585.000 ;
        RECT 754.500 579.600 756.300 584.400 ;
        RECT 757.500 581.400 759.300 585.000 ;
        RECT 754.500 578.400 759.600 579.600 ;
        RECT 754.950 576.450 757.050 577.050 ;
        RECT 739.950 576.000 757.050 576.450 ;
        RECT 740.550 575.550 757.050 576.000 ;
        RECT 731.100 571.050 732.900 572.850 ;
        RECT 734.700 571.050 735.900 575.400 ;
        RECT 754.950 574.950 757.050 575.550 ;
        RECT 744.000 573.450 748.050 574.050 ;
        RECT 737.100 571.050 738.900 572.850 ;
        RECT 743.550 571.950 748.050 573.450 ;
        RECT 694.800 568.950 696.900 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 733.950 568.950 736.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 693.000 563.400 694.800 564.300 ;
        RECT 689.100 562.500 694.800 563.400 ;
        RECT 671.100 560.100 673.500 561.600 ;
        RECT 669.000 557.100 670.800 558.900 ;
        RECT 647.400 555.900 654.000 556.800 ;
        RECT 647.400 555.600 648.900 555.900 ;
        RECT 574.500 549.000 576.300 555.600 ;
        RECT 590.100 549.000 591.900 555.600 ;
        RECT 593.100 549.600 594.900 555.600 ;
        RECT 596.100 549.000 597.900 555.600 ;
        RECT 611.100 549.000 612.900 555.600 ;
        RECT 614.100 549.600 615.900 555.600 ;
        RECT 617.100 549.000 618.900 555.600 ;
        RECT 629.100 549.600 630.900 555.600 ;
        RECT 632.100 549.000 633.900 555.600 ;
        RECT 644.100 549.000 645.900 555.600 ;
        RECT 647.100 549.600 648.900 555.600 ;
        RECT 653.100 555.600 654.000 555.900 ;
        RECT 650.100 549.000 651.900 555.000 ;
        RECT 653.100 549.600 654.900 555.600 ;
        RECT 668.700 549.000 670.500 555.600 ;
        RECT 671.700 549.600 673.500 560.100 ;
        RECT 676.800 549.000 678.600 561.600 ;
        RECT 689.100 555.600 690.300 562.500 ;
        RECT 695.700 561.600 696.900 568.950 ;
        RECT 710.100 567.150 711.900 568.950 ;
        RECT 689.100 549.600 690.900 555.600 ;
        RECT 692.100 549.000 693.900 559.800 ;
        RECT 695.100 549.600 696.900 561.600 ;
        RECT 713.100 555.600 714.300 568.950 ;
        RECT 728.100 567.150 729.900 568.950 ;
        RECT 734.700 561.600 735.900 568.950 ;
        RECT 743.550 568.050 744.450 571.950 ;
        RECT 749.100 571.050 750.900 572.850 ;
        RECT 755.250 571.050 757.050 572.850 ;
        RECT 758.700 571.050 759.600 578.400 ;
        RECT 775.500 576.000 777.300 584.400 ;
        RECT 774.000 574.800 777.300 576.000 ;
        RECT 782.100 575.400 783.900 585.000 ;
        RECT 768.000 573.450 772.050 574.050 ;
        RECT 767.550 571.950 772.050 573.450 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 743.550 566.550 748.050 568.050 ;
        RECT 752.250 567.150 754.050 568.950 ;
        RECT 744.000 565.950 748.050 566.550 ;
        RECT 758.700 561.600 759.600 568.950 ;
        RECT 767.550 568.050 768.450 571.950 ;
        RECT 774.000 571.050 774.900 574.800 ;
        RECT 784.950 573.450 787.050 574.050 ;
        RECT 793.950 573.450 796.050 577.050 ;
        RECT 799.500 576.000 801.300 584.400 ;
        RECT 784.950 573.000 796.050 573.450 ;
        RECT 798.000 574.800 801.300 576.000 ;
        RECT 806.100 575.400 807.900 585.000 ;
        RECT 821.700 577.200 823.500 584.400 ;
        RECT 826.800 578.400 828.600 585.000 ;
        RECT 839.100 579.300 840.900 584.400 ;
        RECT 842.100 580.200 843.900 585.000 ;
        RECT 845.100 579.300 846.900 584.400 ;
        RECT 839.100 577.950 846.900 579.300 ;
        RECT 848.100 578.400 849.900 584.400 ;
        RECT 821.700 576.300 825.900 577.200 ;
        RECT 848.100 576.300 849.300 578.400 ;
        RECT 776.100 571.050 777.900 572.850 ;
        RECT 782.100 571.050 783.900 572.850 ;
        RECT 784.950 572.550 795.450 573.000 ;
        RECT 784.950 571.950 787.050 572.550 ;
        RECT 798.000 571.050 798.900 574.800 ;
        RECT 800.100 571.050 801.900 572.850 ;
        RECT 806.100 571.050 807.900 572.850 ;
        RECT 821.100 571.050 822.900 572.850 ;
        RECT 824.700 571.050 825.900 576.300 ;
        RECT 845.700 575.400 849.300 576.300 ;
        RECT 865.500 576.000 867.300 584.400 ;
        RECT 829.950 573.450 834.000 574.050 ;
        RECT 826.950 571.050 828.750 572.850 ;
        RECT 829.950 571.950 834.450 573.450 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 805.950 568.950 808.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 767.550 566.550 772.050 568.050 ;
        RECT 768.000 565.950 772.050 566.550 ;
        RECT 710.100 549.000 711.900 555.600 ;
        RECT 713.100 549.600 714.900 555.600 ;
        RECT 728.400 549.000 730.200 561.600 ;
        RECT 733.500 560.100 735.900 561.600 ;
        RECT 749.100 560.700 756.900 561.600 ;
        RECT 733.500 549.600 735.300 560.100 ;
        RECT 736.200 557.100 738.000 558.900 ;
        RECT 736.500 549.000 738.300 555.600 ;
        RECT 749.100 549.600 750.900 560.700 ;
        RECT 752.100 549.000 753.900 559.800 ;
        RECT 755.100 549.600 756.900 560.700 ;
        RECT 758.100 549.600 759.900 561.600 ;
        RECT 774.000 556.800 774.900 568.950 ;
        RECT 779.100 567.150 780.900 568.950 ;
        RECT 798.000 556.800 798.900 568.950 ;
        RECT 803.100 567.150 804.900 568.950 ;
        RECT 808.950 564.450 811.050 565.050 ;
        RECT 820.950 564.450 823.050 565.050 ;
        RECT 808.950 563.550 823.050 564.450 ;
        RECT 808.950 562.950 811.050 563.550 ;
        RECT 820.950 562.950 823.050 563.550 ;
        RECT 774.000 555.900 780.600 556.800 ;
        RECT 774.000 555.600 774.900 555.900 ;
        RECT 773.100 549.600 774.900 555.600 ;
        RECT 779.100 555.600 780.600 555.900 ;
        RECT 798.000 555.900 804.600 556.800 ;
        RECT 798.000 555.600 798.900 555.900 ;
        RECT 776.100 549.000 777.900 555.000 ;
        RECT 779.100 549.600 780.900 555.600 ;
        RECT 782.100 549.000 783.900 555.600 ;
        RECT 797.100 549.600 798.900 555.600 ;
        RECT 803.100 555.600 804.600 555.900 ;
        RECT 824.700 555.600 825.900 568.950 ;
        RECT 833.550 568.050 834.450 571.950 ;
        RECT 842.100 571.050 843.900 572.850 ;
        RECT 845.700 571.050 846.900 575.400 ;
        RECT 864.000 574.800 867.300 576.000 ;
        RECT 872.100 575.400 873.900 585.000 ;
        RECT 884.100 581.400 885.900 585.000 ;
        RECT 887.100 581.400 888.900 584.400 ;
        RECT 902.700 581.400 904.500 585.000 ;
        RECT 848.100 571.050 849.900 572.850 ;
        RECT 864.000 571.050 864.900 574.800 ;
        RECT 874.950 573.450 879.000 574.050 ;
        RECT 866.100 571.050 867.900 572.850 ;
        RECT 872.100 571.050 873.900 572.850 ;
        RECT 874.950 571.950 879.450 573.450 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 871.950 568.950 874.050 571.050 ;
        RECT 833.550 566.550 838.050 568.050 ;
        RECT 839.100 567.150 840.900 568.950 ;
        RECT 834.000 565.950 838.050 566.550 ;
        RECT 845.700 561.600 846.900 568.950 ;
        RECT 800.100 549.000 801.900 555.000 ;
        RECT 803.100 549.600 804.900 555.600 ;
        RECT 806.100 549.000 807.900 555.600 ;
        RECT 821.100 549.000 822.900 555.600 ;
        RECT 824.100 549.600 825.900 555.600 ;
        RECT 827.100 549.000 828.900 555.600 ;
        RECT 839.400 549.000 841.200 561.600 ;
        RECT 844.500 560.100 846.900 561.600 ;
        RECT 844.500 549.600 846.300 560.100 ;
        RECT 847.200 557.100 849.000 558.900 ;
        RECT 864.000 556.800 864.900 568.950 ;
        RECT 869.100 567.150 870.900 568.950 ;
        RECT 878.550 568.050 879.450 571.950 ;
        RECT 887.100 571.050 888.300 581.400 ;
        RECT 905.700 579.600 907.500 584.400 ;
        RECT 902.400 578.400 907.500 579.600 ;
        RECT 910.200 578.400 912.000 585.000 ;
        RECT 902.400 571.050 903.300 578.400 ;
        RECT 907.950 576.450 910.050 577.200 ;
        RECT 907.950 575.550 924.450 576.450 ;
        RECT 907.950 575.100 910.050 575.550 ;
        RECT 904.950 571.050 906.750 572.850 ;
        RECT 911.100 571.050 912.900 572.850 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 874.950 566.550 879.450 568.050 ;
        RECT 884.100 567.150 885.900 568.950 ;
        RECT 874.950 565.950 879.000 566.550 ;
        RECT 864.000 555.900 870.600 556.800 ;
        RECT 864.000 555.600 864.900 555.900 ;
        RECT 847.500 549.000 849.300 555.600 ;
        RECT 863.100 549.600 864.900 555.600 ;
        RECT 869.100 555.600 870.600 555.900 ;
        RECT 887.100 555.600 888.300 568.950 ;
        RECT 902.400 561.600 903.300 568.950 ;
        RECT 907.950 567.150 909.750 568.950 ;
        RECT 923.550 567.900 924.450 575.550 ;
        RECT 922.950 565.800 925.050 567.900 ;
        RECT 866.100 549.000 867.900 555.000 ;
        RECT 869.100 549.600 870.900 555.600 ;
        RECT 872.100 549.000 873.900 555.600 ;
        RECT 884.100 549.000 885.900 555.600 ;
        RECT 887.100 549.600 888.900 555.600 ;
        RECT 902.100 549.600 903.900 561.600 ;
        RECT 905.100 560.700 912.900 561.600 ;
        RECT 905.100 549.600 906.900 560.700 ;
        RECT 908.100 549.000 909.900 559.800 ;
        RECT 911.100 549.600 912.900 560.700 ;
        RECT 2.700 539.400 4.500 546.000 ;
        RECT 5.700 540.300 7.500 545.400 ;
        RECT 5.400 539.400 7.500 540.300 ;
        RECT 8.700 539.400 10.500 546.000 ;
        RECT 5.400 538.500 6.300 539.400 ;
        RECT 2.700 537.600 6.300 538.500 ;
        RECT 2.700 521.400 3.900 537.600 ;
        RECT 7.200 536.400 9.000 536.700 ;
        RECT 11.700 536.400 13.500 545.400 ;
        RECT 14.700 539.400 16.500 546.000 ;
        RECT 18.300 542.400 20.100 545.400 ;
        RECT 21.300 542.400 23.100 545.400 ;
        RECT 18.300 540.300 20.400 542.400 ;
        RECT 21.300 540.300 23.400 542.400 ;
        RECT 24.300 539.400 26.100 545.400 ;
        RECT 27.300 539.400 29.100 546.000 ;
        RECT 23.700 537.300 25.800 539.400 ;
        RECT 31.200 537.900 33.000 545.400 ;
        RECT 34.200 539.400 36.000 546.000 ;
        RECT 37.200 539.400 39.000 545.400 ;
        RECT 40.200 542.400 42.000 545.400 ;
        RECT 43.200 542.400 45.000 545.400 ;
        RECT 46.200 542.400 48.000 545.400 ;
        RECT 40.200 540.300 42.300 542.400 ;
        RECT 43.200 540.300 45.300 542.400 ;
        RECT 46.200 540.300 48.300 542.400 ;
        RECT 49.200 539.400 51.000 546.000 ;
        RECT 52.200 539.400 54.000 545.400 ;
        RECT 55.200 539.400 57.000 546.000 ;
        RECT 58.200 539.400 60.000 545.400 ;
        RECT 61.200 539.400 63.000 546.000 ;
        RECT 64.500 539.400 66.300 545.400 ;
        RECT 67.500 539.400 69.300 546.000 ;
        RECT 80.700 539.400 82.500 546.000 ;
        RECT 7.200 535.200 26.400 536.400 ;
        RECT 31.200 535.800 34.500 537.900 ;
        RECT 37.200 535.500 39.900 539.400 ;
        RECT 43.200 538.500 45.300 539.400 ;
        RECT 43.200 537.300 51.300 538.500 ;
        RECT 49.500 536.700 51.300 537.300 ;
        RECT 52.200 536.400 53.400 539.400 ;
        RECT 58.800 538.500 60.000 539.400 ;
        RECT 58.800 537.600 62.700 538.500 ;
        RECT 56.100 536.400 57.900 537.000 ;
        RECT 7.200 534.900 9.000 535.200 ;
        RECT 25.200 534.600 26.400 535.200 ;
        RECT 40.800 534.600 42.900 535.500 ;
        RECT 10.500 533.700 12.300 534.300 ;
        RECT 20.400 533.700 22.500 534.300 ;
        RECT 10.500 532.500 22.500 533.700 ;
        RECT 25.200 533.400 42.900 534.600 ;
        RECT 46.200 534.300 48.300 535.500 ;
        RECT 52.200 535.200 57.900 536.400 ;
        RECT 61.800 534.300 62.700 537.600 ;
        RECT 46.200 533.400 62.700 534.300 ;
        RECT 20.400 532.200 22.500 532.500 ;
        RECT 25.200 531.300 60.900 532.500 ;
        RECT 25.200 530.700 26.400 531.300 ;
        RECT 59.100 530.700 60.900 531.300 ;
        RECT 12.900 529.800 26.400 530.700 ;
        RECT 37.800 529.800 39.900 530.100 ;
        RECT 12.900 529.050 14.700 529.800 ;
        RECT 4.800 526.950 6.900 529.050 ;
        RECT 10.800 527.250 14.700 529.050 ;
        RECT 32.400 528.300 34.500 529.200 ;
        RECT 10.800 526.950 12.900 527.250 ;
        RECT 23.400 527.100 34.500 528.300 ;
        RECT 36.000 528.000 39.900 529.800 ;
        RECT 44.100 528.300 45.900 530.100 ;
        RECT 45.000 527.100 45.900 528.300 ;
        RECT 5.100 525.300 6.900 526.950 ;
        RECT 23.400 526.500 25.200 527.100 ;
        RECT 32.400 526.200 45.900 527.100 ;
        RECT 48.600 526.800 53.700 528.600 ;
        RECT 55.800 526.950 57.900 529.050 ;
        RECT 48.600 525.300 49.500 526.800 ;
        RECT 5.100 524.100 49.500 525.300 ;
        RECT 55.800 524.100 57.300 526.950 ;
        RECT 20.400 521.400 22.200 523.200 ;
        RECT 28.800 522.000 30.900 523.050 ;
        RECT 50.700 522.600 57.300 524.100 ;
        RECT 2.700 520.200 19.500 521.400 ;
        RECT 2.700 516.600 3.900 520.200 ;
        RECT 17.400 519.300 19.500 520.200 ;
        RECT 6.900 518.700 8.700 519.300 ;
        RECT 6.900 517.500 15.300 518.700 ;
        RECT 13.800 516.600 15.300 517.500 ;
        RECT 20.400 518.400 21.300 521.400 ;
        RECT 25.800 521.100 30.900 522.000 ;
        RECT 25.800 520.200 27.600 521.100 ;
        RECT 28.800 520.950 30.900 521.100 ;
        RECT 35.100 521.100 52.200 522.600 ;
        RECT 35.100 520.500 37.200 521.100 ;
        RECT 35.100 518.700 36.900 520.500 ;
        RECT 53.100 519.900 60.900 521.700 ;
        RECT 20.400 517.200 27.600 518.400 ;
        RECT 22.800 516.600 24.600 517.200 ;
        RECT 26.700 516.600 27.600 517.200 ;
        RECT 42.300 516.600 48.900 518.400 ;
        RECT 53.100 516.600 54.600 519.900 ;
        RECT 61.800 516.600 62.700 533.400 ;
        RECT 2.700 510.600 4.500 516.600 ;
        RECT 8.100 510.000 9.900 516.600 ;
        RECT 13.500 510.600 15.300 516.600 ;
        RECT 17.700 513.600 19.800 515.700 ;
        RECT 20.700 513.600 22.800 515.700 ;
        RECT 23.700 513.600 25.800 515.700 ;
        RECT 26.700 515.400 29.400 516.600 ;
        RECT 27.600 514.500 29.400 515.400 ;
        RECT 31.200 514.500 33.900 516.600 ;
        RECT 17.700 510.600 19.500 513.600 ;
        RECT 20.700 510.600 22.500 513.600 ;
        RECT 23.700 510.600 25.500 513.600 ;
        RECT 26.700 510.000 28.500 513.600 ;
        RECT 31.200 510.600 33.000 514.500 ;
        RECT 37.200 513.600 39.300 515.700 ;
        RECT 40.200 513.600 42.300 515.700 ;
        RECT 43.200 513.600 45.300 515.700 ;
        RECT 46.200 513.600 48.300 515.700 ;
        RECT 50.400 515.400 54.600 516.600 ;
        RECT 34.200 510.000 36.000 513.600 ;
        RECT 37.200 510.600 39.000 513.600 ;
        RECT 40.200 510.600 42.000 513.600 ;
        RECT 43.200 510.600 45.000 513.600 ;
        RECT 46.200 510.600 48.000 513.600 ;
        RECT 50.400 510.600 52.200 515.400 ;
        RECT 55.500 510.000 57.300 516.600 ;
        RECT 60.900 510.600 62.700 516.600 ;
        RECT 64.500 529.050 66.000 539.400 ;
        RECT 81.000 536.100 82.800 537.900 ;
        RECT 83.700 534.900 85.500 545.400 ;
        RECT 83.100 533.400 85.500 534.900 ;
        RECT 88.800 533.400 90.600 546.000 ;
        RECT 104.700 539.400 106.500 546.000 ;
        RECT 105.000 536.100 106.800 537.900 ;
        RECT 107.700 534.900 109.500 545.400 ;
        RECT 107.100 533.400 109.500 534.900 ;
        RECT 112.800 533.400 114.600 546.000 ;
        RECT 128.700 539.400 130.500 546.000 ;
        RECT 129.000 536.100 130.800 537.900 ;
        RECT 131.700 534.900 133.500 545.400 ;
        RECT 131.100 533.400 133.500 534.900 ;
        RECT 136.800 533.400 138.600 546.000 ;
        RECT 149.100 533.400 150.900 545.400 ;
        RECT 152.100 534.300 153.900 545.400 ;
        RECT 155.100 535.200 156.900 546.000 ;
        RECT 158.100 534.300 159.900 545.400 ;
        RECT 170.100 539.400 171.900 545.400 ;
        RECT 173.100 539.400 174.900 546.000 ;
        RECT 152.100 533.400 159.900 534.300 ;
        RECT 64.500 526.950 66.900 529.050 ;
        RECT 64.500 513.600 66.000 526.950 ;
        RECT 83.100 526.050 84.300 533.400 ;
        RECT 91.950 528.450 96.000 529.050 ;
        RECT 100.950 528.450 103.050 532.050 ;
        RECT 89.100 526.050 90.900 527.850 ;
        RECT 91.950 526.950 96.450 528.450 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 85.950 523.950 88.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 80.100 522.150 81.900 523.950 ;
        RECT 83.100 519.600 84.300 523.950 ;
        RECT 86.100 522.150 87.900 523.950 ;
        RECT 95.550 520.050 96.450 526.950 ;
        RECT 98.550 528.000 103.050 528.450 ;
        RECT 98.550 527.550 102.450 528.000 ;
        RECT 98.550 523.050 99.450 527.550 ;
        RECT 107.100 526.050 108.300 533.400 ;
        RECT 123.000 528.450 127.050 529.050 ;
        RECT 113.100 526.050 114.900 527.850 ;
        RECT 122.550 526.950 127.050 528.450 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 98.550 521.550 103.050 523.050 ;
        RECT 104.100 522.150 105.900 523.950 ;
        RECT 99.000 520.950 103.050 521.550 ;
        RECT 80.700 518.700 84.300 519.600 ;
        RECT 80.700 516.600 81.900 518.700 ;
        RECT 94.950 517.950 97.050 520.050 ;
        RECT 107.100 519.600 108.300 523.950 ;
        RECT 110.100 522.150 111.900 523.950 ;
        RECT 122.550 523.050 123.450 526.950 ;
        RECT 131.100 526.050 132.300 533.400 ;
        RECT 139.950 528.450 144.000 529.050 ;
        RECT 137.100 526.050 138.900 527.850 ;
        RECT 139.950 526.950 144.450 528.450 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 122.550 521.550 127.050 523.050 ;
        RECT 128.100 522.150 129.900 523.950 ;
        RECT 123.000 520.950 127.050 521.550 ;
        RECT 131.100 519.600 132.300 523.950 ;
        RECT 134.100 522.150 135.900 523.950 ;
        RECT 143.550 523.050 144.450 526.950 ;
        RECT 149.400 526.050 150.300 533.400 ;
        RECT 165.000 528.450 169.050 529.050 ;
        RECT 154.950 526.050 156.750 527.850 ;
        RECT 164.550 526.950 169.050 528.450 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 139.950 521.550 144.450 523.050 ;
        RECT 139.950 520.950 144.000 521.550 ;
        RECT 104.700 518.700 108.300 519.600 ;
        RECT 128.700 518.700 132.300 519.600 ;
        RECT 64.500 510.600 66.300 513.600 ;
        RECT 67.500 510.000 69.300 513.600 ;
        RECT 80.100 510.600 81.900 516.600 ;
        RECT 83.100 515.700 90.900 517.050 ;
        RECT 104.700 516.600 105.900 518.700 ;
        RECT 83.100 510.600 84.900 515.700 ;
        RECT 86.100 510.000 87.900 514.800 ;
        RECT 89.100 510.600 90.900 515.700 ;
        RECT 104.100 510.600 105.900 516.600 ;
        RECT 107.100 515.700 114.900 517.050 ;
        RECT 128.700 516.600 129.900 518.700 ;
        RECT 107.100 510.600 108.900 515.700 ;
        RECT 110.100 510.000 111.900 514.800 ;
        RECT 113.100 510.600 114.900 515.700 ;
        RECT 128.100 510.600 129.900 516.600 ;
        RECT 131.100 515.700 138.900 517.050 ;
        RECT 131.100 510.600 132.900 515.700 ;
        RECT 134.100 510.000 135.900 514.800 ;
        RECT 137.100 510.600 138.900 515.700 ;
        RECT 149.400 516.600 150.300 523.950 ;
        RECT 151.950 522.150 153.750 523.950 ;
        RECT 158.100 522.150 159.900 523.950 ;
        RECT 164.550 523.050 165.450 526.950 ;
        RECT 170.700 526.050 171.900 539.400 ;
        RECT 185.100 533.400 186.900 545.400 ;
        RECT 188.100 534.300 189.900 545.400 ;
        RECT 191.100 535.200 192.900 546.000 ;
        RECT 194.100 534.300 195.900 545.400 ;
        RECT 206.100 539.400 207.900 546.000 ;
        RECT 209.100 539.400 210.900 545.400 ;
        RECT 188.100 533.400 195.900 534.300 ;
        RECT 175.950 528.450 180.000 529.050 ;
        RECT 173.100 526.050 174.900 527.850 ;
        RECT 175.950 526.950 180.450 528.450 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 164.550 521.550 169.050 523.050 ;
        RECT 165.000 520.950 169.050 521.550 ;
        RECT 154.950 519.450 157.050 520.050 ;
        RECT 163.950 519.450 166.050 519.900 ;
        RECT 154.950 518.550 166.050 519.450 ;
        RECT 154.950 517.950 157.050 518.550 ;
        RECT 163.950 517.800 166.050 518.550 ;
        RECT 149.400 515.400 154.500 516.600 ;
        RECT 149.700 510.000 151.500 513.600 ;
        RECT 152.700 510.600 154.500 515.400 ;
        RECT 157.200 510.000 159.000 516.600 ;
        RECT 170.700 513.600 171.900 523.950 ;
        RECT 179.550 523.050 180.450 526.950 ;
        RECT 185.400 526.050 186.300 533.400 ;
        RECT 190.950 526.050 192.750 527.850 ;
        RECT 206.100 526.050 207.900 527.850 ;
        RECT 209.100 526.050 210.300 539.400 ;
        RECT 225.000 534.600 226.800 545.400 ;
        RECT 225.000 533.400 228.600 534.600 ;
        RECT 230.100 533.400 231.900 546.000 ;
        RECT 242.100 533.400 243.900 546.000 ;
        RECT 247.200 534.600 249.000 545.400 ;
        RECT 263.100 539.400 264.900 546.000 ;
        RECT 266.100 539.400 267.900 545.400 ;
        RECT 269.100 539.400 270.900 546.000 ;
        RECT 245.400 533.400 249.000 534.600 ;
        RECT 217.950 529.950 220.050 532.050 ;
        RECT 211.950 528.450 216.000 529.050 ;
        RECT 211.950 526.950 216.450 528.450 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 193.950 523.950 196.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 175.950 521.550 180.450 523.050 ;
        RECT 175.950 520.950 180.000 521.550 ;
        RECT 185.400 516.600 186.300 523.950 ;
        RECT 187.950 522.150 189.750 523.950 ;
        RECT 194.100 522.150 195.900 523.950 ;
        RECT 185.400 515.400 190.500 516.600 ;
        RECT 170.100 510.600 171.900 513.600 ;
        RECT 173.100 510.000 174.900 513.600 ;
        RECT 185.700 510.000 187.500 513.600 ;
        RECT 188.700 510.600 190.500 515.400 ;
        RECT 193.200 510.000 195.000 516.600 ;
        RECT 209.100 513.600 210.300 523.950 ;
        RECT 215.550 523.050 216.450 526.950 ;
        RECT 211.950 521.550 216.450 523.050 ;
        RECT 218.550 523.050 219.450 529.950 ;
        RECT 224.100 526.050 225.900 527.850 ;
        RECT 227.700 526.050 228.600 533.400 ;
        RECT 229.950 526.050 231.750 527.850 ;
        RECT 242.250 526.050 244.050 527.850 ;
        RECT 245.400 526.050 246.300 533.400 ;
        RECT 248.100 526.050 249.900 527.850 ;
        RECT 266.700 526.050 267.900 539.400 ;
        RECT 284.100 533.400 285.900 545.400 ;
        RECT 287.100 535.200 288.900 546.000 ;
        RECT 290.100 539.400 291.900 545.400 ;
        RECT 284.100 526.050 285.300 533.400 ;
        RECT 290.700 532.500 291.900 539.400 ;
        RECT 286.200 531.600 291.900 532.500 ;
        RECT 302.100 533.400 303.900 545.400 ;
        RECT 305.100 535.200 306.900 546.000 ;
        RECT 308.100 539.400 309.900 545.400 ;
        RECT 311.700 539.400 313.500 546.000 ;
        RECT 314.700 540.300 316.500 545.400 ;
        RECT 314.400 539.400 316.500 540.300 ;
        RECT 317.700 539.400 319.500 546.000 ;
        RECT 286.200 530.700 288.000 531.600 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 244.950 523.950 247.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 284.100 523.950 286.200 526.050 ;
        RECT 218.550 521.550 223.050 523.050 ;
        RECT 211.950 520.950 216.000 521.550 ;
        RECT 219.000 520.950 223.050 521.550 ;
        RECT 227.700 513.600 228.600 523.950 ;
        RECT 245.400 513.600 246.300 523.950 ;
        RECT 263.100 522.150 264.900 523.950 ;
        RECT 266.700 518.700 267.900 523.950 ;
        RECT 268.950 522.150 270.750 523.950 ;
        RECT 263.700 517.800 267.900 518.700 ;
        RECT 206.100 510.000 207.900 513.600 ;
        RECT 209.100 510.600 210.900 513.600 ;
        RECT 224.100 510.000 225.900 513.600 ;
        RECT 227.100 510.600 228.900 513.600 ;
        RECT 230.100 510.000 231.900 513.600 ;
        RECT 242.100 510.000 243.900 513.600 ;
        RECT 245.100 510.600 246.900 513.600 ;
        RECT 248.100 510.000 249.900 513.600 ;
        RECT 263.700 510.600 265.500 517.800 ;
        RECT 284.100 516.600 285.300 523.950 ;
        RECT 287.100 519.300 288.000 530.700 ;
        RECT 289.800 526.050 291.600 527.850 ;
        RECT 289.500 523.950 291.600 526.050 ;
        RECT 302.100 526.050 303.300 533.400 ;
        RECT 308.700 532.500 309.900 539.400 ;
        RECT 314.400 538.500 315.300 539.400 ;
        RECT 304.200 531.600 309.900 532.500 ;
        RECT 311.700 537.600 315.300 538.500 ;
        RECT 304.200 530.700 306.000 531.600 ;
        RECT 302.100 523.950 304.200 526.050 ;
        RECT 286.200 518.400 288.000 519.300 ;
        RECT 286.200 517.500 291.900 518.400 ;
        RECT 268.800 510.000 270.600 516.600 ;
        RECT 284.100 510.600 285.900 516.600 ;
        RECT 287.100 510.000 288.900 516.600 ;
        RECT 290.700 513.600 291.900 517.500 ;
        RECT 290.100 510.600 291.900 513.600 ;
        RECT 302.100 516.600 303.300 523.950 ;
        RECT 305.100 519.300 306.000 530.700 ;
        RECT 307.800 526.050 309.600 527.850 ;
        RECT 307.500 523.950 309.600 526.050 ;
        RECT 304.200 518.400 306.000 519.300 ;
        RECT 311.700 521.400 312.900 537.600 ;
        RECT 316.200 536.400 318.000 536.700 ;
        RECT 320.700 536.400 322.500 545.400 ;
        RECT 323.700 539.400 325.500 546.000 ;
        RECT 327.300 542.400 329.100 545.400 ;
        RECT 330.300 542.400 332.100 545.400 ;
        RECT 327.300 540.300 329.400 542.400 ;
        RECT 330.300 540.300 332.400 542.400 ;
        RECT 333.300 539.400 335.100 545.400 ;
        RECT 336.300 539.400 338.100 546.000 ;
        RECT 332.700 537.300 334.800 539.400 ;
        RECT 340.200 537.900 342.000 545.400 ;
        RECT 343.200 539.400 345.000 546.000 ;
        RECT 346.200 539.400 348.000 545.400 ;
        RECT 349.200 542.400 351.000 545.400 ;
        RECT 352.200 542.400 354.000 545.400 ;
        RECT 355.200 542.400 357.000 545.400 ;
        RECT 349.200 540.300 351.300 542.400 ;
        RECT 352.200 540.300 354.300 542.400 ;
        RECT 355.200 540.300 357.300 542.400 ;
        RECT 358.200 539.400 360.000 546.000 ;
        RECT 361.200 539.400 363.000 545.400 ;
        RECT 364.200 539.400 366.000 546.000 ;
        RECT 367.200 539.400 369.000 545.400 ;
        RECT 370.200 539.400 372.000 546.000 ;
        RECT 373.500 539.400 375.300 545.400 ;
        RECT 376.500 539.400 378.300 546.000 ;
        RECT 392.100 539.400 393.900 545.400 ;
        RECT 316.200 535.200 335.400 536.400 ;
        RECT 340.200 535.800 343.500 537.900 ;
        RECT 346.200 535.500 348.900 539.400 ;
        RECT 352.200 538.500 354.300 539.400 ;
        RECT 352.200 537.300 360.300 538.500 ;
        RECT 358.500 536.700 360.300 537.300 ;
        RECT 361.200 536.400 362.400 539.400 ;
        RECT 367.800 538.500 369.000 539.400 ;
        RECT 367.800 537.600 371.700 538.500 ;
        RECT 365.100 536.400 366.900 537.000 ;
        RECT 316.200 534.900 318.000 535.200 ;
        RECT 334.200 534.600 335.400 535.200 ;
        RECT 349.800 534.600 351.900 535.500 ;
        RECT 319.500 533.700 321.300 534.300 ;
        RECT 329.400 533.700 331.500 534.300 ;
        RECT 319.500 532.500 331.500 533.700 ;
        RECT 334.200 533.400 351.900 534.600 ;
        RECT 355.200 534.300 357.300 535.500 ;
        RECT 361.200 535.200 366.900 536.400 ;
        RECT 370.800 534.300 371.700 537.600 ;
        RECT 355.200 533.400 371.700 534.300 ;
        RECT 329.400 532.200 331.500 532.500 ;
        RECT 334.200 531.300 369.900 532.500 ;
        RECT 334.200 530.700 335.400 531.300 ;
        RECT 368.100 530.700 369.900 531.300 ;
        RECT 321.900 529.800 335.400 530.700 ;
        RECT 346.800 529.800 348.900 530.100 ;
        RECT 321.900 529.050 323.700 529.800 ;
        RECT 313.800 526.950 315.900 529.050 ;
        RECT 319.800 527.250 323.700 529.050 ;
        RECT 341.400 528.300 343.500 529.200 ;
        RECT 319.800 526.950 321.900 527.250 ;
        RECT 332.400 527.100 343.500 528.300 ;
        RECT 345.000 528.000 348.900 529.800 ;
        RECT 353.100 528.300 354.900 530.100 ;
        RECT 354.000 527.100 354.900 528.300 ;
        RECT 314.100 525.300 315.900 526.950 ;
        RECT 332.400 526.500 334.200 527.100 ;
        RECT 341.400 526.200 354.900 527.100 ;
        RECT 357.600 526.800 362.700 528.600 ;
        RECT 364.800 526.950 366.900 529.050 ;
        RECT 357.600 525.300 358.500 526.800 ;
        RECT 314.100 524.100 358.500 525.300 ;
        RECT 364.800 524.100 366.300 526.950 ;
        RECT 329.400 521.400 331.200 523.200 ;
        RECT 337.800 522.000 339.900 523.050 ;
        RECT 359.700 522.600 366.300 524.100 ;
        RECT 311.700 520.200 328.500 521.400 ;
        RECT 304.200 517.500 309.900 518.400 ;
        RECT 302.100 510.600 303.900 516.600 ;
        RECT 305.100 510.000 306.900 516.600 ;
        RECT 308.700 513.600 309.900 517.500 ;
        RECT 308.100 510.600 309.900 513.600 ;
        RECT 311.700 516.600 312.900 520.200 ;
        RECT 326.400 519.300 328.500 520.200 ;
        RECT 315.900 518.700 317.700 519.300 ;
        RECT 315.900 517.500 324.300 518.700 ;
        RECT 322.800 516.600 324.300 517.500 ;
        RECT 329.400 518.400 330.300 521.400 ;
        RECT 334.800 521.100 339.900 522.000 ;
        RECT 334.800 520.200 336.600 521.100 ;
        RECT 337.800 520.950 339.900 521.100 ;
        RECT 344.100 521.100 361.200 522.600 ;
        RECT 344.100 520.500 346.200 521.100 ;
        RECT 344.100 518.700 345.900 520.500 ;
        RECT 362.100 519.900 369.900 521.700 ;
        RECT 329.400 517.200 336.600 518.400 ;
        RECT 331.800 516.600 333.600 517.200 ;
        RECT 335.700 516.600 336.600 517.200 ;
        RECT 351.300 516.600 357.900 518.400 ;
        RECT 362.100 516.600 363.600 519.900 ;
        RECT 370.800 516.600 371.700 533.400 ;
        RECT 311.700 510.600 313.500 516.600 ;
        RECT 317.100 510.000 318.900 516.600 ;
        RECT 322.500 510.600 324.300 516.600 ;
        RECT 326.700 513.600 328.800 515.700 ;
        RECT 329.700 513.600 331.800 515.700 ;
        RECT 332.700 513.600 334.800 515.700 ;
        RECT 335.700 515.400 338.400 516.600 ;
        RECT 336.600 514.500 338.400 515.400 ;
        RECT 340.200 514.500 342.900 516.600 ;
        RECT 326.700 510.600 328.500 513.600 ;
        RECT 329.700 510.600 331.500 513.600 ;
        RECT 332.700 510.600 334.500 513.600 ;
        RECT 335.700 510.000 337.500 513.600 ;
        RECT 340.200 510.600 342.000 514.500 ;
        RECT 346.200 513.600 348.300 515.700 ;
        RECT 349.200 513.600 351.300 515.700 ;
        RECT 352.200 513.600 354.300 515.700 ;
        RECT 355.200 513.600 357.300 515.700 ;
        RECT 359.400 515.400 363.600 516.600 ;
        RECT 343.200 510.000 345.000 513.600 ;
        RECT 346.200 510.600 348.000 513.600 ;
        RECT 349.200 510.600 351.000 513.600 ;
        RECT 352.200 510.600 354.000 513.600 ;
        RECT 355.200 510.600 357.000 513.600 ;
        RECT 359.400 510.600 361.200 515.400 ;
        RECT 364.500 510.000 366.300 516.600 ;
        RECT 369.900 510.600 371.700 516.600 ;
        RECT 373.500 529.050 375.000 539.400 ;
        RECT 392.100 532.500 393.300 539.400 ;
        RECT 395.100 535.200 396.900 546.000 ;
        RECT 398.100 533.400 399.900 545.400 ;
        RECT 392.100 531.600 397.800 532.500 ;
        RECT 396.000 530.700 397.800 531.600 ;
        RECT 373.500 526.950 375.900 529.050 ;
        RECT 373.500 513.600 375.000 526.950 ;
        RECT 392.400 526.050 394.200 527.850 ;
        RECT 392.400 523.950 394.500 526.050 ;
        RECT 396.000 519.300 396.900 530.700 ;
        RECT 398.700 526.050 399.900 533.400 ;
        RECT 413.100 539.400 414.900 545.400 ;
        RECT 413.100 532.500 414.300 539.400 ;
        RECT 416.100 535.200 417.900 546.000 ;
        RECT 419.100 533.400 420.900 545.400 ;
        RECT 434.400 533.400 436.200 546.000 ;
        RECT 439.500 534.900 441.300 545.400 ;
        RECT 442.500 539.400 444.300 546.000 ;
        RECT 442.200 536.100 444.000 537.900 ;
        RECT 439.500 533.400 441.900 534.900 ;
        RECT 413.100 531.600 418.800 532.500 ;
        RECT 417.000 530.700 418.800 531.600 ;
        RECT 397.800 523.950 399.900 526.050 ;
        RECT 413.400 526.050 415.200 527.850 ;
        RECT 413.400 523.950 415.500 526.050 ;
        RECT 396.000 518.400 397.800 519.300 ;
        RECT 392.100 517.500 397.800 518.400 ;
        RECT 392.100 513.600 393.300 517.500 ;
        RECT 398.700 516.600 399.900 523.950 ;
        RECT 417.000 519.300 417.900 530.700 ;
        RECT 419.700 526.050 420.900 533.400 ;
        RECT 434.100 526.050 435.900 527.850 ;
        RECT 440.700 526.050 441.900 533.400 ;
        RECT 458.100 533.400 459.900 545.400 ;
        RECT 461.100 535.200 462.900 546.000 ;
        RECT 464.100 539.400 465.900 545.400 ;
        RECT 458.100 526.050 459.300 533.400 ;
        RECT 464.700 532.500 465.900 539.400 ;
        RECT 460.200 531.600 465.900 532.500 ;
        RECT 476.100 539.400 477.900 545.400 ;
        RECT 476.100 532.500 477.300 539.400 ;
        RECT 479.100 535.200 480.900 546.000 ;
        RECT 482.100 533.400 483.900 545.400 ;
        RECT 494.100 539.400 495.900 546.000 ;
        RECT 497.100 539.400 498.900 545.400 ;
        RECT 500.100 539.400 501.900 546.000 ;
        RECT 503.700 539.400 505.500 546.000 ;
        RECT 506.700 540.300 508.500 545.400 ;
        RECT 506.400 539.400 508.500 540.300 ;
        RECT 509.700 539.400 511.500 546.000 ;
        RECT 484.950 537.450 487.050 538.050 ;
        RECT 493.950 537.450 496.050 538.050 ;
        RECT 484.950 536.550 496.050 537.450 ;
        RECT 484.950 535.950 487.050 536.550 ;
        RECT 493.950 535.950 496.050 536.550 ;
        RECT 476.100 531.600 481.800 532.500 ;
        RECT 460.200 530.700 462.000 531.600 ;
        RECT 418.800 523.950 420.900 526.050 ;
        RECT 433.950 523.950 436.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 458.100 523.950 460.200 526.050 ;
        RECT 417.000 518.400 418.800 519.300 ;
        RECT 373.500 510.600 375.300 513.600 ;
        RECT 376.500 510.000 378.300 513.600 ;
        RECT 392.100 510.600 393.900 513.600 ;
        RECT 395.100 510.000 396.900 516.600 ;
        RECT 398.100 510.600 399.900 516.600 ;
        RECT 413.100 517.500 418.800 518.400 ;
        RECT 413.100 513.600 414.300 517.500 ;
        RECT 419.700 516.600 420.900 523.950 ;
        RECT 437.100 522.150 438.900 523.950 ;
        RECT 440.700 519.600 441.900 523.950 ;
        RECT 443.100 522.150 444.900 523.950 ;
        RECT 440.700 518.700 444.300 519.600 ;
        RECT 413.100 510.600 414.900 513.600 ;
        RECT 416.100 510.000 417.900 516.600 ;
        RECT 419.100 510.600 420.900 516.600 ;
        RECT 434.100 515.700 441.900 517.050 ;
        RECT 434.100 510.600 435.900 515.700 ;
        RECT 437.100 510.000 438.900 514.800 ;
        RECT 440.100 510.600 441.900 515.700 ;
        RECT 443.100 516.600 444.300 518.700 ;
        RECT 458.100 516.600 459.300 523.950 ;
        RECT 461.100 519.300 462.000 530.700 ;
        RECT 480.000 530.700 481.800 531.600 ;
        RECT 463.800 526.050 465.600 527.850 ;
        RECT 463.500 523.950 465.600 526.050 ;
        RECT 476.400 526.050 478.200 527.850 ;
        RECT 476.400 523.950 478.500 526.050 ;
        RECT 460.200 518.400 462.000 519.300 ;
        RECT 480.000 519.300 480.900 530.700 ;
        RECT 482.700 526.050 483.900 533.400 ;
        RECT 497.100 526.050 498.300 539.400 ;
        RECT 506.400 538.500 507.300 539.400 ;
        RECT 503.700 537.600 507.300 538.500 ;
        RECT 481.800 523.950 483.900 526.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 480.000 518.400 481.800 519.300 ;
        RECT 460.200 517.500 465.900 518.400 ;
        RECT 443.100 510.600 444.900 516.600 ;
        RECT 458.100 510.600 459.900 516.600 ;
        RECT 461.100 510.000 462.900 516.600 ;
        RECT 464.700 513.600 465.900 517.500 ;
        RECT 464.100 510.600 465.900 513.600 ;
        RECT 476.100 517.500 481.800 518.400 ;
        RECT 476.100 513.600 477.300 517.500 ;
        RECT 482.700 516.600 483.900 523.950 ;
        RECT 494.250 522.150 496.050 523.950 ;
        RECT 497.100 518.700 498.300 523.950 ;
        RECT 500.100 522.150 501.900 523.950 ;
        RECT 503.700 521.400 504.900 537.600 ;
        RECT 508.200 536.400 510.000 536.700 ;
        RECT 512.700 536.400 514.500 545.400 ;
        RECT 515.700 539.400 517.500 546.000 ;
        RECT 519.300 542.400 521.100 545.400 ;
        RECT 522.300 542.400 524.100 545.400 ;
        RECT 519.300 540.300 521.400 542.400 ;
        RECT 522.300 540.300 524.400 542.400 ;
        RECT 525.300 539.400 527.100 545.400 ;
        RECT 528.300 539.400 530.100 546.000 ;
        RECT 524.700 537.300 526.800 539.400 ;
        RECT 532.200 537.900 534.000 545.400 ;
        RECT 535.200 539.400 537.000 546.000 ;
        RECT 538.200 539.400 540.000 545.400 ;
        RECT 541.200 542.400 543.000 545.400 ;
        RECT 544.200 542.400 546.000 545.400 ;
        RECT 547.200 542.400 549.000 545.400 ;
        RECT 541.200 540.300 543.300 542.400 ;
        RECT 544.200 540.300 546.300 542.400 ;
        RECT 547.200 540.300 549.300 542.400 ;
        RECT 550.200 539.400 552.000 546.000 ;
        RECT 553.200 539.400 555.000 545.400 ;
        RECT 556.200 539.400 558.000 546.000 ;
        RECT 559.200 539.400 561.000 545.400 ;
        RECT 562.200 539.400 564.000 546.000 ;
        RECT 565.500 539.400 567.300 545.400 ;
        RECT 568.500 539.400 570.300 546.000 ;
        RECT 581.100 539.400 582.900 545.400 ;
        RECT 508.200 535.200 527.400 536.400 ;
        RECT 532.200 535.800 535.500 537.900 ;
        RECT 538.200 535.500 540.900 539.400 ;
        RECT 544.200 538.500 546.300 539.400 ;
        RECT 544.200 537.300 552.300 538.500 ;
        RECT 550.500 536.700 552.300 537.300 ;
        RECT 553.200 536.400 554.400 539.400 ;
        RECT 559.800 538.500 561.000 539.400 ;
        RECT 559.800 537.600 563.700 538.500 ;
        RECT 557.100 536.400 558.900 537.000 ;
        RECT 508.200 534.900 510.000 535.200 ;
        RECT 526.200 534.600 527.400 535.200 ;
        RECT 541.800 534.600 543.900 535.500 ;
        RECT 511.500 533.700 513.300 534.300 ;
        RECT 521.400 533.700 523.500 534.300 ;
        RECT 511.500 532.500 523.500 533.700 ;
        RECT 526.200 533.400 543.900 534.600 ;
        RECT 547.200 534.300 549.300 535.500 ;
        RECT 553.200 535.200 558.900 536.400 ;
        RECT 562.800 534.300 563.700 537.600 ;
        RECT 547.200 533.400 563.700 534.300 ;
        RECT 521.400 532.200 523.500 532.500 ;
        RECT 526.200 531.300 561.900 532.500 ;
        RECT 526.200 530.700 527.400 531.300 ;
        RECT 560.100 530.700 561.900 531.300 ;
        RECT 513.900 529.800 527.400 530.700 ;
        RECT 538.800 529.800 540.900 530.100 ;
        RECT 513.900 529.050 515.700 529.800 ;
        RECT 505.800 526.950 507.900 529.050 ;
        RECT 511.800 527.250 515.700 529.050 ;
        RECT 533.400 528.300 535.500 529.200 ;
        RECT 511.800 526.950 513.900 527.250 ;
        RECT 524.400 527.100 535.500 528.300 ;
        RECT 537.000 528.000 540.900 529.800 ;
        RECT 545.100 528.300 546.900 530.100 ;
        RECT 546.000 527.100 546.900 528.300 ;
        RECT 506.100 525.300 507.900 526.950 ;
        RECT 524.400 526.500 526.200 527.100 ;
        RECT 533.400 526.200 546.900 527.100 ;
        RECT 549.600 526.800 554.700 528.600 ;
        RECT 556.800 526.950 558.900 529.050 ;
        RECT 549.600 525.300 550.500 526.800 ;
        RECT 506.100 524.100 550.500 525.300 ;
        RECT 556.800 524.100 558.300 526.950 ;
        RECT 521.400 521.400 523.200 523.200 ;
        RECT 529.800 522.000 531.900 523.050 ;
        RECT 551.700 522.600 558.300 524.100 ;
        RECT 503.700 520.200 520.500 521.400 ;
        RECT 497.100 517.800 501.300 518.700 ;
        RECT 476.100 510.600 477.900 513.600 ;
        RECT 479.100 510.000 480.900 516.600 ;
        RECT 482.100 510.600 483.900 516.600 ;
        RECT 494.400 510.000 496.200 516.600 ;
        RECT 499.500 510.600 501.300 517.800 ;
        RECT 503.700 516.600 504.900 520.200 ;
        RECT 518.400 519.300 520.500 520.200 ;
        RECT 507.900 518.700 509.700 519.300 ;
        RECT 507.900 517.500 516.300 518.700 ;
        RECT 514.800 516.600 516.300 517.500 ;
        RECT 521.400 518.400 522.300 521.400 ;
        RECT 526.800 521.100 531.900 522.000 ;
        RECT 526.800 520.200 528.600 521.100 ;
        RECT 529.800 520.950 531.900 521.100 ;
        RECT 536.100 521.100 553.200 522.600 ;
        RECT 536.100 520.500 538.200 521.100 ;
        RECT 536.100 518.700 537.900 520.500 ;
        RECT 554.100 519.900 561.900 521.700 ;
        RECT 521.400 517.200 528.600 518.400 ;
        RECT 523.800 516.600 525.600 517.200 ;
        RECT 527.700 516.600 528.600 517.200 ;
        RECT 543.300 516.600 549.900 518.400 ;
        RECT 554.100 516.600 555.600 519.900 ;
        RECT 562.800 516.600 563.700 533.400 ;
        RECT 503.700 510.600 505.500 516.600 ;
        RECT 509.100 510.000 510.900 516.600 ;
        RECT 514.500 510.600 516.300 516.600 ;
        RECT 518.700 513.600 520.800 515.700 ;
        RECT 521.700 513.600 523.800 515.700 ;
        RECT 524.700 513.600 526.800 515.700 ;
        RECT 527.700 515.400 530.400 516.600 ;
        RECT 528.600 514.500 530.400 515.400 ;
        RECT 532.200 514.500 534.900 516.600 ;
        RECT 518.700 510.600 520.500 513.600 ;
        RECT 521.700 510.600 523.500 513.600 ;
        RECT 524.700 510.600 526.500 513.600 ;
        RECT 527.700 510.000 529.500 513.600 ;
        RECT 532.200 510.600 534.000 514.500 ;
        RECT 538.200 513.600 540.300 515.700 ;
        RECT 541.200 513.600 543.300 515.700 ;
        RECT 544.200 513.600 546.300 515.700 ;
        RECT 547.200 513.600 549.300 515.700 ;
        RECT 551.400 515.400 555.600 516.600 ;
        RECT 535.200 510.000 537.000 513.600 ;
        RECT 538.200 510.600 540.000 513.600 ;
        RECT 541.200 510.600 543.000 513.600 ;
        RECT 544.200 510.600 546.000 513.600 ;
        RECT 547.200 510.600 549.000 513.600 ;
        RECT 551.400 510.600 553.200 515.400 ;
        RECT 556.500 510.000 558.300 516.600 ;
        RECT 561.900 510.600 563.700 516.600 ;
        RECT 565.500 529.050 567.000 539.400 ;
        RECT 581.100 532.500 582.300 539.400 ;
        RECT 584.100 535.200 585.900 546.000 ;
        RECT 587.100 533.400 588.900 545.400 ;
        RECT 581.100 531.600 586.800 532.500 ;
        RECT 585.000 530.700 586.800 531.600 ;
        RECT 565.500 526.950 567.900 529.050 ;
        RECT 565.500 513.600 567.000 526.950 ;
        RECT 581.400 526.050 583.200 527.850 ;
        RECT 581.400 523.950 583.500 526.050 ;
        RECT 585.000 519.300 585.900 530.700 ;
        RECT 587.700 526.050 588.900 533.400 ;
        RECT 586.800 523.950 588.900 526.050 ;
        RECT 585.000 518.400 586.800 519.300 ;
        RECT 581.100 517.500 586.800 518.400 ;
        RECT 581.100 513.600 582.300 517.500 ;
        RECT 587.700 516.600 588.900 523.950 ;
        RECT 565.500 510.600 567.300 513.600 ;
        RECT 568.500 510.000 570.300 513.600 ;
        RECT 581.100 510.600 582.900 513.600 ;
        RECT 584.100 510.000 585.900 516.600 ;
        RECT 587.100 510.600 588.900 516.600 ;
        RECT 602.100 533.400 603.900 545.400 ;
        RECT 605.100 535.200 606.900 546.000 ;
        RECT 608.100 539.400 609.900 545.400 ;
        RECT 620.100 539.400 621.900 546.000 ;
        RECT 623.100 539.400 624.900 545.400 ;
        RECT 602.100 526.050 603.300 533.400 ;
        RECT 608.700 532.500 609.900 539.400 ;
        RECT 604.200 531.600 609.900 532.500 ;
        RECT 604.200 530.700 606.000 531.600 ;
        RECT 602.100 523.950 604.200 526.050 ;
        RECT 602.100 516.600 603.300 523.950 ;
        RECT 605.100 519.300 606.000 530.700 ;
        RECT 607.800 526.050 609.600 527.850 ;
        RECT 607.500 523.950 609.600 526.050 ;
        RECT 620.100 523.950 622.200 526.050 ;
        RECT 620.250 522.150 622.050 523.950 ;
        RECT 623.100 519.300 624.000 539.400 ;
        RECT 626.100 534.000 627.900 546.000 ;
        RECT 629.100 533.400 630.900 545.400 ;
        RECT 641.100 539.400 642.900 546.000 ;
        RECT 644.100 539.400 645.900 545.400 ;
        RECT 647.100 539.400 648.900 546.000 ;
        RECT 625.200 526.050 627.000 527.850 ;
        RECT 629.400 526.050 630.300 533.400 ;
        RECT 644.700 526.050 645.900 539.400 ;
        RECT 662.400 533.400 664.200 546.000 ;
        RECT 667.500 534.900 669.300 545.400 ;
        RECT 670.500 539.400 672.300 546.000 ;
        RECT 683.100 539.400 684.900 545.400 ;
        RECT 686.100 540.000 687.900 546.000 ;
        RECT 684.000 539.100 684.900 539.400 ;
        RECT 689.100 539.400 690.900 545.400 ;
        RECT 692.100 539.400 693.900 546.000 ;
        RECT 707.700 539.400 709.500 546.000 ;
        RECT 689.100 539.100 690.600 539.400 ;
        RECT 684.000 538.200 690.600 539.100 ;
        RECT 670.200 536.100 672.000 537.900 ;
        RECT 667.500 533.400 669.900 534.900 ;
        RECT 662.100 526.050 663.900 527.850 ;
        RECT 668.700 526.050 669.900 533.400 ;
        RECT 673.950 528.450 678.000 529.050 ;
        RECT 673.950 526.950 678.450 528.450 ;
        RECT 625.500 523.950 627.600 526.050 ;
        RECT 628.800 523.950 630.900 526.050 ;
        RECT 640.950 523.950 643.050 526.050 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 604.200 518.400 606.000 519.300 ;
        RECT 620.100 518.400 628.500 519.300 ;
        RECT 604.200 517.500 609.900 518.400 ;
        RECT 602.100 510.600 603.900 516.600 ;
        RECT 605.100 510.000 606.900 516.600 ;
        RECT 608.700 513.600 609.900 517.500 ;
        RECT 608.100 510.600 609.900 513.600 ;
        RECT 620.100 510.600 621.900 518.400 ;
        RECT 626.700 517.500 628.500 518.400 ;
        RECT 629.400 516.600 630.300 523.950 ;
        RECT 641.100 522.150 642.900 523.950 ;
        RECT 644.700 518.700 645.900 523.950 ;
        RECT 646.950 522.150 648.750 523.950 ;
        RECT 665.100 522.150 666.900 523.950 ;
        RECT 668.700 519.600 669.900 523.950 ;
        RECT 671.100 522.150 672.900 523.950 ;
        RECT 677.550 523.050 678.450 526.950 ;
        RECT 684.000 526.050 684.900 538.200 ;
        RECT 708.000 536.100 709.800 537.900 ;
        RECT 685.950 534.450 688.050 535.050 ;
        RECT 703.950 534.450 706.050 535.050 ;
        RECT 710.700 534.900 712.500 545.400 ;
        RECT 685.950 533.550 706.050 534.450 ;
        RECT 685.950 532.950 688.050 533.550 ;
        RECT 703.950 532.950 706.050 533.550 ;
        RECT 710.100 533.400 712.500 534.900 ;
        RECT 715.800 533.400 717.600 546.000 ;
        RECT 731.100 533.400 732.900 545.400 ;
        RECT 734.100 534.300 735.900 545.400 ;
        RECT 737.100 535.200 738.900 546.000 ;
        RECT 740.100 534.300 741.900 545.400 ;
        RECT 755.100 544.500 762.900 545.400 ;
        RECT 755.100 535.200 756.900 544.500 ;
        RECT 758.100 535.800 759.900 543.600 ;
        RECT 734.100 533.400 741.900 534.300 ;
        RECT 685.950 531.450 688.050 531.900 ;
        RECT 685.950 530.550 696.450 531.450 ;
        RECT 685.950 529.800 688.050 530.550 ;
        RECT 695.550 528.450 696.450 530.550 ;
        RECT 689.100 526.050 690.900 527.850 ;
        RECT 695.550 527.550 699.450 528.450 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 673.950 521.550 678.450 523.050 ;
        RECT 673.950 520.950 678.000 521.550 ;
        RECT 684.000 520.200 684.900 523.950 ;
        RECT 686.100 522.150 687.900 523.950 ;
        RECT 692.100 522.150 693.900 523.950 ;
        RECT 698.550 523.050 699.450 527.550 ;
        RECT 710.100 526.050 711.300 533.400 ;
        RECT 715.950 531.450 718.050 532.050 ;
        RECT 715.950 530.550 726.450 531.450 ;
        RECT 715.950 529.950 718.050 530.550 ;
        RECT 718.950 528.450 723.000 529.050 ;
        RECT 716.100 526.050 717.900 527.850 ;
        RECT 718.950 526.950 723.450 528.450 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 694.950 521.550 699.450 523.050 ;
        RECT 707.100 522.150 708.900 523.950 ;
        RECT 694.950 520.950 699.000 521.550 ;
        RECT 668.700 518.700 672.300 519.600 ;
        RECT 684.000 519.000 687.300 520.200 ;
        RECT 710.100 519.600 711.300 523.950 ;
        RECT 713.100 522.150 714.900 523.950 ;
        RECT 722.550 522.900 723.450 526.950 ;
        RECT 721.950 520.800 724.050 522.900 ;
        RECT 624.600 510.000 626.400 516.600 ;
        RECT 627.600 514.800 630.300 516.600 ;
        RECT 641.700 517.800 645.900 518.700 ;
        RECT 627.600 510.600 629.400 514.800 ;
        RECT 641.700 510.600 643.500 517.800 ;
        RECT 646.800 510.000 648.600 516.600 ;
        RECT 662.100 515.700 669.900 517.050 ;
        RECT 662.100 510.600 663.900 515.700 ;
        RECT 665.100 510.000 666.900 514.800 ;
        RECT 668.100 510.600 669.900 515.700 ;
        RECT 671.100 516.600 672.300 518.700 ;
        RECT 671.100 510.600 672.900 516.600 ;
        RECT 685.500 510.600 687.300 519.000 ;
        RECT 692.100 510.000 693.900 519.600 ;
        RECT 707.700 518.700 711.300 519.600 ;
        RECT 718.950 519.450 721.050 519.900 ;
        RECT 725.550 519.450 726.450 530.550 ;
        RECT 731.400 526.050 732.300 533.400 ;
        RECT 736.950 526.050 738.750 527.850 ;
        RECT 758.700 526.050 759.900 535.800 ;
        RECT 761.100 535.800 762.900 544.500 ;
        RECT 764.100 544.500 771.900 545.400 ;
        RECT 764.100 536.700 765.900 544.500 ;
        RECT 767.100 535.800 768.900 543.600 ;
        RECT 761.100 534.900 768.900 535.800 ;
        RECT 770.100 535.500 771.900 544.500 ;
        RECT 773.100 536.400 774.900 546.000 ;
        RECT 776.100 535.500 777.900 545.400 ;
        RECT 788.700 539.400 790.500 546.000 ;
        RECT 789.000 536.100 790.800 537.900 ;
        RECT 770.100 534.600 777.900 535.500 ;
        RECT 791.700 534.900 793.500 545.400 ;
        RECT 791.100 533.400 793.500 534.900 ;
        RECT 796.800 533.400 798.600 546.000 ;
        RECT 809.100 533.400 810.900 545.400 ;
        RECT 812.100 534.300 813.900 545.400 ;
        RECT 815.100 535.200 816.900 546.000 ;
        RECT 818.100 534.300 819.900 545.400 ;
        RECT 830.700 539.400 832.500 546.000 ;
        RECT 831.000 536.100 832.800 537.900 ;
        RECT 833.700 534.900 835.500 545.400 ;
        RECT 812.100 533.400 819.900 534.300 ;
        RECT 833.100 533.400 835.500 534.900 ;
        RECT 838.800 533.400 840.600 546.000 ;
        RECT 854.100 539.400 855.900 545.400 ;
        RECT 857.100 540.000 858.900 546.000 ;
        RECT 855.000 539.100 855.900 539.400 ;
        RECT 860.100 539.400 861.900 545.400 ;
        RECT 863.100 539.400 864.900 546.000 ;
        RECT 860.100 539.100 861.600 539.400 ;
        RECT 855.000 538.200 861.600 539.100 ;
        RECT 784.950 528.450 787.050 529.050 ;
        RECT 763.950 526.050 765.750 527.850 ;
        RECT 773.100 526.050 774.900 527.850 ;
        RECT 779.550 527.550 787.050 528.450 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 733.950 523.950 736.050 526.050 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 758.400 523.950 760.500 526.050 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 773.100 523.950 775.200 526.050 ;
        RECT 707.700 516.600 708.900 518.700 ;
        RECT 718.950 518.550 726.450 519.450 ;
        RECT 718.950 517.800 721.050 518.550 ;
        RECT 707.100 510.600 708.900 516.600 ;
        RECT 710.100 515.700 717.900 517.050 ;
        RECT 710.100 510.600 711.900 515.700 ;
        RECT 713.100 510.000 714.900 514.800 ;
        RECT 716.100 510.600 717.900 515.700 ;
        RECT 731.400 516.600 732.300 523.950 ;
        RECT 733.950 522.150 735.750 523.950 ;
        RECT 740.100 522.150 741.900 523.950 ;
        RECT 736.950 519.450 739.050 520.050 ;
        RECT 754.950 519.450 757.050 520.050 ;
        RECT 736.950 518.550 757.050 519.450 ;
        RECT 736.950 517.950 739.050 518.550 ;
        RECT 754.950 517.950 757.050 518.550 ;
        RECT 731.400 515.400 736.500 516.600 ;
        RECT 731.700 510.000 733.500 513.600 ;
        RECT 734.700 510.600 736.500 515.400 ;
        RECT 739.200 510.000 741.000 516.600 ;
        RECT 758.700 515.400 759.900 523.950 ;
        RECT 767.250 522.150 769.050 523.950 ;
        RECT 760.950 519.450 763.050 520.050 ;
        RECT 779.550 519.450 780.450 527.550 ;
        RECT 784.950 526.950 787.050 527.550 ;
        RECT 791.100 526.050 792.300 533.400 ;
        RECT 797.100 526.050 798.900 527.850 ;
        RECT 809.400 526.050 810.300 533.400 ;
        RECT 820.950 528.450 825.000 529.050 ;
        RECT 814.950 526.050 816.750 527.850 ;
        RECT 820.950 526.950 825.450 528.450 ;
        RECT 787.950 523.950 790.050 526.050 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 808.950 523.950 811.050 526.050 ;
        RECT 811.950 523.950 814.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 788.100 522.150 789.900 523.950 ;
        RECT 791.100 519.600 792.300 523.950 ;
        RECT 794.100 522.150 795.900 523.950 ;
        RECT 760.950 518.550 780.450 519.450 ;
        RECT 788.700 518.700 792.300 519.600 ;
        RECT 760.950 517.950 763.050 518.550 ;
        RECT 788.700 516.600 789.900 518.700 ;
        RECT 758.700 514.500 771.300 515.400 ;
        RECT 763.200 513.600 764.100 514.500 ;
        RECT 770.400 513.600 771.300 514.500 ;
        RECT 763.200 510.600 765.900 513.600 ;
        RECT 767.100 510.000 768.900 513.600 ;
        RECT 770.100 510.600 771.900 513.600 ;
        RECT 773.100 510.000 775.200 513.600 ;
        RECT 788.100 510.600 789.900 516.600 ;
        RECT 791.100 515.700 798.900 517.050 ;
        RECT 791.100 510.600 792.900 515.700 ;
        RECT 794.100 510.000 795.900 514.800 ;
        RECT 797.100 510.600 798.900 515.700 ;
        RECT 809.400 516.600 810.300 523.950 ;
        RECT 811.950 522.150 813.750 523.950 ;
        RECT 818.100 522.150 819.900 523.950 ;
        RECT 824.550 523.050 825.450 526.950 ;
        RECT 833.100 526.050 834.300 533.400 ;
        RECT 850.950 528.450 853.050 529.050 ;
        RECT 839.100 526.050 840.900 527.850 ;
        RECT 845.550 527.550 853.050 528.450 ;
        RECT 829.950 523.950 832.050 526.050 ;
        RECT 832.950 523.950 835.050 526.050 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 824.550 521.550 829.050 523.050 ;
        RECT 830.100 522.150 831.900 523.950 ;
        RECT 825.000 520.950 829.050 521.550 ;
        RECT 833.100 519.600 834.300 523.950 ;
        RECT 836.100 522.150 837.900 523.950 ;
        RECT 845.550 523.050 846.450 527.550 ;
        RECT 850.950 526.950 853.050 527.550 ;
        RECT 855.000 526.050 855.900 538.200 ;
        RECT 875.100 533.400 876.900 545.400 ;
        RECT 878.100 534.300 879.900 545.400 ;
        RECT 881.100 535.200 882.900 546.000 ;
        RECT 884.100 534.300 885.900 545.400 ;
        RECT 878.100 533.400 885.900 534.300 ;
        RECT 896.100 533.400 897.900 545.400 ;
        RECT 899.100 534.300 900.900 545.400 ;
        RECT 902.100 535.200 903.900 546.000 ;
        RECT 905.100 534.300 906.900 545.400 ;
        RECT 920.100 539.400 921.900 545.400 ;
        RECT 923.100 540.000 924.900 546.000 ;
        RECT 899.100 533.400 906.900 534.300 ;
        RECT 921.000 539.100 921.900 539.400 ;
        RECT 926.100 539.400 927.900 545.400 ;
        RECT 929.100 539.400 930.900 546.000 ;
        RECT 926.100 539.100 927.600 539.400 ;
        RECT 921.000 538.200 927.600 539.100 ;
        RECT 865.950 528.450 870.000 529.050 ;
        RECT 860.100 526.050 861.900 527.850 ;
        RECT 865.950 526.950 870.450 528.450 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 841.950 521.550 846.450 523.050 ;
        RECT 841.950 520.950 846.000 521.550 ;
        RECT 830.700 518.700 834.300 519.600 ;
        RECT 855.000 520.200 855.900 523.950 ;
        RECT 857.100 522.150 858.900 523.950 ;
        RECT 863.100 522.150 864.900 523.950 ;
        RECT 869.550 523.050 870.450 526.950 ;
        RECT 875.400 526.050 876.300 533.400 ;
        RECT 880.950 531.450 883.050 532.050 ;
        RECT 880.950 530.550 891.450 531.450 ;
        RECT 880.950 529.950 883.050 530.550 ;
        RECT 880.950 526.050 882.750 527.850 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 880.950 523.950 883.050 526.050 ;
        RECT 883.950 523.950 886.050 526.050 ;
        RECT 865.950 521.550 870.450 523.050 ;
        RECT 865.950 520.950 870.000 521.550 ;
        RECT 855.000 519.000 858.300 520.200 ;
        RECT 830.700 516.600 831.900 518.700 ;
        RECT 809.400 515.400 814.500 516.600 ;
        RECT 809.700 510.000 811.500 513.600 ;
        RECT 812.700 510.600 814.500 515.400 ;
        RECT 817.200 510.000 819.000 516.600 ;
        RECT 830.100 510.600 831.900 516.600 ;
        RECT 833.100 515.700 840.900 517.050 ;
        RECT 833.100 510.600 834.900 515.700 ;
        RECT 836.100 510.000 837.900 514.800 ;
        RECT 839.100 510.600 840.900 515.700 ;
        RECT 856.500 510.600 858.300 519.000 ;
        RECT 863.100 510.000 864.900 519.600 ;
        RECT 875.400 516.600 876.300 523.950 ;
        RECT 877.950 522.150 879.750 523.950 ;
        RECT 884.100 522.150 885.900 523.950 ;
        RECT 890.550 523.050 891.450 530.550 ;
        RECT 896.400 526.050 897.300 533.400 ;
        RECT 910.950 529.950 913.050 532.050 ;
        RECT 901.950 526.050 903.750 527.850 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 890.550 521.550 895.050 523.050 ;
        RECT 891.000 520.950 895.050 521.550 ;
        RECT 896.400 516.600 897.300 523.950 ;
        RECT 898.950 522.150 900.750 523.950 ;
        RECT 905.100 522.150 906.900 523.950 ;
        RECT 911.550 522.450 912.450 529.950 ;
        RECT 921.000 526.050 921.900 538.200 ;
        RECT 926.100 526.050 927.900 527.850 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 922.950 523.950 925.050 526.050 ;
        RECT 925.950 523.950 928.050 526.050 ;
        RECT 928.950 523.950 931.050 526.050 ;
        RECT 916.950 522.450 919.050 523.050 ;
        RECT 911.550 521.550 919.050 522.450 ;
        RECT 916.950 520.950 919.050 521.550 ;
        RECT 921.000 520.200 921.900 523.950 ;
        RECT 923.100 522.150 924.900 523.950 ;
        RECT 929.100 522.150 930.900 523.950 ;
        RECT 904.950 519.450 907.050 520.050 ;
        RECT 910.950 519.450 913.050 520.050 ;
        RECT 904.950 518.550 913.050 519.450 ;
        RECT 921.000 519.000 924.300 520.200 ;
        RECT 904.950 517.950 907.050 518.550 ;
        RECT 910.950 517.950 913.050 518.550 ;
        RECT 875.400 515.400 880.500 516.600 ;
        RECT 875.700 510.000 877.500 513.600 ;
        RECT 878.700 510.600 880.500 515.400 ;
        RECT 883.200 510.000 885.000 516.600 ;
        RECT 896.400 515.400 901.500 516.600 ;
        RECT 896.700 510.000 898.500 513.600 ;
        RECT 899.700 510.600 901.500 515.400 ;
        RECT 904.200 510.000 906.000 516.600 ;
        RECT 922.500 510.600 924.300 519.000 ;
        RECT 929.100 510.000 930.900 519.600 ;
        RECT 14.100 500.400 15.900 506.400 ;
        RECT 17.100 500.400 18.900 507.000 ;
        RECT 20.100 503.400 21.900 506.400 ;
        RECT 14.100 493.050 15.300 500.400 ;
        RECT 20.700 499.500 21.900 503.400 ;
        RECT 16.200 498.600 21.900 499.500 ;
        RECT 23.700 500.400 25.500 506.400 ;
        RECT 29.100 500.400 30.900 507.000 ;
        RECT 34.500 500.400 36.300 506.400 ;
        RECT 38.700 503.400 40.500 506.400 ;
        RECT 41.700 503.400 43.500 506.400 ;
        RECT 44.700 503.400 46.500 506.400 ;
        RECT 47.700 503.400 49.500 507.000 ;
        RECT 38.700 501.300 40.800 503.400 ;
        RECT 41.700 501.300 43.800 503.400 ;
        RECT 44.700 501.300 46.800 503.400 ;
        RECT 52.200 502.500 54.000 506.400 ;
        RECT 55.200 503.400 57.000 507.000 ;
        RECT 58.200 503.400 60.000 506.400 ;
        RECT 61.200 503.400 63.000 506.400 ;
        RECT 64.200 503.400 66.000 506.400 ;
        RECT 67.200 503.400 69.000 506.400 ;
        RECT 48.600 501.600 50.400 502.500 ;
        RECT 47.700 500.400 50.400 501.600 ;
        RECT 52.200 500.400 54.900 502.500 ;
        RECT 58.200 501.300 60.300 503.400 ;
        RECT 61.200 501.300 63.300 503.400 ;
        RECT 64.200 501.300 66.300 503.400 ;
        RECT 67.200 501.300 69.300 503.400 ;
        RECT 71.400 501.600 73.200 506.400 ;
        RECT 71.400 500.400 75.600 501.600 ;
        RECT 76.500 500.400 78.300 507.000 ;
        RECT 81.900 500.400 83.700 506.400 ;
        RECT 16.200 497.700 18.000 498.600 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 14.100 483.600 15.300 490.950 ;
        RECT 17.100 486.300 18.000 497.700 ;
        RECT 23.700 496.800 24.900 500.400 ;
        RECT 34.800 499.500 36.300 500.400 ;
        RECT 43.800 499.800 45.600 500.400 ;
        RECT 47.700 499.800 48.600 500.400 ;
        RECT 27.900 498.300 36.300 499.500 ;
        RECT 41.400 498.600 48.600 499.800 ;
        RECT 63.300 498.600 69.900 500.400 ;
        RECT 27.900 497.700 29.700 498.300 ;
        RECT 38.400 496.800 40.500 497.700 ;
        RECT 23.700 495.600 40.500 496.800 ;
        RECT 41.400 495.600 42.300 498.600 ;
        RECT 46.800 495.900 48.600 496.800 ;
        RECT 56.100 496.500 57.900 498.300 ;
        RECT 74.100 497.100 75.600 500.400 ;
        RECT 49.800 495.900 51.900 496.050 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 19.800 489.150 21.600 490.950 ;
        RECT 16.200 485.400 18.000 486.300 ;
        RECT 16.200 484.500 21.900 485.400 ;
        RECT 14.100 471.600 15.900 483.600 ;
        RECT 17.100 471.000 18.900 481.800 ;
        RECT 20.700 477.600 21.900 484.500 ;
        RECT 23.700 479.400 24.900 495.600 ;
        RECT 41.400 493.800 43.200 495.600 ;
        RECT 46.800 495.000 51.900 495.900 ;
        RECT 49.800 493.950 51.900 495.000 ;
        RECT 56.100 495.900 58.200 496.500 ;
        RECT 56.100 494.400 73.200 495.900 ;
        RECT 74.100 495.300 81.900 497.100 ;
        RECT 71.700 492.900 78.300 494.400 ;
        RECT 26.100 491.700 70.500 492.900 ;
        RECT 26.100 490.050 27.900 491.700 ;
        RECT 25.800 487.950 27.900 490.050 ;
        RECT 31.800 489.750 33.900 490.050 ;
        RECT 44.400 489.900 46.200 490.500 ;
        RECT 53.400 489.900 66.900 490.800 ;
        RECT 31.800 487.950 35.700 489.750 ;
        RECT 44.400 488.700 55.500 489.900 ;
        RECT 33.900 487.200 35.700 487.950 ;
        RECT 53.400 487.800 55.500 488.700 ;
        RECT 57.000 487.200 60.900 489.000 ;
        RECT 66.000 488.700 66.900 489.900 ;
        RECT 33.900 486.300 47.400 487.200 ;
        RECT 58.800 486.900 60.900 487.200 ;
        RECT 65.100 486.900 66.900 488.700 ;
        RECT 69.600 490.200 70.500 491.700 ;
        RECT 69.600 488.400 74.700 490.200 ;
        RECT 76.800 490.050 78.300 492.900 ;
        RECT 76.800 487.950 78.900 490.050 ;
        RECT 46.200 485.700 47.400 486.300 ;
        RECT 80.100 485.700 81.900 486.300 ;
        RECT 41.400 484.500 43.500 484.800 ;
        RECT 46.200 484.500 81.900 485.700 ;
        RECT 31.500 483.300 43.500 484.500 ;
        RECT 82.800 483.600 83.700 500.400 ;
        RECT 31.500 482.700 33.300 483.300 ;
        RECT 41.400 482.700 43.500 483.300 ;
        RECT 46.200 482.400 63.900 483.600 ;
        RECT 28.200 481.800 30.000 482.100 ;
        RECT 46.200 481.800 47.400 482.400 ;
        RECT 28.200 480.600 47.400 481.800 ;
        RECT 61.800 481.500 63.900 482.400 ;
        RECT 67.200 482.700 83.700 483.600 ;
        RECT 67.200 481.500 69.300 482.700 ;
        RECT 28.200 480.300 30.000 480.600 ;
        RECT 23.700 478.500 27.300 479.400 ;
        RECT 26.400 477.600 27.300 478.500 ;
        RECT 20.100 471.600 21.900 477.600 ;
        RECT 23.700 471.000 25.500 477.600 ;
        RECT 26.400 476.700 28.500 477.600 ;
        RECT 26.700 471.600 28.500 476.700 ;
        RECT 29.700 471.000 31.500 477.600 ;
        RECT 32.700 471.600 34.500 480.600 ;
        RECT 44.700 477.600 46.800 479.700 ;
        RECT 52.200 479.100 55.500 481.200 ;
        RECT 35.700 471.000 37.500 477.600 ;
        RECT 39.300 474.600 41.400 476.700 ;
        RECT 42.300 474.600 44.400 476.700 ;
        RECT 39.300 471.600 41.100 474.600 ;
        RECT 42.300 471.600 44.100 474.600 ;
        RECT 45.300 471.600 47.100 477.600 ;
        RECT 48.300 471.000 50.100 477.600 ;
        RECT 52.200 471.600 54.000 479.100 ;
        RECT 58.200 477.600 60.900 481.500 ;
        RECT 73.200 480.600 78.900 481.800 ;
        RECT 70.500 479.700 72.300 480.300 ;
        RECT 64.200 478.500 72.300 479.700 ;
        RECT 64.200 477.600 66.300 478.500 ;
        RECT 73.200 477.600 74.400 480.600 ;
        RECT 77.100 480.000 78.900 480.600 ;
        RECT 82.800 479.400 83.700 482.700 ;
        RECT 79.800 478.500 83.700 479.400 ;
        RECT 85.500 503.400 87.300 506.400 ;
        RECT 88.500 503.400 90.300 507.000 ;
        RECT 104.100 503.400 105.900 507.000 ;
        RECT 107.100 503.400 108.900 506.400 ;
        RECT 110.100 503.400 111.900 507.000 ;
        RECT 85.500 490.050 87.000 503.400 ;
        RECT 107.400 493.050 108.300 503.400 ;
        RECT 113.700 500.400 115.500 506.400 ;
        RECT 119.100 500.400 120.900 507.000 ;
        RECT 124.500 500.400 126.300 506.400 ;
        RECT 128.700 503.400 130.500 506.400 ;
        RECT 131.700 503.400 133.500 506.400 ;
        RECT 134.700 503.400 136.500 506.400 ;
        RECT 137.700 503.400 139.500 507.000 ;
        RECT 128.700 501.300 130.800 503.400 ;
        RECT 131.700 501.300 133.800 503.400 ;
        RECT 134.700 501.300 136.800 503.400 ;
        RECT 142.200 502.500 144.000 506.400 ;
        RECT 145.200 503.400 147.000 507.000 ;
        RECT 148.200 503.400 150.000 506.400 ;
        RECT 151.200 503.400 153.000 506.400 ;
        RECT 154.200 503.400 156.000 506.400 ;
        RECT 157.200 503.400 159.000 506.400 ;
        RECT 138.600 501.600 140.400 502.500 ;
        RECT 137.700 500.400 140.400 501.600 ;
        RECT 142.200 500.400 144.900 502.500 ;
        RECT 148.200 501.300 150.300 503.400 ;
        RECT 151.200 501.300 153.300 503.400 ;
        RECT 154.200 501.300 156.300 503.400 ;
        RECT 157.200 501.300 159.300 503.400 ;
        RECT 161.400 501.600 163.200 506.400 ;
        RECT 161.400 500.400 165.600 501.600 ;
        RECT 166.500 500.400 168.300 507.000 ;
        RECT 171.900 500.400 173.700 506.400 ;
        RECT 113.700 496.800 114.900 500.400 ;
        RECT 124.800 499.500 126.300 500.400 ;
        RECT 133.800 499.800 135.600 500.400 ;
        RECT 137.700 499.800 138.600 500.400 ;
        RECT 117.900 498.300 126.300 499.500 ;
        RECT 131.400 498.600 138.600 499.800 ;
        RECT 153.300 498.600 159.900 500.400 ;
        RECT 117.900 497.700 119.700 498.300 ;
        RECT 128.400 496.800 130.500 497.700 ;
        RECT 113.700 495.600 130.500 496.800 ;
        RECT 131.400 495.600 132.300 498.600 ;
        RECT 136.800 495.900 138.600 496.800 ;
        RECT 146.100 496.500 147.900 498.300 ;
        RECT 164.100 497.100 165.600 500.400 ;
        RECT 139.800 495.900 141.900 496.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 85.500 487.950 87.900 490.050 ;
        RECT 104.250 489.150 106.050 490.950 ;
        RECT 79.800 477.600 81.000 478.500 ;
        RECT 85.500 477.600 87.000 487.950 ;
        RECT 107.400 483.600 108.300 490.950 ;
        RECT 110.100 489.150 111.900 490.950 ;
        RECT 55.200 471.000 57.000 477.600 ;
        RECT 58.200 471.600 60.000 477.600 ;
        RECT 61.200 474.600 63.300 476.700 ;
        RECT 64.200 474.600 66.300 476.700 ;
        RECT 67.200 474.600 69.300 476.700 ;
        RECT 61.200 471.600 63.000 474.600 ;
        RECT 64.200 471.600 66.000 474.600 ;
        RECT 67.200 471.600 69.000 474.600 ;
        RECT 70.200 471.000 72.000 477.600 ;
        RECT 73.200 471.600 75.000 477.600 ;
        RECT 76.200 471.000 78.000 477.600 ;
        RECT 79.200 471.600 81.000 477.600 ;
        RECT 82.200 471.000 84.000 477.600 ;
        RECT 85.500 471.600 87.300 477.600 ;
        RECT 88.500 471.000 90.300 477.600 ;
        RECT 104.100 471.000 105.900 483.600 ;
        RECT 107.400 482.400 111.000 483.600 ;
        RECT 109.200 471.600 111.000 482.400 ;
        RECT 113.700 479.400 114.900 495.600 ;
        RECT 131.400 493.800 133.200 495.600 ;
        RECT 136.800 495.000 141.900 495.900 ;
        RECT 139.800 493.950 141.900 495.000 ;
        RECT 146.100 495.900 148.200 496.500 ;
        RECT 146.100 494.400 163.200 495.900 ;
        RECT 164.100 495.300 171.900 497.100 ;
        RECT 161.700 492.900 168.300 494.400 ;
        RECT 116.100 491.700 160.500 492.900 ;
        RECT 116.100 490.050 117.900 491.700 ;
        RECT 115.800 487.950 117.900 490.050 ;
        RECT 121.800 489.750 123.900 490.050 ;
        RECT 134.400 489.900 136.200 490.500 ;
        RECT 143.400 489.900 156.900 490.800 ;
        RECT 121.800 487.950 125.700 489.750 ;
        RECT 134.400 488.700 145.500 489.900 ;
        RECT 123.900 487.200 125.700 487.950 ;
        RECT 143.400 487.800 145.500 488.700 ;
        RECT 147.000 487.200 150.900 489.000 ;
        RECT 156.000 488.700 156.900 489.900 ;
        RECT 123.900 486.300 137.400 487.200 ;
        RECT 148.800 486.900 150.900 487.200 ;
        RECT 155.100 486.900 156.900 488.700 ;
        RECT 159.600 490.200 160.500 491.700 ;
        RECT 159.600 488.400 164.700 490.200 ;
        RECT 166.800 490.050 168.300 492.900 ;
        RECT 166.800 487.950 168.900 490.050 ;
        RECT 136.200 485.700 137.400 486.300 ;
        RECT 170.100 485.700 171.900 486.300 ;
        RECT 131.400 484.500 133.500 484.800 ;
        RECT 136.200 484.500 171.900 485.700 ;
        RECT 121.500 483.300 133.500 484.500 ;
        RECT 172.800 483.600 173.700 500.400 ;
        RECT 121.500 482.700 123.300 483.300 ;
        RECT 131.400 482.700 133.500 483.300 ;
        RECT 136.200 482.400 153.900 483.600 ;
        RECT 118.200 481.800 120.000 482.100 ;
        RECT 136.200 481.800 137.400 482.400 ;
        RECT 118.200 480.600 137.400 481.800 ;
        RECT 151.800 481.500 153.900 482.400 ;
        RECT 157.200 482.700 173.700 483.600 ;
        RECT 157.200 481.500 159.300 482.700 ;
        RECT 118.200 480.300 120.000 480.600 ;
        RECT 113.700 478.500 117.300 479.400 ;
        RECT 116.400 477.600 117.300 478.500 ;
        RECT 113.700 471.000 115.500 477.600 ;
        RECT 116.400 476.700 118.500 477.600 ;
        RECT 116.700 471.600 118.500 476.700 ;
        RECT 119.700 471.000 121.500 477.600 ;
        RECT 122.700 471.600 124.500 480.600 ;
        RECT 134.700 477.600 136.800 479.700 ;
        RECT 142.200 479.100 145.500 481.200 ;
        RECT 125.700 471.000 127.500 477.600 ;
        RECT 129.300 474.600 131.400 476.700 ;
        RECT 132.300 474.600 134.400 476.700 ;
        RECT 129.300 471.600 131.100 474.600 ;
        RECT 132.300 471.600 134.100 474.600 ;
        RECT 135.300 471.600 137.100 477.600 ;
        RECT 138.300 471.000 140.100 477.600 ;
        RECT 142.200 471.600 144.000 479.100 ;
        RECT 148.200 477.600 150.900 481.500 ;
        RECT 163.200 480.600 168.900 481.800 ;
        RECT 160.500 479.700 162.300 480.300 ;
        RECT 154.200 478.500 162.300 479.700 ;
        RECT 154.200 477.600 156.300 478.500 ;
        RECT 163.200 477.600 164.400 480.600 ;
        RECT 167.100 480.000 168.900 480.600 ;
        RECT 172.800 479.400 173.700 482.700 ;
        RECT 169.800 478.500 173.700 479.400 ;
        RECT 175.500 503.400 177.300 506.400 ;
        RECT 178.500 503.400 180.300 507.000 ;
        RECT 194.700 503.400 196.500 507.000 ;
        RECT 175.500 490.050 177.000 503.400 ;
        RECT 197.700 501.600 199.500 506.400 ;
        RECT 194.400 500.400 199.500 501.600 ;
        RECT 202.200 500.400 204.000 507.000 ;
        RECT 218.400 500.400 220.200 507.000 ;
        RECT 189.000 495.450 193.050 496.050 ;
        RECT 188.550 495.000 193.050 495.450 ;
        RECT 187.950 493.950 193.050 495.000 ;
        RECT 187.950 490.800 190.050 493.950 ;
        RECT 194.400 493.050 195.300 500.400 ;
        RECT 223.500 499.200 225.300 506.400 ;
        RECT 239.100 501.300 240.900 506.400 ;
        RECT 242.100 502.200 243.900 507.000 ;
        RECT 245.100 501.300 246.900 506.400 ;
        RECT 239.100 499.950 246.900 501.300 ;
        RECT 248.100 500.400 249.900 506.400 ;
        RECT 211.950 496.950 214.050 499.050 ;
        RECT 221.100 498.300 225.300 499.200 ;
        RECT 248.100 498.300 249.300 500.400 ;
        RECT 260.700 499.200 262.500 506.400 ;
        RECT 265.800 500.400 267.600 507.000 ;
        RECT 278.100 503.400 279.900 506.400 ;
        RECT 278.100 499.500 279.300 503.400 ;
        RECT 281.100 500.400 282.900 507.000 ;
        RECT 284.100 500.400 285.900 506.400 ;
        RECT 296.100 500.400 297.900 507.000 ;
        RECT 260.700 498.300 264.900 499.200 ;
        RECT 278.100 498.600 283.800 499.500 ;
        RECT 205.950 495.450 210.000 496.050 ;
        RECT 196.950 493.050 198.750 494.850 ;
        RECT 203.100 493.050 204.900 494.850 ;
        RECT 205.950 493.950 210.450 495.450 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 175.500 487.950 177.900 490.050 ;
        RECT 169.800 477.600 171.000 478.500 ;
        RECT 175.500 477.600 177.000 487.950 ;
        RECT 194.400 483.600 195.300 490.950 ;
        RECT 199.950 489.150 201.750 490.950 ;
        RECT 209.550 490.050 210.450 493.950 ;
        RECT 205.950 488.550 210.450 490.050 ;
        RECT 205.950 487.950 210.000 488.550 ;
        RECT 202.950 486.450 205.050 487.050 ;
        RECT 212.550 486.450 213.450 496.950 ;
        RECT 218.250 493.050 220.050 494.850 ;
        RECT 221.100 493.050 222.300 498.300 ;
        RECT 245.700 497.400 249.300 498.300 ;
        RECT 224.100 493.050 225.900 494.850 ;
        RECT 242.100 493.050 243.900 494.850 ;
        RECT 245.700 493.050 246.900 497.400 ;
        RECT 248.100 493.050 249.900 494.850 ;
        RECT 260.100 493.050 261.900 494.850 ;
        RECT 263.700 493.050 264.900 498.300 ;
        RECT 282.000 497.700 283.800 498.600 ;
        RECT 265.950 493.050 267.750 494.850 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 278.400 490.950 280.500 493.050 ;
        RECT 202.950 485.550 213.450 486.450 ;
        RECT 202.950 484.950 205.050 485.550 ;
        RECT 145.200 471.000 147.000 477.600 ;
        RECT 148.200 471.600 150.000 477.600 ;
        RECT 151.200 474.600 153.300 476.700 ;
        RECT 154.200 474.600 156.300 476.700 ;
        RECT 157.200 474.600 159.300 476.700 ;
        RECT 151.200 471.600 153.000 474.600 ;
        RECT 154.200 471.600 156.000 474.600 ;
        RECT 157.200 471.600 159.000 474.600 ;
        RECT 160.200 471.000 162.000 477.600 ;
        RECT 163.200 471.600 165.000 477.600 ;
        RECT 166.200 471.000 168.000 477.600 ;
        RECT 169.200 471.600 171.000 477.600 ;
        RECT 172.200 471.000 174.000 477.600 ;
        RECT 175.500 471.600 177.300 477.600 ;
        RECT 178.500 471.000 180.300 477.600 ;
        RECT 194.100 471.600 195.900 483.600 ;
        RECT 197.100 482.700 204.900 483.600 ;
        RECT 197.100 471.600 198.900 482.700 ;
        RECT 200.100 471.000 201.900 481.800 ;
        RECT 203.100 471.600 204.900 482.700 ;
        RECT 221.100 477.600 222.300 490.950 ;
        RECT 239.100 489.150 240.900 490.950 ;
        RECT 245.700 483.600 246.900 490.950 ;
        RECT 218.100 471.000 219.900 477.600 ;
        RECT 221.100 471.600 222.900 477.600 ;
        RECT 224.100 471.000 225.900 477.600 ;
        RECT 239.400 471.000 241.200 483.600 ;
        RECT 244.500 482.100 246.900 483.600 ;
        RECT 244.500 471.600 246.300 482.100 ;
        RECT 247.200 479.100 249.000 480.900 ;
        RECT 263.700 477.600 264.900 490.950 ;
        RECT 278.400 489.150 280.200 490.950 ;
        RECT 282.000 486.300 282.900 497.700 ;
        RECT 284.700 493.050 285.900 500.400 ;
        RECT 299.100 499.500 300.900 506.400 ;
        RECT 302.100 500.400 303.900 507.000 ;
        RECT 305.100 499.500 306.900 506.400 ;
        RECT 308.100 500.400 309.900 507.000 ;
        RECT 311.100 499.500 312.900 506.400 ;
        RECT 314.100 500.400 315.900 507.000 ;
        RECT 317.100 499.500 318.900 506.400 ;
        RECT 320.100 500.400 321.900 507.000 ;
        RECT 335.100 500.400 336.900 507.000 ;
        RECT 283.800 490.950 285.900 493.050 ;
        RECT 282.000 485.400 283.800 486.300 ;
        RECT 278.100 484.500 283.800 485.400 ;
        RECT 278.100 477.600 279.300 484.500 ;
        RECT 284.700 483.600 285.900 490.950 ;
        RECT 298.050 498.300 300.900 499.500 ;
        RECT 303.000 498.300 306.900 499.500 ;
        RECT 309.000 498.300 312.900 499.500 ;
        RECT 315.000 498.300 318.900 499.500 ;
        RECT 338.100 499.500 339.900 506.400 ;
        RECT 341.100 500.400 342.900 507.000 ;
        RECT 344.100 499.500 345.900 506.400 ;
        RECT 347.100 500.400 348.900 507.000 ;
        RECT 350.100 499.500 351.900 506.400 ;
        RECT 353.100 500.400 354.900 507.000 ;
        RECT 356.100 499.500 357.900 506.400 ;
        RECT 359.100 500.400 360.900 507.000 ;
        RECT 371.100 500.400 372.900 506.400 ;
        RECT 374.100 500.400 375.900 507.000 ;
        RECT 377.100 503.400 378.900 506.400 ;
        RECT 338.100 498.300 342.000 499.500 ;
        RECT 344.100 498.300 348.000 499.500 ;
        RECT 350.100 498.300 354.000 499.500 ;
        RECT 356.100 498.300 358.950 499.500 ;
        RECT 298.050 493.050 299.100 498.300 ;
        RECT 303.000 497.400 304.200 498.300 ;
        RECT 309.000 497.400 310.200 498.300 ;
        RECT 315.000 497.400 316.200 498.300 ;
        RECT 300.000 496.200 304.200 497.400 ;
        RECT 300.000 495.600 301.800 496.200 ;
        RECT 298.050 490.950 301.200 493.050 ;
        RECT 298.050 485.700 299.100 490.950 ;
        RECT 303.000 485.700 304.200 496.200 ;
        RECT 306.000 496.200 310.200 497.400 ;
        RECT 306.000 495.600 307.800 496.200 ;
        RECT 309.000 485.700 310.200 496.200 ;
        RECT 312.000 496.200 316.200 497.400 ;
        RECT 312.000 495.600 313.800 496.200 ;
        RECT 315.000 485.700 316.200 496.200 ;
        RECT 340.800 497.400 342.000 498.300 ;
        RECT 346.800 497.400 348.000 498.300 ;
        RECT 352.800 497.400 354.000 498.300 ;
        RECT 340.800 496.200 345.000 497.400 ;
        RECT 317.400 493.050 319.200 494.850 ;
        RECT 317.100 490.950 319.200 493.050 ;
        RECT 337.800 493.050 339.600 494.850 ;
        RECT 337.800 490.950 339.900 493.050 ;
        RECT 340.800 485.700 342.000 496.200 ;
        RECT 343.200 495.600 345.000 496.200 ;
        RECT 346.800 496.200 351.000 497.400 ;
        RECT 346.800 485.700 348.000 496.200 ;
        RECT 349.200 495.600 351.000 496.200 ;
        RECT 352.800 496.200 357.000 497.400 ;
        RECT 352.800 485.700 354.000 496.200 ;
        RECT 355.200 495.600 357.000 496.200 ;
        RECT 357.900 493.050 358.950 498.300 ;
        RECT 355.800 490.950 358.950 493.050 ;
        RECT 357.900 485.700 358.950 490.950 ;
        RECT 298.050 484.500 300.900 485.700 ;
        RECT 303.000 484.500 306.900 485.700 ;
        RECT 309.000 484.500 312.900 485.700 ;
        RECT 315.000 484.500 318.900 485.700 ;
        RECT 247.500 471.000 249.300 477.600 ;
        RECT 260.100 471.000 261.900 477.600 ;
        RECT 263.100 471.600 264.900 477.600 ;
        RECT 266.100 471.000 267.900 477.600 ;
        RECT 278.100 471.600 279.900 477.600 ;
        RECT 281.100 471.000 282.900 481.800 ;
        RECT 284.100 471.600 285.900 483.600 ;
        RECT 296.100 471.000 297.900 483.600 ;
        RECT 299.100 471.600 300.900 484.500 ;
        RECT 302.100 471.000 303.900 483.600 ;
        RECT 305.100 471.600 306.900 484.500 ;
        RECT 308.100 471.000 309.900 483.600 ;
        RECT 311.100 471.600 312.900 484.500 ;
        RECT 314.100 471.000 315.900 483.600 ;
        RECT 317.100 471.600 318.900 484.500 ;
        RECT 338.100 484.500 342.000 485.700 ;
        RECT 344.100 484.500 348.000 485.700 ;
        RECT 350.100 484.500 354.000 485.700 ;
        RECT 356.100 484.500 358.950 485.700 ;
        RECT 371.100 493.050 372.300 500.400 ;
        RECT 377.700 499.500 378.900 503.400 ;
        RECT 373.200 498.600 378.900 499.500 ;
        RECT 392.100 503.400 393.900 506.400 ;
        RECT 392.100 499.500 393.300 503.400 ;
        RECT 395.100 500.400 396.900 507.000 ;
        RECT 398.100 500.400 399.900 506.400 ;
        RECT 410.400 500.400 412.200 507.000 ;
        RECT 392.100 498.600 397.800 499.500 ;
        RECT 373.200 497.700 375.000 498.600 ;
        RECT 371.100 490.950 373.200 493.050 ;
        RECT 320.100 471.000 321.900 483.600 ;
        RECT 335.100 471.000 336.900 483.600 ;
        RECT 338.100 471.600 339.900 484.500 ;
        RECT 341.100 471.000 342.900 483.600 ;
        RECT 344.100 471.600 345.900 484.500 ;
        RECT 347.100 471.000 348.900 483.600 ;
        RECT 350.100 471.600 351.900 484.500 ;
        RECT 353.100 471.000 354.900 483.600 ;
        RECT 356.100 471.600 357.900 484.500 ;
        RECT 371.100 483.600 372.300 490.950 ;
        RECT 374.100 486.300 375.000 497.700 ;
        RECT 396.000 497.700 397.800 498.600 ;
        RECT 376.500 490.950 378.600 493.050 ;
        RECT 376.800 489.150 378.600 490.950 ;
        RECT 392.400 490.950 394.500 493.050 ;
        RECT 392.400 489.150 394.200 490.950 ;
        RECT 373.200 485.400 375.000 486.300 ;
        RECT 396.000 486.300 396.900 497.700 ;
        RECT 398.700 493.050 399.900 500.400 ;
        RECT 415.500 499.200 417.300 506.400 ;
        RECT 431.100 500.400 432.900 506.400 ;
        RECT 413.100 498.300 417.300 499.200 ;
        RECT 431.700 498.300 432.900 500.400 ;
        RECT 434.100 501.300 435.900 506.400 ;
        RECT 437.100 502.200 438.900 507.000 ;
        RECT 440.100 501.300 441.900 506.400 ;
        RECT 443.700 503.400 445.500 507.000 ;
        RECT 446.700 503.400 448.500 506.400 ;
        RECT 434.100 499.950 441.900 501.300 ;
        RECT 410.250 493.050 412.050 494.850 ;
        RECT 413.100 493.050 414.300 498.300 ;
        RECT 431.700 497.400 435.300 498.300 ;
        RECT 416.100 493.050 417.900 494.850 ;
        RECT 431.100 493.050 432.900 494.850 ;
        RECT 434.100 493.050 435.300 497.400 ;
        RECT 437.100 493.050 438.900 494.850 ;
        RECT 397.800 490.950 399.900 493.050 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 412.950 490.950 415.050 493.050 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 396.000 485.400 397.800 486.300 ;
        RECT 373.200 484.500 378.900 485.400 ;
        RECT 359.100 471.000 360.900 483.600 ;
        RECT 371.100 471.600 372.900 483.600 ;
        RECT 374.100 471.000 375.900 481.800 ;
        RECT 377.700 477.600 378.900 484.500 ;
        RECT 377.100 471.600 378.900 477.600 ;
        RECT 392.100 484.500 397.800 485.400 ;
        RECT 392.100 477.600 393.300 484.500 ;
        RECT 398.700 483.600 399.900 490.950 ;
        RECT 392.100 471.600 393.900 477.600 ;
        RECT 395.100 471.000 396.900 481.800 ;
        RECT 398.100 471.600 399.900 483.600 ;
        RECT 413.100 477.600 414.300 490.950 ;
        RECT 434.100 483.600 435.300 490.950 ;
        RECT 440.100 489.150 441.900 490.950 ;
        RECT 447.000 490.050 448.500 503.400 ;
        RECT 446.100 487.950 448.500 490.050 ;
        RECT 434.100 482.100 436.500 483.600 ;
        RECT 432.000 479.100 433.800 480.900 ;
        RECT 410.100 471.000 411.900 477.600 ;
        RECT 413.100 471.600 414.900 477.600 ;
        RECT 416.100 471.000 417.900 477.600 ;
        RECT 431.700 471.000 433.500 477.600 ;
        RECT 434.700 471.600 436.500 482.100 ;
        RECT 439.800 471.000 441.600 483.600 ;
        RECT 447.000 477.600 448.500 487.950 ;
        RECT 450.300 500.400 452.100 506.400 ;
        RECT 455.700 500.400 457.500 507.000 ;
        RECT 460.800 501.600 462.600 506.400 ;
        RECT 465.000 503.400 466.800 506.400 ;
        RECT 468.000 503.400 469.800 506.400 ;
        RECT 471.000 503.400 472.800 506.400 ;
        RECT 474.000 503.400 475.800 506.400 ;
        RECT 477.000 503.400 478.800 507.000 ;
        RECT 458.400 500.400 462.600 501.600 ;
        RECT 464.700 501.300 466.800 503.400 ;
        RECT 467.700 501.300 469.800 503.400 ;
        RECT 470.700 501.300 472.800 503.400 ;
        RECT 473.700 501.300 475.800 503.400 ;
        RECT 480.000 502.500 481.800 506.400 ;
        RECT 484.500 503.400 486.300 507.000 ;
        RECT 487.500 503.400 489.300 506.400 ;
        RECT 490.500 503.400 492.300 506.400 ;
        RECT 493.500 503.400 495.300 506.400 ;
        RECT 479.100 500.400 481.800 502.500 ;
        RECT 483.600 501.600 485.400 502.500 ;
        RECT 483.600 500.400 486.300 501.600 ;
        RECT 487.200 501.300 489.300 503.400 ;
        RECT 490.200 501.300 492.300 503.400 ;
        RECT 493.200 501.300 495.300 503.400 ;
        RECT 497.700 500.400 499.500 506.400 ;
        RECT 503.100 500.400 504.900 507.000 ;
        RECT 508.500 500.400 510.300 506.400 ;
        RECT 521.100 500.400 522.900 506.400 ;
        RECT 450.300 483.600 451.200 500.400 ;
        RECT 458.400 497.100 459.900 500.400 ;
        RECT 464.100 498.600 470.700 500.400 ;
        RECT 485.400 499.800 486.300 500.400 ;
        RECT 488.400 499.800 490.200 500.400 ;
        RECT 485.400 498.600 492.600 499.800 ;
        RECT 452.100 495.300 459.900 497.100 ;
        RECT 476.100 496.500 477.900 498.300 ;
        RECT 475.800 495.900 477.900 496.500 ;
        RECT 460.800 494.400 477.900 495.900 ;
        RECT 482.100 495.900 484.200 496.050 ;
        RECT 485.400 495.900 487.200 496.800 ;
        RECT 482.100 495.000 487.200 495.900 ;
        RECT 491.700 495.600 492.600 498.600 ;
        RECT 497.700 499.500 499.200 500.400 ;
        RECT 497.700 498.300 506.100 499.500 ;
        RECT 504.300 497.700 506.100 498.300 ;
        RECT 493.500 496.800 495.600 497.700 ;
        RECT 509.100 496.800 510.300 500.400 ;
        RECT 521.700 498.300 522.900 500.400 ;
        RECT 524.100 501.300 525.900 506.400 ;
        RECT 527.100 502.200 528.900 507.000 ;
        RECT 530.100 501.300 531.900 506.400 ;
        RECT 524.100 499.950 531.900 501.300 ;
        RECT 545.700 499.200 547.500 506.400 ;
        RECT 550.800 500.400 552.600 507.000 ;
        RECT 563.100 503.400 564.900 507.000 ;
        RECT 566.100 503.400 567.900 506.400 ;
        RECT 568.950 504.450 571.050 505.050 ;
        RECT 577.950 504.450 580.050 505.050 ;
        RECT 568.950 503.550 580.050 504.450 ;
        RECT 545.700 498.300 549.900 499.200 ;
        RECT 521.700 497.400 525.300 498.300 ;
        RECT 493.500 495.600 510.300 496.800 ;
        RECT 455.700 492.900 462.300 494.400 ;
        RECT 482.100 493.950 484.200 495.000 ;
        RECT 490.800 493.800 492.600 495.600 ;
        RECT 455.700 490.050 457.200 492.900 ;
        RECT 463.500 491.700 507.900 492.900 ;
        RECT 463.500 490.200 464.400 491.700 ;
        RECT 455.100 487.950 457.200 490.050 ;
        RECT 459.300 488.400 464.400 490.200 ;
        RECT 467.100 489.900 480.600 490.800 ;
        RECT 487.800 489.900 489.600 490.500 ;
        RECT 506.100 490.050 507.900 491.700 ;
        RECT 467.100 488.700 468.000 489.900 ;
        RECT 467.100 486.900 468.900 488.700 ;
        RECT 473.100 487.200 477.000 489.000 ;
        RECT 478.500 488.700 489.600 489.900 ;
        RECT 500.100 489.750 502.200 490.050 ;
        RECT 478.500 487.800 480.600 488.700 ;
        RECT 498.300 487.950 502.200 489.750 ;
        RECT 506.100 487.950 508.200 490.050 ;
        RECT 498.300 487.200 500.100 487.950 ;
        RECT 473.100 486.900 475.200 487.200 ;
        RECT 486.600 486.300 500.100 487.200 ;
        RECT 452.100 485.700 453.900 486.300 ;
        RECT 486.600 485.700 487.800 486.300 ;
        RECT 452.100 484.500 487.800 485.700 ;
        RECT 490.500 484.500 492.600 484.800 ;
        RECT 450.300 482.700 466.800 483.600 ;
        RECT 450.300 479.400 451.200 482.700 ;
        RECT 455.100 480.600 460.800 481.800 ;
        RECT 464.700 481.500 466.800 482.700 ;
        RECT 470.100 482.400 487.800 483.600 ;
        RECT 490.500 483.300 502.500 484.500 ;
        RECT 490.500 482.700 492.600 483.300 ;
        RECT 500.700 482.700 502.500 483.300 ;
        RECT 470.100 481.500 472.200 482.400 ;
        RECT 486.600 481.800 487.800 482.400 ;
        RECT 504.000 481.800 505.800 482.100 ;
        RECT 455.100 480.000 456.900 480.600 ;
        RECT 450.300 478.500 454.200 479.400 ;
        RECT 453.000 477.600 454.200 478.500 ;
        RECT 459.600 477.600 460.800 480.600 ;
        RECT 461.700 479.700 463.500 480.300 ;
        RECT 461.700 478.500 469.800 479.700 ;
        RECT 467.700 477.600 469.800 478.500 ;
        RECT 473.100 477.600 475.800 481.500 ;
        RECT 478.500 479.100 481.800 481.200 ;
        RECT 486.600 480.600 505.800 481.800 ;
        RECT 443.700 471.000 445.500 477.600 ;
        RECT 446.700 471.600 448.500 477.600 ;
        RECT 450.000 471.000 451.800 477.600 ;
        RECT 453.000 471.600 454.800 477.600 ;
        RECT 456.000 471.000 457.800 477.600 ;
        RECT 459.000 471.600 460.800 477.600 ;
        RECT 462.000 471.000 463.800 477.600 ;
        RECT 464.700 474.600 466.800 476.700 ;
        RECT 467.700 474.600 469.800 476.700 ;
        RECT 470.700 474.600 472.800 476.700 ;
        RECT 465.000 471.600 466.800 474.600 ;
        RECT 468.000 471.600 469.800 474.600 ;
        RECT 471.000 471.600 472.800 474.600 ;
        RECT 474.000 471.600 475.800 477.600 ;
        RECT 477.000 471.000 478.800 477.600 ;
        RECT 480.000 471.600 481.800 479.100 ;
        RECT 487.200 477.600 489.300 479.700 ;
        RECT 483.900 471.000 485.700 477.600 ;
        RECT 486.900 471.600 488.700 477.600 ;
        RECT 489.600 474.600 491.700 476.700 ;
        RECT 492.600 474.600 494.700 476.700 ;
        RECT 489.900 471.600 491.700 474.600 ;
        RECT 492.900 471.600 494.700 474.600 ;
        RECT 496.500 471.000 498.300 477.600 ;
        RECT 499.500 471.600 501.300 480.600 ;
        RECT 504.000 480.300 505.800 480.600 ;
        RECT 509.100 479.400 510.300 495.600 ;
        RECT 521.100 493.050 522.900 494.850 ;
        RECT 524.100 493.050 525.300 497.400 ;
        RECT 527.100 493.050 528.900 494.850 ;
        RECT 545.100 493.050 546.900 494.850 ;
        RECT 548.700 493.050 549.900 498.300 ;
        RECT 550.950 493.050 552.750 494.850 ;
        RECT 566.100 493.050 567.300 503.400 ;
        RECT 568.950 502.950 571.050 503.550 ;
        RECT 577.950 502.950 580.050 503.550 ;
        RECT 581.100 498.600 582.900 506.400 ;
        RECT 585.600 500.400 587.400 507.000 ;
        RECT 588.600 502.200 590.400 506.400 ;
        RECT 588.600 500.400 591.300 502.200 ;
        RECT 587.700 498.600 589.500 499.500 ;
        RECT 581.100 497.700 589.500 498.600 ;
        RECT 581.250 493.050 583.050 494.850 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 526.950 490.950 529.050 493.050 ;
        RECT 529.950 490.950 532.050 493.050 ;
        RECT 544.950 490.950 547.050 493.050 ;
        RECT 547.950 490.950 550.050 493.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 581.100 490.950 583.200 493.050 ;
        RECT 524.100 483.600 525.300 490.950 ;
        RECT 530.100 489.150 531.900 490.950 ;
        RECT 524.100 482.100 526.500 483.600 ;
        RECT 506.700 478.500 510.300 479.400 ;
        RECT 522.000 479.100 523.800 480.900 ;
        RECT 506.700 477.600 507.600 478.500 ;
        RECT 502.500 471.000 504.300 477.600 ;
        RECT 505.500 476.700 507.600 477.600 ;
        RECT 505.500 471.600 507.300 476.700 ;
        RECT 508.500 471.000 510.300 477.600 ;
        RECT 521.700 471.000 523.500 477.600 ;
        RECT 524.700 471.600 526.500 482.100 ;
        RECT 529.800 471.000 531.600 483.600 ;
        RECT 532.950 480.450 535.050 481.050 ;
        RECT 544.950 480.450 547.050 481.050 ;
        RECT 532.950 479.550 547.050 480.450 ;
        RECT 532.950 478.950 535.050 479.550 ;
        RECT 544.950 478.950 547.050 479.550 ;
        RECT 548.700 477.600 549.900 490.950 ;
        RECT 563.100 489.150 564.900 490.950 ;
        RECT 566.100 477.600 567.300 490.950 ;
        RECT 574.950 486.450 577.050 490.050 ;
        RECT 580.950 486.450 583.050 486.750 ;
        RECT 574.950 486.000 583.050 486.450 ;
        RECT 575.550 485.550 583.050 486.000 ;
        RECT 580.950 484.650 583.050 485.550 ;
        RECT 584.100 477.600 585.000 497.700 ;
        RECT 590.400 493.050 591.300 500.400 ;
        RECT 605.100 501.300 606.900 506.400 ;
        RECT 608.100 502.200 609.900 507.000 ;
        RECT 611.100 501.300 612.900 506.400 ;
        RECT 605.100 499.950 612.900 501.300 ;
        RECT 614.100 500.400 615.900 506.400 ;
        RECT 629.100 503.400 630.900 507.000 ;
        RECT 632.100 503.400 633.900 506.400 ;
        RECT 635.100 503.400 636.900 507.000 ;
        RECT 614.100 498.300 615.300 500.400 ;
        RECT 611.700 497.400 615.300 498.300 ;
        RECT 608.100 493.050 609.900 494.850 ;
        RECT 611.700 493.050 612.900 497.400 ;
        RECT 614.100 493.050 615.900 494.850 ;
        RECT 632.400 493.050 633.300 503.400 ;
        RECT 647.400 500.400 649.200 507.000 ;
        RECT 652.500 499.200 654.300 506.400 ;
        RECT 650.100 498.300 654.300 499.200 ;
        RECT 668.700 499.200 670.500 506.400 ;
        RECT 673.800 500.400 675.600 507.000 ;
        RECT 686.100 501.300 687.900 506.400 ;
        RECT 689.100 502.200 690.900 507.000 ;
        RECT 692.100 501.300 693.900 506.400 ;
        RECT 686.100 499.950 693.900 501.300 ;
        RECT 695.100 500.400 696.900 506.400 ;
        RECT 707.100 503.400 708.900 506.400 ;
        RECT 710.100 503.400 711.900 507.000 ;
        RECT 668.700 498.300 672.900 499.200 ;
        RECT 695.100 498.300 696.300 500.400 ;
        RECT 647.250 493.050 649.050 494.850 ;
        RECT 650.100 493.050 651.300 498.300 ;
        RECT 663.000 495.450 667.050 496.050 ;
        RECT 653.100 493.050 654.900 494.850 ;
        RECT 662.550 493.950 667.050 495.450 ;
        RECT 586.500 490.950 588.600 493.050 ;
        RECT 589.800 490.950 591.900 493.050 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 646.950 490.950 649.050 493.050 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 586.200 489.150 588.000 490.950 ;
        RECT 590.400 483.600 591.300 490.950 ;
        RECT 605.100 489.150 606.900 490.950 ;
        RECT 611.700 483.600 612.900 490.950 ;
        RECT 629.250 489.150 631.050 490.950 ;
        RECT 632.400 483.600 633.300 490.950 ;
        RECT 635.100 489.150 636.900 490.950 ;
        RECT 545.100 471.000 546.900 477.600 ;
        RECT 548.100 471.600 549.900 477.600 ;
        RECT 551.100 471.000 552.900 477.600 ;
        RECT 563.100 471.000 564.900 477.600 ;
        RECT 566.100 471.600 567.900 477.600 ;
        RECT 581.100 471.000 582.900 477.600 ;
        RECT 584.100 471.600 585.900 477.600 ;
        RECT 587.100 471.000 588.900 483.000 ;
        RECT 590.100 471.600 591.900 483.600 ;
        RECT 605.400 471.000 607.200 483.600 ;
        RECT 610.500 482.100 612.900 483.600 ;
        RECT 610.500 471.600 612.300 482.100 ;
        RECT 613.200 479.100 615.000 480.900 ;
        RECT 613.500 471.000 615.300 477.600 ;
        RECT 629.100 471.000 630.900 483.600 ;
        RECT 632.400 482.400 636.000 483.600 ;
        RECT 634.200 471.600 636.000 482.400 ;
        RECT 650.100 477.600 651.300 490.950 ;
        RECT 662.550 490.050 663.450 493.950 ;
        RECT 668.100 493.050 669.900 494.850 ;
        RECT 671.700 493.050 672.900 498.300 ;
        RECT 692.700 497.400 696.300 498.300 ;
        RECT 673.950 493.050 675.750 494.850 ;
        RECT 689.100 493.050 690.900 494.850 ;
        RECT 692.700 493.050 693.900 497.400 ;
        RECT 695.100 493.050 696.900 494.850 ;
        RECT 707.700 493.050 708.900 503.400 ;
        RECT 722.100 501.300 723.900 506.400 ;
        RECT 725.100 502.200 726.900 507.000 ;
        RECT 728.100 501.300 729.900 506.400 ;
        RECT 722.100 499.950 729.900 501.300 ;
        RECT 731.100 500.400 732.900 506.400 ;
        RECT 731.100 498.300 732.300 500.400 ;
        RECT 728.700 497.400 732.300 498.300 ;
        RECT 743.100 497.400 744.900 507.000 ;
        RECT 749.700 498.000 751.500 506.400 ;
        RECT 764.700 499.200 766.500 506.400 ;
        RECT 769.800 500.400 771.600 507.000 ;
        RECT 782.400 500.400 784.200 507.000 ;
        RECT 787.500 499.200 789.300 506.400 ;
        RECT 764.700 498.300 768.900 499.200 ;
        RECT 725.100 493.050 726.900 494.850 ;
        RECT 728.700 493.050 729.900 497.400 ;
        RECT 749.700 496.800 753.000 498.000 ;
        RECT 738.000 495.450 742.050 496.050 ;
        RECT 731.100 493.050 732.900 494.850 ;
        RECT 737.550 493.950 742.050 495.450 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 694.950 490.950 697.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 662.550 488.550 667.050 490.050 ;
        RECT 663.000 487.950 667.050 488.550 ;
        RECT 652.950 480.450 655.050 481.050 ;
        RECT 661.950 480.450 664.050 481.050 ;
        RECT 652.950 479.550 664.050 480.450 ;
        RECT 652.950 478.950 655.050 479.550 ;
        RECT 661.950 478.950 664.050 479.550 ;
        RECT 671.700 477.600 672.900 490.950 ;
        RECT 686.100 489.150 687.900 490.950 ;
        RECT 692.700 483.600 693.900 490.950 ;
        RECT 647.100 471.000 648.900 477.600 ;
        RECT 650.100 471.600 651.900 477.600 ;
        RECT 653.100 471.000 654.900 477.600 ;
        RECT 668.100 471.000 669.900 477.600 ;
        RECT 671.100 471.600 672.900 477.600 ;
        RECT 674.100 471.000 675.900 477.600 ;
        RECT 686.400 471.000 688.200 483.600 ;
        RECT 691.500 482.100 693.900 483.600 ;
        RECT 691.500 471.600 693.300 482.100 ;
        RECT 694.200 479.100 696.000 480.900 ;
        RECT 707.700 477.600 708.900 490.950 ;
        RECT 710.100 489.150 711.900 490.950 ;
        RECT 722.100 489.150 723.900 490.950 ;
        RECT 728.700 483.600 729.900 490.950 ;
        RECT 737.550 490.050 738.450 493.950 ;
        RECT 743.100 493.050 744.900 494.850 ;
        RECT 749.100 493.050 750.900 494.850 ;
        RECT 752.100 493.050 753.000 496.800 ;
        RECT 754.950 495.450 759.000 496.050 ;
        RECT 754.950 493.950 759.450 495.450 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 745.950 490.950 748.050 493.050 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 733.950 488.550 738.450 490.050 ;
        RECT 746.100 489.150 747.900 490.950 ;
        RECT 733.950 487.950 738.000 488.550 ;
        RECT 694.500 471.000 696.300 477.600 ;
        RECT 707.100 471.600 708.900 477.600 ;
        RECT 710.100 471.000 711.900 477.600 ;
        RECT 722.400 471.000 724.200 483.600 ;
        RECT 727.500 482.100 729.900 483.600 ;
        RECT 727.500 471.600 729.300 482.100 ;
        RECT 730.200 479.100 732.000 480.900 ;
        RECT 752.100 478.800 753.000 490.950 ;
        RECT 758.550 490.050 759.450 493.950 ;
        RECT 764.100 493.050 765.900 494.850 ;
        RECT 767.700 493.050 768.900 498.300 ;
        RECT 785.100 498.300 789.300 499.200 ;
        RECT 803.100 500.400 804.900 506.400 ;
        RECT 806.100 501.300 807.900 507.000 ;
        RECT 810.300 501.000 812.100 506.400 ;
        RECT 814.800 501.300 816.600 507.000 ;
        RECT 803.100 499.500 804.600 500.400 ;
        RECT 769.950 493.050 771.750 494.850 ;
        RECT 782.250 493.050 784.050 494.850 ;
        RECT 785.100 493.050 786.300 498.300 ;
        RECT 803.100 498.000 807.600 499.500 ;
        RECT 805.500 497.400 807.600 498.000 ;
        RECT 811.200 498.900 812.100 501.000 ;
        RECT 818.100 500.400 819.900 506.400 ;
        RECT 815.400 499.500 819.900 500.400 ;
        RECT 833.100 501.300 834.900 506.400 ;
        RECT 836.100 502.200 837.900 507.000 ;
        RECT 839.100 501.300 840.900 506.400 ;
        RECT 833.100 499.950 840.900 501.300 ;
        RECT 842.100 500.400 843.900 506.400 ;
        RECT 798.000 495.450 802.050 496.050 ;
        RECT 808.500 495.900 810.300 497.700 ;
        RECT 811.200 496.800 814.200 498.900 ;
        RECT 815.400 497.100 817.500 499.500 ;
        RECT 842.100 498.300 843.300 500.400 ;
        RECT 839.700 497.400 843.300 498.300 ;
        RECT 854.100 497.400 855.900 507.000 ;
        RECT 860.700 498.000 862.500 506.400 ;
        RECT 788.100 493.050 789.900 494.850 ;
        RECT 797.550 493.950 802.050 495.450 ;
        RECT 807.900 495.000 810.000 495.900 ;
        RECT 763.950 490.950 766.050 493.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 797.550 492.450 798.450 493.950 ;
        RECT 803.400 493.800 810.000 495.000 ;
        RECT 803.400 493.200 805.200 493.800 ;
        RECT 794.550 491.550 798.450 492.450 ;
        RECT 758.550 488.550 763.050 490.050 ;
        RECT 759.000 487.950 763.050 488.550 ;
        RECT 754.950 486.450 757.050 487.050 ;
        RECT 763.950 486.450 766.050 487.050 ;
        RECT 754.950 485.550 766.050 486.450 ;
        RECT 754.950 484.950 757.050 485.550 ;
        RECT 763.950 484.950 766.050 485.550 ;
        RECT 746.400 477.900 753.000 478.800 ;
        RECT 746.400 477.600 747.900 477.900 ;
        RECT 730.500 471.000 732.300 477.600 ;
        RECT 743.100 471.000 744.900 477.600 ;
        RECT 746.100 471.600 747.900 477.600 ;
        RECT 752.100 477.600 753.000 477.900 ;
        RECT 767.700 477.600 768.900 490.950 ;
        RECT 785.100 477.600 786.300 490.950 ;
        RECT 794.550 490.050 795.450 491.550 ;
        RECT 803.100 490.950 805.200 493.200 ;
        RECT 790.950 488.550 795.450 490.050 ;
        RECT 807.900 490.800 810.000 492.900 ;
        RECT 807.900 489.000 809.700 490.800 ;
        RECT 811.200 490.050 812.100 496.800 ;
        RECT 813.000 492.900 815.100 495.000 ;
        RECT 836.100 493.050 837.900 494.850 ;
        RECT 839.700 493.050 840.900 497.400 ;
        RECT 860.700 496.800 864.000 498.000 ;
        RECT 878.100 497.400 879.900 507.000 ;
        RECT 884.700 498.000 886.500 506.400 ;
        RECT 899.100 500.400 900.900 506.400 ;
        RECT 899.700 498.300 900.900 500.400 ;
        RECT 902.100 501.300 903.900 506.400 ;
        RECT 905.100 502.200 906.900 507.000 ;
        RECT 908.100 501.300 909.900 506.400 ;
        RECT 902.100 499.950 909.900 501.300 ;
        RECT 920.100 501.300 921.900 506.400 ;
        RECT 923.100 502.200 924.900 507.000 ;
        RECT 926.100 501.300 927.900 506.400 ;
        RECT 920.100 499.950 927.900 501.300 ;
        RECT 929.100 500.400 930.900 506.400 ;
        RECT 929.100 498.300 930.300 500.400 ;
        RECT 884.700 496.800 888.000 498.000 ;
        RECT 899.700 497.400 903.300 498.300 ;
        RECT 842.100 493.050 843.900 494.850 ;
        RECT 854.100 493.050 855.900 494.850 ;
        RECT 860.100 493.050 861.900 494.850 ;
        RECT 863.100 493.050 864.000 496.800 ;
        RECT 878.100 493.050 879.900 494.850 ;
        RECT 884.100 493.050 885.900 494.850 ;
        RECT 887.100 493.050 888.000 496.800 ;
        RECT 899.100 493.050 900.900 494.850 ;
        RECT 902.100 493.050 903.300 497.400 ;
        RECT 926.700 497.400 930.300 498.300 ;
        RECT 905.100 493.050 906.900 494.850 ;
        RECT 923.100 493.050 924.900 494.850 ;
        RECT 926.700 493.050 927.900 497.400 ;
        RECT 929.100 493.050 930.900 494.850 ;
        RECT 813.000 491.100 814.800 492.900 ;
        RECT 817.800 490.950 819.900 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 898.950 490.950 901.050 493.050 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 904.950 490.950 907.050 493.050 ;
        RECT 907.950 490.950 910.050 493.050 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 922.950 490.950 925.050 493.050 ;
        RECT 925.950 490.950 928.050 493.050 ;
        RECT 928.950 490.950 931.050 493.050 ;
        RECT 811.200 488.700 814.200 490.050 ;
        RECT 817.800 489.150 819.600 490.950 ;
        RECT 833.100 489.150 834.900 490.950 ;
        RECT 790.950 487.950 795.000 488.550 ;
        RECT 812.100 487.950 814.200 488.700 ;
        RECT 809.400 485.700 811.200 487.500 ;
        RECT 805.800 484.800 811.200 485.700 ;
        RECT 805.800 483.900 807.900 484.800 ;
        RECT 803.100 482.700 807.900 483.900 ;
        RECT 812.700 483.600 813.900 487.950 ;
        RECT 810.600 482.700 813.900 483.600 ;
        RECT 814.800 483.600 816.900 484.500 ;
        RECT 839.700 483.600 840.900 490.950 ;
        RECT 857.100 489.150 858.900 490.950 ;
        RECT 749.100 471.000 750.900 477.000 ;
        RECT 752.100 471.600 753.900 477.600 ;
        RECT 764.100 471.000 765.900 477.600 ;
        RECT 767.100 471.600 768.900 477.600 ;
        RECT 770.100 471.000 771.900 477.600 ;
        RECT 782.100 471.000 783.900 477.600 ;
        RECT 785.100 471.600 786.900 477.600 ;
        RECT 788.100 471.000 789.900 477.600 ;
        RECT 803.100 471.600 804.900 482.700 ;
        RECT 806.100 471.000 807.900 481.500 ;
        RECT 810.600 471.600 812.400 482.700 ;
        RECT 814.800 482.400 819.900 483.600 ;
        RECT 814.800 471.000 816.900 481.500 ;
        RECT 818.100 471.600 819.900 482.400 ;
        RECT 833.400 471.000 835.200 483.600 ;
        RECT 838.500 482.100 840.900 483.600 ;
        RECT 838.500 471.600 840.300 482.100 ;
        RECT 841.200 479.100 843.000 480.900 ;
        RECT 863.100 478.800 864.000 490.950 ;
        RECT 881.100 489.150 882.900 490.950 ;
        RECT 887.100 478.800 888.000 490.950 ;
        RECT 902.100 483.600 903.300 490.950 ;
        RECT 908.100 489.150 909.900 490.950 ;
        RECT 920.100 489.150 921.900 490.950 ;
        RECT 904.950 486.450 907.050 487.050 ;
        RECT 922.950 486.450 925.050 487.050 ;
        RECT 904.950 485.550 925.050 486.450 ;
        RECT 904.950 484.950 907.050 485.550 ;
        RECT 922.950 484.950 925.050 485.550 ;
        RECT 926.700 483.600 927.900 490.950 ;
        RECT 902.100 482.100 904.500 483.600 ;
        RECT 900.000 479.100 901.800 480.900 ;
        RECT 857.400 477.900 864.000 478.800 ;
        RECT 857.400 477.600 858.900 477.900 ;
        RECT 841.500 471.000 843.300 477.600 ;
        RECT 854.100 471.000 855.900 477.600 ;
        RECT 857.100 471.600 858.900 477.600 ;
        RECT 863.100 477.600 864.000 477.900 ;
        RECT 881.400 477.900 888.000 478.800 ;
        RECT 881.400 477.600 882.900 477.900 ;
        RECT 860.100 471.000 861.900 477.000 ;
        RECT 863.100 471.600 864.900 477.600 ;
        RECT 878.100 471.000 879.900 477.600 ;
        RECT 881.100 471.600 882.900 477.600 ;
        RECT 887.100 477.600 888.000 477.900 ;
        RECT 884.100 471.000 885.900 477.000 ;
        RECT 887.100 471.600 888.900 477.600 ;
        RECT 899.700 471.000 901.500 477.600 ;
        RECT 902.700 471.600 904.500 482.100 ;
        RECT 907.800 471.000 909.600 483.600 ;
        RECT 920.400 471.000 922.200 483.600 ;
        RECT 925.500 482.100 927.900 483.600 ;
        RECT 925.500 471.600 927.300 482.100 ;
        RECT 928.200 479.100 930.000 480.900 ;
        RECT 928.500 471.000 930.300 477.600 ;
        RECT 14.100 461.400 15.900 467.400 ;
        RECT 17.100 461.400 18.900 468.000 ;
        RECT 20.700 461.400 22.500 468.000 ;
        RECT 23.700 461.400 25.500 467.400 ;
        RECT 27.000 461.400 28.800 468.000 ;
        RECT 30.000 461.400 31.800 467.400 ;
        RECT 33.000 461.400 34.800 468.000 ;
        RECT 36.000 461.400 37.800 467.400 ;
        RECT 39.000 461.400 40.800 468.000 ;
        RECT 42.000 464.400 43.800 467.400 ;
        RECT 45.000 464.400 46.800 467.400 ;
        RECT 48.000 464.400 49.800 467.400 ;
        RECT 41.700 462.300 43.800 464.400 ;
        RECT 44.700 462.300 46.800 464.400 ;
        RECT 47.700 462.300 49.800 464.400 ;
        RECT 51.000 461.400 52.800 467.400 ;
        RECT 54.000 461.400 55.800 468.000 ;
        RECT 14.700 448.050 15.900 461.400 ;
        RECT 24.000 451.050 25.500 461.400 ;
        RECT 30.000 460.500 31.200 461.400 ;
        RECT 17.100 448.050 18.900 449.850 ;
        RECT 23.100 448.950 25.500 451.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 14.700 435.600 15.900 445.950 ;
        RECT 24.000 435.600 25.500 448.950 ;
        RECT 14.100 432.600 15.900 435.600 ;
        RECT 17.100 432.000 18.900 435.600 ;
        RECT 20.700 432.000 22.500 435.600 ;
        RECT 23.700 432.600 25.500 435.600 ;
        RECT 27.300 459.600 31.200 460.500 ;
        RECT 27.300 456.300 28.200 459.600 ;
        RECT 32.100 458.400 33.900 459.000 ;
        RECT 36.600 458.400 37.800 461.400 ;
        RECT 44.700 460.500 46.800 461.400 ;
        RECT 38.700 459.300 46.800 460.500 ;
        RECT 38.700 458.700 40.500 459.300 ;
        RECT 32.100 457.200 37.800 458.400 ;
        RECT 50.100 457.500 52.800 461.400 ;
        RECT 57.000 459.900 58.800 467.400 ;
        RECT 60.900 461.400 62.700 468.000 ;
        RECT 63.900 461.400 65.700 467.400 ;
        RECT 66.900 464.400 68.700 467.400 ;
        RECT 69.900 464.400 71.700 467.400 ;
        RECT 66.600 462.300 68.700 464.400 ;
        RECT 69.600 462.300 71.700 464.400 ;
        RECT 73.500 461.400 75.300 468.000 ;
        RECT 55.500 457.800 58.800 459.900 ;
        RECT 64.200 459.300 66.300 461.400 ;
        RECT 76.500 458.400 78.300 467.400 ;
        RECT 79.500 461.400 81.300 468.000 ;
        RECT 82.500 462.300 84.300 467.400 ;
        RECT 82.500 461.400 84.600 462.300 ;
        RECT 85.500 461.400 87.300 468.000 ;
        RECT 83.700 460.500 84.600 461.400 ;
        RECT 83.700 459.600 87.300 460.500 ;
        RECT 81.000 458.400 82.800 458.700 ;
        RECT 41.700 456.300 43.800 457.500 ;
        RECT 27.300 455.400 43.800 456.300 ;
        RECT 47.100 456.600 49.200 457.500 ;
        RECT 63.600 457.200 82.800 458.400 ;
        RECT 63.600 456.600 64.800 457.200 ;
        RECT 81.000 456.900 82.800 457.200 ;
        RECT 47.100 455.400 64.800 456.600 ;
        RECT 67.500 455.700 69.600 456.300 ;
        RECT 77.700 455.700 79.500 456.300 ;
        RECT 27.300 438.600 28.200 455.400 ;
        RECT 67.500 454.500 79.500 455.700 ;
        RECT 29.100 453.300 64.800 454.500 ;
        RECT 67.500 454.200 69.600 454.500 ;
        RECT 29.100 452.700 30.900 453.300 ;
        RECT 63.600 452.700 64.800 453.300 ;
        RECT 32.100 448.950 34.200 451.050 ;
        RECT 32.700 446.100 34.200 448.950 ;
        RECT 36.300 448.800 41.400 450.600 ;
        RECT 40.500 447.300 41.400 448.800 ;
        RECT 44.100 450.300 45.900 452.100 ;
        RECT 50.100 451.800 52.200 452.100 ;
        RECT 63.600 451.800 77.100 452.700 ;
        RECT 44.100 449.100 45.000 450.300 ;
        RECT 50.100 450.000 54.000 451.800 ;
        RECT 55.500 450.300 57.600 451.200 ;
        RECT 75.300 451.050 77.100 451.800 ;
        RECT 55.500 449.100 66.600 450.300 ;
        RECT 75.300 449.250 79.200 451.050 ;
        RECT 44.100 448.200 57.600 449.100 ;
        RECT 64.800 448.500 66.600 449.100 ;
        RECT 77.100 448.950 79.200 449.250 ;
        RECT 83.100 448.950 85.200 451.050 ;
        RECT 83.100 447.300 84.900 448.950 ;
        RECT 40.500 446.100 84.900 447.300 ;
        RECT 32.700 444.600 39.300 446.100 ;
        RECT 29.100 441.900 36.900 443.700 ;
        RECT 37.800 443.100 54.900 444.600 ;
        RECT 52.800 442.500 54.900 443.100 ;
        RECT 59.100 444.000 61.200 445.050 ;
        RECT 59.100 443.100 64.200 444.000 ;
        RECT 67.800 443.400 69.600 445.200 ;
        RECT 86.100 443.400 87.300 459.600 ;
        RECT 98.400 455.400 100.200 468.000 ;
        RECT 103.500 456.900 105.300 467.400 ;
        RECT 106.500 461.400 108.300 468.000 ;
        RECT 122.100 461.400 123.900 468.000 ;
        RECT 125.100 461.400 126.900 467.400 ;
        RECT 128.100 461.400 129.900 468.000 ;
        RECT 131.700 461.400 133.500 468.000 ;
        RECT 134.700 462.300 136.500 467.400 ;
        RECT 134.400 461.400 136.500 462.300 ;
        RECT 137.700 461.400 139.500 468.000 ;
        RECT 106.200 458.100 108.000 459.900 ;
        RECT 103.500 455.400 105.900 456.900 ;
        RECT 98.100 448.050 99.900 449.850 ;
        RECT 104.700 448.050 105.900 455.400 ;
        RECT 106.950 453.450 109.050 454.050 ;
        RECT 106.950 452.550 117.450 453.450 ;
        RECT 106.950 451.950 109.050 452.550 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 101.100 444.150 102.900 445.950 ;
        RECT 59.100 442.950 61.200 443.100 ;
        RECT 35.400 438.600 36.900 441.900 ;
        RECT 53.100 440.700 54.900 442.500 ;
        RECT 62.400 442.200 64.200 443.100 ;
        RECT 68.700 440.400 69.600 443.400 ;
        RECT 70.500 442.200 87.300 443.400 ;
        RECT 70.500 441.300 72.600 442.200 ;
        RECT 81.300 440.700 83.100 441.300 ;
        RECT 41.100 438.600 47.700 440.400 ;
        RECT 62.400 439.200 69.600 440.400 ;
        RECT 74.700 439.500 83.100 440.700 ;
        RECT 62.400 438.600 63.300 439.200 ;
        RECT 65.400 438.600 67.200 439.200 ;
        RECT 74.700 438.600 76.200 439.500 ;
        RECT 86.100 438.600 87.300 442.200 ;
        RECT 104.700 441.600 105.900 445.950 ;
        RECT 107.100 444.150 108.900 445.950 ;
        RECT 116.550 445.050 117.450 452.550 ;
        RECT 125.100 448.050 126.300 461.400 ;
        RECT 134.400 460.500 135.300 461.400 ;
        RECT 131.700 459.600 135.300 460.500 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 127.950 445.950 130.050 448.050 ;
        RECT 116.550 443.550 121.050 445.050 ;
        RECT 122.250 444.150 124.050 445.950 ;
        RECT 117.000 442.950 121.050 443.550 ;
        RECT 104.700 440.700 108.300 441.600 ;
        RECT 27.300 432.600 29.100 438.600 ;
        RECT 32.700 432.000 34.500 438.600 ;
        RECT 35.400 437.400 39.600 438.600 ;
        RECT 37.800 432.600 39.600 437.400 ;
        RECT 41.700 435.600 43.800 437.700 ;
        RECT 44.700 435.600 46.800 437.700 ;
        RECT 47.700 435.600 49.800 437.700 ;
        RECT 50.700 435.600 52.800 437.700 ;
        RECT 56.100 436.500 58.800 438.600 ;
        RECT 60.600 437.400 63.300 438.600 ;
        RECT 60.600 436.500 62.400 437.400 ;
        RECT 42.000 432.600 43.800 435.600 ;
        RECT 45.000 432.600 46.800 435.600 ;
        RECT 48.000 432.600 49.800 435.600 ;
        RECT 51.000 432.600 52.800 435.600 ;
        RECT 54.000 432.000 55.800 435.600 ;
        RECT 57.000 432.600 58.800 436.500 ;
        RECT 64.200 435.600 66.300 437.700 ;
        RECT 67.200 435.600 69.300 437.700 ;
        RECT 70.200 435.600 72.300 437.700 ;
        RECT 61.500 432.000 63.300 435.600 ;
        RECT 64.500 432.600 66.300 435.600 ;
        RECT 67.500 432.600 69.300 435.600 ;
        RECT 70.500 432.600 72.300 435.600 ;
        RECT 74.700 432.600 76.500 438.600 ;
        RECT 80.100 432.000 81.900 438.600 ;
        RECT 85.500 432.600 87.300 438.600 ;
        RECT 98.100 437.700 105.900 439.050 ;
        RECT 98.100 432.600 99.900 437.700 ;
        RECT 101.100 432.000 102.900 436.800 ;
        RECT 104.100 432.600 105.900 437.700 ;
        RECT 107.100 438.600 108.300 440.700 ;
        RECT 125.100 440.700 126.300 445.950 ;
        RECT 128.100 444.150 129.900 445.950 ;
        RECT 131.700 443.400 132.900 459.600 ;
        RECT 136.200 458.400 138.000 458.700 ;
        RECT 140.700 458.400 142.500 467.400 ;
        RECT 143.700 461.400 145.500 468.000 ;
        RECT 147.300 464.400 149.100 467.400 ;
        RECT 150.300 464.400 152.100 467.400 ;
        RECT 147.300 462.300 149.400 464.400 ;
        RECT 150.300 462.300 152.400 464.400 ;
        RECT 153.300 461.400 155.100 467.400 ;
        RECT 156.300 461.400 158.100 468.000 ;
        RECT 152.700 459.300 154.800 461.400 ;
        RECT 160.200 459.900 162.000 467.400 ;
        RECT 163.200 461.400 165.000 468.000 ;
        RECT 166.200 461.400 168.000 467.400 ;
        RECT 169.200 464.400 171.000 467.400 ;
        RECT 172.200 464.400 174.000 467.400 ;
        RECT 175.200 464.400 177.000 467.400 ;
        RECT 169.200 462.300 171.300 464.400 ;
        RECT 172.200 462.300 174.300 464.400 ;
        RECT 175.200 462.300 177.300 464.400 ;
        RECT 178.200 461.400 180.000 468.000 ;
        RECT 181.200 461.400 183.000 467.400 ;
        RECT 184.200 461.400 186.000 468.000 ;
        RECT 187.200 461.400 189.000 467.400 ;
        RECT 190.200 461.400 192.000 468.000 ;
        RECT 193.500 461.400 195.300 467.400 ;
        RECT 196.500 461.400 198.300 468.000 ;
        RECT 200.700 461.400 202.500 468.000 ;
        RECT 203.700 461.400 205.500 467.400 ;
        RECT 207.000 461.400 208.800 468.000 ;
        RECT 210.000 461.400 211.800 467.400 ;
        RECT 213.000 461.400 214.800 468.000 ;
        RECT 216.000 461.400 217.800 467.400 ;
        RECT 219.000 461.400 220.800 468.000 ;
        RECT 222.000 464.400 223.800 467.400 ;
        RECT 225.000 464.400 226.800 467.400 ;
        RECT 228.000 464.400 229.800 467.400 ;
        RECT 221.700 462.300 223.800 464.400 ;
        RECT 224.700 462.300 226.800 464.400 ;
        RECT 227.700 462.300 229.800 464.400 ;
        RECT 231.000 461.400 232.800 467.400 ;
        RECT 234.000 461.400 235.800 468.000 ;
        RECT 136.200 457.200 155.400 458.400 ;
        RECT 160.200 457.800 163.500 459.900 ;
        RECT 166.200 457.500 168.900 461.400 ;
        RECT 172.200 460.500 174.300 461.400 ;
        RECT 172.200 459.300 180.300 460.500 ;
        RECT 178.500 458.700 180.300 459.300 ;
        RECT 181.200 458.400 182.400 461.400 ;
        RECT 187.800 460.500 189.000 461.400 ;
        RECT 187.800 459.600 191.700 460.500 ;
        RECT 185.100 458.400 186.900 459.000 ;
        RECT 136.200 456.900 138.000 457.200 ;
        RECT 154.200 456.600 155.400 457.200 ;
        RECT 169.800 456.600 171.900 457.500 ;
        RECT 139.500 455.700 141.300 456.300 ;
        RECT 149.400 455.700 151.500 456.300 ;
        RECT 139.500 454.500 151.500 455.700 ;
        RECT 154.200 455.400 171.900 456.600 ;
        RECT 175.200 456.300 177.300 457.500 ;
        RECT 181.200 457.200 186.900 458.400 ;
        RECT 190.800 456.300 191.700 459.600 ;
        RECT 175.200 455.400 191.700 456.300 ;
        RECT 149.400 454.200 151.500 454.500 ;
        RECT 154.200 453.300 189.900 454.500 ;
        RECT 154.200 452.700 155.400 453.300 ;
        RECT 188.100 452.700 189.900 453.300 ;
        RECT 141.900 451.800 155.400 452.700 ;
        RECT 166.800 451.800 168.900 452.100 ;
        RECT 141.900 451.050 143.700 451.800 ;
        RECT 133.800 448.950 135.900 451.050 ;
        RECT 139.800 449.250 143.700 451.050 ;
        RECT 161.400 450.300 163.500 451.200 ;
        RECT 139.800 448.950 141.900 449.250 ;
        RECT 152.400 449.100 163.500 450.300 ;
        RECT 165.000 450.000 168.900 451.800 ;
        RECT 173.100 450.300 174.900 452.100 ;
        RECT 174.000 449.100 174.900 450.300 ;
        RECT 134.100 447.300 135.900 448.950 ;
        RECT 152.400 448.500 154.200 449.100 ;
        RECT 161.400 448.200 174.900 449.100 ;
        RECT 177.600 448.800 182.700 450.600 ;
        RECT 184.800 448.950 186.900 451.050 ;
        RECT 177.600 447.300 178.500 448.800 ;
        RECT 134.100 446.100 178.500 447.300 ;
        RECT 184.800 446.100 186.300 448.950 ;
        RECT 149.400 443.400 151.200 445.200 ;
        RECT 157.800 444.000 159.900 445.050 ;
        RECT 179.700 444.600 186.300 446.100 ;
        RECT 131.700 442.200 148.500 443.400 ;
        RECT 125.100 439.800 129.300 440.700 ;
        RECT 107.100 432.600 108.900 438.600 ;
        RECT 122.400 432.000 124.200 438.600 ;
        RECT 127.500 432.600 129.300 439.800 ;
        RECT 131.700 438.600 132.900 442.200 ;
        RECT 146.400 441.300 148.500 442.200 ;
        RECT 135.900 440.700 137.700 441.300 ;
        RECT 135.900 439.500 144.300 440.700 ;
        RECT 142.800 438.600 144.300 439.500 ;
        RECT 149.400 440.400 150.300 443.400 ;
        RECT 154.800 443.100 159.900 444.000 ;
        RECT 154.800 442.200 156.600 443.100 ;
        RECT 157.800 442.950 159.900 443.100 ;
        RECT 164.100 443.100 181.200 444.600 ;
        RECT 164.100 442.500 166.200 443.100 ;
        RECT 164.100 440.700 165.900 442.500 ;
        RECT 182.100 441.900 189.900 443.700 ;
        RECT 149.400 439.200 156.600 440.400 ;
        RECT 151.800 438.600 153.600 439.200 ;
        RECT 155.700 438.600 156.600 439.200 ;
        RECT 171.300 438.600 177.900 440.400 ;
        RECT 182.100 438.600 183.600 441.900 ;
        RECT 190.800 438.600 191.700 455.400 ;
        RECT 131.700 432.600 133.500 438.600 ;
        RECT 137.100 432.000 138.900 438.600 ;
        RECT 142.500 432.600 144.300 438.600 ;
        RECT 146.700 435.600 148.800 437.700 ;
        RECT 149.700 435.600 151.800 437.700 ;
        RECT 152.700 435.600 154.800 437.700 ;
        RECT 155.700 437.400 158.400 438.600 ;
        RECT 156.600 436.500 158.400 437.400 ;
        RECT 160.200 436.500 162.900 438.600 ;
        RECT 146.700 432.600 148.500 435.600 ;
        RECT 149.700 432.600 151.500 435.600 ;
        RECT 152.700 432.600 154.500 435.600 ;
        RECT 155.700 432.000 157.500 435.600 ;
        RECT 160.200 432.600 162.000 436.500 ;
        RECT 166.200 435.600 168.300 437.700 ;
        RECT 169.200 435.600 171.300 437.700 ;
        RECT 172.200 435.600 174.300 437.700 ;
        RECT 175.200 435.600 177.300 437.700 ;
        RECT 179.400 437.400 183.600 438.600 ;
        RECT 163.200 432.000 165.000 435.600 ;
        RECT 166.200 432.600 168.000 435.600 ;
        RECT 169.200 432.600 171.000 435.600 ;
        RECT 172.200 432.600 174.000 435.600 ;
        RECT 175.200 432.600 177.000 435.600 ;
        RECT 179.400 432.600 181.200 437.400 ;
        RECT 184.500 432.000 186.300 438.600 ;
        RECT 189.900 432.600 191.700 438.600 ;
        RECT 193.500 451.050 195.000 461.400 ;
        RECT 204.000 451.050 205.500 461.400 ;
        RECT 210.000 460.500 211.200 461.400 ;
        RECT 193.500 448.950 195.900 451.050 ;
        RECT 203.100 448.950 205.500 451.050 ;
        RECT 193.500 435.600 195.000 448.950 ;
        RECT 204.000 435.600 205.500 448.950 ;
        RECT 193.500 432.600 195.300 435.600 ;
        RECT 196.500 432.000 198.300 435.600 ;
        RECT 200.700 432.000 202.500 435.600 ;
        RECT 203.700 432.600 205.500 435.600 ;
        RECT 207.300 459.600 211.200 460.500 ;
        RECT 207.300 456.300 208.200 459.600 ;
        RECT 212.100 458.400 213.900 459.000 ;
        RECT 216.600 458.400 217.800 461.400 ;
        RECT 224.700 460.500 226.800 461.400 ;
        RECT 218.700 459.300 226.800 460.500 ;
        RECT 218.700 458.700 220.500 459.300 ;
        RECT 212.100 457.200 217.800 458.400 ;
        RECT 230.100 457.500 232.800 461.400 ;
        RECT 237.000 459.900 238.800 467.400 ;
        RECT 240.900 461.400 242.700 468.000 ;
        RECT 243.900 461.400 245.700 467.400 ;
        RECT 246.900 464.400 248.700 467.400 ;
        RECT 249.900 464.400 251.700 467.400 ;
        RECT 246.600 462.300 248.700 464.400 ;
        RECT 249.600 462.300 251.700 464.400 ;
        RECT 253.500 461.400 255.300 468.000 ;
        RECT 235.500 457.800 238.800 459.900 ;
        RECT 244.200 459.300 246.300 461.400 ;
        RECT 256.500 458.400 258.300 467.400 ;
        RECT 259.500 461.400 261.300 468.000 ;
        RECT 262.500 462.300 264.300 467.400 ;
        RECT 262.500 461.400 264.600 462.300 ;
        RECT 265.500 461.400 267.300 468.000 ;
        RECT 269.700 461.400 271.500 468.000 ;
        RECT 272.700 462.300 274.500 467.400 ;
        RECT 272.400 461.400 274.500 462.300 ;
        RECT 275.700 461.400 277.500 468.000 ;
        RECT 263.700 460.500 264.600 461.400 ;
        RECT 272.400 460.500 273.300 461.400 ;
        RECT 263.700 459.600 267.300 460.500 ;
        RECT 261.000 458.400 262.800 458.700 ;
        RECT 221.700 456.300 223.800 457.500 ;
        RECT 207.300 455.400 223.800 456.300 ;
        RECT 227.100 456.600 229.200 457.500 ;
        RECT 243.600 457.200 262.800 458.400 ;
        RECT 243.600 456.600 244.800 457.200 ;
        RECT 261.000 456.900 262.800 457.200 ;
        RECT 227.100 455.400 244.800 456.600 ;
        RECT 247.500 455.700 249.600 456.300 ;
        RECT 257.700 455.700 259.500 456.300 ;
        RECT 207.300 438.600 208.200 455.400 ;
        RECT 247.500 454.500 259.500 455.700 ;
        RECT 209.100 453.300 244.800 454.500 ;
        RECT 247.500 454.200 249.600 454.500 ;
        RECT 209.100 452.700 210.900 453.300 ;
        RECT 243.600 452.700 244.800 453.300 ;
        RECT 212.100 448.950 214.200 451.050 ;
        RECT 212.700 446.100 214.200 448.950 ;
        RECT 216.300 448.800 221.400 450.600 ;
        RECT 220.500 447.300 221.400 448.800 ;
        RECT 224.100 450.300 225.900 452.100 ;
        RECT 230.100 451.800 232.200 452.100 ;
        RECT 243.600 451.800 257.100 452.700 ;
        RECT 224.100 449.100 225.000 450.300 ;
        RECT 230.100 450.000 234.000 451.800 ;
        RECT 235.500 450.300 237.600 451.200 ;
        RECT 255.300 451.050 257.100 451.800 ;
        RECT 235.500 449.100 246.600 450.300 ;
        RECT 255.300 449.250 259.200 451.050 ;
        RECT 224.100 448.200 237.600 449.100 ;
        RECT 244.800 448.500 246.600 449.100 ;
        RECT 257.100 448.950 259.200 449.250 ;
        RECT 263.100 448.950 265.200 451.050 ;
        RECT 263.100 447.300 264.900 448.950 ;
        RECT 220.500 446.100 264.900 447.300 ;
        RECT 212.700 444.600 219.300 446.100 ;
        RECT 209.100 441.900 216.900 443.700 ;
        RECT 217.800 443.100 234.900 444.600 ;
        RECT 232.800 442.500 234.900 443.100 ;
        RECT 239.100 444.000 241.200 445.050 ;
        RECT 239.100 443.100 244.200 444.000 ;
        RECT 247.800 443.400 249.600 445.200 ;
        RECT 266.100 443.400 267.300 459.600 ;
        RECT 239.100 442.950 241.200 443.100 ;
        RECT 215.400 438.600 216.900 441.900 ;
        RECT 233.100 440.700 234.900 442.500 ;
        RECT 242.400 442.200 244.200 443.100 ;
        RECT 248.700 440.400 249.600 443.400 ;
        RECT 250.500 442.200 267.300 443.400 ;
        RECT 250.500 441.300 252.600 442.200 ;
        RECT 261.300 440.700 263.100 441.300 ;
        RECT 221.100 438.600 227.700 440.400 ;
        RECT 242.400 439.200 249.600 440.400 ;
        RECT 254.700 439.500 263.100 440.700 ;
        RECT 242.400 438.600 243.300 439.200 ;
        RECT 245.400 438.600 247.200 439.200 ;
        RECT 254.700 438.600 256.200 439.500 ;
        RECT 266.100 438.600 267.300 442.200 ;
        RECT 207.300 432.600 209.100 438.600 ;
        RECT 212.700 432.000 214.500 438.600 ;
        RECT 215.400 437.400 219.600 438.600 ;
        RECT 217.800 432.600 219.600 437.400 ;
        RECT 221.700 435.600 223.800 437.700 ;
        RECT 224.700 435.600 226.800 437.700 ;
        RECT 227.700 435.600 229.800 437.700 ;
        RECT 230.700 435.600 232.800 437.700 ;
        RECT 236.100 436.500 238.800 438.600 ;
        RECT 240.600 437.400 243.300 438.600 ;
        RECT 240.600 436.500 242.400 437.400 ;
        RECT 222.000 432.600 223.800 435.600 ;
        RECT 225.000 432.600 226.800 435.600 ;
        RECT 228.000 432.600 229.800 435.600 ;
        RECT 231.000 432.600 232.800 435.600 ;
        RECT 234.000 432.000 235.800 435.600 ;
        RECT 237.000 432.600 238.800 436.500 ;
        RECT 244.200 435.600 246.300 437.700 ;
        RECT 247.200 435.600 249.300 437.700 ;
        RECT 250.200 435.600 252.300 437.700 ;
        RECT 241.500 432.000 243.300 435.600 ;
        RECT 244.500 432.600 246.300 435.600 ;
        RECT 247.500 432.600 249.300 435.600 ;
        RECT 250.500 432.600 252.300 435.600 ;
        RECT 254.700 432.600 256.500 438.600 ;
        RECT 260.100 432.000 261.900 438.600 ;
        RECT 265.500 432.600 267.300 438.600 ;
        RECT 269.700 459.600 273.300 460.500 ;
        RECT 269.700 443.400 270.900 459.600 ;
        RECT 274.200 458.400 276.000 458.700 ;
        RECT 278.700 458.400 280.500 467.400 ;
        RECT 281.700 461.400 283.500 468.000 ;
        RECT 285.300 464.400 287.100 467.400 ;
        RECT 288.300 464.400 290.100 467.400 ;
        RECT 285.300 462.300 287.400 464.400 ;
        RECT 288.300 462.300 290.400 464.400 ;
        RECT 291.300 461.400 293.100 467.400 ;
        RECT 294.300 461.400 296.100 468.000 ;
        RECT 290.700 459.300 292.800 461.400 ;
        RECT 298.200 459.900 300.000 467.400 ;
        RECT 301.200 461.400 303.000 468.000 ;
        RECT 304.200 461.400 306.000 467.400 ;
        RECT 307.200 464.400 309.000 467.400 ;
        RECT 310.200 464.400 312.000 467.400 ;
        RECT 313.200 464.400 315.000 467.400 ;
        RECT 307.200 462.300 309.300 464.400 ;
        RECT 310.200 462.300 312.300 464.400 ;
        RECT 313.200 462.300 315.300 464.400 ;
        RECT 316.200 461.400 318.000 468.000 ;
        RECT 319.200 461.400 321.000 467.400 ;
        RECT 322.200 461.400 324.000 468.000 ;
        RECT 325.200 461.400 327.000 467.400 ;
        RECT 328.200 461.400 330.000 468.000 ;
        RECT 331.500 461.400 333.300 467.400 ;
        RECT 334.500 461.400 336.300 468.000 ;
        RECT 338.700 461.400 340.500 468.000 ;
        RECT 341.700 462.300 343.500 467.400 ;
        RECT 341.400 461.400 343.500 462.300 ;
        RECT 344.700 461.400 346.500 468.000 ;
        RECT 274.200 457.200 293.400 458.400 ;
        RECT 298.200 457.800 301.500 459.900 ;
        RECT 304.200 457.500 306.900 461.400 ;
        RECT 310.200 460.500 312.300 461.400 ;
        RECT 310.200 459.300 318.300 460.500 ;
        RECT 316.500 458.700 318.300 459.300 ;
        RECT 319.200 458.400 320.400 461.400 ;
        RECT 325.800 460.500 327.000 461.400 ;
        RECT 325.800 459.600 329.700 460.500 ;
        RECT 323.100 458.400 324.900 459.000 ;
        RECT 274.200 456.900 276.000 457.200 ;
        RECT 292.200 456.600 293.400 457.200 ;
        RECT 307.800 456.600 309.900 457.500 ;
        RECT 277.500 455.700 279.300 456.300 ;
        RECT 287.400 455.700 289.500 456.300 ;
        RECT 277.500 454.500 289.500 455.700 ;
        RECT 292.200 455.400 309.900 456.600 ;
        RECT 313.200 456.300 315.300 457.500 ;
        RECT 319.200 457.200 324.900 458.400 ;
        RECT 328.800 456.300 329.700 459.600 ;
        RECT 313.200 455.400 329.700 456.300 ;
        RECT 287.400 454.200 289.500 454.500 ;
        RECT 292.200 453.300 327.900 454.500 ;
        RECT 292.200 452.700 293.400 453.300 ;
        RECT 326.100 452.700 327.900 453.300 ;
        RECT 279.900 451.800 293.400 452.700 ;
        RECT 304.800 451.800 306.900 452.100 ;
        RECT 279.900 451.050 281.700 451.800 ;
        RECT 271.800 448.950 273.900 451.050 ;
        RECT 277.800 449.250 281.700 451.050 ;
        RECT 299.400 450.300 301.500 451.200 ;
        RECT 277.800 448.950 279.900 449.250 ;
        RECT 290.400 449.100 301.500 450.300 ;
        RECT 303.000 450.000 306.900 451.800 ;
        RECT 311.100 450.300 312.900 452.100 ;
        RECT 312.000 449.100 312.900 450.300 ;
        RECT 272.100 447.300 273.900 448.950 ;
        RECT 290.400 448.500 292.200 449.100 ;
        RECT 299.400 448.200 312.900 449.100 ;
        RECT 315.600 448.800 320.700 450.600 ;
        RECT 322.800 448.950 324.900 451.050 ;
        RECT 315.600 447.300 316.500 448.800 ;
        RECT 272.100 446.100 316.500 447.300 ;
        RECT 322.800 446.100 324.300 448.950 ;
        RECT 287.400 443.400 289.200 445.200 ;
        RECT 295.800 444.000 297.900 445.050 ;
        RECT 317.700 444.600 324.300 446.100 ;
        RECT 269.700 442.200 286.500 443.400 ;
        RECT 269.700 438.600 270.900 442.200 ;
        RECT 284.400 441.300 286.500 442.200 ;
        RECT 273.900 440.700 275.700 441.300 ;
        RECT 273.900 439.500 282.300 440.700 ;
        RECT 280.800 438.600 282.300 439.500 ;
        RECT 287.400 440.400 288.300 443.400 ;
        RECT 292.800 443.100 297.900 444.000 ;
        RECT 292.800 442.200 294.600 443.100 ;
        RECT 295.800 442.950 297.900 443.100 ;
        RECT 302.100 443.100 319.200 444.600 ;
        RECT 302.100 442.500 304.200 443.100 ;
        RECT 302.100 440.700 303.900 442.500 ;
        RECT 320.100 441.900 327.900 443.700 ;
        RECT 287.400 439.200 294.600 440.400 ;
        RECT 289.800 438.600 291.600 439.200 ;
        RECT 293.700 438.600 294.600 439.200 ;
        RECT 309.300 438.600 315.900 440.400 ;
        RECT 320.100 438.600 321.600 441.900 ;
        RECT 328.800 438.600 329.700 455.400 ;
        RECT 269.700 432.600 271.500 438.600 ;
        RECT 275.100 432.000 276.900 438.600 ;
        RECT 280.500 432.600 282.300 438.600 ;
        RECT 284.700 435.600 286.800 437.700 ;
        RECT 287.700 435.600 289.800 437.700 ;
        RECT 290.700 435.600 292.800 437.700 ;
        RECT 293.700 437.400 296.400 438.600 ;
        RECT 294.600 436.500 296.400 437.400 ;
        RECT 298.200 436.500 300.900 438.600 ;
        RECT 284.700 432.600 286.500 435.600 ;
        RECT 287.700 432.600 289.500 435.600 ;
        RECT 290.700 432.600 292.500 435.600 ;
        RECT 293.700 432.000 295.500 435.600 ;
        RECT 298.200 432.600 300.000 436.500 ;
        RECT 304.200 435.600 306.300 437.700 ;
        RECT 307.200 435.600 309.300 437.700 ;
        RECT 310.200 435.600 312.300 437.700 ;
        RECT 313.200 435.600 315.300 437.700 ;
        RECT 317.400 437.400 321.600 438.600 ;
        RECT 301.200 432.000 303.000 435.600 ;
        RECT 304.200 432.600 306.000 435.600 ;
        RECT 307.200 432.600 309.000 435.600 ;
        RECT 310.200 432.600 312.000 435.600 ;
        RECT 313.200 432.600 315.000 435.600 ;
        RECT 317.400 432.600 319.200 437.400 ;
        RECT 322.500 432.000 324.300 438.600 ;
        RECT 327.900 432.600 329.700 438.600 ;
        RECT 331.500 451.050 333.000 461.400 ;
        RECT 341.400 460.500 342.300 461.400 ;
        RECT 338.700 459.600 342.300 460.500 ;
        RECT 331.500 448.950 333.900 451.050 ;
        RECT 331.500 435.600 333.000 448.950 ;
        RECT 338.700 443.400 339.900 459.600 ;
        RECT 343.200 458.400 345.000 458.700 ;
        RECT 347.700 458.400 349.500 467.400 ;
        RECT 350.700 461.400 352.500 468.000 ;
        RECT 354.300 464.400 356.100 467.400 ;
        RECT 357.300 464.400 359.100 467.400 ;
        RECT 354.300 462.300 356.400 464.400 ;
        RECT 357.300 462.300 359.400 464.400 ;
        RECT 360.300 461.400 362.100 467.400 ;
        RECT 363.300 461.400 365.100 468.000 ;
        RECT 359.700 459.300 361.800 461.400 ;
        RECT 367.200 459.900 369.000 467.400 ;
        RECT 370.200 461.400 372.000 468.000 ;
        RECT 373.200 461.400 375.000 467.400 ;
        RECT 376.200 464.400 378.000 467.400 ;
        RECT 379.200 464.400 381.000 467.400 ;
        RECT 382.200 464.400 384.000 467.400 ;
        RECT 376.200 462.300 378.300 464.400 ;
        RECT 379.200 462.300 381.300 464.400 ;
        RECT 382.200 462.300 384.300 464.400 ;
        RECT 385.200 461.400 387.000 468.000 ;
        RECT 388.200 461.400 390.000 467.400 ;
        RECT 391.200 461.400 393.000 468.000 ;
        RECT 394.200 461.400 396.000 467.400 ;
        RECT 397.200 461.400 399.000 468.000 ;
        RECT 400.500 461.400 402.300 467.400 ;
        RECT 403.500 461.400 405.300 468.000 ;
        RECT 343.200 457.200 362.400 458.400 ;
        RECT 367.200 457.800 370.500 459.900 ;
        RECT 373.200 457.500 375.900 461.400 ;
        RECT 379.200 460.500 381.300 461.400 ;
        RECT 379.200 459.300 387.300 460.500 ;
        RECT 385.500 458.700 387.300 459.300 ;
        RECT 388.200 458.400 389.400 461.400 ;
        RECT 394.800 460.500 396.000 461.400 ;
        RECT 394.800 459.600 398.700 460.500 ;
        RECT 392.100 458.400 393.900 459.000 ;
        RECT 343.200 456.900 345.000 457.200 ;
        RECT 361.200 456.600 362.400 457.200 ;
        RECT 376.800 456.600 378.900 457.500 ;
        RECT 346.500 455.700 348.300 456.300 ;
        RECT 356.400 455.700 358.500 456.300 ;
        RECT 346.500 454.500 358.500 455.700 ;
        RECT 361.200 455.400 378.900 456.600 ;
        RECT 382.200 456.300 384.300 457.500 ;
        RECT 388.200 457.200 393.900 458.400 ;
        RECT 397.800 456.300 398.700 459.600 ;
        RECT 382.200 455.400 398.700 456.300 ;
        RECT 356.400 454.200 358.500 454.500 ;
        RECT 361.200 453.300 396.900 454.500 ;
        RECT 361.200 452.700 362.400 453.300 ;
        RECT 395.100 452.700 396.900 453.300 ;
        RECT 348.900 451.800 362.400 452.700 ;
        RECT 373.800 451.800 375.900 452.100 ;
        RECT 348.900 451.050 350.700 451.800 ;
        RECT 340.800 448.950 342.900 451.050 ;
        RECT 346.800 449.250 350.700 451.050 ;
        RECT 368.400 450.300 370.500 451.200 ;
        RECT 346.800 448.950 348.900 449.250 ;
        RECT 359.400 449.100 370.500 450.300 ;
        RECT 372.000 450.000 375.900 451.800 ;
        RECT 380.100 450.300 381.900 452.100 ;
        RECT 381.000 449.100 381.900 450.300 ;
        RECT 341.100 447.300 342.900 448.950 ;
        RECT 359.400 448.500 361.200 449.100 ;
        RECT 368.400 448.200 381.900 449.100 ;
        RECT 384.600 448.800 389.700 450.600 ;
        RECT 391.800 448.950 393.900 451.050 ;
        RECT 384.600 447.300 385.500 448.800 ;
        RECT 341.100 446.100 385.500 447.300 ;
        RECT 391.800 446.100 393.300 448.950 ;
        RECT 356.400 443.400 358.200 445.200 ;
        RECT 364.800 444.000 366.900 445.050 ;
        RECT 386.700 444.600 393.300 446.100 ;
        RECT 338.700 442.200 355.500 443.400 ;
        RECT 338.700 438.600 339.900 442.200 ;
        RECT 353.400 441.300 355.500 442.200 ;
        RECT 342.900 440.700 344.700 441.300 ;
        RECT 342.900 439.500 351.300 440.700 ;
        RECT 349.800 438.600 351.300 439.500 ;
        RECT 356.400 440.400 357.300 443.400 ;
        RECT 361.800 443.100 366.900 444.000 ;
        RECT 361.800 442.200 363.600 443.100 ;
        RECT 364.800 442.950 366.900 443.100 ;
        RECT 371.100 443.100 388.200 444.600 ;
        RECT 371.100 442.500 373.200 443.100 ;
        RECT 371.100 440.700 372.900 442.500 ;
        RECT 389.100 441.900 396.900 443.700 ;
        RECT 356.400 439.200 363.600 440.400 ;
        RECT 358.800 438.600 360.600 439.200 ;
        RECT 362.700 438.600 363.600 439.200 ;
        RECT 378.300 438.600 384.900 440.400 ;
        RECT 389.100 438.600 390.600 441.900 ;
        RECT 397.800 438.600 398.700 455.400 ;
        RECT 331.500 432.600 333.300 435.600 ;
        RECT 334.500 432.000 336.300 435.600 ;
        RECT 338.700 432.600 340.500 438.600 ;
        RECT 344.100 432.000 345.900 438.600 ;
        RECT 349.500 432.600 351.300 438.600 ;
        RECT 353.700 435.600 355.800 437.700 ;
        RECT 356.700 435.600 358.800 437.700 ;
        RECT 359.700 435.600 361.800 437.700 ;
        RECT 362.700 437.400 365.400 438.600 ;
        RECT 363.600 436.500 365.400 437.400 ;
        RECT 367.200 436.500 369.900 438.600 ;
        RECT 353.700 432.600 355.500 435.600 ;
        RECT 356.700 432.600 358.500 435.600 ;
        RECT 359.700 432.600 361.500 435.600 ;
        RECT 362.700 432.000 364.500 435.600 ;
        RECT 367.200 432.600 369.000 436.500 ;
        RECT 373.200 435.600 375.300 437.700 ;
        RECT 376.200 435.600 378.300 437.700 ;
        RECT 379.200 435.600 381.300 437.700 ;
        RECT 382.200 435.600 384.300 437.700 ;
        RECT 386.400 437.400 390.600 438.600 ;
        RECT 370.200 432.000 372.000 435.600 ;
        RECT 373.200 432.600 375.000 435.600 ;
        RECT 376.200 432.600 378.000 435.600 ;
        RECT 379.200 432.600 381.000 435.600 ;
        RECT 382.200 432.600 384.000 435.600 ;
        RECT 386.400 432.600 388.200 437.400 ;
        RECT 391.500 432.000 393.300 438.600 ;
        RECT 396.900 432.600 398.700 438.600 ;
        RECT 400.500 451.050 402.000 461.400 ;
        RECT 416.100 455.400 417.900 467.400 ;
        RECT 419.100 457.200 420.900 468.000 ;
        RECT 422.100 461.400 423.900 467.400 ;
        RECT 425.700 461.400 427.500 468.000 ;
        RECT 428.700 461.400 430.500 467.400 ;
        RECT 432.000 461.400 433.800 468.000 ;
        RECT 435.000 461.400 436.800 467.400 ;
        RECT 438.000 461.400 439.800 468.000 ;
        RECT 441.000 461.400 442.800 467.400 ;
        RECT 444.000 461.400 445.800 468.000 ;
        RECT 447.000 464.400 448.800 467.400 ;
        RECT 450.000 464.400 451.800 467.400 ;
        RECT 453.000 464.400 454.800 467.400 ;
        RECT 446.700 462.300 448.800 464.400 ;
        RECT 449.700 462.300 451.800 464.400 ;
        RECT 452.700 462.300 454.800 464.400 ;
        RECT 456.000 461.400 457.800 467.400 ;
        RECT 459.000 461.400 460.800 468.000 ;
        RECT 400.500 448.950 402.900 451.050 ;
        RECT 400.500 435.600 402.000 448.950 ;
        RECT 416.100 448.050 417.300 455.400 ;
        RECT 422.700 454.500 423.900 461.400 ;
        RECT 418.200 453.600 423.900 454.500 ;
        RECT 418.200 452.700 420.000 453.600 ;
        RECT 416.100 445.950 418.200 448.050 ;
        RECT 416.100 438.600 417.300 445.950 ;
        RECT 419.100 441.300 420.000 452.700 ;
        RECT 429.000 451.050 430.500 461.400 ;
        RECT 435.000 460.500 436.200 461.400 ;
        RECT 421.800 448.050 423.600 449.850 ;
        RECT 428.100 448.950 430.500 451.050 ;
        RECT 421.500 445.950 423.600 448.050 ;
        RECT 418.200 440.400 420.000 441.300 ;
        RECT 418.200 439.500 423.900 440.400 ;
        RECT 400.500 432.600 402.300 435.600 ;
        RECT 403.500 432.000 405.300 435.600 ;
        RECT 416.100 432.600 417.900 438.600 ;
        RECT 419.100 432.000 420.900 438.600 ;
        RECT 422.700 435.600 423.900 439.500 ;
        RECT 429.000 435.600 430.500 448.950 ;
        RECT 422.100 432.600 423.900 435.600 ;
        RECT 425.700 432.000 427.500 435.600 ;
        RECT 428.700 432.600 430.500 435.600 ;
        RECT 432.300 459.600 436.200 460.500 ;
        RECT 432.300 456.300 433.200 459.600 ;
        RECT 437.100 458.400 438.900 459.000 ;
        RECT 441.600 458.400 442.800 461.400 ;
        RECT 449.700 460.500 451.800 461.400 ;
        RECT 443.700 459.300 451.800 460.500 ;
        RECT 443.700 458.700 445.500 459.300 ;
        RECT 437.100 457.200 442.800 458.400 ;
        RECT 455.100 457.500 457.800 461.400 ;
        RECT 462.000 459.900 463.800 467.400 ;
        RECT 465.900 461.400 467.700 468.000 ;
        RECT 468.900 461.400 470.700 467.400 ;
        RECT 471.900 464.400 473.700 467.400 ;
        RECT 474.900 464.400 476.700 467.400 ;
        RECT 471.600 462.300 473.700 464.400 ;
        RECT 474.600 462.300 476.700 464.400 ;
        RECT 478.500 461.400 480.300 468.000 ;
        RECT 460.500 457.800 463.800 459.900 ;
        RECT 469.200 459.300 471.300 461.400 ;
        RECT 481.500 458.400 483.300 467.400 ;
        RECT 484.500 461.400 486.300 468.000 ;
        RECT 487.500 462.300 489.300 467.400 ;
        RECT 487.500 461.400 489.600 462.300 ;
        RECT 490.500 461.400 492.300 468.000 ;
        RECT 506.100 461.400 507.900 467.400 ;
        RECT 488.700 460.500 489.600 461.400 ;
        RECT 488.700 459.600 492.300 460.500 ;
        RECT 486.000 458.400 487.800 458.700 ;
        RECT 446.700 456.300 448.800 457.500 ;
        RECT 432.300 455.400 448.800 456.300 ;
        RECT 452.100 456.600 454.200 457.500 ;
        RECT 468.600 457.200 487.800 458.400 ;
        RECT 468.600 456.600 469.800 457.200 ;
        RECT 486.000 456.900 487.800 457.200 ;
        RECT 452.100 455.400 469.800 456.600 ;
        RECT 472.500 455.700 474.600 456.300 ;
        RECT 482.700 455.700 484.500 456.300 ;
        RECT 432.300 438.600 433.200 455.400 ;
        RECT 472.500 454.500 484.500 455.700 ;
        RECT 434.100 453.300 469.800 454.500 ;
        RECT 472.500 454.200 474.600 454.500 ;
        RECT 434.100 452.700 435.900 453.300 ;
        RECT 468.600 452.700 469.800 453.300 ;
        RECT 437.100 448.950 439.200 451.050 ;
        RECT 437.700 446.100 439.200 448.950 ;
        RECT 441.300 448.800 446.400 450.600 ;
        RECT 445.500 447.300 446.400 448.800 ;
        RECT 449.100 450.300 450.900 452.100 ;
        RECT 455.100 451.800 457.200 452.100 ;
        RECT 468.600 451.800 482.100 452.700 ;
        RECT 449.100 449.100 450.000 450.300 ;
        RECT 455.100 450.000 459.000 451.800 ;
        RECT 460.500 450.300 462.600 451.200 ;
        RECT 480.300 451.050 482.100 451.800 ;
        RECT 460.500 449.100 471.600 450.300 ;
        RECT 480.300 449.250 484.200 451.050 ;
        RECT 449.100 448.200 462.600 449.100 ;
        RECT 469.800 448.500 471.600 449.100 ;
        RECT 482.100 448.950 484.200 449.250 ;
        RECT 488.100 448.950 490.200 451.050 ;
        RECT 488.100 447.300 489.900 448.950 ;
        RECT 445.500 446.100 489.900 447.300 ;
        RECT 437.700 444.600 444.300 446.100 ;
        RECT 434.100 441.900 441.900 443.700 ;
        RECT 442.800 443.100 459.900 444.600 ;
        RECT 457.800 442.500 459.900 443.100 ;
        RECT 464.100 444.000 466.200 445.050 ;
        RECT 464.100 443.100 469.200 444.000 ;
        RECT 472.800 443.400 474.600 445.200 ;
        RECT 491.100 443.400 492.300 459.600 ;
        RECT 506.100 454.500 507.300 461.400 ;
        RECT 509.100 457.200 510.900 468.000 ;
        RECT 512.100 455.400 513.900 467.400 ;
        RECT 506.100 453.600 511.800 454.500 ;
        RECT 510.000 452.700 511.800 453.600 ;
        RECT 506.400 448.050 508.200 449.850 ;
        RECT 506.400 445.950 508.500 448.050 ;
        RECT 464.100 442.950 466.200 443.100 ;
        RECT 440.400 438.600 441.900 441.900 ;
        RECT 458.100 440.700 459.900 442.500 ;
        RECT 467.400 442.200 469.200 443.100 ;
        RECT 473.700 440.400 474.600 443.400 ;
        RECT 475.500 442.200 492.300 443.400 ;
        RECT 475.500 441.300 477.600 442.200 ;
        RECT 486.300 440.700 488.100 441.300 ;
        RECT 446.100 438.600 452.700 440.400 ;
        RECT 467.400 439.200 474.600 440.400 ;
        RECT 479.700 439.500 488.100 440.700 ;
        RECT 467.400 438.600 468.300 439.200 ;
        RECT 470.400 438.600 472.200 439.200 ;
        RECT 479.700 438.600 481.200 439.500 ;
        RECT 491.100 438.600 492.300 442.200 ;
        RECT 510.000 441.300 510.900 452.700 ;
        RECT 512.700 448.050 513.900 455.400 ;
        RECT 527.100 461.400 528.900 467.400 ;
        RECT 527.100 454.500 528.300 461.400 ;
        RECT 530.100 457.200 531.900 468.000 ;
        RECT 533.100 455.400 534.900 467.400 ;
        RECT 548.100 461.400 549.900 468.000 ;
        RECT 551.100 461.400 552.900 467.400 ;
        RECT 527.100 453.600 532.800 454.500 ;
        RECT 531.000 452.700 532.800 453.600 ;
        RECT 511.800 445.950 513.900 448.050 ;
        RECT 527.400 448.050 529.200 449.850 ;
        RECT 527.400 445.950 529.500 448.050 ;
        RECT 510.000 440.400 511.800 441.300 ;
        RECT 432.300 432.600 434.100 438.600 ;
        RECT 437.700 432.000 439.500 438.600 ;
        RECT 440.400 437.400 444.600 438.600 ;
        RECT 442.800 432.600 444.600 437.400 ;
        RECT 446.700 435.600 448.800 437.700 ;
        RECT 449.700 435.600 451.800 437.700 ;
        RECT 452.700 435.600 454.800 437.700 ;
        RECT 455.700 435.600 457.800 437.700 ;
        RECT 461.100 436.500 463.800 438.600 ;
        RECT 465.600 437.400 468.300 438.600 ;
        RECT 465.600 436.500 467.400 437.400 ;
        RECT 447.000 432.600 448.800 435.600 ;
        RECT 450.000 432.600 451.800 435.600 ;
        RECT 453.000 432.600 454.800 435.600 ;
        RECT 456.000 432.600 457.800 435.600 ;
        RECT 459.000 432.000 460.800 435.600 ;
        RECT 462.000 432.600 463.800 436.500 ;
        RECT 469.200 435.600 471.300 437.700 ;
        RECT 472.200 435.600 474.300 437.700 ;
        RECT 475.200 435.600 477.300 437.700 ;
        RECT 466.500 432.000 468.300 435.600 ;
        RECT 469.500 432.600 471.300 435.600 ;
        RECT 472.500 432.600 474.300 435.600 ;
        RECT 475.500 432.600 477.300 435.600 ;
        RECT 479.700 432.600 481.500 438.600 ;
        RECT 485.100 432.000 486.900 438.600 ;
        RECT 490.500 432.600 492.300 438.600 ;
        RECT 506.100 439.500 511.800 440.400 ;
        RECT 506.100 435.600 507.300 439.500 ;
        RECT 512.700 438.600 513.900 445.950 ;
        RECT 531.000 441.300 531.900 452.700 ;
        RECT 533.700 448.050 534.900 455.400 ;
        RECT 532.800 445.950 534.900 448.050 ;
        RECT 548.100 445.950 550.200 448.050 ;
        RECT 531.000 440.400 532.800 441.300 ;
        RECT 506.100 432.600 507.900 435.600 ;
        RECT 509.100 432.000 510.900 438.600 ;
        RECT 512.100 432.600 513.900 438.600 ;
        RECT 527.100 439.500 532.800 440.400 ;
        RECT 527.100 435.600 528.300 439.500 ;
        RECT 533.700 438.600 534.900 445.950 ;
        RECT 548.250 444.150 550.050 445.950 ;
        RECT 551.100 441.300 552.000 461.400 ;
        RECT 554.100 456.000 555.900 468.000 ;
        RECT 557.100 455.400 558.900 467.400 ;
        RECT 569.100 461.400 570.900 468.000 ;
        RECT 572.100 461.400 573.900 467.400 ;
        RECT 575.100 461.400 576.900 468.000 ;
        RECT 590.100 461.400 591.900 467.400 ;
        RECT 593.100 461.400 594.900 468.000 ;
        RECT 553.200 448.050 555.000 449.850 ;
        RECT 557.400 448.050 558.300 455.400 ;
        RECT 562.950 453.450 565.050 454.050 ;
        RECT 568.950 453.450 571.050 454.050 ;
        RECT 562.950 452.550 571.050 453.450 ;
        RECT 562.950 451.950 565.050 452.550 ;
        RECT 568.950 451.950 571.050 452.550 ;
        RECT 572.700 448.050 573.900 461.400 ;
        RECT 574.950 459.450 577.050 460.050 ;
        RECT 586.950 459.450 589.050 460.050 ;
        RECT 574.950 458.550 589.050 459.450 ;
        RECT 574.950 457.950 577.050 458.550 ;
        RECT 586.950 457.950 589.050 458.550 ;
        RECT 586.950 450.450 589.050 451.050 ;
        RECT 581.550 449.550 589.050 450.450 ;
        RECT 553.500 445.950 555.600 448.050 ;
        RECT 556.800 445.950 558.900 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 527.100 432.600 528.900 435.600 ;
        RECT 530.100 432.000 531.900 438.600 ;
        RECT 533.100 432.600 534.900 438.600 ;
        RECT 548.100 440.400 556.500 441.300 ;
        RECT 548.100 432.600 549.900 440.400 ;
        RECT 554.700 439.500 556.500 440.400 ;
        RECT 557.400 438.600 558.300 445.950 ;
        RECT 569.100 444.150 570.900 445.950 ;
        RECT 572.700 440.700 573.900 445.950 ;
        RECT 574.950 444.150 576.750 445.950 ;
        RECT 581.550 445.050 582.450 449.550 ;
        RECT 586.950 448.950 589.050 449.550 ;
        RECT 590.700 448.050 591.900 461.400 ;
        RECT 608.100 456.600 609.900 467.400 ;
        RECT 611.100 457.500 612.900 468.000 ;
        RECT 614.100 466.500 621.900 467.400 ;
        RECT 614.100 456.600 615.900 466.500 ;
        RECT 608.100 455.700 615.900 456.600 ;
        RECT 617.100 454.500 618.900 465.600 ;
        RECT 620.100 455.400 621.900 466.500 ;
        RECT 632.100 461.400 633.900 468.000 ;
        RECT 635.100 461.400 636.900 467.400 ;
        RECT 638.100 462.000 639.900 468.000 ;
        RECT 635.400 461.100 636.900 461.400 ;
        RECT 641.100 461.400 642.900 467.400 ;
        RECT 641.100 461.100 642.000 461.400 ;
        RECT 635.400 460.200 642.000 461.100 ;
        RECT 614.100 453.600 618.900 454.500 ;
        RECT 593.100 448.050 594.900 449.850 ;
        RECT 611.250 448.050 613.050 449.850 ;
        RECT 614.100 448.050 615.000 453.600 ;
        RECT 617.100 448.050 618.900 449.850 ;
        RECT 635.100 448.050 636.900 449.850 ;
        RECT 641.100 448.050 642.000 460.200 ;
        RECT 656.400 455.400 658.200 468.000 ;
        RECT 661.500 456.900 663.300 467.400 ;
        RECT 664.500 461.400 666.300 468.000 ;
        RECT 680.100 461.400 681.900 468.000 ;
        RECT 683.100 461.400 684.900 467.400 ;
        RECT 664.200 458.100 666.000 459.900 ;
        RECT 661.500 455.400 663.900 456.900 ;
        RECT 651.000 450.450 655.050 451.050 ;
        RECT 650.550 448.950 655.050 450.450 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 577.950 443.550 582.450 445.050 ;
        RECT 577.950 442.950 582.000 443.550 ;
        RECT 552.600 432.000 554.400 438.600 ;
        RECT 555.600 436.800 558.300 438.600 ;
        RECT 569.700 439.800 573.900 440.700 ;
        RECT 555.600 432.600 557.400 436.800 ;
        RECT 569.700 432.600 571.500 439.800 ;
        RECT 574.800 432.000 576.600 438.600 ;
        RECT 590.700 435.600 591.900 445.950 ;
        RECT 608.250 444.150 610.050 445.950 ;
        RECT 601.950 441.450 604.050 442.050 ;
        RECT 610.950 441.450 613.050 442.050 ;
        RECT 601.950 440.550 613.050 441.450 ;
        RECT 601.950 439.950 604.050 440.550 ;
        RECT 610.950 439.950 613.050 440.550 ;
        RECT 614.100 438.600 615.300 445.950 ;
        RECT 620.100 444.150 621.900 445.950 ;
        RECT 632.100 444.150 633.900 445.950 ;
        RECT 638.100 444.150 639.900 445.950 ;
        RECT 641.100 442.200 642.000 445.950 ;
        RECT 650.550 445.050 651.450 448.950 ;
        RECT 656.100 448.050 657.900 449.850 ;
        RECT 662.700 448.050 663.900 455.400 ;
        RECT 667.950 456.450 670.050 457.050 ;
        RECT 679.950 456.450 682.050 457.050 ;
        RECT 667.950 455.550 682.050 456.450 ;
        RECT 667.950 454.950 670.050 455.550 ;
        RECT 679.950 454.950 682.050 455.550 ;
        RECT 664.950 453.450 667.050 454.200 ;
        RECT 670.950 453.450 673.050 453.900 ;
        RECT 664.950 452.550 673.050 453.450 ;
        RECT 664.950 452.100 667.050 452.550 ;
        RECT 670.950 451.800 673.050 452.550 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 680.100 445.950 682.200 448.050 ;
        RECT 650.550 443.550 655.050 445.050 ;
        RECT 659.100 444.150 660.900 445.950 ;
        RECT 651.000 442.950 655.050 443.550 ;
        RECT 622.950 441.450 625.050 442.050 ;
        RECT 628.950 441.450 631.050 442.050 ;
        RECT 622.950 440.550 631.050 441.450 ;
        RECT 622.950 439.950 625.050 440.550 ;
        RECT 628.950 439.950 631.050 440.550 ;
        RECT 590.100 432.600 591.900 435.600 ;
        RECT 593.100 432.000 594.900 435.600 ;
        RECT 608.700 432.000 610.500 438.600 ;
        RECT 613.200 432.600 615.000 438.600 ;
        RECT 617.700 432.000 619.500 438.600 ;
        RECT 632.100 432.000 633.900 441.600 ;
        RECT 638.700 441.000 642.000 442.200 ;
        RECT 662.700 441.600 663.900 445.950 ;
        RECT 665.100 444.150 666.900 445.950 ;
        RECT 680.250 444.150 682.050 445.950 ;
        RECT 638.700 432.600 640.500 441.000 ;
        RECT 662.700 440.700 666.300 441.600 ;
        RECT 683.100 441.300 684.000 461.400 ;
        RECT 686.100 456.000 687.900 468.000 ;
        RECT 689.100 455.400 690.900 467.400 ;
        RECT 693.000 456.450 697.050 457.050 ;
        RECT 685.200 448.050 687.000 449.850 ;
        RECT 689.400 448.050 690.300 455.400 ;
        RECT 692.550 454.950 697.050 456.450 ;
        RECT 701.400 455.400 703.200 468.000 ;
        RECT 706.500 456.900 708.300 467.400 ;
        RECT 709.500 461.400 711.300 468.000 ;
        RECT 722.100 461.400 723.900 468.000 ;
        RECT 725.100 461.400 726.900 467.400 ;
        RECT 728.100 462.000 729.900 468.000 ;
        RECT 725.400 461.100 726.900 461.400 ;
        RECT 731.100 461.400 732.900 467.400 ;
        RECT 746.100 461.400 747.900 468.000 ;
        RECT 749.100 461.400 750.900 467.400 ;
        RECT 731.100 461.100 732.000 461.400 ;
        RECT 725.400 460.200 732.000 461.100 ;
        RECT 709.200 458.100 711.000 459.900 ;
        RECT 706.500 455.400 708.900 456.900 ;
        RECT 685.500 445.950 687.600 448.050 ;
        RECT 688.800 445.950 690.900 448.050 ;
        RECT 656.100 437.700 663.900 439.050 ;
        RECT 656.100 432.600 657.900 437.700 ;
        RECT 659.100 432.000 660.900 436.800 ;
        RECT 662.100 432.600 663.900 437.700 ;
        RECT 665.100 438.600 666.300 440.700 ;
        RECT 680.100 440.400 688.500 441.300 ;
        RECT 665.100 432.600 666.900 438.600 ;
        RECT 680.100 432.600 681.900 440.400 ;
        RECT 686.700 439.500 688.500 440.400 ;
        RECT 689.400 438.600 690.300 445.950 ;
        RECT 692.550 442.050 693.450 454.950 ;
        RECT 696.000 450.450 700.050 451.050 ;
        RECT 695.550 448.950 700.050 450.450 ;
        RECT 695.550 445.050 696.450 448.950 ;
        RECT 701.100 448.050 702.900 449.850 ;
        RECT 707.700 448.050 708.900 455.400 ;
        RECT 725.100 448.050 726.900 449.850 ;
        RECT 731.100 448.050 732.000 460.200 ;
        RECT 733.950 450.450 738.000 451.050 ;
        RECT 733.950 448.950 738.450 450.450 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 695.550 443.550 700.050 445.050 ;
        RECT 704.100 444.150 705.900 445.950 ;
        RECT 696.000 442.950 700.050 443.550 ;
        RECT 691.950 439.950 694.050 442.050 ;
        RECT 707.700 441.600 708.900 445.950 ;
        RECT 710.100 444.150 711.900 445.950 ;
        RECT 722.100 444.150 723.900 445.950 ;
        RECT 728.100 444.150 729.900 445.950 ;
        RECT 731.100 442.200 732.000 445.950 ;
        RECT 707.700 440.700 711.300 441.600 ;
        RECT 684.600 432.000 686.400 438.600 ;
        RECT 687.600 436.800 690.300 438.600 ;
        RECT 701.100 437.700 708.900 439.050 ;
        RECT 687.600 432.600 689.400 436.800 ;
        RECT 701.100 432.600 702.900 437.700 ;
        RECT 704.100 432.000 705.900 436.800 ;
        RECT 707.100 432.600 708.900 437.700 ;
        RECT 710.100 438.600 711.300 440.700 ;
        RECT 710.100 432.600 711.900 438.600 ;
        RECT 722.100 432.000 723.900 441.600 ;
        RECT 728.700 441.000 732.000 442.200 ;
        RECT 737.550 441.900 738.450 448.950 ;
        RECT 746.100 445.950 748.200 448.050 ;
        RECT 746.250 444.150 748.050 445.950 ;
        RECT 728.700 432.600 730.500 441.000 ;
        RECT 736.950 439.800 739.050 441.900 ;
        RECT 749.100 441.300 750.000 461.400 ;
        RECT 752.100 456.000 753.900 468.000 ;
        RECT 755.100 455.400 756.900 467.400 ;
        RECT 770.100 461.400 771.900 468.000 ;
        RECT 773.100 461.400 774.900 467.400 ;
        RECT 776.100 461.400 777.900 468.000 ;
        RECT 791.100 461.400 792.900 468.000 ;
        RECT 794.100 461.400 795.900 467.400 ;
        RECT 751.200 448.050 753.000 449.850 ;
        RECT 755.400 448.050 756.300 455.400 ;
        RECT 773.700 448.050 774.900 461.400 ;
        RECT 751.500 445.950 753.600 448.050 ;
        RECT 754.800 445.950 756.900 448.050 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 791.100 445.950 793.200 448.050 ;
        RECT 746.100 440.400 754.500 441.300 ;
        RECT 746.100 432.600 747.900 440.400 ;
        RECT 752.700 439.500 754.500 440.400 ;
        RECT 755.400 438.600 756.300 445.950 ;
        RECT 770.100 444.150 771.900 445.950 ;
        RECT 773.700 440.700 774.900 445.950 ;
        RECT 775.950 444.150 777.750 445.950 ;
        RECT 791.250 444.150 793.050 445.950 ;
        RECT 794.100 441.300 795.000 461.400 ;
        RECT 797.100 456.000 798.900 468.000 ;
        RECT 800.100 455.400 801.900 467.400 ;
        RECT 815.100 461.400 816.900 468.000 ;
        RECT 818.100 461.400 819.900 467.400 ;
        RECT 821.100 461.400 822.900 468.000 ;
        RECT 833.100 461.400 834.900 468.000 ;
        RECT 836.100 461.400 837.900 467.400 ;
        RECT 839.100 462.000 840.900 468.000 ;
        RECT 796.200 448.050 798.000 449.850 ;
        RECT 800.400 448.050 801.300 455.400 ;
        RECT 818.100 448.050 819.300 461.400 ;
        RECT 836.400 461.100 837.900 461.400 ;
        RECT 842.100 461.400 843.900 467.400 ;
        RECT 854.100 461.400 855.900 468.000 ;
        RECT 857.100 461.400 858.900 467.400 ;
        RECT 860.100 462.000 861.900 468.000 ;
        RECT 842.100 461.100 843.000 461.400 ;
        RECT 836.400 460.200 843.000 461.100 ;
        RECT 857.400 461.100 858.900 461.400 ;
        RECT 863.100 461.400 864.900 467.400 ;
        RECT 863.100 461.100 864.000 461.400 ;
        RECT 857.400 460.200 864.000 461.100 ;
        RECT 836.100 448.050 837.900 449.850 ;
        RECT 842.100 448.050 843.000 460.200 ;
        RECT 857.100 448.050 858.900 449.850 ;
        RECT 863.100 448.050 864.000 460.200 ;
        RECT 878.100 456.300 879.900 467.400 ;
        RECT 881.100 457.200 882.900 468.000 ;
        RECT 884.100 456.300 885.900 467.400 ;
        RECT 878.100 455.400 885.900 456.300 ;
        RECT 887.100 455.400 888.900 467.400 ;
        RECT 902.400 455.400 904.200 468.000 ;
        RECT 907.500 456.900 909.300 467.400 ;
        RECT 910.500 461.400 912.300 468.000 ;
        RECT 910.200 458.100 912.000 459.900 ;
        RECT 907.500 455.400 909.900 456.900 ;
        RECT 923.100 456.300 924.900 467.400 ;
        RECT 926.100 457.200 927.900 468.000 ;
        RECT 929.100 456.300 930.900 467.400 ;
        RECT 923.100 455.400 930.900 456.300 ;
        RECT 932.100 455.400 933.900 467.400 ;
        RECT 868.950 453.450 871.050 454.050 ;
        RECT 877.950 453.450 880.050 454.050 ;
        RECT 868.950 452.550 880.050 453.450 ;
        RECT 868.950 451.950 871.050 452.550 ;
        RECT 877.950 451.950 880.050 452.550 ;
        RECT 873.000 450.450 877.050 451.050 ;
        RECT 872.550 448.950 877.050 450.450 ;
        RECT 796.500 445.950 798.600 448.050 ;
        RECT 799.800 445.950 801.900 448.050 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 750.600 432.000 752.400 438.600 ;
        RECT 753.600 436.800 756.300 438.600 ;
        RECT 770.700 439.800 774.900 440.700 ;
        RECT 791.100 440.400 799.500 441.300 ;
        RECT 753.600 432.600 755.400 436.800 ;
        RECT 770.700 432.600 772.500 439.800 ;
        RECT 775.800 432.000 777.600 438.600 ;
        RECT 791.100 432.600 792.900 440.400 ;
        RECT 797.700 439.500 799.500 440.400 ;
        RECT 800.400 438.600 801.300 445.950 ;
        RECT 815.250 444.150 817.050 445.950 ;
        RECT 818.100 440.700 819.300 445.950 ;
        RECT 821.100 444.150 822.900 445.950 ;
        RECT 833.100 444.150 834.900 445.950 ;
        RECT 839.100 444.150 840.900 445.950 ;
        RECT 842.100 442.200 843.000 445.950 ;
        RECT 854.100 444.150 855.900 445.950 ;
        RECT 860.100 444.150 861.900 445.950 ;
        RECT 863.100 442.200 864.000 445.950 ;
        RECT 872.550 444.450 873.450 448.950 ;
        RECT 881.250 448.050 883.050 449.850 ;
        RECT 887.700 448.050 888.600 455.400 ;
        RECT 897.000 450.450 901.050 451.050 ;
        RECT 896.550 448.950 901.050 450.450 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 872.550 443.550 876.450 444.450 ;
        RECT 878.100 444.150 879.900 445.950 ;
        RECT 884.250 444.150 886.050 445.950 ;
        RECT 818.100 439.800 822.300 440.700 ;
        RECT 795.600 432.000 797.400 438.600 ;
        RECT 798.600 436.800 801.300 438.600 ;
        RECT 798.600 432.600 800.400 436.800 ;
        RECT 815.400 432.000 817.200 438.600 ;
        RECT 820.500 432.600 822.300 439.800 ;
        RECT 833.100 432.000 834.900 441.600 ;
        RECT 839.700 441.000 843.000 442.200 ;
        RECT 839.700 432.600 841.500 441.000 ;
        RECT 854.100 432.000 855.900 441.600 ;
        RECT 860.700 441.000 864.000 442.200 ;
        RECT 875.550 441.450 876.450 443.550 ;
        RECT 883.950 441.450 886.050 442.050 ;
        RECT 860.700 432.600 862.500 441.000 ;
        RECT 875.550 440.550 886.050 441.450 ;
        RECT 883.950 439.950 886.050 440.550 ;
        RECT 887.700 438.600 888.600 445.950 ;
        RECT 896.550 445.050 897.450 448.950 ;
        RECT 902.100 448.050 903.900 449.850 ;
        RECT 908.700 448.050 909.900 455.400 ;
        RECT 916.950 453.450 919.050 454.050 ;
        RECT 922.950 453.450 925.050 454.200 ;
        RECT 928.950 453.450 931.050 454.050 ;
        RECT 916.950 452.550 931.050 453.450 ;
        RECT 916.950 451.950 919.050 452.550 ;
        RECT 922.950 452.100 925.050 452.550 ;
        RECT 928.950 451.950 931.050 452.550 ;
        RECT 926.250 448.050 928.050 449.850 ;
        RECT 932.700 448.050 933.600 455.400 ;
        RECT 901.950 445.950 904.050 448.050 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 907.950 445.950 910.050 448.050 ;
        RECT 910.950 445.950 913.050 448.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 925.950 445.950 928.050 448.050 ;
        RECT 928.950 445.950 931.050 448.050 ;
        RECT 931.950 445.950 934.050 448.050 ;
        RECT 896.550 443.550 901.050 445.050 ;
        RECT 905.100 444.150 906.900 445.950 ;
        RECT 897.000 442.950 901.050 443.550 ;
        RECT 908.700 441.600 909.900 445.950 ;
        RECT 911.100 444.150 912.900 445.950 ;
        RECT 923.100 444.150 924.900 445.950 ;
        RECT 929.250 444.150 931.050 445.950 ;
        RECT 908.700 440.700 912.300 441.600 ;
        RECT 879.000 432.000 880.800 438.600 ;
        RECT 883.500 437.400 888.600 438.600 ;
        RECT 902.100 437.700 909.900 439.050 ;
        RECT 883.500 432.600 885.300 437.400 ;
        RECT 886.500 432.000 888.300 435.600 ;
        RECT 902.100 432.600 903.900 437.700 ;
        RECT 905.100 432.000 906.900 436.800 ;
        RECT 908.100 432.600 909.900 437.700 ;
        RECT 911.100 438.600 912.300 440.700 ;
        RECT 932.700 438.600 933.600 445.950 ;
        RECT 911.100 432.600 912.900 438.600 ;
        RECT 924.000 432.000 925.800 438.600 ;
        RECT 928.500 437.400 933.600 438.600 ;
        RECT 928.500 432.600 930.300 437.400 ;
        RECT 931.500 432.000 933.300 435.600 ;
        RECT 11.100 422.400 12.900 428.400 ;
        RECT 14.100 422.400 15.900 429.000 ;
        RECT 17.100 425.400 18.900 428.400 ;
        RECT 11.100 415.050 12.300 422.400 ;
        RECT 17.700 421.500 18.900 425.400 ;
        RECT 13.200 420.600 18.900 421.500 ;
        RECT 32.100 422.400 33.900 428.400 ;
        RECT 35.100 422.400 36.900 429.000 ;
        RECT 38.100 425.400 39.900 428.400 ;
        RECT 13.200 419.700 15.000 420.600 ;
        RECT 11.100 412.950 13.200 415.050 ;
        RECT 11.100 405.600 12.300 412.950 ;
        RECT 14.100 408.300 15.000 419.700 ;
        RECT 32.100 415.050 33.300 422.400 ;
        RECT 38.700 421.500 39.900 425.400 ;
        RECT 34.200 420.600 39.900 421.500 ;
        RECT 34.200 419.700 36.000 420.600 ;
        RECT 16.500 412.950 18.600 415.050 ;
        RECT 16.800 411.150 18.600 412.950 ;
        RECT 32.100 412.950 34.200 415.050 ;
        RECT 13.200 407.400 15.000 408.300 ;
        RECT 13.200 406.500 18.900 407.400 ;
        RECT 11.100 393.600 12.900 405.600 ;
        RECT 14.100 393.000 15.900 403.800 ;
        RECT 17.700 399.600 18.900 406.500 ;
        RECT 17.100 393.600 18.900 399.600 ;
        RECT 32.100 405.600 33.300 412.950 ;
        RECT 35.100 408.300 36.000 419.700 ;
        RECT 50.100 419.400 51.900 429.000 ;
        RECT 56.700 420.000 58.500 428.400 ;
        RECT 71.100 425.400 72.900 428.400 ;
        RECT 71.100 421.500 72.300 425.400 ;
        RECT 74.100 422.400 75.900 429.000 ;
        RECT 77.100 422.400 78.900 428.400 ;
        RECT 89.100 422.400 90.900 429.000 ;
        RECT 92.100 422.400 93.900 428.400 ;
        RECT 95.100 422.400 96.900 429.000 ;
        RECT 71.100 420.600 76.800 421.500 ;
        RECT 56.700 418.800 60.000 420.000 ;
        RECT 50.100 415.050 51.900 416.850 ;
        RECT 56.100 415.050 57.900 416.850 ;
        RECT 59.100 415.050 60.000 418.800 ;
        RECT 75.000 419.700 76.800 420.600 ;
        RECT 37.500 412.950 39.600 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 55.950 412.950 58.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 71.400 412.950 73.500 415.050 ;
        RECT 37.800 411.150 39.600 412.950 ;
        RECT 53.100 411.150 54.900 412.950 ;
        RECT 34.200 407.400 36.000 408.300 ;
        RECT 34.200 406.500 39.900 407.400 ;
        RECT 32.100 393.600 33.900 405.600 ;
        RECT 35.100 393.000 36.900 403.800 ;
        RECT 38.700 399.600 39.900 406.500 ;
        RECT 59.100 400.800 60.000 412.950 ;
        RECT 71.400 411.150 73.200 412.950 ;
        RECT 75.000 408.300 75.900 419.700 ;
        RECT 77.700 415.050 78.900 422.400 ;
        RECT 92.550 415.050 93.600 422.400 ;
        RECT 107.700 421.200 109.500 428.400 ;
        RECT 112.800 422.400 114.600 429.000 ;
        RECT 128.100 425.400 129.900 429.000 ;
        RECT 131.100 425.400 132.900 428.400 ;
        RECT 146.100 425.400 147.900 429.000 ;
        RECT 149.100 425.400 150.900 428.400 ;
        RECT 152.100 425.400 153.900 429.000 ;
        RECT 107.700 420.300 111.900 421.200 ;
        RECT 94.800 415.050 96.600 416.850 ;
        RECT 107.100 415.050 108.900 416.850 ;
        RECT 110.700 415.050 111.900 420.300 ;
        RECT 112.950 420.450 115.050 420.900 ;
        RECT 127.950 420.450 130.050 421.050 ;
        RECT 112.950 419.550 130.050 420.450 ;
        RECT 112.950 418.800 115.050 419.550 ;
        RECT 127.950 418.950 130.050 419.550 ;
        RECT 112.950 415.050 114.750 416.850 ;
        RECT 131.100 415.050 132.300 425.400 ;
        RECT 149.700 415.050 150.600 425.400 ;
        RECT 167.100 422.400 168.900 429.000 ;
        RECT 170.100 422.400 171.900 428.400 ;
        RECT 185.100 423.300 186.900 428.400 ;
        RECT 188.100 424.200 189.900 429.000 ;
        RECT 191.100 423.300 192.900 428.400 ;
        RECT 167.100 415.050 168.900 416.850 ;
        RECT 170.100 415.050 171.300 422.400 ;
        RECT 185.100 421.950 192.900 423.300 ;
        RECT 194.100 422.400 195.900 428.400 ;
        RECT 206.100 422.400 207.900 429.000 ;
        RECT 209.100 422.400 210.900 428.400 ;
        RECT 212.100 422.400 213.900 429.000 ;
        RECT 224.100 422.400 225.900 429.000 ;
        RECT 194.100 420.300 195.300 422.400 ;
        RECT 191.700 419.400 195.300 420.300 ;
        RECT 180.000 417.450 184.050 418.050 ;
        RECT 179.550 415.950 184.050 417.450 ;
        RECT 76.800 412.950 78.900 415.050 ;
        RECT 89.400 412.950 93.600 415.050 ;
        RECT 94.500 412.950 96.600 415.050 ;
        RECT 106.950 412.950 109.050 415.050 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 75.000 407.400 76.800 408.300 ;
        RECT 53.400 399.900 60.000 400.800 ;
        RECT 53.400 399.600 54.900 399.900 ;
        RECT 38.100 393.600 39.900 399.600 ;
        RECT 50.100 393.000 51.900 399.600 ;
        RECT 53.100 393.600 54.900 399.600 ;
        RECT 59.100 399.600 60.000 399.900 ;
        RECT 71.100 406.500 76.800 407.400 ;
        RECT 71.100 399.600 72.300 406.500 ;
        RECT 77.700 405.600 78.900 412.950 ;
        RECT 92.550 405.600 93.600 412.950 ;
        RECT 56.100 393.000 57.900 399.000 ;
        RECT 59.100 393.600 60.900 399.600 ;
        RECT 71.100 393.600 72.900 399.600 ;
        RECT 74.100 393.000 75.900 403.800 ;
        RECT 77.100 393.600 78.900 405.600 ;
        RECT 89.100 393.000 90.900 405.600 ;
        RECT 92.100 393.600 93.900 405.600 ;
        RECT 95.100 393.000 96.900 405.600 ;
        RECT 110.700 399.600 111.900 412.950 ;
        RECT 128.100 411.150 129.900 412.950 ;
        RECT 131.100 399.600 132.300 412.950 ;
        RECT 146.100 411.150 147.900 412.950 ;
        RECT 149.700 405.600 150.600 412.950 ;
        RECT 151.950 411.150 153.750 412.950 ;
        RECT 170.100 405.600 171.300 412.950 ;
        RECT 179.550 412.050 180.450 415.950 ;
        RECT 188.100 415.050 189.900 416.850 ;
        RECT 191.700 415.050 192.900 419.400 ;
        RECT 196.950 417.450 201.000 418.050 ;
        RECT 194.100 415.050 195.900 416.850 ;
        RECT 196.950 415.950 201.450 417.450 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 193.950 412.950 196.050 415.050 ;
        RECT 179.550 410.550 184.050 412.050 ;
        RECT 185.100 411.150 186.900 412.950 ;
        RECT 180.000 409.950 184.050 410.550 ;
        RECT 191.700 405.600 192.900 412.950 ;
        RECT 200.550 412.050 201.450 415.950 ;
        RECT 206.400 415.050 208.200 416.850 ;
        RECT 209.400 415.050 210.450 422.400 ;
        RECT 227.100 421.500 228.900 428.400 ;
        RECT 230.100 422.400 231.900 429.000 ;
        RECT 233.100 421.500 234.900 428.400 ;
        RECT 236.100 422.400 237.900 429.000 ;
        RECT 239.100 421.500 240.900 428.400 ;
        RECT 242.100 422.400 243.900 429.000 ;
        RECT 245.100 421.500 246.900 428.400 ;
        RECT 248.100 422.400 249.900 429.000 ;
        RECT 227.100 420.300 231.000 421.500 ;
        RECT 233.100 420.300 237.000 421.500 ;
        RECT 239.100 420.300 243.000 421.500 ;
        RECT 245.100 420.300 247.950 421.500 ;
        RECT 263.700 421.200 265.500 428.400 ;
        RECT 268.800 422.400 270.600 429.000 ;
        RECT 281.100 422.400 282.900 428.400 ;
        RECT 263.700 420.300 267.900 421.200 ;
        RECT 229.800 419.400 231.000 420.300 ;
        RECT 235.800 419.400 237.000 420.300 ;
        RECT 241.800 419.400 243.000 420.300 ;
        RECT 229.800 418.200 234.000 419.400 ;
        RECT 226.800 415.050 228.600 416.850 ;
        RECT 206.400 412.950 208.500 415.050 ;
        RECT 209.400 412.950 213.600 415.050 ;
        RECT 226.800 412.950 228.900 415.050 ;
        RECT 196.950 410.550 201.450 412.050 ;
        RECT 196.950 409.950 201.000 410.550 ;
        RECT 209.400 405.600 210.450 412.950 ;
        RECT 229.800 407.700 231.000 418.200 ;
        RECT 232.200 417.600 234.000 418.200 ;
        RECT 235.800 418.200 240.000 419.400 ;
        RECT 235.800 407.700 237.000 418.200 ;
        RECT 238.200 417.600 240.000 418.200 ;
        RECT 241.800 418.200 246.000 419.400 ;
        RECT 241.800 407.700 243.000 418.200 ;
        RECT 244.200 417.600 246.000 418.200 ;
        RECT 246.900 415.050 247.950 420.300 ;
        RECT 263.100 415.050 264.900 416.850 ;
        RECT 266.700 415.050 267.900 420.300 ;
        RECT 281.700 420.300 282.900 422.400 ;
        RECT 284.100 423.300 285.900 428.400 ;
        RECT 287.100 424.200 288.900 429.000 ;
        RECT 290.100 423.300 291.900 428.400 ;
        RECT 284.100 421.950 291.900 423.300 ;
        RECT 302.100 425.400 303.900 428.400 ;
        RECT 302.100 421.500 303.300 425.400 ;
        RECT 305.100 422.400 306.900 429.000 ;
        RECT 308.100 422.400 309.900 428.400 ;
        RECT 323.100 422.400 324.900 428.400 ;
        RECT 326.100 422.400 327.900 429.000 ;
        RECT 329.700 422.400 331.500 428.400 ;
        RECT 335.100 422.400 336.900 429.000 ;
        RECT 340.500 422.400 342.300 428.400 ;
        RECT 344.700 425.400 346.500 428.400 ;
        RECT 347.700 425.400 349.500 428.400 ;
        RECT 350.700 425.400 352.500 428.400 ;
        RECT 353.700 425.400 355.500 429.000 ;
        RECT 344.700 423.300 346.800 425.400 ;
        RECT 347.700 423.300 349.800 425.400 ;
        RECT 350.700 423.300 352.800 425.400 ;
        RECT 358.200 424.500 360.000 428.400 ;
        RECT 361.200 425.400 363.000 429.000 ;
        RECT 364.200 425.400 366.000 428.400 ;
        RECT 367.200 425.400 369.000 428.400 ;
        RECT 370.200 425.400 372.000 428.400 ;
        RECT 373.200 425.400 375.000 428.400 ;
        RECT 354.600 423.600 356.400 424.500 ;
        RECT 353.700 422.400 356.400 423.600 ;
        RECT 358.200 422.400 360.900 424.500 ;
        RECT 364.200 423.300 366.300 425.400 ;
        RECT 367.200 423.300 369.300 425.400 ;
        RECT 370.200 423.300 372.300 425.400 ;
        RECT 373.200 423.300 375.300 425.400 ;
        RECT 377.400 423.600 379.200 428.400 ;
        RECT 377.400 422.400 381.600 423.600 ;
        RECT 382.500 422.400 384.300 429.000 ;
        RECT 387.900 422.400 389.700 428.400 ;
        RECT 302.100 420.600 307.800 421.500 ;
        RECT 281.700 419.400 285.300 420.300 ;
        RECT 268.950 415.050 270.750 416.850 ;
        RECT 281.100 415.050 282.900 416.850 ;
        RECT 284.100 415.050 285.300 419.400 ;
        RECT 306.000 419.700 307.800 420.600 ;
        RECT 287.100 415.050 288.900 416.850 ;
        RECT 244.800 412.950 247.950 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 302.400 412.950 304.500 415.050 ;
        RECT 246.900 407.700 247.950 412.950 ;
        RECT 227.100 406.500 231.000 407.700 ;
        RECT 233.100 406.500 237.000 407.700 ;
        RECT 239.100 406.500 243.000 407.700 ;
        RECT 245.100 406.500 247.950 407.700 ;
        RECT 147.000 404.400 150.600 405.600 ;
        RECT 107.100 393.000 108.900 399.600 ;
        RECT 110.100 393.600 111.900 399.600 ;
        RECT 113.100 393.000 114.900 399.600 ;
        RECT 128.100 393.000 129.900 399.600 ;
        RECT 131.100 393.600 132.900 399.600 ;
        RECT 147.000 393.600 148.800 404.400 ;
        RECT 152.100 393.000 153.900 405.600 ;
        RECT 167.100 393.000 168.900 405.600 ;
        RECT 170.100 393.600 171.900 405.600 ;
        RECT 185.400 393.000 187.200 405.600 ;
        RECT 190.500 404.100 192.900 405.600 ;
        RECT 190.500 393.600 192.300 404.100 ;
        RECT 193.200 401.100 195.000 402.900 ;
        RECT 193.500 393.000 195.300 399.600 ;
        RECT 206.100 393.000 207.900 405.600 ;
        RECT 209.100 393.600 210.900 405.600 ;
        RECT 212.100 393.000 213.900 405.600 ;
        RECT 224.100 393.000 225.900 405.600 ;
        RECT 227.100 393.600 228.900 406.500 ;
        RECT 230.100 393.000 231.900 405.600 ;
        RECT 233.100 393.600 234.900 406.500 ;
        RECT 236.100 393.000 237.900 405.600 ;
        RECT 239.100 393.600 240.900 406.500 ;
        RECT 242.100 393.000 243.900 405.600 ;
        RECT 245.100 393.600 246.900 406.500 ;
        RECT 248.100 393.000 249.900 405.600 ;
        RECT 266.700 399.600 267.900 412.950 ;
        RECT 271.950 408.450 274.050 409.050 ;
        RECT 280.950 408.450 283.050 409.050 ;
        RECT 271.950 407.550 283.050 408.450 ;
        RECT 271.950 406.950 274.050 407.550 ;
        RECT 280.950 406.950 283.050 407.550 ;
        RECT 284.100 405.600 285.300 412.950 ;
        RECT 290.100 411.150 291.900 412.950 ;
        RECT 302.400 411.150 304.200 412.950 ;
        RECT 306.000 408.300 306.900 419.700 ;
        RECT 308.700 415.050 309.900 422.400 ;
        RECT 323.700 415.050 324.900 422.400 ;
        RECT 329.700 418.800 330.900 422.400 ;
        RECT 340.800 421.500 342.300 422.400 ;
        RECT 349.800 421.800 351.600 422.400 ;
        RECT 353.700 421.800 354.600 422.400 ;
        RECT 333.900 420.300 342.300 421.500 ;
        RECT 347.400 420.600 354.600 421.800 ;
        RECT 369.300 420.600 375.900 422.400 ;
        RECT 333.900 419.700 335.700 420.300 ;
        RECT 344.400 418.800 346.500 419.700 ;
        RECT 329.700 417.600 346.500 418.800 ;
        RECT 347.400 417.600 348.300 420.600 ;
        RECT 352.800 417.900 354.600 418.800 ;
        RECT 362.100 418.500 363.900 420.300 ;
        RECT 380.100 419.100 381.600 422.400 ;
        RECT 355.800 417.900 357.900 418.050 ;
        RECT 326.100 415.050 327.900 416.850 ;
        RECT 307.800 412.950 309.900 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 306.000 407.400 307.800 408.300 ;
        RECT 302.100 406.500 307.800 407.400 ;
        RECT 284.100 404.100 286.500 405.600 ;
        RECT 282.000 401.100 283.800 402.900 ;
        RECT 263.100 393.000 264.900 399.600 ;
        RECT 266.100 393.600 267.900 399.600 ;
        RECT 269.100 393.000 270.900 399.600 ;
        RECT 281.700 393.000 283.500 399.600 ;
        RECT 284.700 393.600 286.500 404.100 ;
        RECT 289.800 393.000 291.600 405.600 ;
        RECT 302.100 399.600 303.300 406.500 ;
        RECT 308.700 405.600 309.900 412.950 ;
        RECT 323.700 405.600 324.900 412.950 ;
        RECT 302.100 393.600 303.900 399.600 ;
        RECT 305.100 393.000 306.900 403.800 ;
        RECT 308.100 393.600 309.900 405.600 ;
        RECT 323.100 393.600 324.900 405.600 ;
        RECT 326.100 393.000 327.900 405.600 ;
        RECT 329.700 401.400 330.900 417.600 ;
        RECT 347.400 415.800 349.200 417.600 ;
        RECT 352.800 417.000 357.900 417.900 ;
        RECT 355.800 415.950 357.900 417.000 ;
        RECT 362.100 417.900 364.200 418.500 ;
        RECT 362.100 416.400 379.200 417.900 ;
        RECT 380.100 417.300 387.900 419.100 ;
        RECT 377.700 414.900 384.300 416.400 ;
        RECT 332.100 413.700 376.500 414.900 ;
        RECT 332.100 412.050 333.900 413.700 ;
        RECT 331.800 409.950 333.900 412.050 ;
        RECT 337.800 411.750 339.900 412.050 ;
        RECT 350.400 411.900 352.200 412.500 ;
        RECT 359.400 411.900 372.900 412.800 ;
        RECT 337.800 409.950 341.700 411.750 ;
        RECT 350.400 410.700 361.500 411.900 ;
        RECT 339.900 409.200 341.700 409.950 ;
        RECT 359.400 409.800 361.500 410.700 ;
        RECT 363.000 409.200 366.900 411.000 ;
        RECT 372.000 410.700 372.900 411.900 ;
        RECT 339.900 408.300 353.400 409.200 ;
        RECT 364.800 408.900 366.900 409.200 ;
        RECT 371.100 408.900 372.900 410.700 ;
        RECT 375.600 412.200 376.500 413.700 ;
        RECT 375.600 410.400 380.700 412.200 ;
        RECT 382.800 412.050 384.300 414.900 ;
        RECT 382.800 409.950 384.900 412.050 ;
        RECT 352.200 407.700 353.400 408.300 ;
        RECT 386.100 407.700 387.900 408.300 ;
        RECT 347.400 406.500 349.500 406.800 ;
        RECT 352.200 406.500 387.900 407.700 ;
        RECT 337.500 405.300 349.500 406.500 ;
        RECT 388.800 405.600 389.700 422.400 ;
        RECT 337.500 404.700 339.300 405.300 ;
        RECT 347.400 404.700 349.500 405.300 ;
        RECT 352.200 404.400 369.900 405.600 ;
        RECT 334.200 403.800 336.000 404.100 ;
        RECT 352.200 403.800 353.400 404.400 ;
        RECT 334.200 402.600 353.400 403.800 ;
        RECT 367.800 403.500 369.900 404.400 ;
        RECT 373.200 404.700 389.700 405.600 ;
        RECT 373.200 403.500 375.300 404.700 ;
        RECT 334.200 402.300 336.000 402.600 ;
        RECT 329.700 400.500 333.300 401.400 ;
        RECT 332.400 399.600 333.300 400.500 ;
        RECT 329.700 393.000 331.500 399.600 ;
        RECT 332.400 398.700 334.500 399.600 ;
        RECT 332.700 393.600 334.500 398.700 ;
        RECT 335.700 393.000 337.500 399.600 ;
        RECT 338.700 393.600 340.500 402.600 ;
        RECT 350.700 399.600 352.800 401.700 ;
        RECT 358.200 401.100 361.500 403.200 ;
        RECT 341.700 393.000 343.500 399.600 ;
        RECT 345.300 396.600 347.400 398.700 ;
        RECT 348.300 396.600 350.400 398.700 ;
        RECT 345.300 393.600 347.100 396.600 ;
        RECT 348.300 393.600 350.100 396.600 ;
        RECT 351.300 393.600 353.100 399.600 ;
        RECT 354.300 393.000 356.100 399.600 ;
        RECT 358.200 393.600 360.000 401.100 ;
        RECT 364.200 399.600 366.900 403.500 ;
        RECT 379.200 402.600 384.900 403.800 ;
        RECT 376.500 401.700 378.300 402.300 ;
        RECT 370.200 400.500 378.300 401.700 ;
        RECT 370.200 399.600 372.300 400.500 ;
        RECT 379.200 399.600 380.400 402.600 ;
        RECT 383.100 402.000 384.900 402.600 ;
        RECT 388.800 401.400 389.700 404.700 ;
        RECT 385.800 400.500 389.700 401.400 ;
        RECT 391.500 425.400 393.300 428.400 ;
        RECT 394.500 425.400 396.300 429.000 ;
        RECT 391.500 412.050 393.000 425.400 ;
        RECT 407.100 422.400 408.900 429.000 ;
        RECT 410.100 422.400 411.900 428.400 ;
        RECT 425.100 422.400 426.900 428.400 ;
        RECT 428.100 422.400 429.900 429.000 ;
        RECT 431.100 425.400 432.900 428.400 ;
        RECT 407.100 415.050 408.900 416.850 ;
        RECT 410.100 415.050 411.300 422.400 ;
        RECT 425.100 415.050 426.300 422.400 ;
        RECT 431.700 421.500 432.900 425.400 ;
        RECT 427.200 420.600 432.900 421.500 ;
        RECT 446.100 425.400 447.900 428.400 ;
        RECT 446.100 421.500 447.300 425.400 ;
        RECT 449.100 422.400 450.900 429.000 ;
        RECT 452.100 422.400 453.900 428.400 ;
        RECT 464.100 422.400 465.900 429.000 ;
        RECT 467.100 422.400 468.900 428.400 ;
        RECT 446.100 420.600 451.800 421.500 ;
        RECT 427.200 419.700 429.000 420.600 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 425.100 412.950 427.200 415.050 ;
        RECT 391.500 409.950 393.900 412.050 ;
        RECT 385.800 399.600 387.000 400.500 ;
        RECT 391.500 399.600 393.000 409.950 ;
        RECT 410.100 405.600 411.300 412.950 ;
        RECT 425.100 405.600 426.300 412.950 ;
        RECT 428.100 408.300 429.000 419.700 ;
        RECT 450.000 419.700 451.800 420.600 ;
        RECT 430.500 412.950 432.600 415.050 ;
        RECT 430.800 411.150 432.600 412.950 ;
        RECT 446.400 412.950 448.500 415.050 ;
        RECT 446.400 411.150 448.200 412.950 ;
        RECT 427.200 407.400 429.000 408.300 ;
        RECT 450.000 408.300 450.900 419.700 ;
        RECT 452.700 415.050 453.900 422.400 ;
        RECT 464.100 415.050 465.900 416.850 ;
        RECT 467.100 415.050 468.300 422.400 ;
        RECT 479.100 420.600 480.900 428.400 ;
        RECT 483.600 422.400 485.400 429.000 ;
        RECT 486.600 424.200 488.400 428.400 ;
        RECT 500.100 425.400 501.900 429.000 ;
        RECT 503.100 425.400 504.900 428.400 ;
        RECT 515.100 425.400 516.900 428.400 ;
        RECT 486.600 422.400 489.300 424.200 ;
        RECT 485.700 420.600 487.500 421.500 ;
        RECT 479.100 419.700 487.500 420.600 ;
        RECT 479.250 415.050 481.050 416.850 ;
        RECT 451.800 412.950 453.900 415.050 ;
        RECT 463.950 412.950 466.050 415.050 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 479.100 412.950 481.200 415.050 ;
        RECT 450.000 407.400 451.800 408.300 ;
        RECT 427.200 406.500 432.900 407.400 ;
        RECT 361.200 393.000 363.000 399.600 ;
        RECT 364.200 393.600 366.000 399.600 ;
        RECT 367.200 396.600 369.300 398.700 ;
        RECT 370.200 396.600 372.300 398.700 ;
        RECT 373.200 396.600 375.300 398.700 ;
        RECT 367.200 393.600 369.000 396.600 ;
        RECT 370.200 393.600 372.000 396.600 ;
        RECT 373.200 393.600 375.000 396.600 ;
        RECT 376.200 393.000 378.000 399.600 ;
        RECT 379.200 393.600 381.000 399.600 ;
        RECT 382.200 393.000 384.000 399.600 ;
        RECT 385.200 393.600 387.000 399.600 ;
        RECT 388.200 393.000 390.000 399.600 ;
        RECT 391.500 393.600 393.300 399.600 ;
        RECT 394.500 393.000 396.300 399.600 ;
        RECT 407.100 393.000 408.900 405.600 ;
        RECT 410.100 393.600 411.900 405.600 ;
        RECT 425.100 393.600 426.900 405.600 ;
        RECT 428.100 393.000 429.900 403.800 ;
        RECT 431.700 399.600 432.900 406.500 ;
        RECT 431.100 393.600 432.900 399.600 ;
        RECT 446.100 406.500 451.800 407.400 ;
        RECT 446.100 399.600 447.300 406.500 ;
        RECT 452.700 405.600 453.900 412.950 ;
        RECT 467.100 405.600 468.300 412.950 ;
        RECT 446.100 393.600 447.900 399.600 ;
        RECT 449.100 393.000 450.900 403.800 ;
        RECT 452.100 393.600 453.900 405.600 ;
        RECT 464.100 393.000 465.900 405.600 ;
        RECT 467.100 393.600 468.900 405.600 ;
        RECT 482.100 399.600 483.000 419.700 ;
        RECT 488.400 415.050 489.300 422.400 ;
        RECT 503.100 415.050 504.300 425.400 ;
        RECT 515.100 421.500 516.300 425.400 ;
        RECT 518.100 422.400 519.900 429.000 ;
        RECT 521.100 422.400 522.900 428.400 ;
        RECT 515.100 420.600 520.800 421.500 ;
        RECT 519.000 419.700 520.800 420.600 ;
        RECT 484.500 412.950 486.600 415.050 ;
        RECT 487.800 412.950 489.900 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 515.400 412.950 517.500 415.050 ;
        RECT 484.200 411.150 486.000 412.950 ;
        RECT 488.400 405.600 489.300 412.950 ;
        RECT 500.100 411.150 501.900 412.950 ;
        RECT 479.100 393.000 480.900 399.600 ;
        RECT 482.100 393.600 483.900 399.600 ;
        RECT 485.100 393.000 486.900 405.000 ;
        RECT 488.100 393.600 489.900 405.600 ;
        RECT 503.100 399.600 504.300 412.950 ;
        RECT 515.400 411.150 517.200 412.950 ;
        RECT 519.000 408.300 519.900 419.700 ;
        RECT 521.700 415.050 522.900 422.400 ;
        RECT 536.100 425.400 537.900 428.400 ;
        RECT 536.100 421.500 537.300 425.400 ;
        RECT 539.100 422.400 540.900 429.000 ;
        RECT 542.100 422.400 543.900 428.400 ;
        RECT 536.100 420.600 541.800 421.500 ;
        RECT 540.000 419.700 541.800 420.600 ;
        RECT 520.800 412.950 522.900 415.050 ;
        RECT 519.000 407.400 520.800 408.300 ;
        RECT 515.100 406.500 520.800 407.400 ;
        RECT 515.100 399.600 516.300 406.500 ;
        RECT 521.700 405.600 522.900 412.950 ;
        RECT 536.400 412.950 538.500 415.050 ;
        RECT 536.400 411.150 538.200 412.950 ;
        RECT 540.000 408.300 540.900 419.700 ;
        RECT 542.700 415.050 543.900 422.400 ;
        RECT 554.100 420.600 555.900 428.400 ;
        RECT 558.600 422.400 560.400 429.000 ;
        RECT 561.600 424.200 563.400 428.400 ;
        RECT 561.600 422.400 564.300 424.200 ;
        RECT 560.700 420.600 562.500 421.500 ;
        RECT 554.100 419.700 562.500 420.600 ;
        RECT 554.250 415.050 556.050 416.850 ;
        RECT 541.800 412.950 543.900 415.050 ;
        RECT 554.100 412.950 556.200 415.050 ;
        RECT 540.000 407.400 541.800 408.300 ;
        RECT 500.100 393.000 501.900 399.600 ;
        RECT 503.100 393.600 504.900 399.600 ;
        RECT 515.100 393.600 516.900 399.600 ;
        RECT 518.100 393.000 519.900 403.800 ;
        RECT 521.100 393.600 522.900 405.600 ;
        RECT 536.100 406.500 541.800 407.400 ;
        RECT 536.100 399.600 537.300 406.500 ;
        RECT 542.700 405.600 543.900 412.950 ;
        RECT 536.100 393.600 537.900 399.600 ;
        RECT 539.100 393.000 540.900 403.800 ;
        RECT 542.100 393.600 543.900 405.600 ;
        RECT 557.100 399.600 558.000 419.700 ;
        RECT 563.400 415.050 564.300 422.400 ;
        RECT 578.100 422.400 579.900 428.400 ;
        RECT 581.100 422.400 582.900 429.000 ;
        RECT 584.100 425.400 585.900 428.400 ;
        RECT 578.100 415.050 579.300 422.400 ;
        RECT 584.700 421.500 585.900 425.400 ;
        RECT 580.200 420.600 585.900 421.500 ;
        RECT 596.100 420.600 597.900 428.400 ;
        RECT 600.600 422.400 602.400 429.000 ;
        RECT 603.600 424.200 605.400 428.400 ;
        RECT 603.600 422.400 606.300 424.200 ;
        RECT 602.700 420.600 604.500 421.500 ;
        RECT 580.200 419.700 582.000 420.600 ;
        RECT 596.100 419.700 604.500 420.600 ;
        RECT 559.500 412.950 561.600 415.050 ;
        RECT 562.800 412.950 564.900 415.050 ;
        RECT 578.100 412.950 580.200 415.050 ;
        RECT 559.200 411.150 561.000 412.950 ;
        RECT 563.400 405.600 564.300 412.950 ;
        RECT 578.100 405.600 579.300 412.950 ;
        RECT 581.100 408.300 582.000 419.700 ;
        RECT 596.250 415.050 598.050 416.850 ;
        RECT 583.500 412.950 585.600 415.050 ;
        RECT 596.100 412.950 598.200 415.050 ;
        RECT 583.800 411.150 585.600 412.950 ;
        RECT 580.200 407.400 582.000 408.300 ;
        RECT 586.950 408.450 589.050 409.050 ;
        RECT 595.950 408.450 598.050 409.050 ;
        RECT 586.950 407.550 598.050 408.450 ;
        RECT 580.200 406.500 585.900 407.400 ;
        RECT 586.950 406.950 589.050 407.550 ;
        RECT 595.950 406.950 598.050 407.550 ;
        RECT 554.100 393.000 555.900 399.600 ;
        RECT 557.100 393.600 558.900 399.600 ;
        RECT 560.100 393.000 561.900 405.000 ;
        RECT 563.100 393.600 564.900 405.600 ;
        RECT 578.100 393.600 579.900 405.600 ;
        RECT 581.100 393.000 582.900 403.800 ;
        RECT 584.700 399.600 585.900 406.500 ;
        RECT 599.100 399.600 600.000 419.700 ;
        RECT 605.400 415.050 606.300 422.400 ;
        RECT 620.100 423.300 621.900 428.400 ;
        RECT 623.100 424.200 624.900 429.000 ;
        RECT 626.100 423.300 627.900 428.400 ;
        RECT 620.100 421.950 627.900 423.300 ;
        RECT 629.100 422.400 630.900 428.400 ;
        RECT 641.400 422.400 643.200 429.000 ;
        RECT 629.100 420.300 630.300 422.400 ;
        RECT 646.500 421.200 648.300 428.400 ;
        RECT 649.950 426.450 652.050 427.050 ;
        RECT 658.950 426.450 661.050 427.050 ;
        RECT 649.950 425.550 661.050 426.450 ;
        RECT 649.950 424.950 652.050 425.550 ;
        RECT 658.950 424.950 661.050 425.550 ;
        RECT 664.500 422.400 666.300 429.000 ;
        RECT 669.000 422.400 670.800 428.400 ;
        RECT 673.500 422.400 675.300 429.000 ;
        RECT 626.700 419.400 630.300 420.300 ;
        RECT 644.100 420.300 648.300 421.200 ;
        RECT 615.000 417.450 619.050 418.050 ;
        RECT 614.550 415.950 619.050 417.450 ;
        RECT 601.500 412.950 603.600 415.050 ;
        RECT 604.800 412.950 606.900 415.050 ;
        RECT 601.200 411.150 603.000 412.950 ;
        RECT 605.400 405.600 606.300 412.950 ;
        RECT 614.550 412.050 615.450 415.950 ;
        RECT 623.100 415.050 624.900 416.850 ;
        RECT 626.700 415.050 627.900 419.400 ;
        RECT 631.950 417.450 636.000 418.050 ;
        RECT 629.100 415.050 630.900 416.850 ;
        RECT 631.950 415.950 636.450 417.450 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 614.550 410.550 619.050 412.050 ;
        RECT 620.100 411.150 621.900 412.950 ;
        RECT 615.000 409.950 619.050 410.550 ;
        RECT 607.950 408.450 610.050 409.050 ;
        RECT 622.950 408.450 625.050 409.050 ;
        RECT 607.950 407.550 625.050 408.450 ;
        RECT 607.950 406.950 610.050 407.550 ;
        RECT 622.950 406.950 625.050 407.550 ;
        RECT 626.700 405.600 627.900 412.950 ;
        RECT 635.550 412.050 636.450 415.950 ;
        RECT 641.250 415.050 643.050 416.850 ;
        RECT 644.100 415.050 645.300 420.300 ;
        RECT 649.950 417.450 652.050 420.900 ;
        RECT 655.950 417.450 658.050 418.050 ;
        RECT 649.950 417.000 658.050 417.450 ;
        RECT 647.100 415.050 648.900 416.850 ;
        RECT 650.550 416.550 658.050 417.000 ;
        RECT 655.950 415.950 658.050 416.550 ;
        RECT 662.100 415.050 663.900 416.850 ;
        RECT 668.700 415.050 669.900 422.400 ;
        RECT 686.700 421.200 688.500 428.400 ;
        RECT 691.800 422.400 693.600 429.000 ;
        RECT 704.100 423.300 705.900 428.400 ;
        RECT 707.100 424.200 708.900 429.000 ;
        RECT 710.100 423.300 711.900 428.400 ;
        RECT 704.100 421.950 711.900 423.300 ;
        RECT 713.100 422.400 714.900 428.400 ;
        RECT 670.950 420.450 673.050 421.050 ;
        RECT 682.950 420.450 685.050 421.050 ;
        RECT 670.950 419.550 685.050 420.450 ;
        RECT 686.700 420.300 690.900 421.200 ;
        RECT 713.100 420.300 714.300 422.400 ;
        RECT 728.700 421.200 730.500 428.400 ;
        RECT 733.800 422.400 735.600 429.000 ;
        RECT 746.100 425.400 747.900 429.000 ;
        RECT 749.100 425.400 750.900 428.400 ;
        RECT 752.100 425.400 753.900 429.000 ;
        RECT 728.700 420.300 732.900 421.200 ;
        RECT 670.950 418.950 673.050 419.550 ;
        RECT 682.950 418.950 685.050 419.550 ;
        RECT 673.950 415.050 675.750 416.850 ;
        RECT 686.100 415.050 687.900 416.850 ;
        RECT 689.700 415.050 690.900 420.300 ;
        RECT 710.700 419.400 714.300 420.300 ;
        RECT 691.950 415.050 693.750 416.850 ;
        RECT 707.100 415.050 708.900 416.850 ;
        RECT 710.700 415.050 711.900 419.400 ;
        RECT 713.100 415.050 714.900 416.850 ;
        RECT 728.100 415.050 729.900 416.850 ;
        RECT 731.700 415.050 732.900 420.300 ;
        RECT 733.950 415.050 735.750 416.850 ;
        RECT 749.700 415.050 750.600 425.400 ;
        RECT 751.950 423.450 754.050 424.050 ;
        RECT 763.950 423.450 766.050 424.050 ;
        RECT 751.950 422.550 766.050 423.450 ;
        RECT 751.950 421.950 754.050 422.550 ;
        RECT 763.950 421.950 766.050 422.550 ;
        RECT 767.100 419.400 768.900 429.000 ;
        RECT 773.700 420.000 775.500 428.400 ;
        RECT 792.000 422.400 793.800 429.000 ;
        RECT 796.500 423.600 798.300 428.400 ;
        RECT 799.500 425.400 801.300 429.000 ;
        RECT 812.100 425.400 813.900 429.000 ;
        RECT 815.100 425.400 816.900 428.400 ;
        RECT 796.500 422.400 801.600 423.600 ;
        RECT 773.700 418.800 777.000 420.000 ;
        RECT 767.100 415.050 768.900 416.850 ;
        RECT 773.100 415.050 774.900 416.850 ;
        RECT 776.100 415.050 777.000 418.800 ;
        RECT 786.000 417.450 790.050 418.050 ;
        RECT 785.550 415.950 790.050 417.450 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 635.550 410.550 640.050 412.050 ;
        RECT 636.000 409.950 640.050 410.550 ;
        RECT 584.100 393.600 585.900 399.600 ;
        RECT 596.100 393.000 597.900 399.600 ;
        RECT 599.100 393.600 600.900 399.600 ;
        RECT 602.100 393.000 603.900 405.000 ;
        RECT 605.100 393.600 606.900 405.600 ;
        RECT 620.400 393.000 622.200 405.600 ;
        RECT 625.500 404.100 627.900 405.600 ;
        RECT 625.500 393.600 627.300 404.100 ;
        RECT 628.200 401.100 630.000 402.900 ;
        RECT 644.100 399.600 645.300 412.950 ;
        RECT 665.100 411.150 666.900 412.950 ;
        RECT 669.000 407.400 669.900 412.950 ;
        RECT 670.950 411.150 672.750 412.950 ;
        RECT 665.100 406.500 669.900 407.400 ;
        RECT 670.950 408.450 673.050 409.050 ;
        RECT 679.950 408.450 682.050 409.050 ;
        RECT 670.950 407.550 682.050 408.450 ;
        RECT 670.950 406.950 673.050 407.550 ;
        RECT 679.950 406.950 682.050 407.550 ;
        RECT 628.500 393.000 630.300 399.600 ;
        RECT 641.100 393.000 642.900 399.600 ;
        RECT 644.100 393.600 645.900 399.600 ;
        RECT 647.100 393.000 648.900 399.600 ;
        RECT 662.100 394.500 663.900 405.600 ;
        RECT 665.100 395.400 666.900 406.500 ;
        RECT 676.950 405.450 679.050 406.050 ;
        RECT 685.950 405.450 688.050 406.050 ;
        RECT 668.100 404.400 675.900 405.300 ;
        RECT 668.100 394.500 669.900 404.400 ;
        RECT 662.100 393.600 669.900 394.500 ;
        RECT 671.100 393.000 672.900 403.500 ;
        RECT 674.100 393.600 675.900 404.400 ;
        RECT 676.950 404.550 688.050 405.450 ;
        RECT 676.950 403.950 679.050 404.550 ;
        RECT 685.950 403.950 688.050 404.550 ;
        RECT 689.700 399.600 690.900 412.950 ;
        RECT 704.100 411.150 705.900 412.950 ;
        RECT 710.700 405.600 711.900 412.950 ;
        RECT 715.950 408.450 718.050 409.050 ;
        RECT 721.950 408.450 724.050 409.050 ;
        RECT 715.950 407.550 724.050 408.450 ;
        RECT 715.950 406.950 718.050 407.550 ;
        RECT 721.950 406.950 724.050 407.550 ;
        RECT 686.100 393.000 687.900 399.600 ;
        RECT 689.100 393.600 690.900 399.600 ;
        RECT 692.100 393.000 693.900 399.600 ;
        RECT 704.400 393.000 706.200 405.600 ;
        RECT 709.500 404.100 711.900 405.600 ;
        RECT 709.500 393.600 711.300 404.100 ;
        RECT 712.200 401.100 714.000 402.900 ;
        RECT 731.700 399.600 732.900 412.950 ;
        RECT 746.100 411.150 747.900 412.950 ;
        RECT 733.950 408.450 736.050 409.050 ;
        RECT 739.950 408.450 742.050 409.050 ;
        RECT 733.950 407.550 742.050 408.450 ;
        RECT 733.950 406.950 736.050 407.550 ;
        RECT 739.950 406.950 742.050 407.550 ;
        RECT 749.700 405.600 750.600 412.950 ;
        RECT 751.950 411.150 753.750 412.950 ;
        RECT 770.100 411.150 771.900 412.950 ;
        RECT 747.000 404.400 750.600 405.600 ;
        RECT 712.500 393.000 714.300 399.600 ;
        RECT 728.100 393.000 729.900 399.600 ;
        RECT 731.100 393.600 732.900 399.600 ;
        RECT 734.100 393.000 735.900 399.600 ;
        RECT 747.000 393.600 748.800 404.400 ;
        RECT 752.100 393.000 753.900 405.600 ;
        RECT 776.100 400.800 777.000 412.950 ;
        RECT 778.950 411.450 781.050 412.050 ;
        RECT 785.550 411.450 786.450 415.950 ;
        RECT 791.100 415.050 792.900 416.850 ;
        RECT 797.250 415.050 799.050 416.850 ;
        RECT 800.700 415.050 801.600 422.400 ;
        RECT 807.000 417.450 811.050 418.050 ;
        RECT 806.550 415.950 811.050 417.450 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 796.950 412.950 799.050 415.050 ;
        RECT 799.950 412.950 802.050 415.050 ;
        RECT 778.950 410.550 786.450 411.450 ;
        RECT 794.250 411.150 796.050 412.950 ;
        RECT 778.950 409.950 781.050 410.550 ;
        RECT 800.700 405.600 801.600 412.950 ;
        RECT 806.550 411.900 807.450 415.950 ;
        RECT 815.100 415.050 816.300 425.400 ;
        RECT 830.100 422.400 831.900 428.400 ;
        RECT 820.950 418.950 823.050 421.050 ;
        RECT 830.700 420.300 831.900 422.400 ;
        RECT 833.100 423.300 834.900 428.400 ;
        RECT 836.100 424.200 837.900 429.000 ;
        RECT 839.100 423.300 840.900 428.400 ;
        RECT 833.100 421.950 840.900 423.300 ;
        RECT 851.100 423.300 852.900 428.400 ;
        RECT 854.100 424.200 855.900 429.000 ;
        RECT 857.100 423.300 858.900 428.400 ;
        RECT 851.100 421.950 858.900 423.300 ;
        RECT 860.100 422.400 861.900 428.400 ;
        RECT 860.100 420.300 861.300 422.400 ;
        RECT 830.700 419.400 834.300 420.300 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 805.950 409.800 808.050 411.900 ;
        RECT 812.100 411.150 813.900 412.950 ;
        RECT 770.400 399.900 777.000 400.800 ;
        RECT 770.400 399.600 771.900 399.900 ;
        RECT 767.100 393.000 768.900 399.600 ;
        RECT 770.100 393.600 771.900 399.600 ;
        RECT 776.100 399.600 777.000 399.900 ;
        RECT 791.100 404.700 798.900 405.600 ;
        RECT 773.100 393.000 774.900 399.000 ;
        RECT 776.100 393.600 777.900 399.600 ;
        RECT 791.100 393.600 792.900 404.700 ;
        RECT 794.100 393.000 795.900 403.800 ;
        RECT 797.100 393.600 798.900 404.700 ;
        RECT 800.100 393.600 801.900 405.600 ;
        RECT 815.100 399.600 816.300 412.950 ;
        RECT 821.550 412.050 822.450 418.950 ;
        RECT 825.000 417.450 829.050 418.050 ;
        RECT 817.950 410.550 822.450 412.050 ;
        RECT 824.550 415.950 829.050 417.450 ;
        RECT 824.550 412.050 825.450 415.950 ;
        RECT 830.100 415.050 831.900 416.850 ;
        RECT 833.100 415.050 834.300 419.400 ;
        RECT 857.700 419.400 861.300 420.300 ;
        RECT 872.100 419.400 873.900 429.000 ;
        RECT 878.700 420.000 880.500 428.400 ;
        RECT 898.500 420.000 900.300 428.400 ;
        RECT 841.950 417.450 846.000 418.050 ;
        RECT 836.100 415.050 837.900 416.850 ;
        RECT 841.950 415.950 846.450 417.450 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 824.550 410.550 829.050 412.050 ;
        RECT 817.950 409.950 822.000 410.550 ;
        RECT 825.000 409.950 829.050 410.550 ;
        RECT 833.100 405.600 834.300 412.950 ;
        RECT 839.100 411.150 840.900 412.950 ;
        RECT 845.550 412.050 846.450 415.950 ;
        RECT 854.100 415.050 855.900 416.850 ;
        RECT 857.700 415.050 858.900 419.400 ;
        RECT 878.700 418.800 882.000 420.000 ;
        RECT 867.000 417.450 871.050 418.050 ;
        RECT 860.100 415.050 861.900 416.850 ;
        RECT 866.550 415.950 871.050 417.450 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 845.550 410.550 850.050 412.050 ;
        RECT 851.100 411.150 852.900 412.950 ;
        RECT 846.000 409.950 850.050 410.550 ;
        RECT 835.950 408.450 838.050 409.050 ;
        RECT 853.950 408.450 856.050 409.050 ;
        RECT 835.950 407.550 856.050 408.450 ;
        RECT 835.950 406.950 838.050 407.550 ;
        RECT 853.950 406.950 856.050 407.550 ;
        RECT 857.700 405.600 858.900 412.950 ;
        RECT 866.550 412.050 867.450 415.950 ;
        RECT 872.100 415.050 873.900 416.850 ;
        RECT 878.100 415.050 879.900 416.850 ;
        RECT 881.100 415.050 882.000 418.800 ;
        RECT 897.000 418.800 900.300 420.000 ;
        RECT 905.100 419.400 906.900 429.000 ;
        RECT 921.000 422.400 922.800 429.000 ;
        RECT 925.500 423.600 927.300 428.400 ;
        RECT 928.500 425.400 930.300 429.000 ;
        RECT 925.500 422.400 930.600 423.600 ;
        RECT 897.000 415.050 897.900 418.800 ;
        RECT 899.100 415.050 900.900 416.850 ;
        RECT 905.100 415.050 906.900 416.850 ;
        RECT 920.100 415.050 921.900 416.850 ;
        RECT 926.250 415.050 928.050 416.850 ;
        RECT 929.700 415.050 930.600 422.400 ;
        RECT 871.950 412.950 874.050 415.050 ;
        RECT 874.950 412.950 877.050 415.050 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 895.950 412.950 898.050 415.050 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 904.950 412.950 907.050 415.050 ;
        RECT 919.950 412.950 922.050 415.050 ;
        RECT 922.950 412.950 925.050 415.050 ;
        RECT 925.950 412.950 928.050 415.050 ;
        RECT 928.950 412.950 931.050 415.050 ;
        RECT 862.950 410.550 867.450 412.050 ;
        RECT 875.100 411.150 876.900 412.950 ;
        RECT 862.950 409.950 867.000 410.550 ;
        RECT 833.100 404.100 835.500 405.600 ;
        RECT 831.000 401.100 832.800 402.900 ;
        RECT 812.100 393.000 813.900 399.600 ;
        RECT 815.100 393.600 816.900 399.600 ;
        RECT 830.700 393.000 832.500 399.600 ;
        RECT 833.700 393.600 835.500 404.100 ;
        RECT 838.800 393.000 840.600 405.600 ;
        RECT 851.400 393.000 853.200 405.600 ;
        RECT 856.500 404.100 858.900 405.600 ;
        RECT 856.500 393.600 858.300 404.100 ;
        RECT 859.200 401.100 861.000 402.900 ;
        RECT 881.100 400.800 882.000 412.950 ;
        RECT 875.400 399.900 882.000 400.800 ;
        RECT 875.400 399.600 876.900 399.900 ;
        RECT 859.500 393.000 861.300 399.600 ;
        RECT 872.100 393.000 873.900 399.600 ;
        RECT 875.100 393.600 876.900 399.600 ;
        RECT 881.100 399.600 882.000 399.900 ;
        RECT 897.000 400.800 897.900 412.950 ;
        RECT 902.100 411.150 903.900 412.950 ;
        RECT 923.250 411.150 925.050 412.950 ;
        RECT 898.950 408.450 901.050 409.050 ;
        RECT 925.950 408.450 928.050 409.050 ;
        RECT 898.950 407.550 928.050 408.450 ;
        RECT 898.950 406.950 901.050 407.550 ;
        RECT 925.950 406.950 928.050 407.550 ;
        RECT 929.700 405.600 930.600 412.950 ;
        RECT 920.100 404.700 927.900 405.600 ;
        RECT 897.000 399.900 903.600 400.800 ;
        RECT 897.000 399.600 897.900 399.900 ;
        RECT 878.100 393.000 879.900 399.000 ;
        RECT 881.100 393.600 882.900 399.600 ;
        RECT 896.100 393.600 897.900 399.600 ;
        RECT 902.100 399.600 903.600 399.900 ;
        RECT 899.100 393.000 900.900 399.000 ;
        RECT 902.100 393.600 903.900 399.600 ;
        RECT 905.100 393.000 906.900 399.600 ;
        RECT 920.100 393.600 921.900 404.700 ;
        RECT 923.100 393.000 924.900 403.800 ;
        RECT 926.100 393.600 927.900 404.700 ;
        RECT 929.100 393.600 930.900 405.600 ;
        RECT 14.100 377.400 15.900 390.000 ;
        RECT 17.100 376.500 18.900 389.400 ;
        RECT 20.100 377.400 21.900 390.000 ;
        RECT 23.100 376.500 24.900 389.400 ;
        RECT 26.100 377.400 27.900 390.000 ;
        RECT 29.100 376.500 30.900 389.400 ;
        RECT 32.100 377.400 33.900 390.000 ;
        RECT 35.100 376.500 36.900 389.400 ;
        RECT 38.100 377.400 39.900 390.000 ;
        RECT 53.100 378.600 54.900 389.400 ;
        RECT 56.100 379.500 57.900 390.000 ;
        RECT 59.100 388.500 66.900 389.400 ;
        RECT 59.100 378.600 60.900 388.500 ;
        RECT 53.100 377.700 60.900 378.600 ;
        RECT 62.100 376.500 63.900 387.600 ;
        RECT 65.100 377.400 66.900 388.500 ;
        RECT 68.700 383.400 70.500 390.000 ;
        RECT 71.700 383.400 73.500 389.400 ;
        RECT 75.000 383.400 76.800 390.000 ;
        RECT 78.000 383.400 79.800 389.400 ;
        RECT 81.000 383.400 82.800 390.000 ;
        RECT 84.000 383.400 85.800 389.400 ;
        RECT 87.000 383.400 88.800 390.000 ;
        RECT 90.000 386.400 91.800 389.400 ;
        RECT 93.000 386.400 94.800 389.400 ;
        RECT 96.000 386.400 97.800 389.400 ;
        RECT 89.700 384.300 91.800 386.400 ;
        RECT 92.700 384.300 94.800 386.400 ;
        RECT 95.700 384.300 97.800 386.400 ;
        RECT 99.000 383.400 100.800 389.400 ;
        RECT 102.000 383.400 103.800 390.000 ;
        RECT 17.100 375.300 21.000 376.500 ;
        RECT 23.100 375.300 27.000 376.500 ;
        RECT 29.100 375.300 33.000 376.500 ;
        RECT 35.100 375.300 37.950 376.500 ;
        RECT 16.800 367.950 18.900 370.050 ;
        RECT 16.800 366.150 18.600 367.950 ;
        RECT 19.800 364.800 21.000 375.300 ;
        RECT 22.200 364.800 24.000 365.400 ;
        RECT 19.800 363.600 24.000 364.800 ;
        RECT 25.800 364.800 27.000 375.300 ;
        RECT 28.200 364.800 30.000 365.400 ;
        RECT 25.800 363.600 30.000 364.800 ;
        RECT 31.800 364.800 33.000 375.300 ;
        RECT 36.900 370.050 37.950 375.300 ;
        RECT 59.100 375.600 63.900 376.500 ;
        RECT 56.250 370.050 58.050 371.850 ;
        RECT 59.100 370.050 60.000 375.600 ;
        RECT 72.000 373.050 73.500 383.400 ;
        RECT 78.000 382.500 79.200 383.400 ;
        RECT 62.100 370.050 63.900 371.850 ;
        RECT 71.100 370.950 73.500 373.050 ;
        RECT 34.800 367.950 37.950 370.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 34.200 364.800 36.000 365.400 ;
        RECT 31.800 363.600 36.000 364.800 ;
        RECT 19.800 362.700 21.000 363.600 ;
        RECT 25.800 362.700 27.000 363.600 ;
        RECT 31.800 362.700 33.000 363.600 ;
        RECT 36.900 362.700 37.950 367.950 ;
        RECT 53.250 366.150 55.050 367.950 ;
        RECT 17.100 361.500 21.000 362.700 ;
        RECT 23.100 361.500 27.000 362.700 ;
        RECT 29.100 361.500 33.000 362.700 ;
        RECT 35.100 361.500 37.950 362.700 ;
        RECT 14.100 354.000 15.900 360.600 ;
        RECT 17.100 354.600 18.900 361.500 ;
        RECT 20.100 354.000 21.900 360.600 ;
        RECT 23.100 354.600 24.900 361.500 ;
        RECT 26.100 354.000 27.900 360.600 ;
        RECT 29.100 354.600 30.900 361.500 ;
        RECT 32.100 354.000 33.900 360.600 ;
        RECT 35.100 354.600 36.900 361.500 ;
        RECT 59.100 360.600 60.300 367.950 ;
        RECT 65.100 366.150 66.900 367.950 ;
        RECT 38.100 354.000 39.900 360.600 ;
        RECT 53.700 354.000 55.500 360.600 ;
        RECT 58.200 354.600 60.000 360.600 ;
        RECT 62.700 354.000 64.500 360.600 ;
        RECT 72.000 357.600 73.500 370.950 ;
        RECT 68.700 354.000 70.500 357.600 ;
        RECT 71.700 354.600 73.500 357.600 ;
        RECT 75.300 381.600 79.200 382.500 ;
        RECT 75.300 378.300 76.200 381.600 ;
        RECT 80.100 380.400 81.900 381.000 ;
        RECT 84.600 380.400 85.800 383.400 ;
        RECT 92.700 382.500 94.800 383.400 ;
        RECT 86.700 381.300 94.800 382.500 ;
        RECT 86.700 380.700 88.500 381.300 ;
        RECT 80.100 379.200 85.800 380.400 ;
        RECT 98.100 379.500 100.800 383.400 ;
        RECT 105.000 381.900 106.800 389.400 ;
        RECT 108.900 383.400 110.700 390.000 ;
        RECT 111.900 383.400 113.700 389.400 ;
        RECT 114.900 386.400 116.700 389.400 ;
        RECT 117.900 386.400 119.700 389.400 ;
        RECT 114.600 384.300 116.700 386.400 ;
        RECT 117.600 384.300 119.700 386.400 ;
        RECT 121.500 383.400 123.300 390.000 ;
        RECT 103.500 379.800 106.800 381.900 ;
        RECT 112.200 381.300 114.300 383.400 ;
        RECT 124.500 380.400 126.300 389.400 ;
        RECT 127.500 383.400 129.300 390.000 ;
        RECT 130.500 384.300 132.300 389.400 ;
        RECT 130.500 383.400 132.600 384.300 ;
        RECT 133.500 383.400 135.300 390.000 ;
        RECT 131.700 382.500 132.600 383.400 ;
        RECT 131.700 381.600 135.300 382.500 ;
        RECT 129.000 380.400 130.800 380.700 ;
        RECT 89.700 378.300 91.800 379.500 ;
        RECT 75.300 377.400 91.800 378.300 ;
        RECT 95.100 378.600 97.200 379.500 ;
        RECT 111.600 379.200 130.800 380.400 ;
        RECT 111.600 378.600 112.800 379.200 ;
        RECT 129.000 378.900 130.800 379.200 ;
        RECT 95.100 377.400 112.800 378.600 ;
        RECT 115.500 377.700 117.600 378.300 ;
        RECT 125.700 377.700 127.500 378.300 ;
        RECT 75.300 360.600 76.200 377.400 ;
        RECT 115.500 376.500 127.500 377.700 ;
        RECT 77.100 375.300 112.800 376.500 ;
        RECT 115.500 376.200 117.600 376.500 ;
        RECT 77.100 374.700 78.900 375.300 ;
        RECT 111.600 374.700 112.800 375.300 ;
        RECT 80.100 370.950 82.200 373.050 ;
        RECT 80.700 368.100 82.200 370.950 ;
        RECT 84.300 370.800 89.400 372.600 ;
        RECT 88.500 369.300 89.400 370.800 ;
        RECT 92.100 372.300 93.900 374.100 ;
        RECT 98.100 373.800 100.200 374.100 ;
        RECT 111.600 373.800 125.100 374.700 ;
        RECT 92.100 371.100 93.000 372.300 ;
        RECT 98.100 372.000 102.000 373.800 ;
        RECT 103.500 372.300 105.600 373.200 ;
        RECT 123.300 373.050 125.100 373.800 ;
        RECT 103.500 371.100 114.600 372.300 ;
        RECT 123.300 371.250 127.200 373.050 ;
        RECT 92.100 370.200 105.600 371.100 ;
        RECT 112.800 370.500 114.600 371.100 ;
        RECT 125.100 370.950 127.200 371.250 ;
        RECT 131.100 370.950 133.200 373.050 ;
        RECT 131.100 369.300 132.900 370.950 ;
        RECT 88.500 368.100 132.900 369.300 ;
        RECT 80.700 366.600 87.300 368.100 ;
        RECT 77.100 363.900 84.900 365.700 ;
        RECT 85.800 365.100 102.900 366.600 ;
        RECT 100.800 364.500 102.900 365.100 ;
        RECT 107.100 366.000 109.200 367.050 ;
        RECT 107.100 365.100 112.200 366.000 ;
        RECT 115.800 365.400 117.600 367.200 ;
        RECT 134.100 365.400 135.300 381.600 ;
        RECT 146.100 377.400 147.900 389.400 ;
        RECT 149.100 378.300 150.900 389.400 ;
        RECT 152.100 379.200 153.900 390.000 ;
        RECT 155.100 378.300 156.900 389.400 ;
        RECT 170.100 383.400 171.900 390.000 ;
        RECT 173.100 383.400 174.900 389.400 ;
        RECT 149.100 377.400 156.900 378.300 ;
        RECT 146.400 370.050 147.300 377.400 ;
        RECT 151.950 370.050 153.750 371.850 ;
        RECT 170.100 370.050 171.900 371.850 ;
        RECT 173.100 370.050 174.300 383.400 ;
        RECT 185.100 378.600 186.900 389.400 ;
        RECT 188.100 379.500 189.900 390.000 ;
        RECT 191.100 388.500 198.900 389.400 ;
        RECT 191.100 378.600 192.900 388.500 ;
        RECT 185.100 377.700 192.900 378.600 ;
        RECT 194.100 376.500 195.900 387.600 ;
        RECT 197.100 377.400 198.900 388.500 ;
        RECT 212.100 383.400 213.900 389.400 ;
        RECT 215.100 383.400 216.900 390.000 ;
        RECT 230.100 383.400 231.900 390.000 ;
        RECT 233.100 383.400 234.900 389.400 ;
        RECT 236.100 383.400 237.900 390.000 ;
        RECT 248.100 383.400 249.900 389.400 ;
        RECT 251.100 383.400 252.900 390.000 ;
        RECT 191.100 375.600 195.900 376.500 ;
        RECT 180.000 372.450 184.050 373.050 ;
        RECT 179.550 370.950 184.050 372.450 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 148.950 367.950 151.050 370.050 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 107.100 364.950 109.200 365.100 ;
        RECT 83.400 360.600 84.900 363.900 ;
        RECT 101.100 362.700 102.900 364.500 ;
        RECT 110.400 364.200 112.200 365.100 ;
        RECT 116.700 362.400 117.600 365.400 ;
        RECT 118.500 364.200 135.300 365.400 ;
        RECT 118.500 363.300 120.600 364.200 ;
        RECT 129.300 362.700 131.100 363.300 ;
        RECT 89.100 360.600 95.700 362.400 ;
        RECT 110.400 361.200 117.600 362.400 ;
        RECT 122.700 361.500 131.100 362.700 ;
        RECT 110.400 360.600 111.300 361.200 ;
        RECT 113.400 360.600 115.200 361.200 ;
        RECT 122.700 360.600 124.200 361.500 ;
        RECT 134.100 360.600 135.300 364.200 ;
        RECT 75.300 354.600 77.100 360.600 ;
        RECT 80.700 354.000 82.500 360.600 ;
        RECT 83.400 359.400 87.600 360.600 ;
        RECT 85.800 354.600 87.600 359.400 ;
        RECT 89.700 357.600 91.800 359.700 ;
        RECT 92.700 357.600 94.800 359.700 ;
        RECT 95.700 357.600 97.800 359.700 ;
        RECT 98.700 357.600 100.800 359.700 ;
        RECT 104.100 358.500 106.800 360.600 ;
        RECT 108.600 359.400 111.300 360.600 ;
        RECT 108.600 358.500 110.400 359.400 ;
        RECT 90.000 354.600 91.800 357.600 ;
        RECT 93.000 354.600 94.800 357.600 ;
        RECT 96.000 354.600 97.800 357.600 ;
        RECT 99.000 354.600 100.800 357.600 ;
        RECT 102.000 354.000 103.800 357.600 ;
        RECT 105.000 354.600 106.800 358.500 ;
        RECT 112.200 357.600 114.300 359.700 ;
        RECT 115.200 357.600 117.300 359.700 ;
        RECT 118.200 357.600 120.300 359.700 ;
        RECT 109.500 354.000 111.300 357.600 ;
        RECT 112.500 354.600 114.300 357.600 ;
        RECT 115.500 354.600 117.300 357.600 ;
        RECT 118.500 354.600 120.300 357.600 ;
        RECT 122.700 354.600 124.500 360.600 ;
        RECT 128.100 354.000 129.900 360.600 ;
        RECT 133.500 354.600 135.300 360.600 ;
        RECT 146.400 360.600 147.300 367.950 ;
        RECT 148.950 366.150 150.750 367.950 ;
        RECT 155.100 366.150 156.900 367.950 ;
        RECT 146.400 359.400 151.500 360.600 ;
        RECT 146.700 354.000 148.500 357.600 ;
        RECT 149.700 354.600 151.500 359.400 ;
        RECT 154.200 354.000 156.000 360.600 ;
        RECT 173.100 357.600 174.300 367.950 ;
        RECT 179.550 367.050 180.450 370.950 ;
        RECT 188.250 370.050 190.050 371.850 ;
        RECT 191.100 370.050 192.000 375.600 ;
        RECT 196.950 375.450 199.050 376.200 ;
        RECT 196.950 374.550 204.450 375.450 ;
        RECT 196.950 374.100 199.050 374.550 ;
        RECT 194.100 370.050 195.900 371.850 ;
        RECT 184.950 367.950 187.050 370.050 ;
        RECT 187.950 367.950 190.050 370.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 175.950 365.550 180.450 367.050 ;
        RECT 185.250 366.150 187.050 367.950 ;
        RECT 175.950 364.950 180.000 365.550 ;
        RECT 191.100 360.600 192.300 367.950 ;
        RECT 197.100 366.150 198.900 367.950 ;
        RECT 203.550 366.450 204.450 374.550 ;
        RECT 212.700 370.050 213.900 383.400 ;
        RECT 217.950 372.450 222.000 373.050 ;
        RECT 215.100 370.050 216.900 371.850 ;
        RECT 217.950 370.950 222.450 372.450 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 200.550 365.550 204.450 366.450 ;
        RECT 193.950 363.450 196.050 364.050 ;
        RECT 200.550 363.450 201.450 365.550 ;
        RECT 193.950 362.550 201.450 363.450 ;
        RECT 193.950 361.950 196.050 362.550 ;
        RECT 170.100 354.000 171.900 357.600 ;
        RECT 173.100 354.600 174.900 357.600 ;
        RECT 185.700 354.000 187.500 360.600 ;
        RECT 190.200 354.600 192.000 360.600 ;
        RECT 194.700 354.000 196.500 360.600 ;
        RECT 212.700 357.600 213.900 367.950 ;
        RECT 221.550 364.050 222.450 370.950 ;
        RECT 233.700 370.050 234.900 383.400 ;
        RECT 248.700 370.050 249.900 383.400 ;
        RECT 263.400 377.400 265.200 390.000 ;
        RECT 268.500 378.900 270.300 389.400 ;
        RECT 271.500 383.400 273.300 390.000 ;
        RECT 271.200 380.100 273.000 381.900 ;
        RECT 268.500 377.400 270.900 378.900 ;
        RECT 287.400 377.400 289.200 390.000 ;
        RECT 292.500 378.900 294.300 389.400 ;
        RECT 295.500 383.400 297.300 390.000 ;
        RECT 308.100 383.400 309.900 390.000 ;
        RECT 311.100 383.400 312.900 389.400 ;
        RECT 314.100 383.400 315.900 390.000 ;
        RECT 326.700 383.400 328.500 390.000 ;
        RECT 295.200 380.100 297.000 381.900 ;
        RECT 292.500 377.400 294.900 378.900 ;
        RECT 251.100 370.050 252.900 371.850 ;
        RECT 263.100 370.050 264.900 371.850 ;
        RECT 269.700 370.050 270.900 377.400 ;
        RECT 287.100 370.050 288.900 371.850 ;
        RECT 293.700 370.050 294.900 377.400 ;
        RECT 311.700 370.050 312.900 383.400 ;
        RECT 327.000 380.100 328.800 381.900 ;
        RECT 329.700 378.900 331.500 389.400 ;
        RECT 329.100 377.400 331.500 378.900 ;
        RECT 334.800 377.400 336.600 390.000 ;
        RECT 347.100 377.400 348.900 390.000 ;
        RECT 350.100 377.400 351.900 389.400 ;
        RECT 362.100 383.400 363.900 390.000 ;
        RECT 365.100 383.400 366.900 389.400 ;
        RECT 313.950 375.450 316.050 376.050 ;
        RECT 319.950 375.450 322.050 376.050 ;
        RECT 313.950 374.550 322.050 375.450 ;
        RECT 313.950 373.950 316.050 374.550 ;
        RECT 319.950 373.950 322.050 374.550 ;
        RECT 329.100 370.050 330.300 377.400 ;
        RECT 335.100 370.050 336.900 371.850 ;
        RECT 350.100 370.050 351.300 377.400 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 247.950 367.950 250.050 370.050 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 295.950 367.950 298.050 370.050 ;
        RECT 307.950 367.950 310.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 328.950 367.950 331.050 370.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 349.950 367.950 352.050 370.050 ;
        RECT 362.100 367.950 364.200 370.050 ;
        RECT 230.100 366.150 231.900 367.950 ;
        RECT 220.950 361.950 223.050 364.050 ;
        RECT 233.700 362.700 234.900 367.950 ;
        RECT 235.950 366.150 237.750 367.950 ;
        RECT 230.700 361.800 234.900 362.700 ;
        RECT 212.100 354.600 213.900 357.600 ;
        RECT 215.100 354.000 216.900 357.600 ;
        RECT 230.700 354.600 232.500 361.800 ;
        RECT 235.800 354.000 237.600 360.600 ;
        RECT 248.700 357.600 249.900 367.950 ;
        RECT 266.100 366.150 267.900 367.950 ;
        RECT 269.700 363.600 270.900 367.950 ;
        RECT 272.100 366.150 273.900 367.950 ;
        RECT 290.100 366.150 291.900 367.950 ;
        RECT 293.700 363.600 294.900 367.950 ;
        RECT 296.100 366.150 297.900 367.950 ;
        RECT 308.100 366.150 309.900 367.950 ;
        RECT 269.700 362.700 273.300 363.600 ;
        RECT 293.700 362.700 297.300 363.600 ;
        RECT 311.700 362.700 312.900 367.950 ;
        RECT 313.950 366.150 315.750 367.950 ;
        RECT 326.100 366.150 327.900 367.950 ;
        RECT 263.100 359.700 270.900 361.050 ;
        RECT 248.100 354.600 249.900 357.600 ;
        RECT 251.100 354.000 252.900 357.600 ;
        RECT 263.100 354.600 264.900 359.700 ;
        RECT 266.100 354.000 267.900 358.800 ;
        RECT 269.100 354.600 270.900 359.700 ;
        RECT 272.100 360.600 273.300 362.700 ;
        RECT 272.100 354.600 273.900 360.600 ;
        RECT 287.100 359.700 294.900 361.050 ;
        RECT 287.100 354.600 288.900 359.700 ;
        RECT 290.100 354.000 291.900 358.800 ;
        RECT 293.100 354.600 294.900 359.700 ;
        RECT 296.100 360.600 297.300 362.700 ;
        RECT 308.700 361.800 312.900 362.700 ;
        RECT 313.950 363.450 316.050 364.050 ;
        RECT 319.950 363.450 322.050 364.050 ;
        RECT 329.100 363.600 330.300 367.950 ;
        RECT 332.100 366.150 333.900 367.950 ;
        RECT 347.100 366.150 348.900 367.950 ;
        RECT 313.950 362.550 322.050 363.450 ;
        RECT 313.950 361.950 316.050 362.550 ;
        RECT 319.950 361.950 322.050 362.550 ;
        RECT 326.700 362.700 330.300 363.600 ;
        RECT 296.100 354.600 297.900 360.600 ;
        RECT 308.700 354.600 310.500 361.800 ;
        RECT 326.700 360.600 327.900 362.700 ;
        RECT 313.800 354.000 315.600 360.600 ;
        RECT 326.100 354.600 327.900 360.600 ;
        RECT 329.100 359.700 336.900 361.050 ;
        RECT 350.100 360.600 351.300 367.950 ;
        RECT 362.250 366.150 364.050 367.950 ;
        RECT 365.100 363.300 366.000 383.400 ;
        RECT 368.100 378.000 369.900 390.000 ;
        RECT 371.100 377.400 372.900 389.400 ;
        RECT 386.400 377.400 388.200 390.000 ;
        RECT 391.500 378.900 393.300 389.400 ;
        RECT 394.500 383.400 396.300 390.000 ;
        RECT 410.100 383.400 411.900 390.000 ;
        RECT 413.100 383.400 414.900 389.400 ;
        RECT 394.200 380.100 396.000 381.900 ;
        RECT 391.500 377.400 393.900 378.900 ;
        RECT 367.200 370.050 369.000 371.850 ;
        RECT 371.400 370.050 372.300 377.400 ;
        RECT 386.100 370.050 387.900 371.850 ;
        RECT 392.700 370.050 393.900 377.400 ;
        RECT 367.500 367.950 369.600 370.050 ;
        RECT 370.800 367.950 372.900 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 394.950 367.950 397.050 370.050 ;
        RECT 410.100 367.950 412.200 370.050 ;
        RECT 362.100 362.400 370.500 363.300 ;
        RECT 329.100 354.600 330.900 359.700 ;
        RECT 332.100 354.000 333.900 358.800 ;
        RECT 335.100 354.600 336.900 359.700 ;
        RECT 347.100 354.000 348.900 360.600 ;
        RECT 350.100 354.600 351.900 360.600 ;
        RECT 362.100 354.600 363.900 362.400 ;
        RECT 368.700 361.500 370.500 362.400 ;
        RECT 371.400 360.600 372.300 367.950 ;
        RECT 389.100 366.150 390.900 367.950 ;
        RECT 392.700 363.600 393.900 367.950 ;
        RECT 395.100 366.150 396.900 367.950 ;
        RECT 410.250 366.150 412.050 367.950 ;
        RECT 392.700 362.700 396.300 363.600 ;
        RECT 413.100 363.300 414.000 383.400 ;
        RECT 416.100 378.000 417.900 390.000 ;
        RECT 419.100 377.400 420.900 389.400 ;
        RECT 431.100 383.400 432.900 390.000 ;
        RECT 434.100 383.400 435.900 389.400 ;
        RECT 437.100 383.400 438.900 390.000 ;
        RECT 449.700 383.400 451.500 390.000 ;
        RECT 415.200 370.050 417.000 371.850 ;
        RECT 419.400 370.050 420.300 377.400 ;
        RECT 434.100 370.050 435.300 383.400 ;
        RECT 450.000 380.100 451.800 381.900 ;
        RECT 452.700 378.900 454.500 389.400 ;
        RECT 452.100 377.400 454.500 378.900 ;
        RECT 457.800 377.400 459.600 390.000 ;
        RECT 473.400 377.400 475.200 390.000 ;
        RECT 478.500 378.900 480.300 389.400 ;
        RECT 481.500 383.400 483.300 390.000 ;
        RECT 494.100 383.400 495.900 390.000 ;
        RECT 497.100 383.400 498.900 389.400 ;
        RECT 500.100 383.400 501.900 390.000 ;
        RECT 481.200 380.100 483.000 381.900 ;
        RECT 478.500 377.400 480.900 378.900 ;
        RECT 452.100 370.050 453.300 377.400 ;
        RECT 458.100 370.050 459.900 371.850 ;
        RECT 473.100 370.050 474.900 371.850 ;
        RECT 479.700 370.050 480.900 377.400 ;
        RECT 497.100 370.050 498.300 383.400 ;
        RECT 512.100 377.400 513.900 389.400 ;
        RECT 515.100 378.000 516.900 390.000 ;
        RECT 518.100 383.400 519.900 389.400 ;
        RECT 521.100 383.400 522.900 390.000 ;
        RECT 536.700 383.400 538.500 390.000 ;
        RECT 512.700 370.050 513.600 377.400 ;
        RECT 516.000 370.050 517.800 371.850 ;
        RECT 415.500 367.950 417.600 370.050 ;
        RECT 418.800 367.950 420.900 370.050 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 512.100 367.950 514.200 370.050 ;
        RECT 515.400 367.950 517.500 370.050 ;
        RECT 366.600 354.000 368.400 360.600 ;
        RECT 369.600 358.800 372.300 360.600 ;
        RECT 386.100 359.700 393.900 361.050 ;
        RECT 369.600 354.600 371.400 358.800 ;
        RECT 386.100 354.600 387.900 359.700 ;
        RECT 389.100 354.000 390.900 358.800 ;
        RECT 392.100 354.600 393.900 359.700 ;
        RECT 395.100 360.600 396.300 362.700 ;
        RECT 410.100 362.400 418.500 363.300 ;
        RECT 395.100 354.600 396.900 360.600 ;
        RECT 410.100 354.600 411.900 362.400 ;
        RECT 416.700 361.500 418.500 362.400 ;
        RECT 419.400 360.600 420.300 367.950 ;
        RECT 431.250 366.150 433.050 367.950 ;
        RECT 434.100 362.700 435.300 367.950 ;
        RECT 437.100 366.150 438.900 367.950 ;
        RECT 449.100 366.150 450.900 367.950 ;
        RECT 452.100 363.600 453.300 367.950 ;
        RECT 455.100 366.150 456.900 367.950 ;
        RECT 476.100 366.150 477.900 367.950 ;
        RECT 449.700 362.700 453.300 363.600 ;
        RECT 479.700 363.600 480.900 367.950 ;
        RECT 482.100 366.150 483.900 367.950 ;
        RECT 494.250 366.150 496.050 367.950 ;
        RECT 479.700 362.700 483.300 363.600 ;
        RECT 434.100 361.800 438.300 362.700 ;
        RECT 414.600 354.000 416.400 360.600 ;
        RECT 417.600 358.800 420.300 360.600 ;
        RECT 417.600 354.600 419.400 358.800 ;
        RECT 431.400 354.000 433.200 360.600 ;
        RECT 436.500 354.600 438.300 361.800 ;
        RECT 449.700 360.600 450.900 362.700 ;
        RECT 449.100 354.600 450.900 360.600 ;
        RECT 452.100 359.700 459.900 361.050 ;
        RECT 452.100 354.600 453.900 359.700 ;
        RECT 455.100 354.000 456.900 358.800 ;
        RECT 458.100 354.600 459.900 359.700 ;
        RECT 473.100 359.700 480.900 361.050 ;
        RECT 473.100 354.600 474.900 359.700 ;
        RECT 476.100 354.000 477.900 358.800 ;
        RECT 479.100 354.600 480.900 359.700 ;
        RECT 482.100 360.600 483.300 362.700 ;
        RECT 497.100 362.700 498.300 367.950 ;
        RECT 500.100 366.150 501.900 367.950 ;
        RECT 497.100 361.800 501.300 362.700 ;
        RECT 482.100 354.600 483.900 360.600 ;
        RECT 494.400 354.000 496.200 360.600 ;
        RECT 499.500 354.600 501.300 361.800 ;
        RECT 512.700 360.600 513.600 367.950 ;
        RECT 519.000 363.300 519.900 383.400 ;
        RECT 537.000 380.100 538.800 381.900 ;
        RECT 539.700 378.900 541.500 389.400 ;
        RECT 539.100 377.400 541.500 378.900 ;
        RECT 544.800 377.400 546.600 390.000 ;
        RECT 560.100 383.400 561.900 390.000 ;
        RECT 563.100 383.400 564.900 389.400 ;
        RECT 566.100 383.400 567.900 390.000 ;
        RECT 578.100 383.400 579.900 390.000 ;
        RECT 581.100 383.400 582.900 389.400 ;
        RECT 531.000 372.450 535.050 373.050 ;
        RECT 530.550 370.950 535.050 372.450 ;
        RECT 520.800 367.950 522.900 370.050 ;
        RECT 520.950 366.150 522.750 367.950 ;
        RECT 530.550 367.050 531.450 370.950 ;
        RECT 539.100 370.050 540.300 377.400 ;
        RECT 544.950 375.450 547.050 376.050 ;
        RECT 559.950 375.450 562.050 376.200 ;
        RECT 544.950 374.550 562.050 375.450 ;
        RECT 544.950 373.950 547.050 374.550 ;
        RECT 559.950 374.100 562.050 374.550 ;
        RECT 545.100 370.050 546.900 371.850 ;
        RECT 563.700 370.050 564.900 383.400 ;
        RECT 568.950 375.450 571.050 376.050 ;
        RECT 574.950 375.450 577.050 376.050 ;
        RECT 568.950 374.550 577.050 375.450 ;
        RECT 568.950 373.950 571.050 374.550 ;
        RECT 574.950 373.950 577.050 374.550 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 578.100 367.950 580.200 370.050 ;
        RECT 530.550 365.550 535.050 367.050 ;
        RECT 536.100 366.150 537.900 367.950 ;
        RECT 531.000 364.950 535.050 365.550 ;
        RECT 539.100 363.600 540.300 367.950 ;
        RECT 542.100 366.150 543.900 367.950 ;
        RECT 560.100 366.150 561.900 367.950 ;
        RECT 514.500 362.400 522.900 363.300 ;
        RECT 514.500 361.500 516.300 362.400 ;
        RECT 512.700 358.800 515.400 360.600 ;
        RECT 513.600 354.600 515.400 358.800 ;
        RECT 516.600 354.000 518.400 360.600 ;
        RECT 521.100 354.600 522.900 362.400 ;
        RECT 536.700 362.700 540.300 363.600 ;
        RECT 563.700 362.700 564.900 367.950 ;
        RECT 565.950 366.150 567.750 367.950 ;
        RECT 578.250 366.150 580.050 367.950 ;
        RECT 581.100 363.300 582.000 383.400 ;
        RECT 584.100 378.000 585.900 390.000 ;
        RECT 587.100 377.400 588.900 389.400 ;
        RECT 602.400 377.400 604.200 390.000 ;
        RECT 607.500 378.900 609.300 389.400 ;
        RECT 610.500 383.400 612.300 390.000 ;
        RECT 610.200 380.100 612.000 381.900 ;
        RECT 607.500 377.400 609.900 378.900 ;
        RECT 618.000 378.450 622.050 379.050 ;
        RECT 583.200 370.050 585.000 371.850 ;
        RECT 587.400 370.050 588.300 377.400 ;
        RECT 602.100 370.050 603.900 371.850 ;
        RECT 608.700 370.050 609.900 377.400 ;
        RECT 617.550 376.950 622.050 378.450 ;
        RECT 623.400 377.400 625.200 390.000 ;
        RECT 628.500 378.900 630.300 389.400 ;
        RECT 631.500 383.400 633.300 390.000 ;
        RECT 644.100 383.400 645.900 390.000 ;
        RECT 647.100 383.400 648.900 389.400 ;
        RECT 650.100 383.400 651.900 390.000 ;
        RECT 662.100 383.400 663.900 390.000 ;
        RECT 665.100 383.400 666.900 389.400 ;
        RECT 668.100 383.400 669.900 390.000 ;
        RECT 683.100 388.500 690.900 389.400 ;
        RECT 631.200 380.100 633.000 381.900 ;
        RECT 628.500 377.400 630.900 378.900 ;
        RECT 583.500 367.950 585.600 370.050 ;
        RECT 586.800 367.950 588.900 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 610.950 367.950 613.050 370.050 ;
        RECT 536.700 360.600 537.900 362.700 ;
        RECT 560.700 361.800 564.900 362.700 ;
        RECT 578.100 362.400 586.500 363.300 ;
        RECT 536.100 354.600 537.900 360.600 ;
        RECT 539.100 359.700 546.900 361.050 ;
        RECT 539.100 354.600 540.900 359.700 ;
        RECT 542.100 354.000 543.900 358.800 ;
        RECT 545.100 354.600 546.900 359.700 ;
        RECT 560.700 354.600 562.500 361.800 ;
        RECT 565.800 354.000 567.600 360.600 ;
        RECT 578.100 354.600 579.900 362.400 ;
        RECT 584.700 361.500 586.500 362.400 ;
        RECT 587.400 360.600 588.300 367.950 ;
        RECT 605.100 366.150 606.900 367.950 ;
        RECT 608.700 363.600 609.900 367.950 ;
        RECT 611.100 366.150 612.900 367.950 ;
        RECT 617.550 367.050 618.450 376.950 ;
        RECT 623.100 370.050 624.900 371.850 ;
        RECT 629.700 370.050 630.900 377.400 ;
        RECT 631.950 375.450 634.050 375.900 ;
        RECT 631.950 374.550 639.450 375.450 ;
        RECT 631.950 373.800 634.050 374.550 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 617.550 365.550 622.050 367.050 ;
        RECT 626.100 366.150 627.900 367.950 ;
        RECT 618.000 364.950 622.050 365.550 ;
        RECT 629.700 363.600 630.900 367.950 ;
        RECT 632.100 366.150 633.900 367.950 ;
        RECT 638.550 367.050 639.450 374.550 ;
        RECT 647.700 370.050 648.900 383.400 ;
        RECT 665.700 370.050 666.900 383.400 ;
        RECT 683.100 377.400 684.900 388.500 ;
        RECT 686.100 376.500 687.900 387.600 ;
        RECT 689.100 378.600 690.900 388.500 ;
        RECT 692.100 379.500 693.900 390.000 ;
        RECT 695.100 378.600 696.900 389.400 ;
        RECT 707.100 383.400 708.900 390.000 ;
        RECT 710.100 383.400 711.900 389.400 ;
        RECT 713.100 384.000 714.900 390.000 ;
        RECT 710.400 383.100 711.900 383.400 ;
        RECT 716.100 383.400 717.900 389.400 ;
        RECT 718.950 387.450 721.050 387.900 ;
        RECT 724.950 387.450 727.050 388.050 ;
        RECT 718.950 386.550 727.050 387.450 ;
        RECT 718.950 385.800 721.050 386.550 ;
        RECT 724.950 385.950 727.050 386.550 ;
        RECT 716.100 383.100 717.000 383.400 ;
        RECT 710.400 382.200 717.000 383.100 ;
        RECT 689.100 377.700 696.900 378.600 ;
        RECT 686.100 375.600 690.900 376.500 ;
        RECT 670.950 372.450 675.000 373.050 ;
        RECT 670.950 370.950 675.450 372.450 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 638.550 365.550 643.050 367.050 ;
        RECT 644.100 366.150 645.900 367.950 ;
        RECT 639.000 364.950 643.050 365.550 ;
        RECT 608.700 362.700 612.300 363.600 ;
        RECT 629.700 362.700 633.300 363.600 ;
        RECT 647.700 362.700 648.900 367.950 ;
        RECT 649.950 366.150 651.750 367.950 ;
        RECT 662.100 366.150 663.900 367.950 ;
        RECT 665.700 362.700 666.900 367.950 ;
        RECT 667.950 366.150 669.750 367.950 ;
        RECT 674.550 367.050 675.450 370.950 ;
        RECT 686.100 370.050 687.900 371.850 ;
        RECT 690.000 370.050 690.900 375.600 ;
        RECT 697.950 372.450 702.000 373.050 ;
        RECT 691.950 370.050 693.750 371.850 ;
        RECT 697.950 370.950 702.450 372.450 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 670.950 365.550 675.450 367.050 ;
        RECT 683.100 366.150 684.900 367.950 ;
        RECT 670.950 364.950 675.000 365.550 ;
        RECT 582.600 354.000 584.400 360.600 ;
        RECT 585.600 358.800 588.300 360.600 ;
        RECT 602.100 359.700 609.900 361.050 ;
        RECT 585.600 354.600 587.400 358.800 ;
        RECT 602.100 354.600 603.900 359.700 ;
        RECT 605.100 354.000 606.900 358.800 ;
        RECT 608.100 354.600 609.900 359.700 ;
        RECT 611.100 360.600 612.300 362.700 ;
        RECT 611.100 354.600 612.900 360.600 ;
        RECT 623.100 359.700 630.900 361.050 ;
        RECT 623.100 354.600 624.900 359.700 ;
        RECT 626.100 354.000 627.900 358.800 ;
        RECT 629.100 354.600 630.900 359.700 ;
        RECT 632.100 360.600 633.300 362.700 ;
        RECT 644.700 361.800 648.900 362.700 ;
        RECT 662.700 361.800 666.900 362.700 ;
        RECT 632.100 354.600 633.900 360.600 ;
        RECT 644.700 354.600 646.500 361.800 ;
        RECT 649.800 354.000 651.600 360.600 ;
        RECT 662.700 354.600 664.500 361.800 ;
        RECT 689.700 360.600 690.900 367.950 ;
        RECT 694.950 366.150 696.750 367.950 ;
        RECT 701.550 367.050 702.450 370.950 ;
        RECT 710.100 370.050 711.900 371.850 ;
        RECT 716.100 370.050 717.000 382.200 ;
        RECT 732.000 378.600 733.800 389.400 ;
        RECT 732.000 377.400 735.600 378.600 ;
        RECT 737.100 377.400 738.900 390.000 ;
        RECT 749.100 383.400 750.900 389.400 ;
        RECT 752.100 383.400 753.900 390.000 ;
        RECT 767.100 383.400 768.900 390.000 ;
        RECT 770.100 383.400 771.900 389.400 ;
        RECT 773.100 384.000 774.900 390.000 ;
        RECT 731.100 370.050 732.900 371.850 ;
        RECT 734.700 370.050 735.600 377.400 ;
        RECT 736.950 370.050 738.750 371.850 ;
        RECT 749.700 370.050 750.900 383.400 ;
        RECT 770.400 383.100 771.900 383.400 ;
        RECT 776.100 383.400 777.900 389.400 ;
        RECT 788.700 383.400 790.500 390.000 ;
        RECT 776.100 383.100 777.000 383.400 ;
        RECT 770.400 382.200 777.000 383.100 ;
        RECT 752.100 370.050 753.900 371.850 ;
        RECT 770.100 370.050 771.900 371.850 ;
        RECT 776.100 370.050 777.000 382.200 ;
        RECT 789.000 380.100 790.800 381.900 ;
        RECT 791.700 378.900 793.500 389.400 ;
        RECT 791.100 377.400 793.500 378.900 ;
        RECT 796.800 377.400 798.600 390.000 ;
        RECT 809.400 377.400 811.200 390.000 ;
        RECT 814.500 378.900 816.300 389.400 ;
        RECT 817.500 383.400 819.300 390.000 ;
        RECT 830.100 388.500 837.900 389.400 ;
        RECT 817.200 380.100 819.000 381.900 ;
        RECT 814.500 377.400 816.900 378.900 ;
        RECT 830.100 377.400 831.900 388.500 ;
        RECT 791.100 370.050 792.300 377.400 ;
        RECT 807.000 375.450 811.050 376.050 ;
        RECT 806.550 373.950 811.050 375.450 ;
        RECT 806.550 372.450 807.450 373.950 ;
        RECT 797.100 370.050 798.900 371.850 ;
        RECT 803.550 371.550 807.450 372.450 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 709.950 367.950 712.050 370.050 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 769.950 367.950 772.050 370.050 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 790.950 367.950 793.050 370.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 701.550 365.550 706.050 367.050 ;
        RECT 707.100 366.150 708.900 367.950 ;
        RECT 713.100 366.150 714.900 367.950 ;
        RECT 702.000 364.950 706.050 365.550 ;
        RECT 716.100 364.200 717.000 367.950 ;
        RECT 667.800 354.000 669.600 360.600 ;
        RECT 685.500 354.000 687.300 360.600 ;
        RECT 690.000 354.600 691.800 360.600 ;
        RECT 694.500 354.000 696.300 360.600 ;
        RECT 707.100 354.000 708.900 363.600 ;
        RECT 713.700 363.000 717.000 364.200 ;
        RECT 718.950 363.450 721.050 364.050 ;
        RECT 730.950 363.450 733.050 364.050 ;
        RECT 713.700 354.600 715.500 363.000 ;
        RECT 718.950 362.550 733.050 363.450 ;
        RECT 718.950 361.950 721.050 362.550 ;
        RECT 730.950 361.950 733.050 362.550 ;
        RECT 734.700 357.600 735.600 367.950 ;
        RECT 749.700 357.600 750.900 367.950 ;
        RECT 767.100 366.150 768.900 367.950 ;
        RECT 773.100 366.150 774.900 367.950 ;
        RECT 776.100 364.200 777.000 367.950 ;
        RECT 788.100 366.150 789.900 367.950 ;
        RECT 731.100 354.000 732.900 357.600 ;
        RECT 734.100 354.600 735.900 357.600 ;
        RECT 737.100 354.000 738.900 357.600 ;
        RECT 749.100 354.600 750.900 357.600 ;
        RECT 752.100 354.000 753.900 357.600 ;
        RECT 767.100 354.000 768.900 363.600 ;
        RECT 773.700 363.000 777.000 364.200 ;
        RECT 791.100 363.600 792.300 367.950 ;
        RECT 794.100 366.150 795.900 367.950 ;
        RECT 803.550 367.050 804.450 371.550 ;
        RECT 809.100 370.050 810.900 371.850 ;
        RECT 815.700 370.050 816.900 377.400 ;
        RECT 833.100 376.500 834.900 387.600 ;
        RECT 836.100 378.600 837.900 388.500 ;
        RECT 839.100 379.500 840.900 390.000 ;
        RECT 842.100 378.600 843.900 389.400 ;
        RECT 836.100 377.700 843.900 378.600 ;
        RECT 857.400 377.400 859.200 390.000 ;
        RECT 862.500 378.900 864.300 389.400 ;
        RECT 865.500 383.400 867.300 390.000 ;
        RECT 881.100 383.400 882.900 389.400 ;
        RECT 884.100 384.000 885.900 390.000 ;
        RECT 882.000 383.100 882.900 383.400 ;
        RECT 887.100 383.400 888.900 389.400 ;
        RECT 890.100 383.400 891.900 390.000 ;
        RECT 887.100 383.100 888.600 383.400 ;
        RECT 882.000 382.200 888.600 383.100 ;
        RECT 865.200 380.100 867.000 381.900 ;
        RECT 862.500 377.400 864.900 378.900 ;
        RECT 817.950 375.450 820.050 376.200 ;
        RECT 833.100 375.600 837.900 376.500 ;
        RECT 817.950 374.550 825.450 375.450 ;
        RECT 817.950 374.100 820.050 374.550 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 803.550 365.550 808.050 367.050 ;
        RECT 812.100 366.150 813.900 367.950 ;
        RECT 804.000 364.950 808.050 365.550 ;
        RECT 773.700 354.600 775.500 363.000 ;
        RECT 788.700 362.700 792.300 363.600 ;
        RECT 815.700 363.600 816.900 367.950 ;
        RECT 818.100 366.150 819.900 367.950 ;
        RECT 824.550 366.450 825.450 374.550 ;
        RECT 833.100 370.050 834.900 371.850 ;
        RECT 837.000 370.050 837.900 375.600 ;
        RECT 838.950 370.050 840.750 371.850 ;
        RECT 857.100 370.050 858.900 371.850 ;
        RECT 863.700 370.050 864.900 377.400 ;
        RECT 868.950 372.450 871.050 373.050 ;
        RECT 874.950 372.450 877.050 373.050 ;
        RECT 868.950 371.550 877.050 372.450 ;
        RECT 868.950 370.950 871.050 371.550 ;
        RECT 874.950 370.950 877.050 371.550 ;
        RECT 882.000 370.050 882.900 382.200 ;
        RECT 905.100 378.300 906.900 389.400 ;
        RECT 908.100 379.200 909.900 390.000 ;
        RECT 911.100 378.300 912.900 389.400 ;
        RECT 905.100 377.400 912.900 378.300 ;
        RECT 914.100 377.400 915.900 389.400 ;
        RECT 895.950 375.450 898.050 376.050 ;
        RECT 910.950 375.450 913.050 376.050 ;
        RECT 895.950 374.550 913.050 375.450 ;
        RECT 895.950 373.950 898.050 374.550 ;
        RECT 910.950 373.950 913.050 374.550 ;
        RECT 887.100 370.050 888.900 371.850 ;
        RECT 908.250 370.050 910.050 371.850 ;
        RECT 914.700 370.050 915.600 377.400 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 835.950 367.950 838.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 880.950 367.950 883.050 370.050 ;
        RECT 883.950 367.950 886.050 370.050 ;
        RECT 886.950 367.950 889.050 370.050 ;
        RECT 889.950 367.950 892.050 370.050 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 907.950 367.950 910.050 370.050 ;
        RECT 910.950 367.950 913.050 370.050 ;
        RECT 913.950 367.950 916.050 370.050 ;
        RECT 824.550 365.550 828.450 366.450 ;
        RECT 830.100 366.150 831.900 367.950 ;
        RECT 815.700 362.700 819.300 363.600 ;
        RECT 788.700 360.600 789.900 362.700 ;
        RECT 788.100 354.600 789.900 360.600 ;
        RECT 791.100 359.700 798.900 361.050 ;
        RECT 791.100 354.600 792.900 359.700 ;
        RECT 794.100 354.000 795.900 358.800 ;
        RECT 797.100 354.600 798.900 359.700 ;
        RECT 809.100 359.700 816.900 361.050 ;
        RECT 809.100 354.600 810.900 359.700 ;
        RECT 812.100 354.000 813.900 358.800 ;
        RECT 815.100 354.600 816.900 359.700 ;
        RECT 818.100 360.600 819.300 362.700 ;
        RECT 827.550 363.450 828.450 365.550 ;
        RECT 832.950 363.450 835.050 364.050 ;
        RECT 827.550 362.550 835.050 363.450 ;
        RECT 832.950 361.950 835.050 362.550 ;
        RECT 836.700 360.600 837.900 367.950 ;
        RECT 841.950 366.150 843.750 367.950 ;
        RECT 860.100 366.150 861.900 367.950 ;
        RECT 863.700 363.600 864.900 367.950 ;
        RECT 866.100 366.150 867.900 367.950 ;
        RECT 882.000 364.200 882.900 367.950 ;
        RECT 884.100 366.150 885.900 367.950 ;
        RECT 890.100 366.150 891.900 367.950 ;
        RECT 905.100 366.150 906.900 367.950 ;
        RECT 911.250 366.150 913.050 367.950 ;
        RECT 863.700 362.700 867.300 363.600 ;
        RECT 882.000 363.000 885.300 364.200 ;
        RECT 818.100 354.600 819.900 360.600 ;
        RECT 832.500 354.000 834.300 360.600 ;
        RECT 837.000 354.600 838.800 360.600 ;
        RECT 841.500 354.000 843.300 360.600 ;
        RECT 857.100 359.700 864.900 361.050 ;
        RECT 857.100 354.600 858.900 359.700 ;
        RECT 860.100 354.000 861.900 358.800 ;
        RECT 863.100 354.600 864.900 359.700 ;
        RECT 866.100 360.600 867.300 362.700 ;
        RECT 866.100 354.600 867.900 360.600 ;
        RECT 883.500 354.600 885.300 363.000 ;
        RECT 890.100 354.000 891.900 363.600 ;
        RECT 914.700 360.600 915.600 367.950 ;
        RECT 906.000 354.000 907.800 360.600 ;
        RECT 910.500 359.400 915.600 360.600 ;
        RECT 910.500 354.600 912.300 359.400 ;
        RECT 913.500 354.000 915.300 357.600 ;
        RECT 14.100 344.400 15.900 351.000 ;
        RECT 17.100 343.500 18.900 350.400 ;
        RECT 20.100 344.400 21.900 351.000 ;
        RECT 23.100 343.500 24.900 350.400 ;
        RECT 26.100 344.400 27.900 351.000 ;
        RECT 29.100 343.500 30.900 350.400 ;
        RECT 32.100 344.400 33.900 351.000 ;
        RECT 35.100 343.500 36.900 350.400 ;
        RECT 38.100 344.400 39.900 351.000 ;
        RECT 53.100 347.400 54.900 350.400 ;
        RECT 56.100 347.400 57.900 351.000 ;
        RECT 59.700 347.400 61.500 351.000 ;
        RECT 62.700 347.400 64.500 350.400 ;
        RECT 17.100 342.300 21.000 343.500 ;
        RECT 23.100 342.300 27.000 343.500 ;
        RECT 29.100 342.300 33.000 343.500 ;
        RECT 35.100 342.300 37.950 343.500 ;
        RECT 19.800 341.400 21.000 342.300 ;
        RECT 25.800 341.400 27.000 342.300 ;
        RECT 31.800 341.400 33.000 342.300 ;
        RECT 19.800 340.200 24.000 341.400 ;
        RECT 16.800 337.050 18.600 338.850 ;
        RECT 16.800 334.950 18.900 337.050 ;
        RECT 19.800 329.700 21.000 340.200 ;
        RECT 22.200 339.600 24.000 340.200 ;
        RECT 25.800 340.200 30.000 341.400 ;
        RECT 25.800 329.700 27.000 340.200 ;
        RECT 28.200 339.600 30.000 340.200 ;
        RECT 31.800 340.200 36.000 341.400 ;
        RECT 31.800 329.700 33.000 340.200 ;
        RECT 34.200 339.600 36.000 340.200 ;
        RECT 36.900 337.050 37.950 342.300 ;
        RECT 53.700 337.050 54.900 347.400 ;
        RECT 34.800 334.950 37.950 337.050 ;
        RECT 52.950 334.950 55.050 337.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 36.900 329.700 37.950 334.950 ;
        RECT 17.100 328.500 21.000 329.700 ;
        RECT 23.100 328.500 27.000 329.700 ;
        RECT 29.100 328.500 33.000 329.700 ;
        RECT 35.100 328.500 37.950 329.700 ;
        RECT 14.100 315.000 15.900 327.600 ;
        RECT 17.100 315.600 18.900 328.500 ;
        RECT 20.100 315.000 21.900 327.600 ;
        RECT 23.100 315.600 24.900 328.500 ;
        RECT 26.100 315.000 27.900 327.600 ;
        RECT 29.100 315.600 30.900 328.500 ;
        RECT 32.100 315.000 33.900 327.600 ;
        RECT 35.100 315.600 36.900 328.500 ;
        RECT 38.100 315.000 39.900 327.600 ;
        RECT 53.700 321.600 54.900 334.950 ;
        RECT 56.100 333.150 57.900 334.950 ;
        RECT 63.000 334.050 64.500 347.400 ;
        RECT 62.100 331.950 64.500 334.050 ;
        RECT 63.000 321.600 64.500 331.950 ;
        RECT 66.300 344.400 68.100 350.400 ;
        RECT 71.700 344.400 73.500 351.000 ;
        RECT 76.800 345.600 78.600 350.400 ;
        RECT 81.000 347.400 82.800 350.400 ;
        RECT 84.000 347.400 85.800 350.400 ;
        RECT 87.000 347.400 88.800 350.400 ;
        RECT 90.000 347.400 91.800 350.400 ;
        RECT 93.000 347.400 94.800 351.000 ;
        RECT 74.400 344.400 78.600 345.600 ;
        RECT 80.700 345.300 82.800 347.400 ;
        RECT 83.700 345.300 85.800 347.400 ;
        RECT 86.700 345.300 88.800 347.400 ;
        RECT 89.700 345.300 91.800 347.400 ;
        RECT 96.000 346.500 97.800 350.400 ;
        RECT 100.500 347.400 102.300 351.000 ;
        RECT 103.500 347.400 105.300 350.400 ;
        RECT 106.500 347.400 108.300 350.400 ;
        RECT 109.500 347.400 111.300 350.400 ;
        RECT 95.100 344.400 97.800 346.500 ;
        RECT 99.600 345.600 101.400 346.500 ;
        RECT 99.600 344.400 102.300 345.600 ;
        RECT 103.200 345.300 105.300 347.400 ;
        RECT 106.200 345.300 108.300 347.400 ;
        RECT 109.200 345.300 111.300 347.400 ;
        RECT 113.700 344.400 115.500 350.400 ;
        RECT 119.100 344.400 120.900 351.000 ;
        RECT 124.500 344.400 126.300 350.400 ;
        RECT 140.700 347.400 142.500 351.000 ;
        RECT 143.700 345.600 145.500 350.400 ;
        RECT 66.300 327.600 67.200 344.400 ;
        RECT 74.400 341.100 75.900 344.400 ;
        RECT 80.100 342.600 86.700 344.400 ;
        RECT 101.400 343.800 102.300 344.400 ;
        RECT 104.400 343.800 106.200 344.400 ;
        RECT 101.400 342.600 108.600 343.800 ;
        RECT 68.100 339.300 75.900 341.100 ;
        RECT 92.100 340.500 93.900 342.300 ;
        RECT 91.800 339.900 93.900 340.500 ;
        RECT 76.800 338.400 93.900 339.900 ;
        RECT 98.100 339.900 100.200 340.050 ;
        RECT 101.400 339.900 103.200 340.800 ;
        RECT 98.100 339.000 103.200 339.900 ;
        RECT 107.700 339.600 108.600 342.600 ;
        RECT 113.700 343.500 115.200 344.400 ;
        RECT 113.700 342.300 122.100 343.500 ;
        RECT 120.300 341.700 122.100 342.300 ;
        RECT 109.500 340.800 111.600 341.700 ;
        RECT 125.100 340.800 126.300 344.400 ;
        RECT 109.500 339.600 126.300 340.800 ;
        RECT 140.400 344.400 145.500 345.600 ;
        RECT 148.200 344.400 150.000 351.000 ;
        RECT 161.700 347.400 163.500 351.000 ;
        RECT 164.700 345.600 166.500 350.400 ;
        RECT 161.400 344.400 166.500 345.600 ;
        RECT 169.200 344.400 171.000 351.000 ;
        RECT 182.100 344.400 183.900 350.400 ;
        RECT 71.700 336.900 78.300 338.400 ;
        RECT 98.100 337.950 100.200 339.000 ;
        RECT 106.800 337.800 108.600 339.600 ;
        RECT 71.700 334.050 73.200 336.900 ;
        RECT 79.500 335.700 123.900 336.900 ;
        RECT 79.500 334.200 80.400 335.700 ;
        RECT 71.100 331.950 73.200 334.050 ;
        RECT 75.300 332.400 80.400 334.200 ;
        RECT 83.100 333.900 96.600 334.800 ;
        RECT 103.800 333.900 105.600 334.500 ;
        RECT 122.100 334.050 123.900 335.700 ;
        RECT 83.100 332.700 84.000 333.900 ;
        RECT 83.100 330.900 84.900 332.700 ;
        RECT 89.100 331.200 93.000 333.000 ;
        RECT 94.500 332.700 105.600 333.900 ;
        RECT 116.100 333.750 118.200 334.050 ;
        RECT 94.500 331.800 96.600 332.700 ;
        RECT 114.300 331.950 118.200 333.750 ;
        RECT 122.100 331.950 124.200 334.050 ;
        RECT 114.300 331.200 116.100 331.950 ;
        RECT 89.100 330.900 91.200 331.200 ;
        RECT 102.600 330.300 116.100 331.200 ;
        RECT 68.100 329.700 69.900 330.300 ;
        RECT 102.600 329.700 103.800 330.300 ;
        RECT 68.100 328.500 103.800 329.700 ;
        RECT 106.500 328.500 108.600 328.800 ;
        RECT 66.300 326.700 82.800 327.600 ;
        RECT 66.300 323.400 67.200 326.700 ;
        RECT 71.100 324.600 76.800 325.800 ;
        RECT 80.700 325.500 82.800 326.700 ;
        RECT 86.100 326.400 103.800 327.600 ;
        RECT 106.500 327.300 118.500 328.500 ;
        RECT 106.500 326.700 108.600 327.300 ;
        RECT 116.700 326.700 118.500 327.300 ;
        RECT 86.100 325.500 88.200 326.400 ;
        RECT 102.600 325.800 103.800 326.400 ;
        RECT 120.000 325.800 121.800 326.100 ;
        RECT 71.100 324.000 72.900 324.600 ;
        RECT 66.300 322.500 70.200 323.400 ;
        RECT 69.000 321.600 70.200 322.500 ;
        RECT 75.600 321.600 76.800 324.600 ;
        RECT 77.700 323.700 79.500 324.300 ;
        RECT 77.700 322.500 85.800 323.700 ;
        RECT 83.700 321.600 85.800 322.500 ;
        RECT 89.100 321.600 91.800 325.500 ;
        RECT 94.500 323.100 97.800 325.200 ;
        RECT 102.600 324.600 121.800 325.800 ;
        RECT 53.100 315.600 54.900 321.600 ;
        RECT 56.100 315.000 57.900 321.600 ;
        RECT 59.700 315.000 61.500 321.600 ;
        RECT 62.700 315.600 64.500 321.600 ;
        RECT 66.000 315.000 67.800 321.600 ;
        RECT 69.000 315.600 70.800 321.600 ;
        RECT 72.000 315.000 73.800 321.600 ;
        RECT 75.000 315.600 76.800 321.600 ;
        RECT 78.000 315.000 79.800 321.600 ;
        RECT 80.700 318.600 82.800 320.700 ;
        RECT 83.700 318.600 85.800 320.700 ;
        RECT 86.700 318.600 88.800 320.700 ;
        RECT 81.000 315.600 82.800 318.600 ;
        RECT 84.000 315.600 85.800 318.600 ;
        RECT 87.000 315.600 88.800 318.600 ;
        RECT 90.000 315.600 91.800 321.600 ;
        RECT 93.000 315.000 94.800 321.600 ;
        RECT 96.000 315.600 97.800 323.100 ;
        RECT 103.200 321.600 105.300 323.700 ;
        RECT 99.900 315.000 101.700 321.600 ;
        RECT 102.900 315.600 104.700 321.600 ;
        RECT 105.600 318.600 107.700 320.700 ;
        RECT 108.600 318.600 110.700 320.700 ;
        RECT 105.900 315.600 107.700 318.600 ;
        RECT 108.900 315.600 110.700 318.600 ;
        RECT 112.500 315.000 114.300 321.600 ;
        RECT 115.500 315.600 117.300 324.600 ;
        RECT 120.000 324.300 121.800 324.600 ;
        RECT 125.100 323.400 126.300 339.600 ;
        RECT 135.000 339.450 139.050 340.050 ;
        RECT 134.550 337.950 139.050 339.450 ;
        RECT 134.550 334.050 135.450 337.950 ;
        RECT 140.400 337.050 141.300 344.400 ;
        RECT 142.950 337.050 144.750 338.850 ;
        RECT 149.100 337.050 150.900 338.850 ;
        RECT 161.400 337.050 162.300 344.400 ;
        RECT 182.700 342.300 183.900 344.400 ;
        RECT 185.100 345.300 186.900 350.400 ;
        RECT 188.100 346.200 189.900 351.000 ;
        RECT 191.100 345.300 192.900 350.400 ;
        RECT 185.100 343.950 192.900 345.300 ;
        RECT 206.400 344.400 208.200 351.000 ;
        RECT 211.500 343.200 213.300 350.400 ;
        RECT 227.100 347.400 228.900 350.400 ;
        RECT 230.100 347.400 231.900 351.000 ;
        RECT 242.100 347.400 243.900 351.000 ;
        RECT 245.100 347.400 246.900 350.400 ;
        RECT 260.100 347.400 261.900 351.000 ;
        RECT 263.100 347.400 264.900 350.400 ;
        RECT 209.100 342.300 213.300 343.200 ;
        RECT 182.700 341.400 186.300 342.300 ;
        RECT 172.950 339.450 177.000 340.050 ;
        RECT 163.950 337.050 165.750 338.850 ;
        RECT 170.100 337.050 171.900 338.850 ;
        RECT 172.950 337.950 177.450 339.450 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 134.550 332.550 139.050 334.050 ;
        RECT 135.000 331.950 139.050 332.550 ;
        RECT 140.400 327.600 141.300 334.950 ;
        RECT 145.950 333.150 147.750 334.950 ;
        RECT 142.950 330.450 145.050 331.050 ;
        RECT 151.950 330.450 154.050 331.050 ;
        RECT 157.950 330.450 160.050 331.050 ;
        RECT 142.950 329.550 160.050 330.450 ;
        RECT 142.950 328.950 145.050 329.550 ;
        RECT 151.950 328.950 154.050 329.550 ;
        RECT 157.950 328.950 160.050 329.550 ;
        RECT 161.400 327.600 162.300 334.950 ;
        RECT 166.950 333.150 168.750 334.950 ;
        RECT 176.550 334.050 177.450 337.950 ;
        RECT 182.100 337.050 183.900 338.850 ;
        RECT 185.100 337.050 186.300 341.400 ;
        RECT 188.100 337.050 189.900 338.850 ;
        RECT 206.250 337.050 208.050 338.850 ;
        RECT 209.100 337.050 210.300 342.300 ;
        RECT 212.100 337.050 213.900 338.850 ;
        RECT 227.700 337.050 228.900 347.400 ;
        RECT 245.100 337.050 246.300 347.400 ;
        RECT 263.100 337.050 264.300 347.400 ;
        RECT 275.100 344.400 276.900 350.400 ;
        RECT 278.100 345.000 279.900 351.000 ;
        RECT 284.700 350.400 285.900 351.000 ;
        RECT 281.100 347.400 282.900 350.400 ;
        RECT 284.100 347.400 285.900 350.400 ;
        RECT 275.100 337.050 276.000 344.400 ;
        RECT 281.700 343.200 282.600 347.400 ;
        RECT 296.400 344.400 298.200 351.000 ;
        RECT 301.500 343.200 303.300 350.400 ;
        RECT 317.400 344.400 319.200 351.000 ;
        RECT 322.500 343.200 324.300 350.400 ;
        RECT 338.700 344.400 340.500 351.000 ;
        RECT 343.200 344.400 345.000 350.400 ;
        RECT 347.700 344.400 349.500 351.000 ;
        RECT 367.500 344.400 369.300 351.000 ;
        RECT 372.000 344.400 373.800 350.400 ;
        RECT 376.500 344.400 378.300 351.000 ;
        RECT 389.100 347.400 390.900 351.000 ;
        RECT 392.100 347.400 393.900 350.400 ;
        RECT 277.200 342.300 282.600 343.200 ;
        RECT 299.100 342.300 303.300 343.200 ;
        RECT 310.950 342.450 313.050 343.050 ;
        RECT 316.950 342.450 319.050 343.050 ;
        RECT 277.200 341.400 279.300 342.300 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 275.100 334.950 277.200 337.050 ;
        RECT 172.950 332.550 177.450 334.050 ;
        RECT 172.950 331.950 177.000 332.550 ;
        RECT 185.100 327.600 186.300 334.950 ;
        RECT 191.100 333.150 192.900 334.950 ;
        RECT 122.700 322.500 126.300 323.400 ;
        RECT 122.700 321.600 123.600 322.500 ;
        RECT 118.500 315.000 120.300 321.600 ;
        RECT 121.500 320.700 123.600 321.600 ;
        RECT 121.500 315.600 123.300 320.700 ;
        RECT 124.500 315.000 126.300 321.600 ;
        RECT 140.100 315.600 141.900 327.600 ;
        RECT 143.100 326.700 150.900 327.600 ;
        RECT 143.100 315.600 144.900 326.700 ;
        RECT 146.100 315.000 147.900 325.800 ;
        RECT 149.100 315.600 150.900 326.700 ;
        RECT 161.100 315.600 162.900 327.600 ;
        RECT 164.100 326.700 171.900 327.600 ;
        RECT 164.100 315.600 165.900 326.700 ;
        RECT 167.100 315.000 168.900 325.800 ;
        RECT 170.100 315.600 171.900 326.700 ;
        RECT 185.100 326.100 187.500 327.600 ;
        RECT 183.000 323.100 184.800 324.900 ;
        RECT 182.700 315.000 184.500 321.600 ;
        RECT 185.700 315.600 187.500 326.100 ;
        RECT 190.800 315.000 192.600 327.600 ;
        RECT 209.100 321.600 210.300 334.950 ;
        RECT 227.700 321.600 228.900 334.950 ;
        RECT 230.100 333.150 231.900 334.950 ;
        RECT 242.100 333.150 243.900 334.950 ;
        RECT 245.100 321.600 246.300 334.950 ;
        RECT 260.100 333.150 261.900 334.950 ;
        RECT 263.100 321.600 264.300 334.950 ;
        RECT 276.000 327.600 277.200 334.950 ;
        RECT 278.400 330.900 279.300 341.400 ;
        RECT 283.800 337.050 285.600 338.850 ;
        RECT 296.250 337.050 298.050 338.850 ;
        RECT 299.100 337.050 300.300 342.300 ;
        RECT 310.950 341.550 319.050 342.450 ;
        RECT 310.950 340.950 313.050 341.550 ;
        RECT 316.950 340.950 319.050 341.550 ;
        RECT 320.100 342.300 324.300 343.200 ;
        RECT 312.000 339.450 316.050 340.050 ;
        RECT 302.100 337.050 303.900 338.850 ;
        RECT 311.550 337.950 316.050 339.450 ;
        RECT 280.500 334.950 282.600 337.050 ;
        RECT 283.800 334.950 285.900 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 280.200 333.150 282.000 334.950 ;
        RECT 278.100 330.300 279.900 330.900 ;
        RECT 278.100 329.100 285.900 330.300 ;
        RECT 284.700 327.600 285.900 329.100 ;
        RECT 276.000 326.100 278.400 327.600 ;
        RECT 206.100 315.000 207.900 321.600 ;
        RECT 209.100 315.600 210.900 321.600 ;
        RECT 212.100 315.000 213.900 321.600 ;
        RECT 227.100 315.600 228.900 321.600 ;
        RECT 230.100 315.000 231.900 321.600 ;
        RECT 242.100 315.000 243.900 321.600 ;
        RECT 245.100 315.600 246.900 321.600 ;
        RECT 260.100 315.000 261.900 321.600 ;
        RECT 263.100 315.600 264.900 321.600 ;
        RECT 276.600 315.600 278.400 326.100 ;
        RECT 279.600 315.000 281.400 327.600 ;
        RECT 284.100 315.600 285.900 327.600 ;
        RECT 299.100 321.600 300.300 334.950 ;
        RECT 311.550 333.450 312.450 337.950 ;
        RECT 317.250 337.050 319.050 338.850 ;
        RECT 320.100 337.050 321.300 342.300 ;
        RECT 323.100 337.050 324.900 338.850 ;
        RECT 338.250 337.050 340.050 338.850 ;
        RECT 344.100 337.050 345.300 344.400 ;
        RECT 352.950 339.450 357.000 340.050 ;
        RECT 350.100 337.050 351.900 338.850 ;
        RECT 352.950 337.950 357.450 339.450 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 311.550 332.550 315.450 333.450 ;
        RECT 314.550 331.050 315.450 332.550 ;
        RECT 314.550 329.550 319.050 331.050 ;
        RECT 315.000 328.950 319.050 329.550 ;
        RECT 320.100 321.600 321.300 334.950 ;
        RECT 341.250 333.150 343.050 334.950 ;
        RECT 336.000 330.450 340.050 331.050 ;
        RECT 335.550 328.950 340.050 330.450 ;
        RECT 344.100 329.400 345.000 334.950 ;
        RECT 347.100 333.150 348.900 334.950 ;
        RECT 356.550 333.450 357.450 337.950 ;
        RECT 365.100 337.050 366.900 338.850 ;
        RECT 371.700 337.050 372.900 344.400 ;
        RECT 379.950 339.450 384.000 340.050 ;
        RECT 376.950 337.050 378.750 338.850 ;
        RECT 379.950 337.950 384.450 339.450 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 361.950 333.450 364.050 334.050 ;
        RECT 356.550 332.550 364.050 333.450 ;
        RECT 368.100 333.150 369.900 334.950 ;
        RECT 361.950 331.950 364.050 332.550 ;
        RECT 372.000 329.400 372.900 334.950 ;
        RECT 373.950 333.150 375.750 334.950 ;
        RECT 322.950 327.450 325.050 328.050 ;
        RECT 335.550 327.450 336.450 328.950 ;
        RECT 344.100 328.500 348.900 329.400 ;
        RECT 322.950 326.550 336.450 327.450 ;
        RECT 322.950 325.950 325.050 326.550 ;
        RECT 338.100 326.400 345.900 327.300 ;
        RECT 296.100 315.000 297.900 321.600 ;
        RECT 299.100 315.600 300.900 321.600 ;
        RECT 302.100 315.000 303.900 321.600 ;
        RECT 317.100 315.000 318.900 321.600 ;
        RECT 320.100 315.600 321.900 321.600 ;
        RECT 323.100 315.000 324.900 321.600 ;
        RECT 325.950 321.450 328.050 325.050 ;
        RECT 334.950 321.450 337.050 322.050 ;
        RECT 325.950 321.000 337.050 321.450 ;
        RECT 326.550 320.550 337.050 321.000 ;
        RECT 334.950 319.950 337.050 320.550 ;
        RECT 338.100 315.600 339.900 326.400 ;
        RECT 341.100 315.000 342.900 325.500 ;
        RECT 344.100 316.500 345.900 326.400 ;
        RECT 347.100 317.400 348.900 328.500 ;
        RECT 368.100 328.500 372.900 329.400 ;
        RECT 373.950 330.450 376.050 331.050 ;
        RECT 383.550 330.450 384.450 337.950 ;
        RECT 392.100 337.050 393.300 347.400 ;
        RECT 404.100 341.400 405.900 351.000 ;
        RECT 410.700 342.000 412.500 350.400 ;
        RECT 426.000 344.400 427.800 351.000 ;
        RECT 430.500 345.600 432.300 350.400 ;
        RECT 433.500 347.400 435.300 351.000 ;
        RECT 430.500 344.400 435.600 345.600 ;
        RECT 410.700 340.800 414.000 342.000 ;
        RECT 404.100 337.050 405.900 338.850 ;
        RECT 410.100 337.050 411.900 338.850 ;
        RECT 413.100 337.050 414.000 340.800 ;
        RECT 420.000 339.450 424.050 340.050 ;
        RECT 419.550 337.950 424.050 339.450 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 403.950 334.950 406.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 389.100 333.150 390.900 334.950 ;
        RECT 373.950 329.550 384.450 330.450 ;
        RECT 373.950 328.950 376.050 329.550 ;
        RECT 350.100 316.500 351.900 327.600 ;
        RECT 344.100 315.600 351.900 316.500 ;
        RECT 365.100 316.500 366.900 327.600 ;
        RECT 368.100 317.400 369.900 328.500 ;
        RECT 371.100 326.400 378.900 327.300 ;
        RECT 371.100 316.500 372.900 326.400 ;
        RECT 365.100 315.600 372.900 316.500 ;
        RECT 374.100 315.000 375.900 325.500 ;
        RECT 377.100 315.600 378.900 326.400 ;
        RECT 392.100 321.600 393.300 334.950 ;
        RECT 407.100 333.150 408.900 334.950 ;
        RECT 397.950 330.450 400.050 331.050 ;
        RECT 409.950 330.450 412.050 331.050 ;
        RECT 397.950 329.550 412.050 330.450 ;
        RECT 397.950 328.950 400.050 329.550 ;
        RECT 409.950 328.950 412.050 329.550 ;
        RECT 413.100 322.800 414.000 334.950 ;
        RECT 419.550 334.050 420.450 337.950 ;
        RECT 425.100 337.050 426.900 338.850 ;
        RECT 431.250 337.050 433.050 338.850 ;
        RECT 434.700 337.050 435.600 344.400 ;
        RECT 451.500 342.000 453.300 350.400 ;
        RECT 450.000 340.800 453.300 342.000 ;
        RECT 458.100 341.400 459.900 351.000 ;
        RECT 475.500 342.000 477.300 350.400 ;
        RECT 474.000 340.800 477.300 342.000 ;
        RECT 482.100 341.400 483.900 351.000 ;
        RECT 494.100 347.400 495.900 351.000 ;
        RECT 497.100 347.400 498.900 350.400 ;
        RECT 500.100 347.400 501.900 351.000 ;
        RECT 450.000 337.050 450.900 340.800 ;
        RECT 452.100 337.050 453.900 338.850 ;
        RECT 458.100 337.050 459.900 338.850 ;
        RECT 474.000 337.050 474.900 340.800 ;
        RECT 476.100 337.050 477.900 338.850 ;
        RECT 482.100 337.050 483.900 338.850 ;
        RECT 497.700 337.050 498.600 347.400 ;
        RECT 515.700 343.200 517.500 350.400 ;
        RECT 520.800 344.400 522.600 351.000 ;
        RECT 515.700 342.300 519.900 343.200 ;
        RECT 502.950 339.450 505.050 340.050 ;
        RECT 502.950 338.550 510.450 339.450 ;
        RECT 502.950 337.950 505.050 338.550 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 415.950 332.550 420.450 334.050 ;
        RECT 428.250 333.150 430.050 334.950 ;
        RECT 415.950 331.950 420.000 332.550 ;
        RECT 434.700 327.600 435.600 334.950 ;
        RECT 407.400 321.900 414.000 322.800 ;
        RECT 407.400 321.600 408.900 321.900 ;
        RECT 389.100 315.000 390.900 321.600 ;
        RECT 392.100 315.600 393.900 321.600 ;
        RECT 404.100 315.000 405.900 321.600 ;
        RECT 407.100 315.600 408.900 321.600 ;
        RECT 413.100 321.600 414.000 321.900 ;
        RECT 425.100 326.700 432.900 327.600 ;
        RECT 410.100 315.000 411.900 321.000 ;
        RECT 413.100 315.600 414.900 321.600 ;
        RECT 425.100 315.600 426.900 326.700 ;
        RECT 428.100 315.000 429.900 325.800 ;
        RECT 431.100 315.600 432.900 326.700 ;
        RECT 434.100 315.600 435.900 327.600 ;
        RECT 450.000 322.800 450.900 334.950 ;
        RECT 455.100 333.150 456.900 334.950 ;
        RECT 457.950 330.450 460.050 331.050 ;
        RECT 466.950 330.450 469.050 331.050 ;
        RECT 457.950 329.550 469.050 330.450 ;
        RECT 457.950 328.950 460.050 329.550 ;
        RECT 466.950 328.950 469.050 329.550 ;
        RECT 474.000 322.800 474.900 334.950 ;
        RECT 479.100 333.150 480.900 334.950 ;
        RECT 494.100 333.150 495.900 334.950 ;
        RECT 497.700 327.600 498.600 334.950 ;
        RECT 499.950 333.150 501.750 334.950 ;
        RECT 509.550 333.900 510.450 338.550 ;
        RECT 515.100 337.050 516.900 338.850 ;
        RECT 518.700 337.050 519.900 342.300 ;
        RECT 535.500 342.000 537.300 350.400 ;
        RECT 534.000 340.800 537.300 342.000 ;
        RECT 542.100 341.400 543.900 351.000 ;
        RECT 556.500 344.400 558.300 351.000 ;
        RECT 561.000 344.400 562.800 350.400 ;
        RECT 565.500 344.400 567.300 351.000 ;
        RECT 581.700 344.400 583.500 351.000 ;
        RECT 586.200 344.400 588.000 350.400 ;
        RECT 590.700 344.400 592.500 351.000 ;
        RECT 553.950 342.450 556.050 343.050 ;
        RECT 548.550 341.550 556.050 342.450 ;
        RECT 528.000 339.450 532.050 340.050 ;
        RECT 520.950 337.050 522.750 338.850 ;
        RECT 527.550 337.950 532.050 339.450 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 508.950 331.800 511.050 333.900 ;
        RECT 495.000 326.400 498.600 327.600 ;
        RECT 450.000 321.900 456.600 322.800 ;
        RECT 450.000 321.600 450.900 321.900 ;
        RECT 449.100 315.600 450.900 321.600 ;
        RECT 455.100 321.600 456.600 321.900 ;
        RECT 474.000 321.900 480.600 322.800 ;
        RECT 474.000 321.600 474.900 321.900 ;
        RECT 452.100 315.000 453.900 321.000 ;
        RECT 455.100 315.600 456.900 321.600 ;
        RECT 458.100 315.000 459.900 321.600 ;
        RECT 473.100 315.600 474.900 321.600 ;
        RECT 479.100 321.600 480.600 321.900 ;
        RECT 476.100 315.000 477.900 321.000 ;
        RECT 479.100 315.600 480.900 321.600 ;
        RECT 482.100 315.000 483.900 321.600 ;
        RECT 495.000 315.600 496.800 326.400 ;
        RECT 500.100 315.000 501.900 327.600 ;
        RECT 518.700 321.600 519.900 334.950 ;
        RECT 527.550 334.050 528.450 337.950 ;
        RECT 534.000 337.050 534.900 340.800 ;
        RECT 536.100 337.050 537.900 338.850 ;
        RECT 542.100 337.050 543.900 338.850 ;
        RECT 532.950 334.950 535.050 337.050 ;
        RECT 535.950 334.950 538.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 523.950 332.550 528.450 334.050 ;
        RECT 523.950 331.950 528.000 332.550 ;
        RECT 534.000 322.800 534.900 334.950 ;
        RECT 539.100 333.150 540.900 334.950 ;
        RECT 548.550 334.050 549.450 341.550 ;
        RECT 553.950 340.950 556.050 341.550 ;
        RECT 554.100 337.050 555.900 338.850 ;
        RECT 560.700 337.050 561.900 344.400 ;
        RECT 565.950 337.050 567.750 338.850 ;
        RECT 581.250 337.050 583.050 338.850 ;
        RECT 587.100 337.050 588.300 344.400 ;
        RECT 608.700 343.200 610.500 350.400 ;
        RECT 613.800 344.400 615.600 351.000 ;
        RECT 592.950 342.450 595.050 343.050 ;
        RECT 601.950 342.450 604.050 343.050 ;
        RECT 592.950 341.550 604.050 342.450 ;
        RECT 608.700 342.300 612.900 343.200 ;
        RECT 592.950 340.950 595.050 341.550 ;
        RECT 601.950 340.950 604.050 341.550 ;
        RECT 593.100 337.050 594.900 338.850 ;
        RECT 608.100 337.050 609.900 338.850 ;
        RECT 611.700 337.050 612.900 342.300 ;
        RECT 613.950 342.450 616.050 343.050 ;
        RECT 613.950 341.550 621.450 342.450 ;
        RECT 613.950 340.950 616.050 341.550 ;
        RECT 613.950 337.050 615.750 338.850 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 544.950 332.550 549.450 334.050 ;
        RECT 557.100 333.150 558.900 334.950 ;
        RECT 544.950 331.950 549.000 332.550 ;
        RECT 561.000 329.400 561.900 334.950 ;
        RECT 562.950 333.150 564.750 334.950 ;
        RECT 584.250 333.150 586.050 334.950 ;
        RECT 557.100 328.500 561.900 329.400 ;
        RECT 587.100 329.400 588.000 334.950 ;
        RECT 590.100 333.150 591.900 334.950 ;
        RECT 587.100 328.500 591.900 329.400 ;
        RECT 534.000 321.900 540.600 322.800 ;
        RECT 534.000 321.600 534.900 321.900 ;
        RECT 515.100 315.000 516.900 321.600 ;
        RECT 518.100 315.600 519.900 321.600 ;
        RECT 521.100 315.000 522.900 321.600 ;
        RECT 533.100 315.600 534.900 321.600 ;
        RECT 539.100 321.600 540.600 321.900 ;
        RECT 536.100 315.000 537.900 321.000 ;
        RECT 539.100 315.600 540.900 321.600 ;
        RECT 542.100 315.000 543.900 321.600 ;
        RECT 554.100 316.500 555.900 327.600 ;
        RECT 557.100 317.400 558.900 328.500 ;
        RECT 560.100 326.400 567.900 327.300 ;
        RECT 560.100 316.500 561.900 326.400 ;
        RECT 554.100 315.600 561.900 316.500 ;
        RECT 563.100 315.000 564.900 325.500 ;
        RECT 566.100 315.600 567.900 326.400 ;
        RECT 581.100 326.400 588.900 327.300 ;
        RECT 581.100 315.600 582.900 326.400 ;
        RECT 584.100 315.000 585.900 325.500 ;
        RECT 587.100 316.500 588.900 326.400 ;
        RECT 590.100 317.400 591.900 328.500 ;
        RECT 593.100 316.500 594.900 327.600 ;
        RECT 611.700 321.600 612.900 334.950 ;
        RECT 620.550 333.450 621.450 341.550 ;
        RECT 626.100 341.400 627.900 351.000 ;
        RECT 632.700 342.000 634.500 350.400 ;
        RECT 647.100 347.400 648.900 351.000 ;
        RECT 650.100 347.400 651.900 350.400 ;
        RECT 632.700 340.800 636.000 342.000 ;
        RECT 626.100 337.050 627.900 338.850 ;
        RECT 632.100 337.050 633.900 338.850 ;
        RECT 635.100 337.050 636.000 340.800 ;
        RECT 650.100 337.050 651.300 347.400 ;
        RECT 665.100 341.400 666.900 351.000 ;
        RECT 671.700 342.000 673.500 350.400 ;
        RECT 689.700 343.200 691.500 350.400 ;
        RECT 694.800 344.400 696.600 351.000 ;
        RECT 707.100 347.400 708.900 351.000 ;
        RECT 710.100 347.400 711.900 350.400 ;
        RECT 689.700 342.300 693.900 343.200 ;
        RECT 671.700 340.800 675.000 342.000 ;
        RECT 652.950 339.450 657.000 340.050 ;
        RECT 652.950 337.950 657.450 339.450 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 631.950 334.950 634.050 337.050 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 620.550 332.550 624.450 333.450 ;
        RECT 629.100 333.150 630.900 334.950 ;
        RECT 623.550 330.450 624.450 332.550 ;
        RECT 631.950 330.450 634.050 331.050 ;
        RECT 623.550 329.550 634.050 330.450 ;
        RECT 631.950 328.950 634.050 329.550 ;
        RECT 635.100 322.800 636.000 334.950 ;
        RECT 647.100 333.150 648.900 334.950 ;
        RECT 629.400 321.900 636.000 322.800 ;
        RECT 629.400 321.600 630.900 321.900 ;
        RECT 587.100 315.600 594.900 316.500 ;
        RECT 608.100 315.000 609.900 321.600 ;
        RECT 611.100 315.600 612.900 321.600 ;
        RECT 614.100 315.000 615.900 321.600 ;
        RECT 626.100 315.000 627.900 321.600 ;
        RECT 629.100 315.600 630.900 321.600 ;
        RECT 635.100 321.600 636.000 321.900 ;
        RECT 650.100 321.600 651.300 334.950 ;
        RECT 656.550 334.050 657.450 337.950 ;
        RECT 665.100 337.050 666.900 338.850 ;
        RECT 671.100 337.050 672.900 338.850 ;
        RECT 674.100 337.050 675.000 340.800 ;
        RECT 676.950 339.450 681.000 340.050 ;
        RECT 676.950 337.950 681.450 339.450 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 652.950 332.550 657.450 334.050 ;
        RECT 668.100 333.150 669.900 334.950 ;
        RECT 652.950 331.950 657.000 332.550 ;
        RECT 674.100 322.800 675.000 334.950 ;
        RECT 680.550 333.450 681.450 337.950 ;
        RECT 689.100 337.050 690.900 338.850 ;
        RECT 692.700 337.050 693.900 342.300 ;
        RECT 694.950 337.050 696.750 338.850 ;
        RECT 710.100 337.050 711.300 347.400 ;
        RECT 722.100 345.300 723.900 350.400 ;
        RECT 725.100 346.200 726.900 351.000 ;
        RECT 728.100 345.300 729.900 350.400 ;
        RECT 722.100 343.950 729.900 345.300 ;
        RECT 731.100 344.400 732.900 350.400 ;
        RECT 743.700 347.400 745.500 351.000 ;
        RECT 746.700 345.600 748.500 350.400 ;
        RECT 743.400 344.400 748.500 345.600 ;
        RECT 751.200 344.400 753.000 351.000 ;
        RECT 764.100 347.400 765.900 350.400 ;
        RECT 767.100 347.400 768.900 351.000 ;
        RECT 731.100 342.300 732.300 344.400 ;
        RECT 728.700 341.400 732.300 342.300 ;
        RECT 712.950 339.450 717.000 340.050 ;
        RECT 712.950 337.950 717.450 339.450 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 706.950 334.950 709.050 337.050 ;
        RECT 709.950 334.950 712.050 337.050 ;
        RECT 685.950 333.450 688.050 334.050 ;
        RECT 680.550 332.550 688.050 333.450 ;
        RECT 685.950 331.950 688.050 332.550 ;
        RECT 679.950 324.450 682.050 325.050 ;
        RECT 688.950 324.450 691.050 325.050 ;
        RECT 679.950 323.550 691.050 324.450 ;
        RECT 679.950 322.950 682.050 323.550 ;
        RECT 688.950 322.950 691.050 323.550 ;
        RECT 668.400 321.900 675.000 322.800 ;
        RECT 668.400 321.600 669.900 321.900 ;
        RECT 632.100 315.000 633.900 321.000 ;
        RECT 635.100 315.600 636.900 321.600 ;
        RECT 647.100 315.000 648.900 321.600 ;
        RECT 650.100 315.600 651.900 321.600 ;
        RECT 665.100 315.000 666.900 321.600 ;
        RECT 668.100 315.600 669.900 321.600 ;
        RECT 674.100 321.600 675.000 321.900 ;
        RECT 692.700 321.600 693.900 334.950 ;
        RECT 707.100 333.150 708.900 334.950 ;
        RECT 710.100 321.600 711.300 334.950 ;
        RECT 716.550 334.050 717.450 337.950 ;
        RECT 725.100 337.050 726.900 338.850 ;
        RECT 728.700 337.050 729.900 341.400 ;
        RECT 738.000 339.450 742.050 340.050 ;
        RECT 731.100 337.050 732.900 338.850 ;
        RECT 737.550 337.950 742.050 339.450 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 727.950 334.950 730.050 337.050 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 716.550 332.550 721.050 334.050 ;
        RECT 722.100 333.150 723.900 334.950 ;
        RECT 717.000 331.950 721.050 332.550 ;
        RECT 728.700 327.600 729.900 334.950 ;
        RECT 737.550 334.050 738.450 337.950 ;
        RECT 743.400 337.050 744.300 344.400 ;
        RECT 754.950 339.450 759.000 340.050 ;
        RECT 745.950 337.050 747.750 338.850 ;
        RECT 752.100 337.050 753.900 338.850 ;
        RECT 754.950 337.950 759.450 339.450 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 733.950 332.550 738.450 334.050 ;
        RECT 733.950 331.950 738.000 332.550 ;
        RECT 743.400 327.600 744.300 334.950 ;
        RECT 748.950 333.150 750.750 334.950 ;
        RECT 758.550 334.050 759.450 337.950 ;
        RECT 764.700 337.050 765.900 347.400 ;
        RECT 782.100 341.400 783.900 351.000 ;
        RECT 788.700 342.000 790.500 350.400 ;
        RECT 803.400 344.400 805.200 351.000 ;
        RECT 808.500 343.200 810.300 350.400 ;
        RECT 806.100 342.300 810.300 343.200 ;
        RECT 824.100 342.600 825.900 350.400 ;
        RECT 828.600 344.400 830.400 351.000 ;
        RECT 831.600 346.200 833.400 350.400 ;
        RECT 831.600 344.400 834.300 346.200 ;
        RECT 830.700 342.600 832.500 343.500 ;
        RECT 788.700 340.800 792.000 342.000 ;
        RECT 782.100 337.050 783.900 338.850 ;
        RECT 788.100 337.050 789.900 338.850 ;
        RECT 791.100 337.050 792.000 340.800 ;
        RECT 803.250 337.050 805.050 338.850 ;
        RECT 806.100 337.050 807.300 342.300 ;
        RECT 824.100 341.700 832.500 342.600 ;
        RECT 809.100 337.050 810.900 338.850 ;
        RECT 824.250 337.050 826.050 338.850 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 824.100 334.950 826.200 337.050 ;
        RECT 754.950 332.550 759.450 334.050 ;
        RECT 754.950 331.950 759.000 332.550 ;
        RECT 671.100 315.000 672.900 321.000 ;
        RECT 674.100 315.600 675.900 321.600 ;
        RECT 689.100 315.000 690.900 321.600 ;
        RECT 692.100 315.600 693.900 321.600 ;
        RECT 695.100 315.000 696.900 321.600 ;
        RECT 697.950 318.900 702.000 319.050 ;
        RECT 697.950 316.950 703.050 318.900 ;
        RECT 700.950 316.800 703.050 316.950 ;
        RECT 707.100 315.000 708.900 321.600 ;
        RECT 710.100 315.600 711.900 321.600 ;
        RECT 722.400 315.000 724.200 327.600 ;
        RECT 727.500 326.100 729.900 327.600 ;
        RECT 727.500 315.600 729.300 326.100 ;
        RECT 730.200 323.100 732.000 324.900 ;
        RECT 730.500 315.000 732.300 321.600 ;
        RECT 743.100 315.600 744.900 327.600 ;
        RECT 746.100 326.700 753.900 327.600 ;
        RECT 746.100 315.600 747.900 326.700 ;
        RECT 749.100 315.000 750.900 325.800 ;
        RECT 752.100 315.600 753.900 326.700 ;
        RECT 764.700 321.600 765.900 334.950 ;
        RECT 767.100 333.150 768.900 334.950 ;
        RECT 785.100 333.150 786.900 334.950 ;
        RECT 791.100 322.800 792.000 334.950 ;
        RECT 785.400 321.900 792.000 322.800 ;
        RECT 785.400 321.600 786.900 321.900 ;
        RECT 764.100 315.600 765.900 321.600 ;
        RECT 767.100 315.000 768.900 321.600 ;
        RECT 782.100 315.000 783.900 321.600 ;
        RECT 785.100 315.600 786.900 321.600 ;
        RECT 791.100 321.600 792.000 321.900 ;
        RECT 806.100 321.600 807.300 334.950 ;
        RECT 808.950 330.450 811.050 331.050 ;
        RECT 823.950 330.450 826.050 331.050 ;
        RECT 808.950 329.550 826.050 330.450 ;
        RECT 808.950 328.950 811.050 329.550 ;
        RECT 823.950 328.950 826.050 329.550 ;
        RECT 827.100 321.600 828.000 341.700 ;
        RECT 833.400 337.050 834.300 344.400 ;
        RECT 848.100 345.300 849.900 350.400 ;
        RECT 851.100 346.200 852.900 351.000 ;
        RECT 854.100 345.300 855.900 350.400 ;
        RECT 848.100 343.950 855.900 345.300 ;
        RECT 857.100 344.400 858.900 350.400 ;
        RECT 857.100 342.300 858.300 344.400 ;
        RECT 854.700 341.400 858.300 342.300 ;
        RECT 872.100 341.400 873.900 351.000 ;
        RECT 878.700 342.000 880.500 350.400 ;
        RECT 883.950 348.450 886.050 349.050 ;
        RECT 889.950 348.450 892.050 349.050 ;
        RECT 883.950 347.550 892.050 348.450 ;
        RECT 883.950 346.950 886.050 347.550 ;
        RECT 889.950 346.950 892.050 347.550 ;
        RECT 893.100 344.400 894.900 350.400 ;
        RECT 893.700 342.300 894.900 344.400 ;
        RECT 896.100 345.300 897.900 350.400 ;
        RECT 899.100 346.200 900.900 351.000 ;
        RECT 902.100 345.300 903.900 350.400 ;
        RECT 896.100 343.950 903.900 345.300 ;
        RECT 917.100 344.400 918.900 350.400 ;
        RECT 917.700 342.300 918.900 344.400 ;
        RECT 920.100 345.300 921.900 350.400 ;
        RECT 923.100 346.200 924.900 351.000 ;
        RECT 926.100 345.300 927.900 350.400 ;
        RECT 920.100 343.950 927.900 345.300 ;
        RECT 851.100 337.050 852.900 338.850 ;
        RECT 854.700 337.050 855.900 341.400 ;
        RECT 878.700 340.800 882.000 342.000 ;
        RECT 893.700 341.400 897.300 342.300 ;
        RECT 917.700 341.400 921.300 342.300 ;
        RECT 868.950 339.450 871.050 340.050 ;
        RECT 857.100 337.050 858.900 338.850 ;
        RECT 863.550 338.550 871.050 339.450 ;
        RECT 829.500 334.950 831.600 337.050 ;
        RECT 832.800 334.950 834.900 337.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 829.200 333.150 831.000 334.950 ;
        RECT 833.400 327.600 834.300 334.950 ;
        RECT 848.100 333.150 849.900 334.950 ;
        RECT 854.700 327.600 855.900 334.950 ;
        RECT 863.550 334.050 864.450 338.550 ;
        RECT 868.950 337.950 871.050 338.550 ;
        RECT 872.100 337.050 873.900 338.850 ;
        RECT 878.100 337.050 879.900 338.850 ;
        RECT 881.100 337.050 882.000 340.800 ;
        RECT 893.100 337.050 894.900 338.850 ;
        RECT 896.100 337.050 897.300 341.400 ;
        RECT 912.000 339.450 916.050 340.050 ;
        RECT 899.100 337.050 900.900 338.850 ;
        RECT 911.550 337.950 916.050 339.450 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 859.950 332.550 864.450 334.050 ;
        RECT 875.100 333.150 876.900 334.950 ;
        RECT 859.950 331.950 864.000 332.550 ;
        RECT 788.100 315.000 789.900 321.000 ;
        RECT 791.100 315.600 792.900 321.600 ;
        RECT 803.100 315.000 804.900 321.600 ;
        RECT 806.100 315.600 807.900 321.600 ;
        RECT 809.100 315.000 810.900 321.600 ;
        RECT 824.100 315.000 825.900 321.600 ;
        RECT 827.100 315.600 828.900 321.600 ;
        RECT 830.100 315.000 831.900 327.000 ;
        RECT 833.100 315.600 834.900 327.600 ;
        RECT 848.400 315.000 850.200 327.600 ;
        RECT 853.500 326.100 855.900 327.600 ;
        RECT 853.500 315.600 855.300 326.100 ;
        RECT 856.200 323.100 858.000 324.900 ;
        RECT 881.100 322.800 882.000 334.950 ;
        RECT 896.100 327.600 897.300 334.950 ;
        RECT 902.100 333.150 903.900 334.950 ;
        RECT 911.550 334.050 912.450 337.950 ;
        RECT 917.100 337.050 918.900 338.850 ;
        RECT 920.100 337.050 921.300 341.400 ;
        RECT 923.100 337.050 924.900 338.850 ;
        RECT 916.950 334.950 919.050 337.050 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 911.550 332.550 916.050 334.050 ;
        RECT 912.000 331.950 916.050 332.550 ;
        RECT 920.100 327.600 921.300 334.950 ;
        RECT 926.100 333.150 927.900 334.950 ;
        RECT 896.100 326.100 898.500 327.600 ;
        RECT 894.000 323.100 895.800 324.900 ;
        RECT 875.400 321.900 882.000 322.800 ;
        RECT 875.400 321.600 876.900 321.900 ;
        RECT 856.500 315.000 858.300 321.600 ;
        RECT 872.100 315.000 873.900 321.600 ;
        RECT 875.100 315.600 876.900 321.600 ;
        RECT 881.100 321.600 882.000 321.900 ;
        RECT 878.100 315.000 879.900 321.000 ;
        RECT 881.100 315.600 882.900 321.600 ;
        RECT 893.700 315.000 895.500 321.600 ;
        RECT 896.700 315.600 898.500 326.100 ;
        RECT 901.800 315.000 903.600 327.600 ;
        RECT 920.100 326.100 922.500 327.600 ;
        RECT 918.000 323.100 919.800 324.900 ;
        RECT 917.700 315.000 919.500 321.600 ;
        RECT 920.700 315.600 922.500 326.100 ;
        RECT 925.800 315.000 927.600 327.600 ;
        RECT 11.100 305.400 12.900 312.000 ;
        RECT 14.100 305.400 15.900 311.400 ;
        RECT 11.100 292.050 12.900 293.850 ;
        RECT 14.100 292.050 15.300 305.400 ;
        RECT 29.100 300.600 30.900 311.400 ;
        RECT 32.100 301.500 33.900 312.000 ;
        RECT 35.100 310.500 42.900 311.400 ;
        RECT 35.100 300.600 36.900 310.500 ;
        RECT 29.100 299.700 36.900 300.600 ;
        RECT 38.100 298.500 39.900 309.600 ;
        RECT 41.100 299.400 42.900 310.500 ;
        RECT 53.100 305.400 54.900 312.000 ;
        RECT 56.100 305.400 57.900 311.400 ;
        RECT 59.700 305.400 61.500 312.000 ;
        RECT 62.700 305.400 64.500 311.400 ;
        RECT 66.000 305.400 67.800 312.000 ;
        RECT 69.000 305.400 70.800 311.400 ;
        RECT 72.000 305.400 73.800 312.000 ;
        RECT 75.000 305.400 76.800 311.400 ;
        RECT 78.000 305.400 79.800 312.000 ;
        RECT 81.000 308.400 82.800 311.400 ;
        RECT 84.000 308.400 85.800 311.400 ;
        RECT 87.000 308.400 88.800 311.400 ;
        RECT 80.700 306.300 82.800 308.400 ;
        RECT 83.700 306.300 85.800 308.400 ;
        RECT 86.700 306.300 88.800 308.400 ;
        RECT 90.000 305.400 91.800 311.400 ;
        RECT 93.000 305.400 94.800 312.000 ;
        RECT 35.100 297.600 39.900 298.500 ;
        RECT 32.250 292.050 34.050 293.850 ;
        RECT 35.100 292.050 36.000 297.600 ;
        RECT 48.000 294.450 52.050 295.050 ;
        RECT 38.100 292.050 39.900 293.850 ;
        RECT 47.550 292.950 52.050 294.450 ;
        RECT 10.950 289.950 13.050 292.050 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 28.950 289.950 31.050 292.050 ;
        RECT 31.950 289.950 34.050 292.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 14.100 279.600 15.300 289.950 ;
        RECT 29.250 288.150 31.050 289.950 ;
        RECT 35.100 282.600 36.300 289.950 ;
        RECT 41.100 288.150 42.900 289.950 ;
        RECT 47.550 289.050 48.450 292.950 ;
        RECT 53.100 292.050 54.900 293.850 ;
        RECT 56.100 292.050 57.300 305.400 ;
        RECT 63.000 295.050 64.500 305.400 ;
        RECT 69.000 304.500 70.200 305.400 ;
        RECT 62.100 292.950 64.500 295.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 47.550 287.550 52.050 289.050 ;
        RECT 48.000 286.950 52.050 287.550 ;
        RECT 11.100 276.000 12.900 279.600 ;
        RECT 14.100 276.600 15.900 279.600 ;
        RECT 29.700 276.000 31.500 282.600 ;
        RECT 34.200 276.600 36.000 282.600 ;
        RECT 38.700 276.000 40.500 282.600 ;
        RECT 56.100 279.600 57.300 289.950 ;
        RECT 63.000 279.600 64.500 292.950 ;
        RECT 53.100 276.000 54.900 279.600 ;
        RECT 56.100 276.600 57.900 279.600 ;
        RECT 59.700 276.000 61.500 279.600 ;
        RECT 62.700 276.600 64.500 279.600 ;
        RECT 66.300 303.600 70.200 304.500 ;
        RECT 66.300 300.300 67.200 303.600 ;
        RECT 71.100 302.400 72.900 303.000 ;
        RECT 75.600 302.400 76.800 305.400 ;
        RECT 83.700 304.500 85.800 305.400 ;
        RECT 77.700 303.300 85.800 304.500 ;
        RECT 77.700 302.700 79.500 303.300 ;
        RECT 71.100 301.200 76.800 302.400 ;
        RECT 89.100 301.500 91.800 305.400 ;
        RECT 96.000 303.900 97.800 311.400 ;
        RECT 99.900 305.400 101.700 312.000 ;
        RECT 102.900 305.400 104.700 311.400 ;
        RECT 105.900 308.400 107.700 311.400 ;
        RECT 108.900 308.400 110.700 311.400 ;
        RECT 105.600 306.300 107.700 308.400 ;
        RECT 108.600 306.300 110.700 308.400 ;
        RECT 112.500 305.400 114.300 312.000 ;
        RECT 94.500 301.800 97.800 303.900 ;
        RECT 103.200 303.300 105.300 305.400 ;
        RECT 115.500 302.400 117.300 311.400 ;
        RECT 118.500 305.400 120.300 312.000 ;
        RECT 121.500 306.300 123.300 311.400 ;
        RECT 121.500 305.400 123.600 306.300 ;
        RECT 124.500 305.400 126.300 312.000 ;
        RECT 122.700 304.500 123.600 305.400 ;
        RECT 122.700 303.600 126.300 304.500 ;
        RECT 120.000 302.400 121.800 302.700 ;
        RECT 80.700 300.300 82.800 301.500 ;
        RECT 66.300 299.400 82.800 300.300 ;
        RECT 86.100 300.600 88.200 301.500 ;
        RECT 102.600 301.200 121.800 302.400 ;
        RECT 102.600 300.600 103.800 301.200 ;
        RECT 120.000 300.900 121.800 301.200 ;
        RECT 86.100 299.400 103.800 300.600 ;
        RECT 106.500 299.700 108.600 300.300 ;
        RECT 116.700 299.700 118.500 300.300 ;
        RECT 66.300 282.600 67.200 299.400 ;
        RECT 106.500 298.500 118.500 299.700 ;
        RECT 68.100 297.300 103.800 298.500 ;
        RECT 106.500 298.200 108.600 298.500 ;
        RECT 68.100 296.700 69.900 297.300 ;
        RECT 102.600 296.700 103.800 297.300 ;
        RECT 71.100 292.950 73.200 295.050 ;
        RECT 71.700 290.100 73.200 292.950 ;
        RECT 75.300 292.800 80.400 294.600 ;
        RECT 79.500 291.300 80.400 292.800 ;
        RECT 83.100 294.300 84.900 296.100 ;
        RECT 89.100 295.800 91.200 296.100 ;
        RECT 102.600 295.800 116.100 296.700 ;
        RECT 83.100 293.100 84.000 294.300 ;
        RECT 89.100 294.000 93.000 295.800 ;
        RECT 94.500 294.300 96.600 295.200 ;
        RECT 114.300 295.050 116.100 295.800 ;
        RECT 94.500 293.100 105.600 294.300 ;
        RECT 114.300 293.250 118.200 295.050 ;
        RECT 83.100 292.200 96.600 293.100 ;
        RECT 103.800 292.500 105.600 293.100 ;
        RECT 116.100 292.950 118.200 293.250 ;
        RECT 122.100 292.950 124.200 295.050 ;
        RECT 122.100 291.300 123.900 292.950 ;
        RECT 79.500 290.100 123.900 291.300 ;
        RECT 71.700 288.600 78.300 290.100 ;
        RECT 68.100 285.900 75.900 287.700 ;
        RECT 76.800 287.100 93.900 288.600 ;
        RECT 91.800 286.500 93.900 287.100 ;
        RECT 98.100 288.000 100.200 289.050 ;
        RECT 98.100 287.100 103.200 288.000 ;
        RECT 106.800 287.400 108.600 289.200 ;
        RECT 125.100 287.400 126.300 303.600 ;
        RECT 140.100 300.600 141.900 311.400 ;
        RECT 143.100 301.500 144.900 312.000 ;
        RECT 146.100 310.500 153.900 311.400 ;
        RECT 146.100 300.600 147.900 310.500 ;
        RECT 140.100 299.700 147.900 300.600 ;
        RECT 149.100 298.500 150.900 309.600 ;
        RECT 152.100 299.400 153.900 310.500 ;
        RECT 167.100 305.400 168.900 311.400 ;
        RECT 170.100 306.000 171.900 312.000 ;
        RECT 168.000 305.100 168.900 305.400 ;
        RECT 173.100 305.400 174.900 311.400 ;
        RECT 176.100 305.400 177.900 312.000 ;
        RECT 173.100 305.100 174.600 305.400 ;
        RECT 168.000 304.200 174.600 305.100 ;
        RECT 146.100 297.600 150.900 298.500 ;
        RECT 136.950 294.450 139.050 295.050 ;
        RECT 98.100 286.950 100.200 287.100 ;
        RECT 74.400 282.600 75.900 285.900 ;
        RECT 92.100 284.700 93.900 286.500 ;
        RECT 101.400 286.200 103.200 287.100 ;
        RECT 107.700 284.400 108.600 287.400 ;
        RECT 109.500 286.200 126.300 287.400 ;
        RECT 109.500 285.300 111.600 286.200 ;
        RECT 120.300 284.700 122.100 285.300 ;
        RECT 80.100 282.600 86.700 284.400 ;
        RECT 101.400 283.200 108.600 284.400 ;
        RECT 113.700 283.500 122.100 284.700 ;
        RECT 101.400 282.600 102.300 283.200 ;
        RECT 104.400 282.600 106.200 283.200 ;
        RECT 113.700 282.600 115.200 283.500 ;
        RECT 125.100 282.600 126.300 286.200 ;
        RECT 128.550 293.550 139.050 294.450 ;
        RECT 128.550 285.900 129.450 293.550 ;
        RECT 136.950 292.950 139.050 293.550 ;
        RECT 143.250 292.050 145.050 293.850 ;
        RECT 146.100 292.050 147.000 297.600 ;
        RECT 149.100 292.050 150.900 293.850 ;
        RECT 168.000 292.050 168.900 304.200 ;
        RECT 188.100 299.400 189.900 312.000 ;
        RECT 193.200 300.600 195.000 311.400 ;
        RECT 209.100 305.400 210.900 312.000 ;
        RECT 212.100 305.400 213.900 311.400 ;
        RECT 224.100 305.400 225.900 312.000 ;
        RECT 227.100 305.400 228.900 311.400 ;
        RECT 230.100 306.000 231.900 312.000 ;
        RECT 191.400 299.400 195.000 300.600 ;
        RECT 169.950 297.450 172.050 298.050 ;
        RECT 181.950 297.450 184.050 298.050 ;
        RECT 187.950 297.450 190.050 298.050 ;
        RECT 169.950 296.550 190.050 297.450 ;
        RECT 169.950 295.950 172.050 296.550 ;
        RECT 181.950 295.950 184.050 296.550 ;
        RECT 187.950 295.950 190.050 296.550 ;
        RECT 173.100 292.050 174.900 293.850 ;
        RECT 188.250 292.050 190.050 293.850 ;
        RECT 191.400 292.050 192.300 299.400 ;
        RECT 194.100 292.050 195.900 293.850 ;
        RECT 209.100 292.050 210.900 293.850 ;
        RECT 212.100 292.050 213.300 305.400 ;
        RECT 227.400 305.100 228.900 305.400 ;
        RECT 233.100 305.400 234.900 311.400 ;
        RECT 233.100 305.100 234.000 305.400 ;
        RECT 227.400 304.200 234.000 305.100 ;
        RECT 214.950 294.450 219.000 295.050 ;
        RECT 214.950 292.950 219.450 294.450 ;
        RECT 139.950 289.950 142.050 292.050 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 140.250 288.150 142.050 289.950 ;
        RECT 127.950 283.800 130.050 285.900 ;
        RECT 133.950 285.450 136.050 286.050 ;
        RECT 139.950 285.450 142.050 286.050 ;
        RECT 133.950 284.550 142.050 285.450 ;
        RECT 133.950 283.950 136.050 284.550 ;
        RECT 139.950 283.950 142.050 284.550 ;
        RECT 146.100 282.600 147.300 289.950 ;
        RECT 152.100 288.150 153.900 289.950 ;
        RECT 168.000 286.200 168.900 289.950 ;
        RECT 170.100 288.150 171.900 289.950 ;
        RECT 176.100 288.150 177.900 289.950 ;
        RECT 168.000 285.000 171.300 286.200 ;
        RECT 66.300 276.600 68.100 282.600 ;
        RECT 71.700 276.000 73.500 282.600 ;
        RECT 74.400 281.400 78.600 282.600 ;
        RECT 76.800 276.600 78.600 281.400 ;
        RECT 80.700 279.600 82.800 281.700 ;
        RECT 83.700 279.600 85.800 281.700 ;
        RECT 86.700 279.600 88.800 281.700 ;
        RECT 89.700 279.600 91.800 281.700 ;
        RECT 95.100 280.500 97.800 282.600 ;
        RECT 99.600 281.400 102.300 282.600 ;
        RECT 99.600 280.500 101.400 281.400 ;
        RECT 81.000 276.600 82.800 279.600 ;
        RECT 84.000 276.600 85.800 279.600 ;
        RECT 87.000 276.600 88.800 279.600 ;
        RECT 90.000 276.600 91.800 279.600 ;
        RECT 93.000 276.000 94.800 279.600 ;
        RECT 96.000 276.600 97.800 280.500 ;
        RECT 103.200 279.600 105.300 281.700 ;
        RECT 106.200 279.600 108.300 281.700 ;
        RECT 109.200 279.600 111.300 281.700 ;
        RECT 100.500 276.000 102.300 279.600 ;
        RECT 103.500 276.600 105.300 279.600 ;
        RECT 106.500 276.600 108.300 279.600 ;
        RECT 109.500 276.600 111.300 279.600 ;
        RECT 113.700 276.600 115.500 282.600 ;
        RECT 119.100 276.000 120.900 282.600 ;
        RECT 124.500 276.600 126.300 282.600 ;
        RECT 140.700 276.000 142.500 282.600 ;
        RECT 145.200 276.600 147.000 282.600 ;
        RECT 149.700 276.000 151.500 282.600 ;
        RECT 169.500 276.600 171.300 285.000 ;
        RECT 176.100 276.000 177.900 285.600 ;
        RECT 191.400 279.600 192.300 289.950 ;
        RECT 212.100 279.600 213.300 289.950 ;
        RECT 218.550 289.050 219.450 292.950 ;
        RECT 227.100 292.050 228.900 293.850 ;
        RECT 233.100 292.050 234.000 304.200 ;
        RECT 245.400 299.400 247.200 312.000 ;
        RECT 250.500 300.900 252.300 311.400 ;
        RECT 253.500 305.400 255.300 312.000 ;
        RECT 253.200 302.100 255.000 303.900 ;
        RECT 267.600 300.900 269.400 311.400 ;
        RECT 250.500 299.400 252.900 300.900 ;
        RECT 245.100 292.050 246.900 293.850 ;
        RECT 251.700 292.050 252.900 299.400 ;
        RECT 267.000 299.400 269.400 300.900 ;
        RECT 270.600 299.400 272.400 312.000 ;
        RECT 275.100 299.400 276.900 311.400 ;
        RECT 290.400 299.400 292.200 312.000 ;
        RECT 295.500 300.900 297.300 311.400 ;
        RECT 298.500 305.400 300.300 312.000 ;
        RECT 311.700 305.400 313.500 312.000 ;
        RECT 298.200 302.100 300.000 303.900 ;
        RECT 312.000 302.100 313.800 303.900 ;
        RECT 314.700 300.900 316.500 311.400 ;
        RECT 295.500 299.400 297.900 300.900 ;
        RECT 267.000 292.050 268.200 299.400 ;
        RECT 275.700 297.900 276.900 299.400 ;
        RECT 269.100 296.700 276.900 297.900 ;
        RECT 292.950 297.450 295.050 298.050 ;
        RECT 269.100 296.100 270.900 296.700 ;
        RECT 284.550 296.550 295.050 297.450 ;
        RECT 223.950 289.950 226.050 292.050 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 266.100 289.950 268.200 292.050 ;
        RECT 218.550 287.550 223.050 289.050 ;
        RECT 224.100 288.150 225.900 289.950 ;
        RECT 230.100 288.150 231.900 289.950 ;
        RECT 219.000 286.950 223.050 287.550 ;
        RECT 233.100 286.200 234.000 289.950 ;
        RECT 248.100 288.150 249.900 289.950 ;
        RECT 188.100 276.000 189.900 279.600 ;
        RECT 191.100 276.600 192.900 279.600 ;
        RECT 194.100 276.000 195.900 279.600 ;
        RECT 209.100 276.000 210.900 279.600 ;
        RECT 212.100 276.600 213.900 279.600 ;
        RECT 224.100 276.000 225.900 285.600 ;
        RECT 230.700 285.000 234.000 286.200 ;
        RECT 251.700 285.600 252.900 289.950 ;
        RECT 254.100 288.150 255.900 289.950 ;
        RECT 230.700 276.600 232.500 285.000 ;
        RECT 251.700 284.700 255.300 285.600 ;
        RECT 245.100 281.700 252.900 283.050 ;
        RECT 245.100 276.600 246.900 281.700 ;
        RECT 248.100 276.000 249.900 280.800 ;
        RECT 251.100 276.600 252.900 281.700 ;
        RECT 254.100 282.600 255.300 284.700 ;
        RECT 266.100 282.600 267.000 289.950 ;
        RECT 269.400 285.600 270.300 296.100 ;
        RECT 271.200 292.050 273.000 293.850 ;
        RECT 271.500 289.950 273.600 292.050 ;
        RECT 274.800 289.950 276.900 292.050 ;
        RECT 274.800 288.150 276.600 289.950 ;
        RECT 284.550 289.050 285.450 296.550 ;
        RECT 292.950 295.950 295.050 296.550 ;
        RECT 290.100 292.050 291.900 293.850 ;
        RECT 296.700 292.050 297.900 299.400 ;
        RECT 314.100 299.400 316.500 300.900 ;
        RECT 319.800 299.400 321.600 312.000 ;
        RECT 335.100 305.400 336.900 312.000 ;
        RECT 338.100 305.400 339.900 311.400 ;
        RECT 341.100 305.400 342.900 312.000 ;
        RECT 301.950 297.450 304.050 298.050 ;
        RECT 310.950 297.450 313.050 298.050 ;
        RECT 301.950 296.550 313.050 297.450 ;
        RECT 301.950 295.950 304.050 296.550 ;
        RECT 310.950 295.950 313.050 296.550 ;
        RECT 314.100 292.050 315.300 299.400 ;
        RECT 322.950 294.450 327.000 295.050 ;
        RECT 320.100 292.050 321.900 293.850 ;
        RECT 322.950 292.950 327.450 294.450 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 298.950 289.950 301.050 292.050 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 284.550 287.550 289.050 289.050 ;
        RECT 293.100 288.150 294.900 289.950 ;
        RECT 285.000 286.950 289.050 287.550 ;
        RECT 268.200 284.700 270.300 285.600 ;
        RECT 296.700 285.600 297.900 289.950 ;
        RECT 299.100 288.150 300.900 289.950 ;
        RECT 311.100 288.150 312.900 289.950 ;
        RECT 314.100 285.600 315.300 289.950 ;
        RECT 317.100 288.150 318.900 289.950 ;
        RECT 326.550 289.050 327.450 292.950 ;
        RECT 338.100 292.050 339.300 305.400 ;
        RECT 353.100 300.300 354.900 311.400 ;
        RECT 356.100 301.500 357.900 312.000 ;
        RECT 360.600 300.300 362.400 311.400 ;
        RECT 364.800 301.500 366.900 312.000 ;
        RECT 368.100 300.600 369.900 311.400 ;
        RECT 380.100 305.400 381.900 312.000 ;
        RECT 383.100 305.400 384.900 311.400 ;
        RECT 386.100 305.400 387.900 312.000 ;
        RECT 398.100 305.400 399.900 312.000 ;
        RECT 401.100 305.400 402.900 311.400 ;
        RECT 404.100 305.400 405.900 312.000 ;
        RECT 353.100 299.100 357.900 300.300 ;
        RECT 360.600 299.400 363.900 300.300 ;
        RECT 355.800 298.200 357.900 299.100 ;
        RECT 355.800 297.300 361.200 298.200 ;
        RECT 359.400 295.500 361.200 297.300 ;
        RECT 362.700 295.050 363.900 299.400 ;
        RECT 364.800 299.400 369.900 300.600 ;
        RECT 364.800 298.500 366.900 299.400 ;
        RECT 362.100 294.300 364.200 295.050 ;
        RECT 375.000 294.450 379.050 295.050 ;
        RECT 357.900 292.200 359.700 294.000 ;
        RECT 361.200 292.950 364.200 294.300 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 322.950 287.550 327.450 289.050 ;
        RECT 335.250 288.150 337.050 289.950 ;
        RECT 322.950 286.950 327.000 287.550 ;
        RECT 296.700 284.700 300.300 285.600 ;
        RECT 268.200 283.800 273.600 284.700 ;
        RECT 254.100 276.600 255.900 282.600 ;
        RECT 266.100 276.600 267.900 282.600 ;
        RECT 269.100 276.000 270.900 282.000 ;
        RECT 272.700 279.600 273.600 283.800 ;
        RECT 290.100 281.700 297.900 283.050 ;
        RECT 272.100 276.600 273.900 279.600 ;
        RECT 275.100 276.600 276.900 279.600 ;
        RECT 290.100 276.600 291.900 281.700 ;
        RECT 275.700 276.000 276.900 276.600 ;
        RECT 293.100 276.000 294.900 280.800 ;
        RECT 296.100 276.600 297.900 281.700 ;
        RECT 299.100 282.600 300.300 284.700 ;
        RECT 311.700 284.700 315.300 285.600 ;
        RECT 338.100 284.700 339.300 289.950 ;
        RECT 341.100 288.150 342.900 289.950 ;
        RECT 353.100 289.800 355.200 292.050 ;
        RECT 357.900 290.100 360.000 292.200 ;
        RECT 353.400 289.200 355.200 289.800 ;
        RECT 353.400 288.000 360.000 289.200 ;
        RECT 357.900 287.100 360.000 288.000 ;
        RECT 355.500 285.000 357.600 285.600 ;
        RECT 358.500 285.300 360.300 287.100 ;
        RECT 361.200 286.200 362.100 292.950 ;
        RECT 367.800 292.050 369.600 293.850 ;
        RECT 374.550 292.950 379.050 294.450 ;
        RECT 363.000 290.100 364.800 291.900 ;
        RECT 363.000 288.000 365.100 290.100 ;
        RECT 367.800 289.950 369.900 292.050 ;
        RECT 374.550 289.050 375.450 292.950 ;
        RECT 383.100 292.050 384.300 305.400 ;
        RECT 401.100 292.050 402.300 305.400 ;
        RECT 416.400 299.400 418.200 312.000 ;
        RECT 421.500 300.900 423.300 311.400 ;
        RECT 424.500 305.400 426.300 312.000 ;
        RECT 440.100 305.400 441.900 312.000 ;
        RECT 443.100 305.400 444.900 311.400 ;
        RECT 458.100 305.400 459.900 312.000 ;
        RECT 461.100 305.400 462.900 311.400 ;
        RECT 464.100 305.400 465.900 312.000 ;
        RECT 424.200 302.100 426.000 303.900 ;
        RECT 421.500 299.400 423.900 300.900 ;
        RECT 403.950 297.450 406.050 298.050 ;
        RECT 415.950 297.450 418.050 298.050 ;
        RECT 403.950 296.550 418.050 297.450 ;
        RECT 403.950 295.950 406.050 296.550 ;
        RECT 415.950 295.950 418.050 296.550 ;
        RECT 416.100 292.050 417.900 293.850 ;
        RECT 422.700 292.050 423.900 299.400 ;
        RECT 440.100 292.050 441.900 293.850 ;
        RECT 443.100 292.050 444.300 305.400 ;
        RECT 461.700 292.050 462.900 305.400 ;
        RECT 479.100 300.300 480.900 311.400 ;
        RECT 482.100 301.200 483.900 312.000 ;
        RECT 485.100 300.300 486.900 311.400 ;
        RECT 479.100 299.400 486.900 300.300 ;
        RECT 488.100 299.400 489.900 311.400 ;
        RECT 503.100 299.400 504.900 312.000 ;
        RECT 507.600 299.400 510.900 311.400 ;
        RECT 513.600 299.400 515.400 312.000 ;
        RECT 530.100 305.400 531.900 312.000 ;
        RECT 533.100 305.400 534.900 311.400 ;
        RECT 536.100 305.400 537.900 312.000 ;
        RECT 482.250 292.050 484.050 293.850 ;
        RECT 488.700 292.050 489.600 299.400 ;
        RECT 499.950 294.450 502.050 298.050 ;
        RECT 497.550 294.000 502.050 294.450 ;
        RECT 497.550 293.550 501.450 294.000 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 374.550 287.550 379.050 289.050 ;
        RECT 380.250 288.150 382.050 289.950 ;
        RECT 375.000 286.950 379.050 287.550 ;
        RECT 311.700 282.600 312.900 284.700 ;
        RECT 338.100 283.800 342.300 284.700 ;
        RECT 299.100 276.600 300.900 282.600 ;
        RECT 311.100 276.600 312.900 282.600 ;
        RECT 314.100 281.700 321.900 283.050 ;
        RECT 314.100 276.600 315.900 281.700 ;
        RECT 317.100 276.000 318.900 280.800 ;
        RECT 320.100 276.600 321.900 281.700 ;
        RECT 335.400 276.000 337.200 282.600 ;
        RECT 340.500 276.600 342.300 283.800 ;
        RECT 353.100 283.500 357.600 285.000 ;
        RECT 361.200 284.100 364.200 286.200 ;
        RECT 353.100 282.600 354.600 283.500 ;
        RECT 353.100 276.600 354.900 282.600 ;
        RECT 361.200 282.000 362.100 284.100 ;
        RECT 365.400 283.500 367.500 285.900 ;
        RECT 383.100 284.700 384.300 289.950 ;
        RECT 386.100 288.150 387.900 289.950 ;
        RECT 398.250 288.150 400.050 289.950 ;
        RECT 401.100 284.700 402.300 289.950 ;
        RECT 404.100 288.150 405.900 289.950 ;
        RECT 419.100 288.150 420.900 289.950 ;
        RECT 422.700 285.600 423.900 289.950 ;
        RECT 425.100 288.150 426.900 289.950 ;
        RECT 422.700 284.700 426.300 285.600 ;
        RECT 383.100 283.800 387.300 284.700 ;
        RECT 401.100 283.800 405.300 284.700 ;
        RECT 365.400 282.600 369.900 283.500 ;
        RECT 356.100 276.000 357.900 281.700 ;
        RECT 360.300 276.600 362.100 282.000 ;
        RECT 364.800 276.000 366.600 281.700 ;
        RECT 368.100 276.600 369.900 282.600 ;
        RECT 380.400 276.000 382.200 282.600 ;
        RECT 385.500 276.600 387.300 283.800 ;
        RECT 398.400 276.000 400.200 282.600 ;
        RECT 403.500 276.600 405.300 283.800 ;
        RECT 416.100 281.700 423.900 283.050 ;
        RECT 416.100 276.600 417.900 281.700 ;
        RECT 419.100 276.000 420.900 280.800 ;
        RECT 422.100 276.600 423.900 281.700 ;
        RECT 425.100 282.600 426.300 284.700 ;
        RECT 425.100 276.600 426.900 282.600 ;
        RECT 443.100 279.600 444.300 289.950 ;
        RECT 458.100 288.150 459.900 289.950 ;
        RECT 461.700 284.700 462.900 289.950 ;
        RECT 463.950 288.150 465.750 289.950 ;
        RECT 479.100 288.150 480.900 289.950 ;
        RECT 485.250 288.150 487.050 289.950 ;
        RECT 458.700 283.800 462.900 284.700 ;
        RECT 440.100 276.000 441.900 279.600 ;
        RECT 443.100 276.600 444.900 279.600 ;
        RECT 458.700 276.600 460.500 283.800 ;
        RECT 488.700 282.600 489.600 289.950 ;
        RECT 490.950 288.450 493.050 289.050 ;
        RECT 497.550 288.450 498.450 293.550 ;
        RECT 503.100 292.050 504.900 293.850 ;
        RECT 508.950 292.050 510.000 299.400 ;
        RECT 526.950 294.450 529.050 295.050 ;
        RECT 514.950 292.050 516.750 293.850 ;
        RECT 521.550 293.550 529.050 294.450 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 490.950 287.550 498.450 288.450 ;
        RECT 506.250 288.150 508.050 289.950 ;
        RECT 508.950 289.950 511.050 292.050 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 514.950 289.950 517.050 292.050 ;
        RECT 490.950 286.950 493.050 287.550 ;
        RECT 508.950 285.300 510.000 289.950 ;
        RECT 511.950 288.150 513.750 289.950 ;
        RECT 521.550 289.050 522.450 293.550 ;
        RECT 526.950 292.950 529.050 293.550 ;
        RECT 533.700 292.050 534.900 305.400 ;
        RECT 549.600 299.400 551.400 312.000 ;
        RECT 554.100 299.400 557.400 311.400 ;
        RECT 560.100 299.400 561.900 312.000 ;
        RECT 572.100 305.400 573.900 312.000 ;
        RECT 575.100 305.400 576.900 311.400 ;
        RECT 578.100 305.400 579.900 312.000 ;
        RECT 593.100 305.400 594.900 312.000 ;
        RECT 596.100 305.400 597.900 311.400 ;
        RECT 599.100 305.400 600.900 312.000 ;
        RECT 614.100 305.400 615.900 312.000 ;
        RECT 617.100 305.400 618.900 311.400 ;
        RECT 620.100 305.400 621.900 312.000 ;
        RECT 635.700 305.400 637.500 312.000 ;
        RECT 565.950 303.450 568.050 303.900 ;
        RECT 571.950 303.450 574.050 304.050 ;
        RECT 565.950 302.550 574.050 303.450 ;
        RECT 565.950 301.800 568.050 302.550 ;
        RECT 571.950 301.950 574.050 302.550 ;
        RECT 548.250 292.050 550.050 293.850 ;
        RECT 555.000 292.050 556.050 299.400 ;
        RECT 559.950 297.450 562.050 298.050 ;
        RECT 571.950 297.450 574.050 298.050 ;
        RECT 559.950 296.550 574.050 297.450 ;
        RECT 559.950 295.950 562.050 296.550 ;
        RECT 571.950 295.950 574.050 296.550 ;
        RECT 560.100 292.050 561.900 293.850 ;
        RECT 575.700 292.050 576.900 305.400 ;
        RECT 580.950 294.450 585.000 295.050 ;
        RECT 580.950 292.950 585.450 294.450 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 535.950 289.950 538.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 517.950 287.550 522.450 289.050 ;
        RECT 530.100 288.150 531.900 289.950 ;
        RECT 517.950 286.950 522.000 287.550 ;
        RECT 508.950 284.100 513.300 285.300 ;
        RECT 533.700 284.700 534.900 289.950 ;
        RECT 535.950 288.150 537.750 289.950 ;
        RECT 551.250 288.150 553.050 289.950 ;
        RECT 555.000 285.300 556.050 289.950 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 559.950 289.950 562.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 556.950 288.150 558.750 289.950 ;
        RECT 572.100 288.150 573.900 289.950 ;
        RECT 463.800 276.000 465.600 282.600 ;
        RECT 480.000 276.000 481.800 282.600 ;
        RECT 484.500 281.400 489.600 282.600 ;
        RECT 503.100 282.000 510.900 282.900 ;
        RECT 512.400 282.600 513.300 284.100 ;
        RECT 530.700 283.800 534.900 284.700 ;
        RECT 551.700 284.100 556.050 285.300 ;
        RECT 575.700 284.700 576.900 289.950 ;
        RECT 577.950 288.150 579.750 289.950 ;
        RECT 584.550 288.450 585.450 292.950 ;
        RECT 596.700 292.050 597.900 305.400 ;
        RECT 598.950 297.450 601.050 298.200 ;
        RECT 607.950 297.450 610.050 298.050 ;
        RECT 598.950 296.550 610.050 297.450 ;
        RECT 598.950 296.100 601.050 296.550 ;
        RECT 607.950 295.950 610.050 296.550 ;
        RECT 617.700 292.050 618.900 305.400 ;
        RECT 636.000 302.100 637.800 303.900 ;
        RECT 638.700 300.900 640.500 311.400 ;
        RECT 638.100 299.400 640.500 300.900 ;
        RECT 643.800 299.400 645.600 312.000 ;
        RECT 656.100 305.400 657.900 312.000 ;
        RECT 659.100 305.400 660.900 311.400 ;
        RECT 671.700 305.400 673.500 312.000 ;
        RECT 625.950 297.450 628.050 298.050 ;
        RECT 634.950 297.450 637.050 298.050 ;
        RECT 625.950 296.550 637.050 297.450 ;
        RECT 625.950 295.950 628.050 296.550 ;
        RECT 634.950 295.950 637.050 296.550 ;
        RECT 638.100 292.050 639.300 299.400 ;
        RECT 644.100 292.050 645.900 293.850 ;
        RECT 656.100 292.050 657.900 293.850 ;
        RECT 659.100 292.050 660.300 305.400 ;
        RECT 672.000 302.100 673.800 303.900 ;
        RECT 674.700 300.900 676.500 311.400 ;
        RECT 674.100 299.400 676.500 300.900 ;
        RECT 679.800 299.400 681.600 312.000 ;
        RECT 692.100 305.400 693.900 312.000 ;
        RECT 695.100 305.400 696.900 311.400 ;
        RECT 674.100 292.050 675.300 299.400 ;
        RECT 687.000 294.450 691.050 295.050 ;
        RECT 680.100 292.050 681.900 293.850 ;
        RECT 686.550 292.950 691.050 294.450 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 673.950 289.950 676.050 292.050 ;
        RECT 676.950 289.950 679.050 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 589.950 288.450 592.050 289.050 ;
        RECT 584.550 287.550 592.050 288.450 ;
        RECT 593.100 288.150 594.900 289.950 ;
        RECT 589.950 286.950 592.050 287.550 ;
        RECT 596.700 284.700 597.900 289.950 ;
        RECT 598.950 288.150 600.750 289.950 ;
        RECT 614.100 288.150 615.900 289.950 ;
        RECT 617.700 284.700 618.900 289.950 ;
        RECT 619.950 288.150 621.750 289.950 ;
        RECT 635.100 288.150 636.900 289.950 ;
        RECT 638.100 285.600 639.300 289.950 ;
        RECT 641.100 288.150 642.900 289.950 ;
        RECT 484.500 276.600 486.300 281.400 ;
        RECT 487.500 276.000 489.300 279.600 ;
        RECT 503.100 276.600 504.900 282.000 ;
        RECT 506.100 276.000 507.900 281.100 ;
        RECT 509.100 277.500 510.900 282.000 ;
        RECT 512.100 278.400 513.900 282.600 ;
        RECT 515.100 277.500 516.900 282.600 ;
        RECT 509.100 276.600 516.900 277.500 ;
        RECT 530.700 276.600 532.500 283.800 ;
        RECT 551.700 282.600 552.600 284.100 ;
        RECT 572.700 283.800 576.900 284.700 ;
        RECT 593.700 283.800 597.900 284.700 ;
        RECT 614.700 283.800 618.900 284.700 ;
        RECT 635.700 284.700 639.300 285.600 ;
        RECT 535.800 276.000 537.600 282.600 ;
        RECT 548.100 277.500 549.900 282.600 ;
        RECT 551.100 278.400 552.900 282.600 ;
        RECT 554.100 282.000 561.900 282.900 ;
        RECT 554.100 277.500 555.900 282.000 ;
        RECT 548.100 276.600 555.900 277.500 ;
        RECT 557.100 276.000 558.900 281.100 ;
        RECT 560.100 276.600 561.900 282.000 ;
        RECT 572.700 276.600 574.500 283.800 ;
        RECT 577.800 276.000 579.600 282.600 ;
        RECT 593.700 276.600 595.500 283.800 ;
        RECT 598.800 276.000 600.600 282.600 ;
        RECT 614.700 276.600 616.500 283.800 ;
        RECT 635.700 282.600 636.900 284.700 ;
        RECT 619.800 276.000 621.600 282.600 ;
        RECT 635.100 276.600 636.900 282.600 ;
        RECT 638.100 281.700 645.900 283.050 ;
        RECT 638.100 276.600 639.900 281.700 ;
        RECT 641.100 276.000 642.900 280.800 ;
        RECT 644.100 276.600 645.900 281.700 ;
        RECT 659.100 279.600 660.300 289.950 ;
        RECT 671.100 288.150 672.900 289.950 ;
        RECT 674.100 285.600 675.300 289.950 ;
        RECT 677.100 288.150 678.900 289.950 ;
        RECT 686.550 289.050 687.450 292.950 ;
        RECT 692.100 292.050 693.900 293.850 ;
        RECT 695.100 292.050 696.300 305.400 ;
        RECT 707.100 300.600 708.900 311.400 ;
        RECT 710.100 301.500 712.200 312.000 ;
        RECT 707.100 299.400 712.200 300.600 ;
        RECT 714.600 300.300 716.400 311.400 ;
        RECT 719.100 301.500 720.900 312.000 ;
        RECT 722.100 300.300 723.900 311.400 ;
        RECT 737.100 305.400 738.900 312.000 ;
        RECT 740.100 305.400 741.900 311.400 ;
        RECT 743.100 305.400 744.900 312.000 ;
        RECT 710.100 298.500 712.200 299.400 ;
        RECT 713.100 299.400 716.400 300.300 ;
        RECT 713.100 295.050 714.300 299.400 ;
        RECT 719.100 299.100 723.900 300.300 ;
        RECT 719.100 298.200 721.200 299.100 ;
        RECT 715.800 297.300 721.200 298.200 ;
        RECT 715.800 295.500 717.600 297.300 ;
        RECT 712.800 294.300 714.900 295.050 ;
        RECT 707.400 292.050 709.200 293.850 ;
        RECT 712.800 292.950 715.800 294.300 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 707.100 289.950 709.200 292.050 ;
        RECT 712.200 290.100 714.000 291.900 ;
        RECT 686.550 287.550 691.050 289.050 ;
        RECT 687.000 286.950 691.050 287.550 ;
        RECT 671.700 284.700 675.300 285.600 ;
        RECT 671.700 282.600 672.900 284.700 ;
        RECT 656.100 276.000 657.900 279.600 ;
        RECT 659.100 276.600 660.900 279.600 ;
        RECT 671.100 276.600 672.900 282.600 ;
        RECT 674.100 281.700 681.900 283.050 ;
        RECT 674.100 276.600 675.900 281.700 ;
        RECT 677.100 276.000 678.900 280.800 ;
        RECT 680.100 276.600 681.900 281.700 ;
        RECT 695.100 279.600 696.300 289.950 ;
        RECT 711.900 288.000 714.000 290.100 ;
        RECT 714.900 286.200 715.800 292.950 ;
        RECT 717.300 292.200 719.100 294.000 ;
        RECT 717.000 290.100 719.100 292.200 ;
        RECT 740.700 292.050 741.900 305.400 ;
        RECT 755.100 300.300 756.900 311.400 ;
        RECT 758.100 301.200 759.900 312.000 ;
        RECT 761.100 300.300 762.900 311.400 ;
        RECT 755.100 299.400 762.900 300.300 ;
        RECT 764.100 299.400 765.900 311.400 ;
        RECT 776.100 305.400 777.900 311.400 ;
        RECT 779.100 305.400 780.900 312.000 ;
        RECT 758.250 292.050 760.050 293.850 ;
        RECT 764.700 292.050 765.600 299.400 ;
        RECT 771.000 294.450 775.050 295.050 ;
        RECT 770.550 292.950 775.050 294.450 ;
        RECT 721.800 289.800 723.900 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 754.950 289.950 757.050 292.050 ;
        RECT 757.950 289.950 760.050 292.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 721.800 289.200 723.600 289.800 ;
        RECT 717.000 288.000 723.600 289.200 ;
        RECT 737.100 288.150 738.900 289.950 ;
        RECT 717.000 287.100 719.100 288.000 ;
        RECT 709.500 283.500 711.600 285.900 ;
        RECT 712.800 284.100 715.800 286.200 ;
        RECT 716.700 285.300 718.500 287.100 ;
        RECT 707.100 282.600 711.600 283.500 ;
        RECT 692.100 276.000 693.900 279.600 ;
        RECT 695.100 276.600 696.900 279.600 ;
        RECT 707.100 276.600 708.900 282.600 ;
        RECT 714.900 282.000 715.800 284.100 ;
        RECT 719.400 285.000 721.500 285.600 ;
        RECT 719.400 283.500 723.900 285.000 ;
        RECT 740.700 284.700 741.900 289.950 ;
        RECT 742.950 288.150 744.750 289.950 ;
        RECT 755.100 288.150 756.900 289.950 ;
        RECT 761.250 288.150 763.050 289.950 ;
        RECT 722.400 282.600 723.900 283.500 ;
        RECT 710.400 276.000 712.200 281.700 ;
        RECT 714.900 276.600 716.700 282.000 ;
        RECT 719.100 276.000 720.900 281.700 ;
        RECT 722.100 276.600 723.900 282.600 ;
        RECT 737.700 283.800 741.900 284.700 ;
        RECT 737.700 276.600 739.500 283.800 ;
        RECT 764.700 282.600 765.600 289.950 ;
        RECT 770.550 289.050 771.450 292.950 ;
        RECT 776.700 292.050 777.900 305.400 ;
        RECT 794.100 299.400 795.900 311.400 ;
        RECT 797.100 300.300 798.900 311.400 ;
        RECT 800.100 301.200 801.900 312.000 ;
        RECT 803.100 300.300 804.900 311.400 ;
        RECT 818.100 305.400 819.900 312.000 ;
        RECT 821.100 305.400 822.900 311.400 ;
        RECT 824.100 306.000 825.900 312.000 ;
        RECT 821.400 305.100 822.900 305.400 ;
        RECT 827.100 305.400 828.900 311.400 ;
        RECT 827.100 305.100 828.000 305.400 ;
        RECT 821.400 304.200 828.000 305.100 ;
        RECT 797.100 299.400 804.900 300.300 ;
        RECT 779.100 292.050 780.900 293.850 ;
        RECT 794.400 292.050 795.300 299.400 ;
        RECT 796.950 297.450 799.050 297.900 ;
        RECT 817.950 297.450 820.050 298.050 ;
        RECT 796.950 296.550 820.050 297.450 ;
        RECT 796.950 295.800 799.050 296.550 ;
        RECT 817.950 295.950 820.050 296.550 ;
        RECT 799.950 292.050 801.750 293.850 ;
        RECT 821.100 292.050 822.900 293.850 ;
        RECT 827.100 292.050 828.000 304.200 ;
        RECT 839.100 299.400 840.900 311.400 ;
        RECT 842.100 300.300 843.900 311.400 ;
        RECT 845.100 301.200 846.900 312.000 ;
        RECT 848.100 300.300 849.900 311.400 ;
        RECT 860.100 305.400 861.900 312.000 ;
        RECT 863.100 305.400 864.900 311.400 ;
        RECT 866.100 306.000 867.900 312.000 ;
        RECT 863.400 305.100 864.900 305.400 ;
        RECT 869.100 305.400 870.900 311.400 ;
        RECT 869.100 305.100 870.000 305.400 ;
        RECT 863.400 304.200 870.000 305.100 ;
        RECT 842.100 299.400 849.900 300.300 ;
        RECT 839.400 292.050 840.300 299.400 ;
        RECT 847.950 297.450 850.050 298.050 ;
        RECT 865.950 297.450 868.050 298.050 ;
        RECT 847.950 296.550 868.050 297.450 ;
        RECT 847.950 295.950 850.050 296.550 ;
        RECT 865.950 295.950 868.050 296.550 ;
        RECT 844.950 292.050 846.750 293.850 ;
        RECT 863.100 292.050 864.900 293.850 ;
        RECT 869.100 292.050 870.000 304.200 ;
        RECT 881.100 299.400 882.900 311.400 ;
        RECT 884.100 300.300 885.900 311.400 ;
        RECT 887.100 301.200 888.900 312.000 ;
        RECT 890.100 300.300 891.900 311.400 ;
        RECT 902.100 305.400 903.900 312.000 ;
        RECT 905.100 305.400 906.900 311.400 ;
        RECT 908.100 306.000 909.900 312.000 ;
        RECT 905.400 305.100 906.900 305.400 ;
        RECT 911.100 305.400 912.900 311.400 ;
        RECT 911.100 305.100 912.000 305.400 ;
        RECT 905.400 304.200 912.000 305.100 ;
        RECT 884.100 299.400 891.900 300.300 ;
        RECT 881.400 292.050 882.300 299.400 ;
        RECT 883.950 297.450 886.050 298.050 ;
        RECT 907.950 297.450 910.050 298.050 ;
        RECT 883.950 296.550 910.050 297.450 ;
        RECT 883.950 295.950 886.050 296.550 ;
        RECT 907.950 295.950 910.050 296.550 ;
        RECT 886.950 292.050 888.750 293.850 ;
        RECT 905.100 292.050 906.900 293.850 ;
        RECT 911.100 292.050 912.000 304.200 ;
        RECT 925.950 297.450 928.050 298.050 ;
        RECT 931.950 297.450 934.050 298.050 ;
        RECT 925.950 296.550 934.050 297.450 ;
        RECT 925.950 295.950 928.050 296.550 ;
        RECT 931.950 295.950 934.050 296.550 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 841.950 289.950 844.050 292.050 ;
        RECT 844.950 289.950 847.050 292.050 ;
        RECT 847.950 289.950 850.050 292.050 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 865.950 289.950 868.050 292.050 ;
        RECT 868.950 289.950 871.050 292.050 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 901.950 289.950 904.050 292.050 ;
        RECT 904.950 289.950 907.050 292.050 ;
        RECT 907.950 289.950 910.050 292.050 ;
        RECT 910.950 289.950 913.050 292.050 ;
        RECT 766.950 287.550 771.450 289.050 ;
        RECT 766.950 286.950 771.000 287.550 ;
        RECT 742.800 276.000 744.600 282.600 ;
        RECT 756.000 276.000 757.800 282.600 ;
        RECT 760.500 281.400 765.600 282.600 ;
        RECT 760.500 276.600 762.300 281.400 ;
        RECT 776.700 279.600 777.900 289.950 ;
        RECT 794.400 282.600 795.300 289.950 ;
        RECT 796.950 288.150 798.750 289.950 ;
        RECT 803.100 288.150 804.900 289.950 ;
        RECT 818.100 288.150 819.900 289.950 ;
        RECT 824.100 288.150 825.900 289.950 ;
        RECT 827.100 286.200 828.000 289.950 ;
        RECT 794.400 281.400 799.500 282.600 ;
        RECT 763.500 276.000 765.300 279.600 ;
        RECT 776.100 276.600 777.900 279.600 ;
        RECT 779.100 276.000 780.900 279.600 ;
        RECT 794.700 276.000 796.500 279.600 ;
        RECT 797.700 276.600 799.500 281.400 ;
        RECT 802.200 276.000 804.000 282.600 ;
        RECT 818.100 276.000 819.900 285.600 ;
        RECT 824.700 285.000 828.000 286.200 ;
        RECT 824.700 276.600 826.500 285.000 ;
        RECT 839.400 282.600 840.300 289.950 ;
        RECT 841.950 288.150 843.750 289.950 ;
        RECT 848.100 288.150 849.900 289.950 ;
        RECT 860.100 288.150 861.900 289.950 ;
        RECT 866.100 288.150 867.900 289.950 ;
        RECT 869.100 286.200 870.000 289.950 ;
        RECT 839.400 281.400 844.500 282.600 ;
        RECT 839.700 276.000 841.500 279.600 ;
        RECT 842.700 276.600 844.500 281.400 ;
        RECT 847.200 276.000 849.000 282.600 ;
        RECT 860.100 276.000 861.900 285.600 ;
        RECT 866.700 285.000 870.000 286.200 ;
        RECT 866.700 276.600 868.500 285.000 ;
        RECT 881.400 282.600 882.300 289.950 ;
        RECT 883.950 288.150 885.750 289.950 ;
        RECT 890.100 288.150 891.900 289.950 ;
        RECT 902.100 288.150 903.900 289.950 ;
        RECT 908.100 288.150 909.900 289.950 ;
        RECT 911.100 286.200 912.000 289.950 ;
        RECT 881.400 281.400 886.500 282.600 ;
        RECT 881.700 276.000 883.500 279.600 ;
        RECT 884.700 276.600 886.500 281.400 ;
        RECT 889.200 276.000 891.000 282.600 ;
        RECT 902.100 276.000 903.900 285.600 ;
        RECT 908.700 285.000 912.000 286.200 ;
        RECT 908.700 276.600 910.500 285.000 ;
        RECT 2.700 269.400 4.500 273.000 ;
        RECT 5.700 269.400 7.500 272.400 ;
        RECT 6.000 256.050 7.500 269.400 ;
        RECT 5.100 253.950 7.500 256.050 ;
        RECT 6.000 243.600 7.500 253.950 ;
        RECT 9.300 266.400 11.100 272.400 ;
        RECT 14.700 266.400 16.500 273.000 ;
        RECT 19.800 267.600 21.600 272.400 ;
        RECT 24.000 269.400 25.800 272.400 ;
        RECT 27.000 269.400 28.800 272.400 ;
        RECT 30.000 269.400 31.800 272.400 ;
        RECT 33.000 269.400 34.800 272.400 ;
        RECT 36.000 269.400 37.800 273.000 ;
        RECT 17.400 266.400 21.600 267.600 ;
        RECT 23.700 267.300 25.800 269.400 ;
        RECT 26.700 267.300 28.800 269.400 ;
        RECT 29.700 267.300 31.800 269.400 ;
        RECT 32.700 267.300 34.800 269.400 ;
        RECT 39.000 268.500 40.800 272.400 ;
        RECT 43.500 269.400 45.300 273.000 ;
        RECT 46.500 269.400 48.300 272.400 ;
        RECT 49.500 269.400 51.300 272.400 ;
        RECT 52.500 269.400 54.300 272.400 ;
        RECT 38.100 266.400 40.800 268.500 ;
        RECT 42.600 267.600 44.400 268.500 ;
        RECT 42.600 266.400 45.300 267.600 ;
        RECT 46.200 267.300 48.300 269.400 ;
        RECT 49.200 267.300 51.300 269.400 ;
        RECT 52.200 267.300 54.300 269.400 ;
        RECT 56.700 266.400 58.500 272.400 ;
        RECT 62.100 266.400 63.900 273.000 ;
        RECT 67.500 266.400 69.300 272.400 ;
        RECT 80.100 266.400 81.900 272.400 ;
        RECT 9.300 249.600 10.200 266.400 ;
        RECT 17.400 263.100 18.900 266.400 ;
        RECT 23.100 264.600 29.700 266.400 ;
        RECT 44.400 265.800 45.300 266.400 ;
        RECT 47.400 265.800 49.200 266.400 ;
        RECT 44.400 264.600 51.600 265.800 ;
        RECT 11.100 261.300 18.900 263.100 ;
        RECT 35.100 262.500 36.900 264.300 ;
        RECT 34.800 261.900 36.900 262.500 ;
        RECT 19.800 260.400 36.900 261.900 ;
        RECT 41.100 261.900 43.200 262.050 ;
        RECT 44.400 261.900 46.200 262.800 ;
        RECT 41.100 261.000 46.200 261.900 ;
        RECT 50.700 261.600 51.600 264.600 ;
        RECT 56.700 265.500 58.200 266.400 ;
        RECT 56.700 264.300 65.100 265.500 ;
        RECT 63.300 263.700 65.100 264.300 ;
        RECT 52.500 262.800 54.600 263.700 ;
        RECT 68.100 262.800 69.300 266.400 ;
        RECT 80.700 264.300 81.900 266.400 ;
        RECT 83.100 267.300 84.900 272.400 ;
        RECT 86.100 268.200 87.900 273.000 ;
        RECT 89.100 267.300 90.900 272.400 ;
        RECT 83.100 265.950 90.900 267.300 ;
        RECT 104.700 265.200 106.500 272.400 ;
        RECT 109.800 266.400 111.600 273.000 ;
        RECT 122.700 266.400 124.500 273.000 ;
        RECT 127.200 266.400 129.000 272.400 ;
        RECT 131.700 266.400 133.500 273.000 ;
        RECT 104.700 264.300 108.900 265.200 ;
        RECT 80.700 263.400 84.300 264.300 ;
        RECT 52.500 261.600 69.300 262.800 ;
        RECT 14.700 258.900 21.300 260.400 ;
        RECT 41.100 259.950 43.200 261.000 ;
        RECT 49.800 259.800 51.600 261.600 ;
        RECT 14.700 256.050 16.200 258.900 ;
        RECT 22.500 257.700 66.900 258.900 ;
        RECT 22.500 256.200 23.400 257.700 ;
        RECT 14.100 253.950 16.200 256.050 ;
        RECT 18.300 254.400 23.400 256.200 ;
        RECT 26.100 255.900 39.600 256.800 ;
        RECT 46.800 255.900 48.600 256.500 ;
        RECT 65.100 256.050 66.900 257.700 ;
        RECT 26.100 254.700 27.000 255.900 ;
        RECT 26.100 252.900 27.900 254.700 ;
        RECT 32.100 253.200 36.000 255.000 ;
        RECT 37.500 254.700 48.600 255.900 ;
        RECT 59.100 255.750 61.200 256.050 ;
        RECT 37.500 253.800 39.600 254.700 ;
        RECT 57.300 253.950 61.200 255.750 ;
        RECT 65.100 253.950 67.200 256.050 ;
        RECT 57.300 253.200 59.100 253.950 ;
        RECT 32.100 252.900 34.200 253.200 ;
        RECT 45.600 252.300 59.100 253.200 ;
        RECT 11.100 251.700 12.900 252.300 ;
        RECT 45.600 251.700 46.800 252.300 ;
        RECT 11.100 250.500 46.800 251.700 ;
        RECT 49.500 250.500 51.600 250.800 ;
        RECT 9.300 248.700 25.800 249.600 ;
        RECT 9.300 245.400 10.200 248.700 ;
        RECT 14.100 246.600 19.800 247.800 ;
        RECT 23.700 247.500 25.800 248.700 ;
        RECT 29.100 248.400 46.800 249.600 ;
        RECT 49.500 249.300 61.500 250.500 ;
        RECT 49.500 248.700 51.600 249.300 ;
        RECT 59.700 248.700 61.500 249.300 ;
        RECT 29.100 247.500 31.200 248.400 ;
        RECT 45.600 247.800 46.800 248.400 ;
        RECT 63.000 247.800 64.800 248.100 ;
        RECT 14.100 246.000 15.900 246.600 ;
        RECT 9.300 244.500 13.200 245.400 ;
        RECT 12.000 243.600 13.200 244.500 ;
        RECT 18.600 243.600 19.800 246.600 ;
        RECT 20.700 245.700 22.500 246.300 ;
        RECT 20.700 244.500 28.800 245.700 ;
        RECT 26.700 243.600 28.800 244.500 ;
        RECT 32.100 243.600 34.800 247.500 ;
        RECT 37.500 245.100 40.800 247.200 ;
        RECT 45.600 246.600 64.800 247.800 ;
        RECT 2.700 237.000 4.500 243.600 ;
        RECT 5.700 237.600 7.500 243.600 ;
        RECT 9.000 237.000 10.800 243.600 ;
        RECT 12.000 237.600 13.800 243.600 ;
        RECT 15.000 237.000 16.800 243.600 ;
        RECT 18.000 237.600 19.800 243.600 ;
        RECT 21.000 237.000 22.800 243.600 ;
        RECT 23.700 240.600 25.800 242.700 ;
        RECT 26.700 240.600 28.800 242.700 ;
        RECT 29.700 240.600 31.800 242.700 ;
        RECT 24.000 237.600 25.800 240.600 ;
        RECT 27.000 237.600 28.800 240.600 ;
        RECT 30.000 237.600 31.800 240.600 ;
        RECT 33.000 237.600 34.800 243.600 ;
        RECT 36.000 237.000 37.800 243.600 ;
        RECT 39.000 237.600 40.800 245.100 ;
        RECT 46.200 243.600 48.300 245.700 ;
        RECT 42.900 237.000 44.700 243.600 ;
        RECT 45.900 237.600 47.700 243.600 ;
        RECT 48.600 240.600 50.700 242.700 ;
        RECT 51.600 240.600 53.700 242.700 ;
        RECT 48.900 237.600 50.700 240.600 ;
        RECT 51.900 237.600 53.700 240.600 ;
        RECT 55.500 237.000 57.300 243.600 ;
        RECT 58.500 237.600 60.300 246.600 ;
        RECT 63.000 246.300 64.800 246.600 ;
        RECT 68.100 245.400 69.300 261.600 ;
        RECT 80.100 259.050 81.900 260.850 ;
        RECT 83.100 259.050 84.300 263.400 ;
        RECT 86.100 259.050 87.900 260.850 ;
        RECT 104.100 259.050 105.900 260.850 ;
        RECT 107.700 259.050 108.900 264.300 ;
        RECT 109.950 259.050 111.750 260.850 ;
        RECT 122.250 259.050 124.050 260.850 ;
        RECT 128.100 259.050 129.300 266.400 ;
        RECT 148.500 264.000 150.300 272.400 ;
        RECT 147.000 262.800 150.300 264.000 ;
        RECT 155.100 263.400 156.900 273.000 ;
        RECT 170.700 265.200 172.500 272.400 ;
        RECT 175.800 266.400 177.600 273.000 ;
        RECT 188.100 266.400 189.900 272.400 ;
        RECT 170.700 264.300 174.900 265.200 ;
        RECT 134.100 259.050 135.900 260.850 ;
        RECT 147.000 259.050 147.900 262.800 ;
        RECT 149.100 259.050 150.900 260.850 ;
        RECT 155.100 259.050 156.900 260.850 ;
        RECT 170.100 259.050 171.900 260.850 ;
        RECT 173.700 259.050 174.900 264.300 ;
        RECT 188.700 264.300 189.900 266.400 ;
        RECT 191.100 267.300 192.900 272.400 ;
        RECT 194.100 268.200 195.900 273.000 ;
        RECT 197.100 267.300 198.900 272.400 ;
        RECT 191.100 265.950 198.900 267.300 ;
        RECT 209.100 271.500 216.900 272.400 ;
        RECT 209.100 266.400 210.900 271.500 ;
        RECT 212.100 266.400 213.900 270.600 ;
        RECT 215.100 267.000 216.900 271.500 ;
        RECT 218.100 267.900 219.900 273.000 ;
        RECT 221.100 267.000 222.900 272.400 ;
        RECT 212.700 264.900 213.600 266.400 ;
        RECT 215.100 266.100 222.900 267.000 ;
        RECT 236.400 266.400 238.200 273.000 ;
        RECT 241.500 265.200 243.300 272.400 ;
        RECT 254.100 266.400 255.900 272.400 ;
        RECT 188.700 263.400 192.300 264.300 ;
        RECT 212.700 263.700 217.050 264.900 ;
        RECT 175.950 259.050 177.750 260.850 ;
        RECT 188.100 259.050 189.900 260.850 ;
        RECT 191.100 259.050 192.300 263.400 ;
        RECT 194.100 259.050 195.900 260.850 ;
        RECT 212.250 259.050 214.050 260.850 ;
        RECT 216.000 259.050 217.050 263.700 ;
        RECT 239.100 264.300 243.300 265.200 ;
        RECT 254.700 264.300 255.900 266.400 ;
        RECT 257.100 267.300 258.900 272.400 ;
        RECT 260.100 268.200 261.900 273.000 ;
        RECT 263.100 267.300 264.900 272.400 ;
        RECT 257.100 265.950 264.900 267.300 ;
        RECT 275.100 267.300 276.900 272.400 ;
        RECT 278.100 268.200 279.900 273.000 ;
        RECT 281.100 267.300 282.900 272.400 ;
        RECT 275.100 265.950 282.900 267.300 ;
        RECT 284.100 266.400 285.900 272.400 ;
        RECT 284.100 264.300 285.300 266.400 ;
        RECT 296.700 265.200 298.500 272.400 ;
        RECT 301.800 266.400 303.600 273.000 ;
        RECT 317.100 267.000 318.900 272.400 ;
        RECT 320.100 267.900 321.900 273.000 ;
        RECT 323.100 271.500 330.900 272.400 ;
        RECT 323.100 267.000 324.900 271.500 ;
        RECT 317.100 266.100 324.900 267.000 ;
        RECT 326.100 266.400 327.900 270.600 ;
        RECT 329.100 266.400 330.900 271.500 ;
        RECT 344.100 267.300 345.900 272.400 ;
        RECT 347.100 268.200 348.900 273.000 ;
        RECT 350.100 267.300 351.900 272.400 ;
        RECT 296.700 264.300 300.900 265.200 ;
        RECT 70.950 258.450 75.000 259.050 ;
        RECT 70.950 256.950 75.450 258.450 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 133.950 256.950 136.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 196.950 256.950 199.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 217.950 259.050 219.750 260.850 ;
        RECT 236.250 259.050 238.050 260.850 ;
        RECT 239.100 259.050 240.300 264.300 ;
        RECT 254.700 263.400 258.300 264.300 ;
        RECT 242.100 259.050 243.900 260.850 ;
        RECT 254.100 259.050 255.900 260.850 ;
        RECT 257.100 259.050 258.300 263.400 ;
        RECT 281.700 263.400 285.300 264.300 ;
        RECT 270.000 261.450 274.050 262.050 ;
        RECT 260.100 259.050 261.900 260.850 ;
        RECT 269.550 259.950 274.050 261.450 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 238.950 256.950 241.050 259.050 ;
        RECT 241.950 256.950 244.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 259.950 256.950 262.050 259.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 74.550 256.050 75.450 256.950 ;
        RECT 74.550 254.550 79.050 256.050 ;
        RECT 75.000 253.950 79.050 254.550 ;
        RECT 83.100 249.600 84.300 256.950 ;
        RECT 89.100 255.150 90.900 256.950 ;
        RECT 83.100 248.100 85.500 249.600 ;
        RECT 65.700 244.500 69.300 245.400 ;
        RECT 81.000 245.100 82.800 246.900 ;
        RECT 65.700 243.600 66.600 244.500 ;
        RECT 61.500 237.000 63.300 243.600 ;
        RECT 64.500 242.700 66.600 243.600 ;
        RECT 64.500 237.600 66.300 242.700 ;
        RECT 67.500 237.000 69.300 243.600 ;
        RECT 80.700 237.000 82.500 243.600 ;
        RECT 83.700 237.600 85.500 248.100 ;
        RECT 88.800 237.000 90.600 249.600 ;
        RECT 107.700 243.600 108.900 256.950 ;
        RECT 125.250 255.150 127.050 256.950 ;
        RECT 128.100 251.400 129.000 256.950 ;
        RECT 131.100 255.150 132.900 256.950 ;
        RECT 128.100 250.500 132.900 251.400 ;
        RECT 122.100 248.400 129.900 249.300 ;
        RECT 104.100 237.000 105.900 243.600 ;
        RECT 107.100 237.600 108.900 243.600 ;
        RECT 110.100 237.000 111.900 243.600 ;
        RECT 122.100 237.600 123.900 248.400 ;
        RECT 125.100 237.000 126.900 247.500 ;
        RECT 128.100 238.500 129.900 248.400 ;
        RECT 131.100 239.400 132.900 250.500 ;
        RECT 134.100 238.500 135.900 249.600 ;
        RECT 147.000 244.800 147.900 256.950 ;
        RECT 152.100 255.150 153.900 256.950 ;
        RECT 147.000 243.900 153.600 244.800 ;
        RECT 147.000 243.600 147.900 243.900 ;
        RECT 128.100 237.600 135.900 238.500 ;
        RECT 146.100 237.600 147.900 243.600 ;
        RECT 152.100 243.600 153.600 243.900 ;
        RECT 173.700 243.600 174.900 256.950 ;
        RECT 191.100 249.600 192.300 256.950 ;
        RECT 197.100 255.150 198.900 256.950 ;
        RECT 209.250 255.150 211.050 256.950 ;
        RECT 216.000 249.600 217.050 256.950 ;
        RECT 221.100 255.150 222.900 256.950 ;
        RECT 191.100 248.100 193.500 249.600 ;
        RECT 189.000 245.100 190.800 246.900 ;
        RECT 149.100 237.000 150.900 243.000 ;
        RECT 152.100 237.600 153.900 243.600 ;
        RECT 155.100 237.000 156.900 243.600 ;
        RECT 170.100 237.000 171.900 243.600 ;
        RECT 173.100 237.600 174.900 243.600 ;
        RECT 176.100 237.000 177.900 243.600 ;
        RECT 188.700 237.000 190.500 243.600 ;
        RECT 191.700 237.600 193.500 248.100 ;
        RECT 196.800 237.000 198.600 249.600 ;
        RECT 210.600 237.000 212.400 249.600 ;
        RECT 215.100 237.600 218.400 249.600 ;
        RECT 221.100 237.000 222.900 249.600 ;
        RECT 239.100 243.600 240.300 256.950 ;
        RECT 241.950 252.450 244.050 253.050 ;
        RECT 247.950 252.450 250.050 253.050 ;
        RECT 241.950 251.550 250.050 252.450 ;
        RECT 241.950 250.950 244.050 251.550 ;
        RECT 247.950 250.950 250.050 251.550 ;
        RECT 257.100 249.600 258.300 256.950 ;
        RECT 263.100 255.150 264.900 256.950 ;
        RECT 269.550 256.050 270.450 259.950 ;
        RECT 278.100 259.050 279.900 260.850 ;
        RECT 281.700 259.050 282.900 263.400 ;
        RECT 286.950 261.450 291.000 262.050 ;
        RECT 284.100 259.050 285.900 260.850 ;
        RECT 286.950 259.950 291.450 261.450 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 269.550 254.550 274.050 256.050 ;
        RECT 275.100 255.150 276.900 256.950 ;
        RECT 270.000 253.950 274.050 254.550 ;
        RECT 281.700 249.600 282.900 256.950 ;
        RECT 290.550 256.050 291.450 259.950 ;
        RECT 296.100 259.050 297.900 260.850 ;
        RECT 299.700 259.050 300.900 264.300 ;
        RECT 301.950 264.450 304.050 265.050 ;
        RECT 316.950 264.450 319.050 265.050 ;
        RECT 326.400 264.900 327.300 266.400 ;
        RECT 344.100 265.950 351.900 267.300 ;
        RECT 353.100 266.400 354.900 272.400 ;
        RECT 365.100 269.400 366.900 272.400 ;
        RECT 368.100 269.400 369.900 273.000 ;
        RECT 301.950 263.550 319.050 264.450 ;
        RECT 301.950 262.950 304.050 263.550 ;
        RECT 316.950 262.950 319.050 263.550 ;
        RECT 322.950 263.700 327.300 264.900 ;
        RECT 353.100 264.300 354.300 266.400 ;
        RECT 313.950 261.450 316.050 262.050 ;
        RECT 301.950 259.050 303.750 260.850 ;
        RECT 308.550 260.550 316.050 261.450 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 290.550 254.550 295.050 256.050 ;
        RECT 291.000 253.950 295.050 254.550 ;
        RECT 257.100 248.100 259.500 249.600 ;
        RECT 255.000 245.100 256.800 246.900 ;
        RECT 236.100 237.000 237.900 243.600 ;
        RECT 239.100 237.600 240.900 243.600 ;
        RECT 242.100 237.000 243.900 243.600 ;
        RECT 254.700 237.000 256.500 243.600 ;
        RECT 257.700 237.600 259.500 248.100 ;
        RECT 262.800 237.000 264.600 249.600 ;
        RECT 275.400 237.000 277.200 249.600 ;
        RECT 280.500 248.100 282.900 249.600 ;
        RECT 280.500 237.600 282.300 248.100 ;
        RECT 283.200 245.100 285.000 246.900 ;
        RECT 299.700 243.600 300.900 256.950 ;
        RECT 308.550 256.050 309.450 260.550 ;
        RECT 313.950 259.950 316.050 260.550 ;
        RECT 320.250 259.050 322.050 260.850 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 322.950 259.050 324.000 263.700 ;
        RECT 350.700 263.400 354.300 264.300 ;
        RECT 325.950 259.050 327.750 260.850 ;
        RECT 347.100 259.050 348.900 260.850 ;
        RECT 350.700 259.050 351.900 263.400 ;
        RECT 353.100 259.050 354.900 260.850 ;
        RECT 365.700 259.050 366.900 269.400 ;
        RECT 383.100 266.400 384.900 272.400 ;
        RECT 386.100 267.300 387.900 273.000 ;
        RECT 390.600 266.400 392.400 272.400 ;
        RECT 395.100 267.300 396.900 273.000 ;
        RECT 398.100 266.400 399.900 272.400 ;
        RECT 413.100 266.400 414.900 272.400 ;
        RECT 383.700 264.600 384.900 266.400 ;
        RECT 390.900 264.900 392.100 266.400 ;
        RECT 395.100 265.500 399.900 266.400 ;
        RECT 383.700 263.700 390.000 264.600 ;
        RECT 387.900 261.600 390.000 263.700 ;
        RECT 383.400 259.050 385.200 260.850 ;
        RECT 388.200 259.800 390.000 261.600 ;
        RECT 390.900 262.800 393.900 264.900 ;
        RECT 395.100 264.300 397.200 265.500 ;
        RECT 413.700 264.300 414.900 266.400 ;
        RECT 416.100 267.300 417.900 272.400 ;
        RECT 419.100 268.200 420.900 273.000 ;
        RECT 422.100 267.300 423.900 272.400 ;
        RECT 435.600 268.200 437.400 272.400 ;
        RECT 416.100 265.950 423.900 267.300 ;
        RECT 434.700 266.400 437.400 268.200 ;
        RECT 438.600 266.400 440.400 273.000 ;
        RECT 413.700 263.400 417.300 264.300 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 383.100 258.300 385.200 259.050 ;
        RECT 383.100 256.950 390.000 258.300 ;
        RECT 304.950 254.550 309.450 256.050 ;
        RECT 317.100 255.150 318.900 256.950 ;
        RECT 304.950 253.950 309.000 254.550 ;
        RECT 322.950 249.600 324.000 256.950 ;
        RECT 328.950 255.150 330.750 256.950 ;
        RECT 344.100 255.150 345.900 256.950 ;
        RECT 350.700 249.600 351.900 256.950 ;
        RECT 352.950 252.450 355.050 253.050 ;
        RECT 361.950 252.450 364.050 253.050 ;
        RECT 352.950 251.550 364.050 252.450 ;
        RECT 352.950 250.950 355.050 251.550 ;
        RECT 361.950 250.950 364.050 251.550 ;
        RECT 283.500 237.000 285.300 243.600 ;
        RECT 296.100 237.000 297.900 243.600 ;
        RECT 299.100 237.600 300.900 243.600 ;
        RECT 302.100 237.000 303.900 243.600 ;
        RECT 317.100 237.000 318.900 249.600 ;
        RECT 321.600 237.600 324.900 249.600 ;
        RECT 327.600 237.000 329.400 249.600 ;
        RECT 344.400 237.000 346.200 249.600 ;
        RECT 349.500 248.100 351.900 249.600 ;
        RECT 349.500 237.600 351.300 248.100 ;
        RECT 352.200 245.100 354.000 246.900 ;
        RECT 365.700 243.600 366.900 256.950 ;
        RECT 368.100 255.150 369.900 256.950 ;
        RECT 388.200 256.500 390.000 256.950 ;
        RECT 390.900 257.100 392.100 262.800 ;
        RECT 393.000 259.800 395.100 261.900 ;
        RECT 393.300 258.000 395.100 259.800 ;
        RECT 413.100 259.050 414.900 260.850 ;
        RECT 416.100 259.050 417.300 263.400 ;
        RECT 419.100 259.050 420.900 260.850 ;
        RECT 434.700 259.050 435.600 266.400 ;
        RECT 436.500 264.600 438.300 265.500 ;
        RECT 443.100 264.600 444.900 272.400 ;
        RECT 456.600 268.200 458.400 272.400 ;
        RECT 436.500 263.700 444.900 264.600 ;
        RECT 455.700 266.400 458.400 268.200 ;
        RECT 459.600 266.400 461.400 273.000 ;
        RECT 390.900 256.200 393.300 257.100 ;
        RECT 391.800 256.050 393.300 256.200 ;
        RECT 397.800 256.950 399.900 259.050 ;
        RECT 412.950 256.950 415.050 259.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 434.100 256.950 436.200 259.050 ;
        RECT 437.400 256.950 439.500 259.050 ;
        RECT 387.000 253.500 390.900 255.300 ;
        RECT 388.800 253.200 390.900 253.500 ;
        RECT 391.800 253.950 393.900 256.050 ;
        RECT 397.800 255.150 399.600 256.950 ;
        RECT 391.800 252.000 392.700 253.950 ;
        RECT 385.500 249.600 387.600 251.700 ;
        RECT 391.200 250.950 392.700 252.000 ;
        RECT 391.200 249.600 392.400 250.950 ;
        RECT 383.100 248.700 387.600 249.600 ;
        RECT 352.500 237.000 354.300 243.600 ;
        RECT 365.100 237.600 366.900 243.600 ;
        RECT 368.100 237.000 369.900 243.600 ;
        RECT 383.100 237.600 384.900 248.700 ;
        RECT 386.100 237.000 387.900 247.500 ;
        RECT 390.600 237.600 392.400 249.600 ;
        RECT 395.100 249.600 397.200 250.500 ;
        RECT 416.100 249.600 417.300 256.950 ;
        RECT 422.100 255.150 423.900 256.950 ;
        RECT 434.700 249.600 435.600 256.950 ;
        RECT 438.000 255.150 439.800 256.950 ;
        RECT 395.100 248.400 399.900 249.600 ;
        RECT 395.100 237.000 396.900 247.500 ;
        RECT 398.100 237.600 399.900 248.400 ;
        RECT 416.100 248.100 418.500 249.600 ;
        RECT 414.000 245.100 415.800 246.900 ;
        RECT 413.700 237.000 415.500 243.600 ;
        RECT 416.700 237.600 418.500 248.100 ;
        RECT 421.800 237.000 423.600 249.600 ;
        RECT 434.100 237.600 435.900 249.600 ;
        RECT 437.100 237.000 438.900 249.000 ;
        RECT 441.000 243.600 441.900 263.700 ;
        RECT 442.950 259.050 444.750 260.850 ;
        RECT 455.700 259.050 456.600 266.400 ;
        RECT 457.500 264.600 459.300 265.500 ;
        RECT 464.100 264.600 465.900 272.400 ;
        RECT 479.100 269.400 480.900 273.000 ;
        RECT 482.100 269.400 483.900 272.400 ;
        RECT 485.100 269.400 486.900 273.000 ;
        RECT 457.500 263.700 465.900 264.600 ;
        RECT 442.800 256.950 444.900 259.050 ;
        RECT 455.100 256.950 457.200 259.050 ;
        RECT 458.400 256.950 460.500 259.050 ;
        RECT 455.700 249.600 456.600 256.950 ;
        RECT 459.000 255.150 460.800 256.950 ;
        RECT 440.100 237.600 441.900 243.600 ;
        RECT 443.100 237.000 444.900 243.600 ;
        RECT 455.100 237.600 456.900 249.600 ;
        RECT 458.100 237.000 459.900 249.000 ;
        RECT 462.000 243.600 462.900 263.700 ;
        RECT 463.950 259.050 465.750 260.850 ;
        RECT 482.700 259.050 483.600 269.400 ;
        RECT 499.500 264.000 501.300 272.400 ;
        RECT 498.000 262.800 501.300 264.000 ;
        RECT 506.100 263.400 507.900 273.000 ;
        RECT 521.100 269.400 522.900 272.400 ;
        RECT 524.100 269.400 525.900 273.000 ;
        RECT 539.100 269.400 540.900 272.400 ;
        RECT 542.100 269.400 543.900 273.000 ;
        RECT 557.100 269.400 558.900 273.000 ;
        RECT 560.100 269.400 561.900 272.400 ;
        RECT 563.100 269.400 564.900 273.000 ;
        RECT 498.000 259.050 498.900 262.800 ;
        RECT 500.100 259.050 501.900 260.850 ;
        RECT 506.100 259.050 507.900 260.850 ;
        RECT 521.700 259.050 522.900 269.400 ;
        RECT 523.950 264.450 526.050 265.050 ;
        RECT 532.950 264.450 535.050 265.050 ;
        RECT 523.950 263.550 535.050 264.450 ;
        RECT 523.950 262.950 526.050 263.550 ;
        RECT 532.950 262.950 535.050 263.550 ;
        RECT 539.700 259.050 540.900 269.400 ;
        RECT 560.400 259.050 561.300 269.400 ;
        RECT 575.100 267.300 576.900 272.400 ;
        RECT 578.100 268.200 579.900 273.000 ;
        RECT 581.100 267.300 582.900 272.400 ;
        RECT 575.100 265.950 582.900 267.300 ;
        RECT 584.100 266.400 585.900 272.400 ;
        RECT 596.100 269.400 597.900 272.400 ;
        RECT 599.100 269.400 600.900 273.000 ;
        RECT 584.100 264.300 585.300 266.400 ;
        RECT 581.700 263.400 585.300 264.300 ;
        RECT 578.100 259.050 579.900 260.850 ;
        RECT 581.700 259.050 582.900 263.400 ;
        RECT 586.950 261.450 589.050 265.050 ;
        RECT 586.950 261.000 591.450 261.450 ;
        RECT 584.100 259.050 585.900 260.850 ;
        RECT 587.550 260.550 591.450 261.000 ;
        RECT 463.800 256.950 465.900 259.050 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 479.100 255.150 480.900 256.950 ;
        RECT 482.700 249.600 483.600 256.950 ;
        RECT 484.950 255.150 486.750 256.950 ;
        RECT 480.000 248.400 483.600 249.600 ;
        RECT 461.100 237.600 462.900 243.600 ;
        RECT 464.100 237.000 465.900 243.600 ;
        RECT 480.000 237.600 481.800 248.400 ;
        RECT 485.100 237.000 486.900 249.600 ;
        RECT 498.000 244.800 498.900 256.950 ;
        RECT 503.100 255.150 504.900 256.950 ;
        RECT 498.000 243.900 504.600 244.800 ;
        RECT 498.000 243.600 498.900 243.900 ;
        RECT 497.100 237.600 498.900 243.600 ;
        RECT 503.100 243.600 504.600 243.900 ;
        RECT 521.700 243.600 522.900 256.950 ;
        RECT 524.100 255.150 525.900 256.950 ;
        RECT 539.700 243.600 540.900 256.950 ;
        RECT 542.100 255.150 543.900 256.950 ;
        RECT 557.250 255.150 559.050 256.950 ;
        RECT 560.400 249.600 561.300 256.950 ;
        RECT 563.100 255.150 564.900 256.950 ;
        RECT 575.100 255.150 576.900 256.950 ;
        RECT 581.700 249.600 582.900 256.950 ;
        RECT 590.550 256.050 591.450 260.550 ;
        RECT 596.700 259.050 597.900 269.400 ;
        RECT 611.700 265.200 613.500 272.400 ;
        RECT 616.800 266.400 618.600 273.000 ;
        RECT 629.400 266.400 631.200 273.000 ;
        RECT 634.500 265.200 636.300 272.400 ;
        RECT 611.700 264.300 615.900 265.200 ;
        RECT 628.950 264.450 631.050 265.050 ;
        RECT 611.100 259.050 612.900 260.850 ;
        RECT 614.700 259.050 615.900 264.300 ;
        RECT 623.550 263.550 631.050 264.450 ;
        RECT 616.950 259.050 618.750 260.850 ;
        RECT 595.950 256.950 598.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 590.550 254.550 595.050 256.050 ;
        RECT 591.000 253.950 595.050 254.550 ;
        RECT 500.100 237.000 501.900 243.000 ;
        RECT 503.100 237.600 504.900 243.600 ;
        RECT 506.100 237.000 507.900 243.600 ;
        RECT 521.100 237.600 522.900 243.600 ;
        RECT 524.100 237.000 525.900 243.600 ;
        RECT 539.100 237.600 540.900 243.600 ;
        RECT 542.100 237.000 543.900 243.600 ;
        RECT 557.100 237.000 558.900 249.600 ;
        RECT 560.400 248.400 564.000 249.600 ;
        RECT 562.200 237.600 564.000 248.400 ;
        RECT 575.400 237.000 577.200 249.600 ;
        RECT 580.500 248.100 582.900 249.600 ;
        RECT 580.500 237.600 582.300 248.100 ;
        RECT 583.200 245.100 585.000 246.900 ;
        RECT 596.700 243.600 597.900 256.950 ;
        RECT 599.100 255.150 600.900 256.950 ;
        RECT 601.950 252.450 604.050 253.050 ;
        RECT 610.950 252.450 613.050 253.050 ;
        RECT 601.950 251.550 613.050 252.450 ;
        RECT 601.950 250.950 604.050 251.550 ;
        RECT 610.950 250.950 613.050 251.550 ;
        RECT 614.700 243.600 615.900 256.950 ;
        RECT 623.550 256.050 624.450 263.550 ;
        RECT 628.950 262.950 631.050 263.550 ;
        RECT 632.100 264.300 636.300 265.200 ;
        RECT 629.250 259.050 631.050 260.850 ;
        RECT 632.100 259.050 633.300 264.300 ;
        RECT 647.100 263.400 648.900 273.000 ;
        RECT 653.700 264.000 655.500 272.400 ;
        RECT 673.500 264.000 675.300 272.400 ;
        RECT 653.700 262.800 657.000 264.000 ;
        RECT 637.950 261.450 642.000 262.050 ;
        RECT 635.100 259.050 636.900 260.850 ;
        RECT 637.950 259.950 642.450 261.450 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 623.550 254.550 628.050 256.050 ;
        RECT 624.000 253.950 628.050 254.550 ;
        RECT 632.100 243.600 633.300 256.950 ;
        RECT 641.550 256.050 642.450 259.950 ;
        RECT 647.100 259.050 648.900 260.850 ;
        RECT 653.100 259.050 654.900 260.850 ;
        RECT 656.100 259.050 657.000 262.800 ;
        RECT 672.000 262.800 675.300 264.000 ;
        RECT 680.100 263.400 681.900 273.000 ;
        RECT 692.100 263.400 693.900 273.000 ;
        RECT 698.700 264.000 700.500 272.400 ;
        RECT 713.100 266.400 714.900 272.400 ;
        RECT 713.700 264.300 714.900 266.400 ;
        RECT 716.100 267.300 717.900 272.400 ;
        RECT 719.100 268.200 720.900 273.000 ;
        RECT 722.100 267.300 723.900 272.400 ;
        RECT 734.700 269.400 736.500 273.000 ;
        RECT 737.700 267.600 739.500 272.400 ;
        RECT 716.100 265.950 723.900 267.300 ;
        RECT 734.400 266.400 739.500 267.600 ;
        RECT 742.200 266.400 744.000 273.000 ;
        RECT 698.700 262.800 702.000 264.000 ;
        RECT 713.700 263.400 717.300 264.300 ;
        RECT 658.950 261.450 663.000 262.050 ;
        RECT 658.950 259.950 663.450 261.450 ;
        RECT 646.950 256.950 649.050 259.050 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 641.550 254.550 646.050 256.050 ;
        RECT 650.100 255.150 651.900 256.950 ;
        RECT 642.000 253.950 646.050 254.550 ;
        RECT 656.100 244.800 657.000 256.950 ;
        RECT 662.550 255.450 663.450 259.950 ;
        RECT 672.000 259.050 672.900 262.800 ;
        RECT 674.100 259.050 675.900 260.850 ;
        RECT 680.100 259.050 681.900 260.850 ;
        RECT 692.100 259.050 693.900 260.850 ;
        RECT 698.100 259.050 699.900 260.850 ;
        RECT 701.100 259.050 702.000 262.800 ;
        RECT 713.100 259.050 714.900 260.850 ;
        RECT 716.100 259.050 717.300 263.400 ;
        RECT 724.950 261.450 729.000 262.050 ;
        RECT 719.100 259.050 720.900 260.850 ;
        RECT 724.950 259.950 729.450 261.450 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 667.950 255.450 670.050 256.050 ;
        RECT 662.550 254.550 670.050 255.450 ;
        RECT 667.950 253.950 670.050 254.550 ;
        RECT 650.400 243.900 657.000 244.800 ;
        RECT 650.400 243.600 651.900 243.900 ;
        RECT 583.500 237.000 585.300 243.600 ;
        RECT 596.100 237.600 597.900 243.600 ;
        RECT 599.100 237.000 600.900 243.600 ;
        RECT 611.100 237.000 612.900 243.600 ;
        RECT 614.100 237.600 615.900 243.600 ;
        RECT 617.100 237.000 618.900 243.600 ;
        RECT 629.100 237.000 630.900 243.600 ;
        RECT 632.100 237.600 633.900 243.600 ;
        RECT 635.100 237.000 636.900 243.600 ;
        RECT 647.100 237.000 648.900 243.600 ;
        RECT 650.100 237.600 651.900 243.600 ;
        RECT 656.100 243.600 657.000 243.900 ;
        RECT 672.000 244.800 672.900 256.950 ;
        RECT 677.100 255.150 678.900 256.950 ;
        RECT 695.100 255.150 696.900 256.950 ;
        RECT 673.950 252.450 676.050 253.050 ;
        RECT 697.950 252.450 700.050 253.050 ;
        RECT 673.950 251.550 700.050 252.450 ;
        RECT 673.950 250.950 676.050 251.550 ;
        RECT 697.950 250.950 700.050 251.550 ;
        RECT 701.100 244.800 702.000 256.950 ;
        RECT 716.100 249.600 717.300 256.950 ;
        RECT 722.100 255.150 723.900 256.950 ;
        RECT 728.550 252.900 729.450 259.950 ;
        RECT 734.400 259.050 735.300 266.400 ;
        RECT 760.500 264.000 762.300 272.400 ;
        RECT 759.000 262.800 762.300 264.000 ;
        RECT 767.100 263.400 768.900 273.000 ;
        RECT 779.100 263.400 780.900 273.000 ;
        RECT 785.700 264.000 787.500 272.400 ;
        RECT 800.100 266.400 801.900 272.400 ;
        RECT 800.700 264.300 801.900 266.400 ;
        RECT 803.100 267.300 804.900 272.400 ;
        RECT 806.100 268.200 807.900 273.000 ;
        RECT 809.100 267.300 810.900 272.400 ;
        RECT 803.100 265.950 810.900 267.300 ;
        RECT 821.100 266.400 822.900 272.400 ;
        RECT 821.700 264.300 822.900 266.400 ;
        RECT 824.100 267.300 825.900 272.400 ;
        RECT 827.100 268.200 828.900 273.000 ;
        RECT 830.100 267.300 831.900 272.400 ;
        RECT 824.100 265.950 831.900 267.300 ;
        RECT 785.700 262.800 789.000 264.000 ;
        RECT 800.700 263.400 804.300 264.300 ;
        RECT 821.700 263.400 825.300 264.300 ;
        RECT 847.500 264.000 849.300 272.400 ;
        RECT 736.950 259.050 738.750 260.850 ;
        RECT 743.100 259.050 744.900 260.850 ;
        RECT 759.000 259.050 759.900 262.800 ;
        RECT 769.950 261.450 774.000 262.050 ;
        RECT 761.100 259.050 762.900 260.850 ;
        RECT 767.100 259.050 768.900 260.850 ;
        RECT 769.950 259.950 774.450 261.450 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 736.950 256.950 739.050 259.050 ;
        RECT 739.950 256.950 742.050 259.050 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 727.950 250.800 730.050 252.900 ;
        RECT 734.400 249.600 735.300 256.950 ;
        RECT 739.950 255.150 741.750 256.950 ;
        RECT 716.100 248.100 718.500 249.600 ;
        RECT 714.000 245.100 715.800 246.900 ;
        RECT 672.000 243.900 678.600 244.800 ;
        RECT 672.000 243.600 672.900 243.900 ;
        RECT 653.100 237.000 654.900 243.000 ;
        RECT 656.100 237.600 657.900 243.600 ;
        RECT 671.100 237.600 672.900 243.600 ;
        RECT 677.100 243.600 678.600 243.900 ;
        RECT 695.400 243.900 702.000 244.800 ;
        RECT 695.400 243.600 696.900 243.900 ;
        RECT 674.100 237.000 675.900 243.000 ;
        RECT 677.100 237.600 678.900 243.600 ;
        RECT 680.100 237.000 681.900 243.600 ;
        RECT 692.100 237.000 693.900 243.600 ;
        RECT 695.100 237.600 696.900 243.600 ;
        RECT 701.100 243.600 702.000 243.900 ;
        RECT 698.100 237.000 699.900 243.000 ;
        RECT 701.100 237.600 702.900 243.600 ;
        RECT 713.700 237.000 715.500 243.600 ;
        RECT 716.700 237.600 718.500 248.100 ;
        RECT 721.800 237.000 723.600 249.600 ;
        RECT 734.100 237.600 735.900 249.600 ;
        RECT 737.100 248.700 744.900 249.600 ;
        RECT 737.100 237.600 738.900 248.700 ;
        RECT 740.100 237.000 741.900 247.800 ;
        RECT 743.100 237.600 744.900 248.700 ;
        RECT 759.000 244.800 759.900 256.950 ;
        RECT 764.100 255.150 765.900 256.950 ;
        RECT 773.550 256.050 774.450 259.950 ;
        RECT 779.100 259.050 780.900 260.850 ;
        RECT 785.100 259.050 786.900 260.850 ;
        RECT 788.100 259.050 789.000 262.800 ;
        RECT 800.100 259.050 801.900 260.850 ;
        RECT 803.100 259.050 804.300 263.400 ;
        RECT 806.100 259.050 807.900 260.850 ;
        RECT 821.100 259.050 822.900 260.850 ;
        RECT 824.100 259.050 825.300 263.400 ;
        RECT 846.000 262.800 849.300 264.000 ;
        RECT 854.100 263.400 855.900 273.000 ;
        RECT 869.700 269.400 871.500 273.000 ;
        RECT 872.700 267.600 874.500 272.400 ;
        RECT 869.400 266.400 874.500 267.600 ;
        RECT 877.200 266.400 879.000 273.000 ;
        RECT 893.700 269.400 895.500 273.000 ;
        RECT 896.700 267.600 898.500 272.400 ;
        RECT 893.400 266.400 898.500 267.600 ;
        RECT 901.200 266.400 903.000 273.000 ;
        RECT 827.100 259.050 828.900 260.850 ;
        RECT 846.000 259.050 846.900 262.800 ;
        RECT 848.100 259.050 849.900 260.850 ;
        RECT 854.100 259.050 855.900 260.850 ;
        RECT 869.400 259.050 870.300 266.400 ;
        RECT 874.950 264.450 877.050 264.900 ;
        RECT 874.950 263.550 882.450 264.450 ;
        RECT 874.950 262.800 877.050 263.550 ;
        RECT 881.550 261.450 882.450 263.550 ;
        RECT 871.950 259.050 873.750 260.850 ;
        RECT 878.100 259.050 879.900 260.850 ;
        RECT 881.550 260.550 885.450 261.450 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 769.950 254.550 774.450 256.050 ;
        RECT 782.100 255.150 783.900 256.950 ;
        RECT 769.950 253.950 774.000 254.550 ;
        RECT 760.950 252.450 763.050 253.050 ;
        RECT 784.950 252.450 787.050 253.050 ;
        RECT 760.950 251.550 787.050 252.450 ;
        RECT 760.950 250.950 763.050 251.550 ;
        RECT 784.950 250.950 787.050 251.550 ;
        RECT 788.100 244.800 789.000 256.950 ;
        RECT 803.100 249.600 804.300 256.950 ;
        RECT 809.100 255.150 810.900 256.950 ;
        RECT 824.100 249.600 825.300 256.950 ;
        RECT 830.100 255.150 831.900 256.950 ;
        RECT 803.100 248.100 805.500 249.600 ;
        RECT 801.000 245.100 802.800 246.900 ;
        RECT 759.000 243.900 765.600 244.800 ;
        RECT 759.000 243.600 759.900 243.900 ;
        RECT 758.100 237.600 759.900 243.600 ;
        RECT 764.100 243.600 765.600 243.900 ;
        RECT 782.400 243.900 789.000 244.800 ;
        RECT 782.400 243.600 783.900 243.900 ;
        RECT 761.100 237.000 762.900 243.000 ;
        RECT 764.100 237.600 765.900 243.600 ;
        RECT 767.100 237.000 768.900 243.600 ;
        RECT 779.100 237.000 780.900 243.600 ;
        RECT 782.100 237.600 783.900 243.600 ;
        RECT 788.100 243.600 789.000 243.900 ;
        RECT 785.100 237.000 786.900 243.000 ;
        RECT 788.100 237.600 789.900 243.600 ;
        RECT 800.700 237.000 802.500 243.600 ;
        RECT 803.700 237.600 805.500 248.100 ;
        RECT 808.800 237.000 810.600 249.600 ;
        RECT 824.100 248.100 826.500 249.600 ;
        RECT 822.000 245.100 823.800 246.900 ;
        RECT 821.700 237.000 823.500 243.600 ;
        RECT 824.700 237.600 826.500 248.100 ;
        RECT 829.800 237.000 831.600 249.600 ;
        RECT 846.000 244.800 846.900 256.950 ;
        RECT 851.100 255.150 852.900 256.950 ;
        RECT 853.950 252.450 856.050 253.050 ;
        RECT 865.950 252.450 868.050 253.050 ;
        RECT 853.950 251.550 868.050 252.450 ;
        RECT 853.950 250.950 856.050 251.550 ;
        RECT 865.950 250.950 868.050 251.550 ;
        RECT 869.400 249.600 870.300 256.950 ;
        RECT 874.950 255.150 876.750 256.950 ;
        RECT 884.550 255.450 885.450 260.550 ;
        RECT 893.400 259.050 894.300 266.400 ;
        RECT 914.100 263.400 915.900 273.000 ;
        RECT 920.700 264.000 922.500 272.400 ;
        RECT 920.700 262.800 924.000 264.000 ;
        RECT 895.950 259.050 897.750 260.850 ;
        RECT 902.100 259.050 903.900 260.850 ;
        RECT 914.100 259.050 915.900 260.850 ;
        RECT 920.100 259.050 921.900 260.850 ;
        RECT 923.100 259.050 924.000 262.800 ;
        RECT 925.950 261.450 930.000 262.050 ;
        RECT 925.950 259.950 930.450 261.450 ;
        RECT 892.950 256.950 895.050 259.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 901.950 256.950 904.050 259.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 916.950 256.950 919.050 259.050 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 922.950 256.950 925.050 259.050 ;
        RECT 889.950 255.450 892.050 256.050 ;
        RECT 884.550 254.550 892.050 255.450 ;
        RECT 889.950 253.950 892.050 254.550 ;
        RECT 871.950 252.450 874.050 252.750 ;
        RECT 890.550 252.450 891.450 253.950 ;
        RECT 871.950 251.550 891.450 252.450 ;
        RECT 871.950 250.650 874.050 251.550 ;
        RECT 893.400 249.600 894.300 256.950 ;
        RECT 898.950 255.150 900.750 256.950 ;
        RECT 917.100 255.150 918.900 256.950 ;
        RECT 846.000 243.900 852.600 244.800 ;
        RECT 846.000 243.600 846.900 243.900 ;
        RECT 845.100 237.600 846.900 243.600 ;
        RECT 851.100 243.600 852.600 243.900 ;
        RECT 848.100 237.000 849.900 243.000 ;
        RECT 851.100 237.600 852.900 243.600 ;
        RECT 854.100 237.000 855.900 243.600 ;
        RECT 869.100 237.600 870.900 249.600 ;
        RECT 872.100 248.700 879.900 249.600 ;
        RECT 872.100 237.600 873.900 248.700 ;
        RECT 875.100 237.000 876.900 247.800 ;
        RECT 878.100 237.600 879.900 248.700 ;
        RECT 893.100 237.600 894.900 249.600 ;
        RECT 896.100 248.700 903.900 249.600 ;
        RECT 896.100 237.600 897.900 248.700 ;
        RECT 899.100 237.000 900.900 247.800 ;
        RECT 902.100 237.600 903.900 248.700 ;
        RECT 923.100 244.800 924.000 256.950 ;
        RECT 929.550 255.450 930.450 259.950 ;
        RECT 926.550 255.000 930.450 255.450 ;
        RECT 925.950 254.550 930.450 255.000 ;
        RECT 925.950 250.950 928.050 254.550 ;
        RECT 917.400 243.900 924.000 244.800 ;
        RECT 917.400 243.600 918.900 243.900 ;
        RECT 914.100 237.000 915.900 243.600 ;
        RECT 917.100 237.600 918.900 243.600 ;
        RECT 923.100 243.600 924.000 243.900 ;
        RECT 920.100 237.000 921.900 243.000 ;
        RECT 923.100 237.600 924.900 243.600 ;
        RECT 2.700 227.400 4.500 234.000 ;
        RECT 5.700 227.400 7.500 233.400 ;
        RECT 9.000 227.400 10.800 234.000 ;
        RECT 12.000 227.400 13.800 233.400 ;
        RECT 15.000 227.400 16.800 234.000 ;
        RECT 18.000 227.400 19.800 233.400 ;
        RECT 21.000 227.400 22.800 234.000 ;
        RECT 24.000 230.400 25.800 233.400 ;
        RECT 27.000 230.400 28.800 233.400 ;
        RECT 30.000 230.400 31.800 233.400 ;
        RECT 23.700 228.300 25.800 230.400 ;
        RECT 26.700 228.300 28.800 230.400 ;
        RECT 29.700 228.300 31.800 230.400 ;
        RECT 33.000 227.400 34.800 233.400 ;
        RECT 36.000 227.400 37.800 234.000 ;
        RECT 6.000 217.050 7.500 227.400 ;
        RECT 12.000 226.500 13.200 227.400 ;
        RECT 5.100 214.950 7.500 217.050 ;
        RECT 6.000 201.600 7.500 214.950 ;
        RECT 2.700 198.000 4.500 201.600 ;
        RECT 5.700 198.600 7.500 201.600 ;
        RECT 9.300 225.600 13.200 226.500 ;
        RECT 9.300 222.300 10.200 225.600 ;
        RECT 14.100 224.400 15.900 225.000 ;
        RECT 18.600 224.400 19.800 227.400 ;
        RECT 26.700 226.500 28.800 227.400 ;
        RECT 20.700 225.300 28.800 226.500 ;
        RECT 20.700 224.700 22.500 225.300 ;
        RECT 14.100 223.200 19.800 224.400 ;
        RECT 32.100 223.500 34.800 227.400 ;
        RECT 39.000 225.900 40.800 233.400 ;
        RECT 42.900 227.400 44.700 234.000 ;
        RECT 45.900 227.400 47.700 233.400 ;
        RECT 48.900 230.400 50.700 233.400 ;
        RECT 51.900 230.400 53.700 233.400 ;
        RECT 48.600 228.300 50.700 230.400 ;
        RECT 51.600 228.300 53.700 230.400 ;
        RECT 55.500 227.400 57.300 234.000 ;
        RECT 37.500 223.800 40.800 225.900 ;
        RECT 46.200 225.300 48.300 227.400 ;
        RECT 58.500 224.400 60.300 233.400 ;
        RECT 61.500 227.400 63.300 234.000 ;
        RECT 64.500 228.300 66.300 233.400 ;
        RECT 64.500 227.400 66.600 228.300 ;
        RECT 67.500 227.400 69.300 234.000 ;
        RECT 83.100 227.400 84.900 233.400 ;
        RECT 86.100 227.400 87.900 234.000 ;
        RECT 89.700 227.400 91.500 234.000 ;
        RECT 92.700 227.400 94.500 233.400 ;
        RECT 96.000 227.400 97.800 234.000 ;
        RECT 99.000 227.400 100.800 233.400 ;
        RECT 102.000 227.400 103.800 234.000 ;
        RECT 105.000 227.400 106.800 233.400 ;
        RECT 108.000 227.400 109.800 234.000 ;
        RECT 111.000 230.400 112.800 233.400 ;
        RECT 114.000 230.400 115.800 233.400 ;
        RECT 117.000 230.400 118.800 233.400 ;
        RECT 110.700 228.300 112.800 230.400 ;
        RECT 113.700 228.300 115.800 230.400 ;
        RECT 116.700 228.300 118.800 230.400 ;
        RECT 120.000 227.400 121.800 233.400 ;
        RECT 123.000 227.400 124.800 234.000 ;
        RECT 65.700 226.500 66.600 227.400 ;
        RECT 65.700 225.600 69.300 226.500 ;
        RECT 63.000 224.400 64.800 224.700 ;
        RECT 23.700 222.300 25.800 223.500 ;
        RECT 9.300 221.400 25.800 222.300 ;
        RECT 29.100 222.600 31.200 223.500 ;
        RECT 45.600 223.200 64.800 224.400 ;
        RECT 45.600 222.600 46.800 223.200 ;
        RECT 63.000 222.900 64.800 223.200 ;
        RECT 29.100 221.400 46.800 222.600 ;
        RECT 49.500 221.700 51.600 222.300 ;
        RECT 59.700 221.700 61.500 222.300 ;
        RECT 9.300 204.600 10.200 221.400 ;
        RECT 49.500 220.500 61.500 221.700 ;
        RECT 11.100 219.300 46.800 220.500 ;
        RECT 49.500 220.200 51.600 220.500 ;
        RECT 11.100 218.700 12.900 219.300 ;
        RECT 45.600 218.700 46.800 219.300 ;
        RECT 14.100 214.950 16.200 217.050 ;
        RECT 14.700 212.100 16.200 214.950 ;
        RECT 18.300 214.800 23.400 216.600 ;
        RECT 22.500 213.300 23.400 214.800 ;
        RECT 26.100 216.300 27.900 218.100 ;
        RECT 32.100 217.800 34.200 218.100 ;
        RECT 45.600 217.800 59.100 218.700 ;
        RECT 26.100 215.100 27.000 216.300 ;
        RECT 32.100 216.000 36.000 217.800 ;
        RECT 37.500 216.300 39.600 217.200 ;
        RECT 57.300 217.050 59.100 217.800 ;
        RECT 37.500 215.100 48.600 216.300 ;
        RECT 57.300 215.250 61.200 217.050 ;
        RECT 26.100 214.200 39.600 215.100 ;
        RECT 46.800 214.500 48.600 215.100 ;
        RECT 59.100 214.950 61.200 215.250 ;
        RECT 65.100 214.950 67.200 217.050 ;
        RECT 65.100 213.300 66.900 214.950 ;
        RECT 22.500 212.100 66.900 213.300 ;
        RECT 14.700 210.600 21.300 212.100 ;
        RECT 11.100 207.900 18.900 209.700 ;
        RECT 19.800 209.100 36.900 210.600 ;
        RECT 34.800 208.500 36.900 209.100 ;
        RECT 41.100 210.000 43.200 211.050 ;
        RECT 41.100 209.100 46.200 210.000 ;
        RECT 49.800 209.400 51.600 211.200 ;
        RECT 68.100 209.400 69.300 225.600 ;
        RECT 83.700 214.050 84.900 227.400 ;
        RECT 93.000 217.050 94.500 227.400 ;
        RECT 99.000 226.500 100.200 227.400 ;
        RECT 86.100 214.050 87.900 215.850 ;
        RECT 92.100 214.950 94.500 217.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 41.100 208.950 43.200 209.100 ;
        RECT 17.400 204.600 18.900 207.900 ;
        RECT 35.100 206.700 36.900 208.500 ;
        RECT 44.400 208.200 46.200 209.100 ;
        RECT 50.700 206.400 51.600 209.400 ;
        RECT 52.500 208.200 69.300 209.400 ;
        RECT 52.500 207.300 54.600 208.200 ;
        RECT 63.300 206.700 65.100 207.300 ;
        RECT 23.100 204.600 29.700 206.400 ;
        RECT 44.400 205.200 51.600 206.400 ;
        RECT 56.700 205.500 65.100 206.700 ;
        RECT 44.400 204.600 45.300 205.200 ;
        RECT 47.400 204.600 49.200 205.200 ;
        RECT 56.700 204.600 58.200 205.500 ;
        RECT 68.100 204.600 69.300 208.200 ;
        RECT 9.300 198.600 11.100 204.600 ;
        RECT 14.700 198.000 16.500 204.600 ;
        RECT 17.400 203.400 21.600 204.600 ;
        RECT 19.800 198.600 21.600 203.400 ;
        RECT 23.700 201.600 25.800 203.700 ;
        RECT 26.700 201.600 28.800 203.700 ;
        RECT 29.700 201.600 31.800 203.700 ;
        RECT 32.700 201.600 34.800 203.700 ;
        RECT 38.100 202.500 40.800 204.600 ;
        RECT 42.600 203.400 45.300 204.600 ;
        RECT 42.600 202.500 44.400 203.400 ;
        RECT 24.000 198.600 25.800 201.600 ;
        RECT 27.000 198.600 28.800 201.600 ;
        RECT 30.000 198.600 31.800 201.600 ;
        RECT 33.000 198.600 34.800 201.600 ;
        RECT 36.000 198.000 37.800 201.600 ;
        RECT 39.000 198.600 40.800 202.500 ;
        RECT 46.200 201.600 48.300 203.700 ;
        RECT 49.200 201.600 51.300 203.700 ;
        RECT 52.200 201.600 54.300 203.700 ;
        RECT 43.500 198.000 45.300 201.600 ;
        RECT 46.500 198.600 48.300 201.600 ;
        RECT 49.500 198.600 51.300 201.600 ;
        RECT 52.500 198.600 54.300 201.600 ;
        RECT 56.700 198.600 58.500 204.600 ;
        RECT 62.100 198.000 63.900 204.600 ;
        RECT 67.500 198.600 69.300 204.600 ;
        RECT 83.700 201.600 84.900 211.950 ;
        RECT 93.000 201.600 94.500 214.950 ;
        RECT 83.100 198.600 84.900 201.600 ;
        RECT 86.100 198.000 87.900 201.600 ;
        RECT 89.700 198.000 91.500 201.600 ;
        RECT 92.700 198.600 94.500 201.600 ;
        RECT 96.300 225.600 100.200 226.500 ;
        RECT 96.300 222.300 97.200 225.600 ;
        RECT 101.100 224.400 102.900 225.000 ;
        RECT 105.600 224.400 106.800 227.400 ;
        RECT 113.700 226.500 115.800 227.400 ;
        RECT 107.700 225.300 115.800 226.500 ;
        RECT 107.700 224.700 109.500 225.300 ;
        RECT 101.100 223.200 106.800 224.400 ;
        RECT 119.100 223.500 121.800 227.400 ;
        RECT 126.000 225.900 127.800 233.400 ;
        RECT 129.900 227.400 131.700 234.000 ;
        RECT 132.900 227.400 134.700 233.400 ;
        RECT 135.900 230.400 137.700 233.400 ;
        RECT 138.900 230.400 140.700 233.400 ;
        RECT 135.600 228.300 137.700 230.400 ;
        RECT 138.600 228.300 140.700 230.400 ;
        RECT 142.500 227.400 144.300 234.000 ;
        RECT 124.500 223.800 127.800 225.900 ;
        RECT 133.200 225.300 135.300 227.400 ;
        RECT 145.500 224.400 147.300 233.400 ;
        RECT 148.500 227.400 150.300 234.000 ;
        RECT 151.500 228.300 153.300 233.400 ;
        RECT 151.500 227.400 153.600 228.300 ;
        RECT 154.500 227.400 156.300 234.000 ;
        RECT 170.100 227.400 171.900 233.400 ;
        RECT 152.700 226.500 153.600 227.400 ;
        RECT 152.700 225.600 156.300 226.500 ;
        RECT 150.000 224.400 151.800 224.700 ;
        RECT 110.700 222.300 112.800 223.500 ;
        RECT 96.300 221.400 112.800 222.300 ;
        RECT 116.100 222.600 118.200 223.500 ;
        RECT 132.600 223.200 151.800 224.400 ;
        RECT 132.600 222.600 133.800 223.200 ;
        RECT 150.000 222.900 151.800 223.200 ;
        RECT 116.100 221.400 133.800 222.600 ;
        RECT 136.500 221.700 138.600 222.300 ;
        RECT 146.700 221.700 148.500 222.300 ;
        RECT 96.300 204.600 97.200 221.400 ;
        RECT 136.500 220.500 148.500 221.700 ;
        RECT 98.100 219.300 133.800 220.500 ;
        RECT 136.500 220.200 138.600 220.500 ;
        RECT 98.100 218.700 99.900 219.300 ;
        RECT 132.600 218.700 133.800 219.300 ;
        RECT 101.100 214.950 103.200 217.050 ;
        RECT 101.700 212.100 103.200 214.950 ;
        RECT 105.300 214.800 110.400 216.600 ;
        RECT 109.500 213.300 110.400 214.800 ;
        RECT 113.100 216.300 114.900 218.100 ;
        RECT 119.100 217.800 121.200 218.100 ;
        RECT 132.600 217.800 146.100 218.700 ;
        RECT 113.100 215.100 114.000 216.300 ;
        RECT 119.100 216.000 123.000 217.800 ;
        RECT 124.500 216.300 126.600 217.200 ;
        RECT 144.300 217.050 146.100 217.800 ;
        RECT 124.500 215.100 135.600 216.300 ;
        RECT 144.300 215.250 148.200 217.050 ;
        RECT 113.100 214.200 126.600 215.100 ;
        RECT 133.800 214.500 135.600 215.100 ;
        RECT 146.100 214.950 148.200 215.250 ;
        RECT 152.100 214.950 154.200 217.050 ;
        RECT 152.100 213.300 153.900 214.950 ;
        RECT 109.500 212.100 153.900 213.300 ;
        RECT 101.700 210.600 108.300 212.100 ;
        RECT 98.100 207.900 105.900 209.700 ;
        RECT 106.800 209.100 123.900 210.600 ;
        RECT 121.800 208.500 123.900 209.100 ;
        RECT 128.100 210.000 130.200 211.050 ;
        RECT 128.100 209.100 133.200 210.000 ;
        RECT 136.800 209.400 138.600 211.200 ;
        RECT 155.100 209.400 156.300 225.600 ;
        RECT 170.100 220.500 171.300 227.400 ;
        RECT 173.100 223.200 174.900 234.000 ;
        RECT 176.100 221.400 177.900 233.400 ;
        RECT 191.100 222.600 192.900 233.400 ;
        RECT 194.100 223.500 195.900 234.000 ;
        RECT 191.100 221.400 195.900 222.600 ;
        RECT 170.100 219.600 175.800 220.500 ;
        RECT 174.000 218.700 175.800 219.600 ;
        RECT 170.400 214.050 172.200 215.850 ;
        RECT 170.400 211.950 172.500 214.050 ;
        RECT 128.100 208.950 130.200 209.100 ;
        RECT 104.400 204.600 105.900 207.900 ;
        RECT 122.100 206.700 123.900 208.500 ;
        RECT 131.400 208.200 133.200 209.100 ;
        RECT 137.700 206.400 138.600 209.400 ;
        RECT 139.500 208.200 156.300 209.400 ;
        RECT 139.500 207.300 141.600 208.200 ;
        RECT 150.300 206.700 152.100 207.300 ;
        RECT 110.100 204.600 116.700 206.400 ;
        RECT 131.400 205.200 138.600 206.400 ;
        RECT 143.700 205.500 152.100 206.700 ;
        RECT 131.400 204.600 132.300 205.200 ;
        RECT 134.400 204.600 136.200 205.200 ;
        RECT 143.700 204.600 145.200 205.500 ;
        RECT 155.100 204.600 156.300 208.200 ;
        RECT 174.000 207.300 174.900 218.700 ;
        RECT 176.700 214.050 177.900 221.400 ;
        RECT 193.800 220.500 195.900 221.400 ;
        RECT 198.600 221.400 200.400 233.400 ;
        RECT 203.100 223.500 204.900 234.000 ;
        RECT 206.100 222.300 207.900 233.400 ;
        RECT 203.400 221.400 207.900 222.300 ;
        RECT 218.100 222.600 219.900 233.400 ;
        RECT 221.100 223.500 223.200 234.000 ;
        RECT 218.100 221.400 223.200 222.600 ;
        RECT 225.600 222.300 227.400 233.400 ;
        RECT 230.100 223.500 231.900 234.000 ;
        RECT 233.100 222.300 234.900 233.400 ;
        RECT 245.100 227.400 246.900 234.000 ;
        RECT 248.100 227.400 249.900 233.400 ;
        RECT 251.100 227.400 252.900 234.000 ;
        RECT 266.700 227.400 268.500 234.000 ;
        RECT 198.600 220.050 199.800 221.400 ;
        RECT 198.300 219.000 199.800 220.050 ;
        RECT 203.400 219.300 205.500 221.400 ;
        RECT 221.100 220.500 223.200 221.400 ;
        RECT 224.100 221.400 227.400 222.300 ;
        RECT 198.300 217.050 199.200 219.000 ;
        RECT 191.400 214.050 193.200 215.850 ;
        RECT 197.100 214.950 199.200 217.050 ;
        RECT 200.100 217.500 202.200 217.800 ;
        RECT 200.100 215.700 204.000 217.500 ;
        RECT 224.100 217.050 225.300 221.400 ;
        RECT 230.100 221.100 234.900 222.300 ;
        RECT 230.100 220.200 232.200 221.100 ;
        RECT 226.800 219.300 232.200 220.200 ;
        RECT 238.950 219.450 241.050 220.050 ;
        RECT 244.950 219.450 247.050 220.050 ;
        RECT 226.800 217.500 228.600 219.300 ;
        RECT 238.950 218.550 247.050 219.450 ;
        RECT 238.950 217.950 241.050 218.550 ;
        RECT 244.950 217.950 247.050 218.550 ;
        RECT 223.800 216.300 225.900 217.050 ;
        RECT 175.800 211.950 177.900 214.050 ;
        RECT 191.100 211.950 193.200 214.050 ;
        RECT 197.700 214.800 199.200 214.950 ;
        RECT 197.700 213.900 200.100 214.800 ;
        RECT 174.000 206.400 175.800 207.300 ;
        RECT 96.300 198.600 98.100 204.600 ;
        RECT 101.700 198.000 103.500 204.600 ;
        RECT 104.400 203.400 108.600 204.600 ;
        RECT 106.800 198.600 108.600 203.400 ;
        RECT 110.700 201.600 112.800 203.700 ;
        RECT 113.700 201.600 115.800 203.700 ;
        RECT 116.700 201.600 118.800 203.700 ;
        RECT 119.700 201.600 121.800 203.700 ;
        RECT 125.100 202.500 127.800 204.600 ;
        RECT 129.600 203.400 132.300 204.600 ;
        RECT 129.600 202.500 131.400 203.400 ;
        RECT 111.000 198.600 112.800 201.600 ;
        RECT 114.000 198.600 115.800 201.600 ;
        RECT 117.000 198.600 118.800 201.600 ;
        RECT 120.000 198.600 121.800 201.600 ;
        RECT 123.000 198.000 124.800 201.600 ;
        RECT 126.000 198.600 127.800 202.500 ;
        RECT 133.200 201.600 135.300 203.700 ;
        RECT 136.200 201.600 138.300 203.700 ;
        RECT 139.200 201.600 141.300 203.700 ;
        RECT 130.500 198.000 132.300 201.600 ;
        RECT 133.500 198.600 135.300 201.600 ;
        RECT 136.500 198.600 138.300 201.600 ;
        RECT 139.500 198.600 141.300 201.600 ;
        RECT 143.700 198.600 145.500 204.600 ;
        RECT 149.100 198.000 150.900 204.600 ;
        RECT 154.500 198.600 156.300 204.600 ;
        RECT 170.100 205.500 175.800 206.400 ;
        RECT 170.100 201.600 171.300 205.500 ;
        RECT 176.700 204.600 177.900 211.950 ;
        RECT 195.900 211.200 197.700 213.000 ;
        RECT 195.900 209.100 198.000 211.200 ;
        RECT 198.900 208.200 200.100 213.900 ;
        RECT 201.000 214.050 202.800 214.500 ;
        RECT 218.400 214.050 220.200 215.850 ;
        RECT 223.800 214.950 226.800 216.300 ;
        RECT 201.000 212.700 207.900 214.050 ;
        RECT 205.800 211.950 207.900 212.700 ;
        RECT 218.100 211.950 220.200 214.050 ;
        RECT 223.200 212.100 225.000 213.900 ;
        RECT 193.800 205.500 195.900 206.700 ;
        RECT 197.100 206.100 200.100 208.200 ;
        RECT 201.000 209.400 202.800 211.200 ;
        RECT 205.800 210.150 207.600 211.950 ;
        RECT 222.900 210.000 225.000 212.100 ;
        RECT 201.000 207.300 203.100 209.400 ;
        RECT 225.900 208.200 226.800 214.950 ;
        RECT 228.300 214.200 230.100 216.000 ;
        RECT 228.000 212.100 230.100 214.200 ;
        RECT 248.100 214.050 249.300 227.400 ;
        RECT 267.000 224.100 268.800 225.900 ;
        RECT 269.700 222.900 271.500 233.400 ;
        RECT 269.100 221.400 271.500 222.900 ;
        RECT 274.800 221.400 276.600 234.000 ;
        RECT 287.100 221.400 288.900 233.400 ;
        RECT 290.100 222.000 291.900 234.000 ;
        RECT 293.100 227.400 294.900 233.400 ;
        RECT 296.100 227.400 297.900 234.000 ;
        RECT 311.700 227.400 313.500 234.000 ;
        RECT 269.100 214.050 270.300 221.400 ;
        RECT 271.950 219.450 274.050 219.900 ;
        RECT 283.950 219.450 286.050 220.050 ;
        RECT 271.950 218.550 286.050 219.450 ;
        RECT 271.950 217.800 274.050 218.550 ;
        RECT 283.950 217.950 286.050 218.550 ;
        RECT 275.100 214.050 276.900 215.850 ;
        RECT 287.700 214.050 288.600 221.400 ;
        RECT 291.000 214.050 292.800 215.850 ;
        RECT 232.800 211.800 234.900 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 287.100 211.950 289.200 214.050 ;
        RECT 290.400 211.950 292.500 214.050 ;
        RECT 232.800 211.200 234.600 211.800 ;
        RECT 228.000 210.000 234.600 211.200 ;
        RECT 245.250 210.150 247.050 211.950 ;
        RECT 228.000 209.100 230.100 210.000 ;
        RECT 201.000 206.400 207.300 207.300 ;
        RECT 170.100 198.600 171.900 201.600 ;
        RECT 173.100 198.000 174.900 204.600 ;
        RECT 176.100 198.600 177.900 204.600 ;
        RECT 191.100 204.600 195.900 205.500 ;
        RECT 198.900 204.600 200.100 206.100 ;
        RECT 206.100 204.600 207.300 206.400 ;
        RECT 220.500 205.500 222.600 207.900 ;
        RECT 223.800 206.100 226.800 208.200 ;
        RECT 227.700 207.300 229.500 209.100 ;
        RECT 218.100 204.600 222.600 205.500 ;
        RECT 191.100 198.600 192.900 204.600 ;
        RECT 194.100 198.000 195.900 203.700 ;
        RECT 198.600 198.600 200.400 204.600 ;
        RECT 203.100 198.000 204.900 203.700 ;
        RECT 206.100 198.600 207.900 204.600 ;
        RECT 218.100 198.600 219.900 204.600 ;
        RECT 225.900 204.000 226.800 206.100 ;
        RECT 230.400 207.000 232.500 207.600 ;
        RECT 230.400 205.500 234.900 207.000 ;
        RECT 248.100 206.700 249.300 211.950 ;
        RECT 251.100 210.150 252.900 211.950 ;
        RECT 266.100 210.150 267.900 211.950 ;
        RECT 269.100 207.600 270.300 211.950 ;
        RECT 272.100 210.150 273.900 211.950 ;
        RECT 266.700 206.700 270.300 207.600 ;
        RECT 248.100 205.800 252.300 206.700 ;
        RECT 233.400 204.600 234.900 205.500 ;
        RECT 221.400 198.000 223.200 203.700 ;
        RECT 225.900 198.600 227.700 204.000 ;
        RECT 230.100 198.000 231.900 203.700 ;
        RECT 233.100 198.600 234.900 204.600 ;
        RECT 245.400 198.000 247.200 204.600 ;
        RECT 250.500 198.600 252.300 205.800 ;
        RECT 266.700 204.600 267.900 206.700 ;
        RECT 266.100 198.600 267.900 204.600 ;
        RECT 269.100 203.700 276.900 205.050 ;
        RECT 269.100 198.600 270.900 203.700 ;
        RECT 272.100 198.000 273.900 202.800 ;
        RECT 275.100 198.600 276.900 203.700 ;
        RECT 287.700 204.600 288.600 211.950 ;
        RECT 294.000 207.300 294.900 227.400 ;
        RECT 312.000 224.100 313.800 225.900 ;
        RECT 314.700 222.900 316.500 233.400 ;
        RECT 314.100 221.400 316.500 222.900 ;
        RECT 319.800 221.400 321.600 234.000 ;
        RECT 332.100 227.400 333.900 233.400 ;
        RECT 335.100 228.000 336.900 234.000 ;
        RECT 333.000 227.100 333.900 227.400 ;
        RECT 338.100 227.400 339.900 233.400 ;
        RECT 341.100 227.400 342.900 234.000 ;
        RECT 356.700 227.400 358.500 234.000 ;
        RECT 338.100 227.100 339.600 227.400 ;
        RECT 333.000 226.200 339.600 227.100 ;
        RECT 314.100 214.050 315.300 221.400 ;
        RECT 320.100 214.050 321.900 215.850 ;
        RECT 333.000 214.050 333.900 226.200 ;
        RECT 357.000 224.100 358.800 225.900 ;
        RECT 359.700 222.900 361.500 233.400 ;
        RECT 359.100 221.400 361.500 222.900 ;
        RECT 364.800 221.400 366.600 234.000 ;
        RECT 378.000 222.600 379.800 233.400 ;
        RECT 378.000 221.400 381.600 222.600 ;
        RECT 383.100 221.400 384.900 234.000 ;
        RECT 395.100 221.400 396.900 233.400 ;
        RECT 398.100 222.300 399.900 233.400 ;
        RECT 401.100 223.200 402.900 234.000 ;
        RECT 404.100 222.300 405.900 233.400 ;
        RECT 416.100 227.400 417.900 233.400 ;
        RECT 419.100 228.000 420.900 234.000 ;
        RECT 398.100 221.400 405.900 222.300 ;
        RECT 417.000 227.100 417.900 227.400 ;
        RECT 422.100 227.400 423.900 233.400 ;
        RECT 425.100 227.400 426.900 234.000 ;
        RECT 422.100 227.100 423.600 227.400 ;
        RECT 417.000 226.200 423.600 227.100 ;
        RECT 338.100 214.050 339.900 215.850 ;
        RECT 359.100 214.050 360.300 221.400 ;
        RECT 365.100 214.050 366.900 215.850 ;
        RECT 377.100 214.050 378.900 215.850 ;
        RECT 380.700 214.050 381.600 221.400 ;
        RECT 382.950 214.050 384.750 215.850 ;
        RECT 395.400 214.050 396.300 221.400 ;
        RECT 400.950 214.050 402.750 215.850 ;
        RECT 417.000 214.050 417.900 226.200 ;
        RECT 437.400 221.400 439.200 234.000 ;
        RECT 442.500 222.900 444.300 233.400 ;
        RECT 445.500 227.400 447.300 234.000 ;
        RECT 458.100 227.400 459.900 233.400 ;
        RECT 461.100 227.400 462.900 234.000 ;
        RECT 445.200 224.100 447.000 225.900 ;
        RECT 442.500 221.400 444.900 222.900 ;
        RECT 422.100 214.050 423.900 215.850 ;
        RECT 437.100 214.050 438.900 215.850 ;
        RECT 443.700 214.050 444.900 221.400 ;
        RECT 453.000 216.450 457.050 217.050 ;
        RECT 452.550 214.950 457.050 216.450 ;
        RECT 295.800 211.950 297.900 214.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 400.950 211.950 403.050 214.050 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 436.950 211.950 439.050 214.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 295.950 210.150 297.750 211.950 ;
        RECT 311.100 210.150 312.900 211.950 ;
        RECT 314.100 207.600 315.300 211.950 ;
        RECT 317.100 210.150 318.900 211.950 ;
        RECT 289.500 206.400 297.900 207.300 ;
        RECT 289.500 205.500 291.300 206.400 ;
        RECT 287.700 202.800 290.400 204.600 ;
        RECT 288.600 198.600 290.400 202.800 ;
        RECT 291.600 198.000 293.400 204.600 ;
        RECT 296.100 198.600 297.900 206.400 ;
        RECT 311.700 206.700 315.300 207.600 ;
        RECT 333.000 208.200 333.900 211.950 ;
        RECT 335.100 210.150 336.900 211.950 ;
        RECT 341.100 210.150 342.900 211.950 ;
        RECT 356.100 210.150 357.900 211.950 ;
        RECT 333.000 207.000 336.300 208.200 ;
        RECT 359.100 207.600 360.300 211.950 ;
        RECT 362.100 210.150 363.900 211.950 ;
        RECT 311.700 204.600 312.900 206.700 ;
        RECT 311.100 198.600 312.900 204.600 ;
        RECT 314.100 203.700 321.900 205.050 ;
        RECT 314.100 198.600 315.900 203.700 ;
        RECT 317.100 198.000 318.900 202.800 ;
        RECT 320.100 198.600 321.900 203.700 ;
        RECT 334.500 198.600 336.300 207.000 ;
        RECT 341.100 198.000 342.900 207.600 ;
        RECT 356.700 206.700 360.300 207.600 ;
        RECT 356.700 204.600 357.900 206.700 ;
        RECT 356.100 198.600 357.900 204.600 ;
        RECT 359.100 203.700 366.900 205.050 ;
        RECT 359.100 198.600 360.900 203.700 ;
        RECT 362.100 198.000 363.900 202.800 ;
        RECT 365.100 198.600 366.900 203.700 ;
        RECT 380.700 201.600 381.600 211.950 ;
        RECT 395.400 204.600 396.300 211.950 ;
        RECT 397.950 210.150 399.750 211.950 ;
        RECT 404.100 210.150 405.900 211.950 ;
        RECT 417.000 208.200 417.900 211.950 ;
        RECT 419.100 210.150 420.900 211.950 ;
        RECT 425.100 210.150 426.900 211.950 ;
        RECT 440.100 210.150 441.900 211.950 ;
        RECT 417.000 207.000 420.300 208.200 ;
        RECT 443.700 207.600 444.900 211.950 ;
        RECT 446.100 210.150 447.900 211.950 ;
        RECT 452.550 211.050 453.450 214.950 ;
        RECT 458.700 214.050 459.900 227.400 ;
        RECT 476.400 221.400 478.200 234.000 ;
        RECT 481.500 222.900 483.300 233.400 ;
        RECT 484.500 227.400 486.300 234.000 ;
        RECT 484.200 224.100 486.000 225.900 ;
        RECT 481.500 221.400 483.900 222.900 ;
        RECT 500.100 221.400 501.900 234.000 ;
        RECT 505.200 222.600 507.000 233.400 ;
        RECT 503.400 221.400 507.000 222.600 ;
        RECT 519.000 222.600 520.800 233.400 ;
        RECT 519.000 221.400 522.600 222.600 ;
        RECT 524.100 221.400 525.900 234.000 ;
        RECT 536.700 227.400 538.500 234.000 ;
        RECT 537.000 224.100 538.800 225.900 ;
        RECT 539.700 222.900 541.500 233.400 ;
        RECT 539.100 221.400 541.500 222.900 ;
        RECT 544.800 221.400 546.600 234.000 ;
        RECT 557.100 227.400 558.900 234.000 ;
        RECT 560.100 227.400 561.900 233.400 ;
        RECT 563.100 227.400 564.900 234.000 ;
        RECT 578.100 227.400 579.900 234.000 ;
        RECT 581.100 227.400 582.900 233.400 ;
        RECT 584.100 227.400 585.900 234.000 ;
        RECT 472.950 216.450 475.050 220.050 ;
        RECT 470.550 216.000 475.050 216.450 ;
        RECT 461.100 214.050 462.900 215.850 ;
        RECT 470.550 215.550 474.450 216.000 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 452.550 209.550 457.050 211.050 ;
        RECT 453.000 208.950 457.050 209.550 ;
        RECT 395.400 203.400 400.500 204.600 ;
        RECT 377.100 198.000 378.900 201.600 ;
        RECT 380.100 198.600 381.900 201.600 ;
        RECT 383.100 198.000 384.900 201.600 ;
        RECT 395.700 198.000 397.500 201.600 ;
        RECT 398.700 198.600 400.500 203.400 ;
        RECT 403.200 198.000 405.000 204.600 ;
        RECT 418.500 198.600 420.300 207.000 ;
        RECT 425.100 198.000 426.900 207.600 ;
        RECT 443.700 206.700 447.300 207.600 ;
        RECT 437.100 203.700 444.900 205.050 ;
        RECT 437.100 198.600 438.900 203.700 ;
        RECT 440.100 198.000 441.900 202.800 ;
        RECT 443.100 198.600 444.900 203.700 ;
        RECT 446.100 204.600 447.300 206.700 ;
        RECT 446.100 198.600 447.900 204.600 ;
        RECT 458.700 201.600 459.900 211.950 ;
        RECT 470.550 211.050 471.450 215.550 ;
        RECT 476.100 214.050 477.900 215.850 ;
        RECT 482.700 214.050 483.900 221.400 ;
        RECT 500.250 214.050 502.050 215.850 ;
        RECT 503.400 214.050 504.300 221.400 ;
        RECT 513.000 216.450 517.050 217.050 ;
        RECT 506.100 214.050 507.900 215.850 ;
        RECT 512.550 214.950 517.050 216.450 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 481.950 211.950 484.050 214.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 505.950 211.950 508.050 214.050 ;
        RECT 470.550 209.550 475.050 211.050 ;
        RECT 479.100 210.150 480.900 211.950 ;
        RECT 471.000 208.950 475.050 209.550 ;
        RECT 482.700 207.600 483.900 211.950 ;
        RECT 485.100 210.150 486.900 211.950 ;
        RECT 482.700 206.700 486.300 207.600 ;
        RECT 476.100 203.700 483.900 205.050 ;
        RECT 458.100 198.600 459.900 201.600 ;
        RECT 461.100 198.000 462.900 201.600 ;
        RECT 476.100 198.600 477.900 203.700 ;
        RECT 479.100 198.000 480.900 202.800 ;
        RECT 482.100 198.600 483.900 203.700 ;
        RECT 485.100 204.600 486.300 206.700 ;
        RECT 485.100 198.600 486.900 204.600 ;
        RECT 487.950 201.450 490.050 202.050 ;
        RECT 496.950 201.450 499.050 202.050 ;
        RECT 503.400 201.600 504.300 211.950 ;
        RECT 512.550 211.050 513.450 214.950 ;
        RECT 518.100 214.050 519.900 215.850 ;
        RECT 521.700 214.050 522.600 221.400 ;
        RECT 531.000 216.450 535.050 217.050 ;
        RECT 523.950 214.050 525.750 215.850 ;
        RECT 530.550 214.950 535.050 216.450 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 523.950 211.950 526.050 214.050 ;
        RECT 508.950 209.550 513.450 211.050 ;
        RECT 508.950 208.950 513.000 209.550 ;
        RECT 521.700 201.600 522.600 211.950 ;
        RECT 530.550 211.050 531.450 214.950 ;
        RECT 539.100 214.050 540.300 221.400 ;
        RECT 545.100 214.050 546.900 215.850 ;
        RECT 560.100 214.050 561.300 227.400 ;
        RECT 581.700 214.050 582.900 227.400 ;
        RECT 600.000 222.600 601.800 233.400 ;
        RECT 600.000 221.400 603.600 222.600 ;
        RECT 605.100 221.400 606.900 234.000 ;
        RECT 620.100 227.400 621.900 234.000 ;
        RECT 623.100 227.400 624.900 233.400 ;
        RECT 626.100 227.400 627.900 234.000 ;
        RECT 589.950 219.450 592.050 220.050 ;
        RECT 598.950 219.450 601.050 220.050 ;
        RECT 589.950 218.550 601.050 219.450 ;
        RECT 589.950 217.950 592.050 218.550 ;
        RECT 598.950 217.950 601.050 218.550 ;
        RECT 599.100 214.050 600.900 215.850 ;
        RECT 602.700 214.050 603.600 221.400 ;
        RECT 604.950 214.050 606.750 215.850 ;
        RECT 623.100 214.050 624.300 227.400 ;
        RECT 639.600 222.900 641.400 233.400 ;
        RECT 639.000 221.400 641.400 222.900 ;
        RECT 642.600 221.400 644.400 234.000 ;
        RECT 647.100 221.400 648.900 233.400 ;
        RECT 662.100 227.400 663.900 234.000 ;
        RECT 665.100 227.400 666.900 233.400 ;
        RECT 668.100 227.400 669.900 234.000 ;
        RECT 639.000 214.050 640.200 221.400 ;
        RECT 647.700 219.900 648.900 221.400 ;
        RECT 641.100 218.700 648.900 219.900 ;
        RECT 641.100 218.100 642.900 218.700 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 556.950 211.950 559.050 214.050 ;
        RECT 559.950 211.950 562.050 214.050 ;
        RECT 562.950 211.950 565.050 214.050 ;
        RECT 577.950 211.950 580.050 214.050 ;
        RECT 580.950 211.950 583.050 214.050 ;
        RECT 583.950 211.950 586.050 214.050 ;
        RECT 598.950 211.950 601.050 214.050 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 619.950 211.950 622.050 214.050 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 625.950 211.950 628.050 214.050 ;
        RECT 638.100 211.950 640.200 214.050 ;
        RECT 530.550 209.550 535.050 211.050 ;
        RECT 536.100 210.150 537.900 211.950 ;
        RECT 531.000 208.950 535.050 209.550 ;
        RECT 539.100 207.600 540.300 211.950 ;
        RECT 542.100 210.150 543.900 211.950 ;
        RECT 557.250 210.150 559.050 211.950 ;
        RECT 536.700 206.700 540.300 207.600 ;
        RECT 560.100 206.700 561.300 211.950 ;
        RECT 563.100 210.150 564.900 211.950 ;
        RECT 578.100 210.150 579.900 211.950 ;
        RECT 581.700 206.700 582.900 211.950 ;
        RECT 583.950 210.150 585.750 211.950 ;
        RECT 536.700 204.600 537.900 206.700 ;
        RECT 560.100 205.800 564.300 206.700 ;
        RECT 487.950 200.550 499.050 201.450 ;
        RECT 487.950 199.950 490.050 200.550 ;
        RECT 496.950 199.950 499.050 200.550 ;
        RECT 500.100 198.000 501.900 201.600 ;
        RECT 503.100 198.600 504.900 201.600 ;
        RECT 506.100 198.000 507.900 201.600 ;
        RECT 518.100 198.000 519.900 201.600 ;
        RECT 521.100 198.600 522.900 201.600 ;
        RECT 524.100 198.000 525.900 201.600 ;
        RECT 536.100 198.600 537.900 204.600 ;
        RECT 539.100 203.700 546.900 205.050 ;
        RECT 539.100 198.600 540.900 203.700 ;
        RECT 542.100 198.000 543.900 202.800 ;
        RECT 545.100 198.600 546.900 203.700 ;
        RECT 557.400 198.000 559.200 204.600 ;
        RECT 562.500 198.600 564.300 205.800 ;
        RECT 578.700 205.800 582.900 206.700 ;
        RECT 565.950 201.450 568.050 202.050 ;
        RECT 571.950 201.450 574.050 202.050 ;
        RECT 565.950 200.550 574.050 201.450 ;
        RECT 565.950 199.950 568.050 200.550 ;
        RECT 571.950 199.950 574.050 200.550 ;
        RECT 578.700 198.600 580.500 205.800 ;
        RECT 583.800 198.000 585.600 204.600 ;
        RECT 602.700 201.600 603.600 211.950 ;
        RECT 620.250 210.150 622.050 211.950 ;
        RECT 623.100 206.700 624.300 211.950 ;
        RECT 626.100 210.150 627.900 211.950 ;
        RECT 623.100 205.800 627.300 206.700 ;
        RECT 599.100 198.000 600.900 201.600 ;
        RECT 602.100 198.600 603.900 201.600 ;
        RECT 605.100 198.000 606.900 201.600 ;
        RECT 620.400 198.000 622.200 204.600 ;
        RECT 625.500 198.600 627.300 205.800 ;
        RECT 638.100 204.600 639.000 211.950 ;
        RECT 641.400 207.600 642.300 218.100 ;
        RECT 643.200 214.050 645.000 215.850 ;
        RECT 665.100 214.050 666.300 227.400 ;
        RECT 683.100 222.600 684.900 233.400 ;
        RECT 686.100 223.500 688.200 234.000 ;
        RECT 683.100 221.400 688.200 222.600 ;
        RECT 690.600 222.300 692.400 233.400 ;
        RECT 695.100 223.500 696.900 234.000 ;
        RECT 698.100 222.300 699.900 233.400 ;
        RECT 686.100 220.500 688.200 221.400 ;
        RECT 689.100 221.400 692.400 222.300 ;
        RECT 689.100 217.050 690.300 221.400 ;
        RECT 695.100 221.100 699.900 222.300 ;
        RECT 710.100 222.600 711.900 233.400 ;
        RECT 713.100 223.500 714.900 234.000 ;
        RECT 710.100 221.400 714.900 222.600 ;
        RECT 695.100 220.200 697.200 221.100 ;
        RECT 712.800 220.500 714.900 221.400 ;
        RECT 717.600 221.400 719.400 233.400 ;
        RECT 722.100 223.500 723.900 234.000 ;
        RECT 725.100 222.300 726.900 233.400 ;
        RECT 740.100 227.400 741.900 234.000 ;
        RECT 743.100 227.400 744.900 233.400 ;
        RECT 746.100 228.000 747.900 234.000 ;
        RECT 743.400 227.100 744.900 227.400 ;
        RECT 749.100 227.400 750.900 233.400 ;
        RECT 761.100 227.400 762.900 234.000 ;
        RECT 764.100 227.400 765.900 233.400 ;
        RECT 767.100 227.400 768.900 234.000 ;
        RECT 782.100 227.400 783.900 234.000 ;
        RECT 785.100 227.400 786.900 233.400 ;
        RECT 788.100 227.400 789.900 234.000 ;
        RECT 800.700 227.400 802.500 234.000 ;
        RECT 749.100 227.100 750.000 227.400 ;
        RECT 743.400 226.200 750.000 227.100 ;
        RECT 722.400 221.400 726.900 222.300 ;
        RECT 691.800 219.300 697.200 220.200 ;
        RECT 717.600 220.050 718.800 221.400 ;
        RECT 691.800 217.500 693.600 219.300 ;
        RECT 717.300 219.000 718.800 220.050 ;
        RECT 722.400 219.300 724.500 221.400 ;
        RECT 717.300 217.050 718.200 219.000 ;
        RECT 688.800 216.300 690.900 217.050 ;
        RECT 683.400 214.050 685.200 215.850 ;
        RECT 688.800 214.950 691.800 216.300 ;
        RECT 643.500 211.950 645.600 214.050 ;
        RECT 646.800 211.950 648.900 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 683.100 211.950 685.200 214.050 ;
        RECT 688.200 212.100 690.000 213.900 ;
        RECT 646.800 210.150 648.600 211.950 ;
        RECT 662.250 210.150 664.050 211.950 ;
        RECT 640.200 206.700 642.300 207.600 ;
        RECT 646.950 207.450 649.050 208.050 ;
        RECT 661.950 207.450 664.050 208.050 ;
        RECT 640.200 205.800 645.600 206.700 ;
        RECT 646.950 206.550 664.050 207.450 ;
        RECT 646.950 205.950 649.050 206.550 ;
        RECT 661.950 205.950 664.050 206.550 ;
        RECT 665.100 206.700 666.300 211.950 ;
        RECT 668.100 210.150 669.900 211.950 ;
        RECT 687.900 210.000 690.000 212.100 ;
        RECT 690.900 208.200 691.800 214.950 ;
        RECT 693.300 214.200 695.100 216.000 ;
        RECT 693.000 212.100 695.100 214.200 ;
        RECT 710.400 214.050 712.200 215.850 ;
        RECT 716.100 214.950 718.200 217.050 ;
        RECT 719.100 217.500 721.200 217.800 ;
        RECT 719.100 215.700 723.000 217.500 ;
        RECT 697.800 211.800 699.900 214.050 ;
        RECT 710.100 211.950 712.200 214.050 ;
        RECT 716.700 214.800 718.200 214.950 ;
        RECT 716.700 213.900 719.100 214.800 ;
        RECT 697.800 211.200 699.600 211.800 ;
        RECT 693.000 210.000 699.600 211.200 ;
        RECT 714.900 211.200 716.700 213.000 ;
        RECT 693.000 209.100 695.100 210.000 ;
        RECT 714.900 209.100 717.000 211.200 ;
        RECT 665.100 205.800 669.300 206.700 ;
        RECT 638.100 198.600 639.900 204.600 ;
        RECT 641.100 198.000 642.900 204.000 ;
        RECT 644.700 201.600 645.600 205.800 ;
        RECT 644.100 198.600 645.900 201.600 ;
        RECT 647.100 198.600 648.900 201.600 ;
        RECT 647.700 198.000 648.900 198.600 ;
        RECT 662.400 198.000 664.200 204.600 ;
        RECT 667.500 198.600 669.300 205.800 ;
        RECT 685.500 205.500 687.600 207.900 ;
        RECT 688.800 206.100 691.800 208.200 ;
        RECT 692.700 207.300 694.500 209.100 ;
        RECT 717.900 208.200 719.100 213.900 ;
        RECT 720.000 214.050 721.800 214.500 ;
        RECT 743.100 214.050 744.900 215.850 ;
        RECT 749.100 214.050 750.000 226.200 ;
        RECT 764.100 214.050 765.300 227.400 ;
        RECT 785.100 214.050 786.300 227.400 ;
        RECT 801.000 224.100 802.800 225.900 ;
        RECT 803.700 222.900 805.500 233.400 ;
        RECT 803.100 221.400 805.500 222.900 ;
        RECT 808.800 221.400 810.600 234.000 ;
        RECT 821.100 227.400 822.900 234.000 ;
        RECT 824.100 227.400 825.900 233.400 ;
        RECT 803.100 214.050 804.300 221.400 ;
        RECT 809.100 214.050 810.900 215.850 ;
        RECT 821.100 214.050 822.900 215.850 ;
        RECT 824.100 214.050 825.300 227.400 ;
        RECT 839.100 221.400 840.900 233.400 ;
        RECT 842.100 222.300 843.900 233.400 ;
        RECT 845.100 223.200 846.900 234.000 ;
        RECT 848.100 222.300 849.900 233.400 ;
        RECT 842.100 221.400 849.900 222.300 ;
        RECT 863.100 221.400 864.900 233.400 ;
        RECT 866.100 222.300 867.900 233.400 ;
        RECT 869.100 223.200 870.900 234.000 ;
        RECT 872.100 222.300 873.900 233.400 ;
        RECT 884.100 227.400 885.900 233.400 ;
        RECT 887.100 228.000 888.900 234.000 ;
        RECT 866.100 221.400 873.900 222.300 ;
        RECT 885.000 227.100 885.900 227.400 ;
        RECT 890.100 227.400 891.900 233.400 ;
        RECT 893.100 227.400 894.900 234.000 ;
        RECT 905.100 227.400 906.900 234.000 ;
        RECT 908.100 227.400 909.900 233.400 ;
        RECT 911.100 228.000 912.900 234.000 ;
        RECT 890.100 227.100 891.600 227.400 ;
        RECT 885.000 226.200 891.600 227.100 ;
        RECT 908.400 227.100 909.900 227.400 ;
        RECT 914.100 227.400 915.900 233.400 ;
        RECT 914.100 227.100 915.000 227.400 ;
        RECT 908.400 226.200 915.000 227.100 ;
        RECT 839.400 214.050 840.300 221.400 ;
        RECT 844.950 214.050 846.750 215.850 ;
        RECT 863.400 214.050 864.300 221.400 ;
        RECT 874.950 216.450 879.000 217.050 ;
        RECT 868.950 214.050 870.750 215.850 ;
        RECT 874.950 214.950 879.450 216.450 ;
        RECT 720.000 212.700 726.900 214.050 ;
        RECT 724.800 211.950 726.900 212.700 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 742.950 211.950 745.050 214.050 ;
        RECT 745.950 211.950 748.050 214.050 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 787.950 211.950 790.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 683.100 204.600 687.600 205.500 ;
        RECT 683.100 198.600 684.900 204.600 ;
        RECT 690.900 204.000 691.800 206.100 ;
        RECT 695.400 207.000 697.500 207.600 ;
        RECT 695.400 205.500 699.900 207.000 ;
        RECT 712.800 205.500 714.900 206.700 ;
        RECT 716.100 206.100 719.100 208.200 ;
        RECT 720.000 209.400 721.800 211.200 ;
        RECT 724.800 210.150 726.600 211.950 ;
        RECT 740.100 210.150 741.900 211.950 ;
        RECT 746.100 210.150 747.900 211.950 ;
        RECT 720.000 207.300 722.100 209.400 ;
        RECT 749.100 208.200 750.000 211.950 ;
        RECT 761.250 210.150 763.050 211.950 ;
        RECT 720.000 206.400 726.300 207.300 ;
        RECT 698.400 204.600 699.900 205.500 ;
        RECT 686.400 198.000 688.200 203.700 ;
        RECT 690.900 198.600 692.700 204.000 ;
        RECT 695.100 198.000 696.900 203.700 ;
        RECT 698.100 198.600 699.900 204.600 ;
        RECT 710.100 204.600 714.900 205.500 ;
        RECT 717.900 204.600 719.100 206.100 ;
        RECT 725.100 204.600 726.300 206.400 ;
        RECT 710.100 198.600 711.900 204.600 ;
        RECT 713.100 198.000 714.900 203.700 ;
        RECT 717.600 198.600 719.400 204.600 ;
        RECT 722.100 198.000 723.900 203.700 ;
        RECT 725.100 198.600 726.900 204.600 ;
        RECT 740.100 198.000 741.900 207.600 ;
        RECT 746.700 207.000 750.000 208.200 ;
        RECT 746.700 198.600 748.500 207.000 ;
        RECT 764.100 206.700 765.300 211.950 ;
        RECT 767.100 210.150 768.900 211.950 ;
        RECT 782.250 210.150 784.050 211.950 ;
        RECT 769.950 207.450 772.050 208.050 ;
        RECT 781.950 207.450 784.050 208.050 ;
        RECT 764.100 205.800 768.300 206.700 ;
        RECT 769.950 206.550 784.050 207.450 ;
        RECT 769.950 205.950 772.050 206.550 ;
        RECT 781.950 205.950 784.050 206.550 ;
        RECT 785.100 206.700 786.300 211.950 ;
        RECT 788.100 210.150 789.900 211.950 ;
        RECT 800.100 210.150 801.900 211.950 ;
        RECT 803.100 207.600 804.300 211.950 ;
        RECT 806.100 210.150 807.900 211.950 ;
        RECT 800.700 206.700 804.300 207.600 ;
        RECT 785.100 205.800 789.300 206.700 ;
        RECT 761.400 198.000 763.200 204.600 ;
        RECT 766.500 198.600 768.300 205.800 ;
        RECT 782.400 198.000 784.200 204.600 ;
        RECT 787.500 198.600 789.300 205.800 ;
        RECT 800.700 204.600 801.900 206.700 ;
        RECT 800.100 198.600 801.900 204.600 ;
        RECT 803.100 203.700 810.900 205.050 ;
        RECT 803.100 198.600 804.900 203.700 ;
        RECT 806.100 198.000 807.900 202.800 ;
        RECT 809.100 198.600 810.900 203.700 ;
        RECT 824.100 201.600 825.300 211.950 ;
        RECT 829.950 204.450 832.050 205.050 ;
        RECT 835.950 204.450 838.050 205.050 ;
        RECT 829.950 203.550 838.050 204.450 ;
        RECT 829.950 202.950 832.050 203.550 ;
        RECT 835.950 202.950 838.050 203.550 ;
        RECT 839.400 204.600 840.300 211.950 ;
        RECT 841.950 210.150 843.750 211.950 ;
        RECT 848.100 210.150 849.900 211.950 ;
        RECT 863.400 204.600 864.300 211.950 ;
        RECT 865.950 210.150 867.750 211.950 ;
        RECT 872.100 210.150 873.900 211.950 ;
        RECT 871.950 207.450 874.050 208.050 ;
        RECT 878.550 207.450 879.450 214.950 ;
        RECT 885.000 214.050 885.900 226.200 ;
        RECT 886.950 219.450 889.050 219.900 ;
        RECT 892.950 219.450 895.050 220.200 ;
        RECT 886.950 218.550 895.050 219.450 ;
        RECT 886.950 217.800 889.050 218.550 ;
        RECT 892.950 218.100 895.050 218.550 ;
        RECT 890.100 214.050 891.900 215.850 ;
        RECT 908.100 214.050 909.900 215.850 ;
        RECT 914.100 214.050 915.000 226.200 ;
        RECT 883.950 211.950 886.050 214.050 ;
        RECT 886.950 211.950 889.050 214.050 ;
        RECT 889.950 211.950 892.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 904.950 211.950 907.050 214.050 ;
        RECT 907.950 211.950 910.050 214.050 ;
        RECT 910.950 211.950 913.050 214.050 ;
        RECT 913.950 211.950 916.050 214.050 ;
        RECT 871.950 206.550 879.450 207.450 ;
        RECT 885.000 208.200 885.900 211.950 ;
        RECT 887.100 210.150 888.900 211.950 ;
        RECT 893.100 210.150 894.900 211.950 ;
        RECT 905.100 210.150 906.900 211.950 ;
        RECT 911.100 210.150 912.900 211.950 ;
        RECT 914.100 208.200 915.000 211.950 ;
        RECT 885.000 207.000 888.300 208.200 ;
        RECT 871.950 205.950 874.050 206.550 ;
        RECT 839.400 203.400 844.500 204.600 ;
        RECT 821.100 198.000 822.900 201.600 ;
        RECT 824.100 198.600 825.900 201.600 ;
        RECT 839.700 198.000 841.500 201.600 ;
        RECT 842.700 198.600 844.500 203.400 ;
        RECT 847.200 198.000 849.000 204.600 ;
        RECT 863.400 203.400 868.500 204.600 ;
        RECT 863.700 198.000 865.500 201.600 ;
        RECT 866.700 198.600 868.500 203.400 ;
        RECT 871.200 198.000 873.000 204.600 ;
        RECT 886.500 198.600 888.300 207.000 ;
        RECT 893.100 198.000 894.900 207.600 ;
        RECT 905.100 198.000 906.900 207.600 ;
        RECT 911.700 207.000 915.000 208.200 ;
        RECT 911.700 198.600 913.500 207.000 ;
        RECT 11.100 191.400 12.900 195.000 ;
        RECT 14.100 191.400 15.900 194.400 ;
        RECT 14.100 181.050 15.300 191.400 ;
        RECT 29.700 188.400 31.500 195.000 ;
        RECT 34.200 188.400 36.000 194.400 ;
        RECT 38.700 188.400 40.500 195.000 ;
        RECT 53.100 191.400 54.900 194.400 ;
        RECT 56.100 191.400 57.900 195.000 ;
        RECT 49.950 189.450 52.050 190.050 ;
        RECT 44.550 188.550 52.050 189.450 ;
        RECT 29.250 181.050 31.050 182.850 ;
        RECT 35.100 181.050 36.300 188.400 ;
        RECT 37.950 186.450 40.050 187.200 ;
        RECT 44.550 186.450 45.450 188.550 ;
        RECT 49.950 187.950 52.050 188.550 ;
        RECT 37.950 185.550 45.450 186.450 ;
        RECT 37.950 185.100 40.050 185.550 ;
        RECT 41.100 181.050 42.900 182.850 ;
        RECT 53.700 181.050 54.900 191.400 ;
        RECT 73.500 186.000 75.300 194.400 ;
        RECT 72.000 184.800 75.300 186.000 ;
        RECT 80.100 185.400 81.900 195.000 ;
        RECT 92.100 189.300 93.900 194.400 ;
        RECT 95.100 190.200 96.900 195.000 ;
        RECT 98.100 189.300 99.900 194.400 ;
        RECT 92.100 187.950 99.900 189.300 ;
        RECT 101.100 188.400 102.900 194.400 ;
        RECT 112.950 192.450 115.050 193.050 ;
        RECT 104.550 192.000 115.050 192.450 ;
        RECT 103.950 191.550 115.050 192.000 ;
        RECT 101.100 186.300 102.300 188.400 ;
        RECT 103.950 187.950 106.050 191.550 ;
        RECT 112.950 190.950 115.050 191.550 ;
        RECT 116.100 191.400 117.900 194.400 ;
        RECT 119.100 191.400 120.900 195.000 ;
        RECT 134.700 191.400 136.500 195.000 ;
        RECT 98.700 185.400 102.300 186.300 ;
        RECT 58.950 183.450 63.000 184.050 ;
        RECT 58.950 181.950 63.450 183.450 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 28.950 178.950 31.050 181.050 ;
        RECT 31.950 178.950 34.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 52.950 178.950 55.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 11.100 177.150 12.900 178.950 ;
        RECT 14.100 165.600 15.300 178.950 ;
        RECT 32.250 177.150 34.050 178.950 ;
        RECT 35.100 173.400 36.000 178.950 ;
        RECT 38.100 177.150 39.900 178.950 ;
        RECT 35.100 172.500 39.900 173.400 ;
        RECT 29.100 170.400 36.900 171.300 ;
        RECT 11.100 159.000 12.900 165.600 ;
        RECT 14.100 159.600 15.900 165.600 ;
        RECT 29.100 159.600 30.900 170.400 ;
        RECT 32.100 159.000 33.900 169.500 ;
        RECT 35.100 160.500 36.900 170.400 ;
        RECT 38.100 161.400 39.900 172.500 ;
        RECT 41.100 160.500 42.900 171.600 ;
        RECT 53.700 165.600 54.900 178.950 ;
        RECT 56.100 177.150 57.900 178.950 ;
        RECT 62.550 178.050 63.450 181.950 ;
        RECT 72.000 181.050 72.900 184.800 ;
        RECT 87.000 183.450 91.050 184.050 ;
        RECT 74.100 181.050 75.900 182.850 ;
        RECT 80.100 181.050 81.900 182.850 ;
        RECT 86.550 181.950 91.050 183.450 ;
        RECT 70.950 178.950 73.050 181.050 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 58.950 176.550 63.450 178.050 ;
        RECT 58.950 175.950 63.000 176.550 ;
        RECT 72.000 166.800 72.900 178.950 ;
        RECT 77.100 177.150 78.900 178.950 ;
        RECT 86.550 177.450 87.450 181.950 ;
        RECT 95.100 181.050 96.900 182.850 ;
        RECT 98.700 181.050 99.900 185.400 ;
        RECT 101.100 181.050 102.900 182.850 ;
        RECT 116.700 181.050 117.900 191.400 ;
        RECT 137.700 189.600 139.500 194.400 ;
        RECT 134.400 188.400 139.500 189.600 ;
        RECT 142.200 188.400 144.000 195.000 ;
        RECT 134.400 181.050 135.300 188.400 ;
        RECT 157.500 186.000 159.300 194.400 ;
        RECT 156.000 184.800 159.300 186.000 ;
        RECT 164.100 185.400 165.900 195.000 ;
        RECT 179.100 191.400 180.900 194.400 ;
        RECT 182.100 191.400 183.900 195.000 ;
        RECT 136.950 181.050 138.750 182.850 ;
        RECT 143.100 181.050 144.900 182.850 ;
        RECT 156.000 181.050 156.900 184.800 ;
        RECT 158.100 181.050 159.900 182.850 ;
        RECT 164.100 181.050 165.900 182.850 ;
        RECT 179.700 181.050 180.900 191.400 ;
        RECT 194.700 187.200 196.500 194.400 ;
        RECT 199.800 188.400 201.600 195.000 ;
        RECT 215.100 188.400 216.900 194.400 ;
        RECT 194.700 186.300 198.900 187.200 ;
        RECT 194.100 181.050 195.900 182.850 ;
        RECT 197.700 181.050 198.900 186.300 ;
        RECT 215.700 186.300 216.900 188.400 ;
        RECT 218.100 189.300 219.900 194.400 ;
        RECT 221.100 190.200 222.900 195.000 ;
        RECT 224.100 189.300 225.900 194.400 ;
        RECT 236.100 191.400 237.900 195.000 ;
        RECT 239.100 191.400 240.900 194.400 ;
        RECT 242.100 191.400 243.900 195.000 ;
        RECT 257.100 191.400 258.900 195.000 ;
        RECT 260.100 191.400 261.900 194.400 ;
        RECT 263.100 191.400 264.900 195.000 ;
        RECT 218.100 187.950 225.900 189.300 ;
        RECT 215.700 185.400 219.300 186.300 ;
        RECT 199.950 181.050 201.750 182.850 ;
        RECT 215.100 181.050 216.900 182.850 ;
        RECT 218.100 181.050 219.300 185.400 ;
        RECT 221.100 181.050 222.900 182.850 ;
        RECT 239.700 181.050 240.600 191.400 ;
        RECT 260.400 181.050 261.300 191.400 ;
        RECT 275.400 188.400 277.200 195.000 ;
        RECT 280.500 187.200 282.300 194.400 ;
        RECT 293.100 191.400 294.900 195.000 ;
        RECT 296.100 191.400 297.900 194.400 ;
        RECT 278.100 186.300 282.300 187.200 ;
        RECT 268.950 181.950 271.050 184.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 160.950 178.950 163.050 181.050 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 181.950 178.950 184.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 83.550 177.000 87.450 177.450 ;
        RECT 92.100 177.150 93.900 178.950 ;
        RECT 82.950 176.550 87.450 177.000 ;
        RECT 82.950 172.950 85.050 176.550 ;
        RECT 98.700 171.600 99.900 178.950 ;
        RECT 72.000 165.900 78.600 166.800 ;
        RECT 72.000 165.600 72.900 165.900 ;
        RECT 35.100 159.600 42.900 160.500 ;
        RECT 53.100 159.600 54.900 165.600 ;
        RECT 56.100 159.000 57.900 165.600 ;
        RECT 71.100 159.600 72.900 165.600 ;
        RECT 77.100 165.600 78.600 165.900 ;
        RECT 74.100 159.000 75.900 165.000 ;
        RECT 77.100 159.600 78.900 165.600 ;
        RECT 80.100 159.000 81.900 165.600 ;
        RECT 92.400 159.000 94.200 171.600 ;
        RECT 97.500 170.100 99.900 171.600 ;
        RECT 97.500 159.600 99.300 170.100 ;
        RECT 100.200 167.100 102.000 168.900 ;
        RECT 116.700 165.600 117.900 178.950 ;
        RECT 119.100 177.150 120.900 178.950 ;
        RECT 134.400 171.600 135.300 178.950 ;
        RECT 139.950 177.150 141.750 178.950 ;
        RECT 136.950 174.450 139.050 175.050 ;
        RECT 148.950 174.450 151.050 175.050 ;
        RECT 136.950 173.550 151.050 174.450 ;
        RECT 136.950 172.950 139.050 173.550 ;
        RECT 148.950 172.950 151.050 173.550 ;
        RECT 100.500 159.000 102.300 165.600 ;
        RECT 116.100 159.600 117.900 165.600 ;
        RECT 119.100 159.000 120.900 165.600 ;
        RECT 134.100 159.600 135.900 171.600 ;
        RECT 137.100 170.700 144.900 171.600 ;
        RECT 137.100 159.600 138.900 170.700 ;
        RECT 140.100 159.000 141.900 169.800 ;
        RECT 143.100 159.600 144.900 170.700 ;
        RECT 156.000 166.800 156.900 178.950 ;
        RECT 161.100 177.150 162.900 178.950 ;
        RECT 163.950 174.450 166.050 175.050 ;
        RECT 169.950 174.450 172.050 175.050 ;
        RECT 163.950 173.550 172.050 174.450 ;
        RECT 163.950 172.950 166.050 173.550 ;
        RECT 169.950 172.950 172.050 173.550 ;
        RECT 156.000 165.900 162.600 166.800 ;
        RECT 156.000 165.600 156.900 165.900 ;
        RECT 155.100 159.600 156.900 165.600 ;
        RECT 161.100 165.600 162.600 165.900 ;
        RECT 179.700 165.600 180.900 178.950 ;
        RECT 182.100 177.150 183.900 178.950 ;
        RECT 197.700 165.600 198.900 178.950 ;
        RECT 218.100 171.600 219.300 178.950 ;
        RECT 224.100 177.150 225.900 178.950 ;
        RECT 236.100 177.150 237.900 178.950 ;
        RECT 239.700 171.600 240.600 178.950 ;
        RECT 241.950 177.150 243.750 178.950 ;
        RECT 257.250 177.150 259.050 178.950 ;
        RECT 260.400 171.600 261.300 178.950 ;
        RECT 263.100 177.150 264.900 178.950 ;
        RECT 269.550 178.050 270.450 181.950 ;
        RECT 275.250 181.050 277.050 182.850 ;
        RECT 278.100 181.050 279.300 186.300 ;
        RECT 281.100 181.050 282.900 182.850 ;
        RECT 296.100 181.050 297.300 191.400 ;
        RECT 308.100 189.300 309.900 194.400 ;
        RECT 311.100 190.200 312.900 195.000 ;
        RECT 314.100 189.300 315.900 194.400 ;
        RECT 308.100 187.950 315.900 189.300 ;
        RECT 317.100 188.400 318.900 194.400 ;
        RECT 337.200 191.400 339.900 194.400 ;
        RECT 341.100 191.400 342.900 195.000 ;
        RECT 344.100 191.400 345.900 194.400 ;
        RECT 347.100 191.400 349.200 195.000 ;
        RECT 365.700 191.400 367.500 195.000 ;
        RECT 337.200 190.500 338.100 191.400 ;
        RECT 344.400 190.500 345.300 191.400 ;
        RECT 332.700 189.600 345.300 190.500 ;
        RECT 368.700 189.600 370.500 194.400 ;
        RECT 317.100 186.300 318.300 188.400 ;
        RECT 314.700 185.400 318.300 186.300 ;
        RECT 303.000 183.450 307.050 184.050 ;
        RECT 302.550 181.950 307.050 183.450 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 277.950 178.950 280.050 181.050 ;
        RECT 280.950 178.950 283.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 265.950 176.550 270.450 178.050 ;
        RECT 265.950 175.950 270.000 176.550 ;
        RECT 218.100 170.100 220.500 171.600 ;
        RECT 216.000 167.100 217.800 168.900 ;
        RECT 158.100 159.000 159.900 165.000 ;
        RECT 161.100 159.600 162.900 165.600 ;
        RECT 164.100 159.000 165.900 165.600 ;
        RECT 179.100 159.600 180.900 165.600 ;
        RECT 182.100 159.000 183.900 165.600 ;
        RECT 194.100 159.000 195.900 165.600 ;
        RECT 197.100 159.600 198.900 165.600 ;
        RECT 200.100 159.000 201.900 165.600 ;
        RECT 215.700 159.000 217.500 165.600 ;
        RECT 218.700 159.600 220.500 170.100 ;
        RECT 223.800 159.000 225.600 171.600 ;
        RECT 237.000 170.400 240.600 171.600 ;
        RECT 237.000 159.600 238.800 170.400 ;
        RECT 242.100 159.000 243.900 171.600 ;
        RECT 257.100 159.000 258.900 171.600 ;
        RECT 260.400 170.400 264.000 171.600 ;
        RECT 262.200 159.600 264.000 170.400 ;
        RECT 278.100 165.600 279.300 178.950 ;
        RECT 293.100 177.150 294.900 178.950 ;
        RECT 296.100 165.600 297.300 178.950 ;
        RECT 302.550 178.050 303.450 181.950 ;
        RECT 311.100 181.050 312.900 182.850 ;
        RECT 314.700 181.050 315.900 185.400 ;
        RECT 317.100 181.050 318.900 182.850 ;
        RECT 332.700 181.050 333.900 189.600 ;
        RECT 365.400 188.400 370.500 189.600 ;
        RECT 373.200 188.400 375.000 195.000 ;
        RECT 389.100 191.400 390.900 194.400 ;
        RECT 392.100 191.400 393.900 195.000 ;
        RECT 341.250 181.050 343.050 182.850 ;
        RECT 365.400 181.050 366.300 188.400 ;
        RECT 367.950 181.050 369.750 182.850 ;
        RECT 374.100 181.050 375.900 182.850 ;
        RECT 389.700 181.050 390.900 191.400 ;
        RECT 404.100 188.400 405.900 194.400 ;
        RECT 404.700 186.300 405.900 188.400 ;
        RECT 407.100 189.300 408.900 194.400 ;
        RECT 410.100 190.200 411.900 195.000 ;
        RECT 413.100 189.300 414.900 194.400 ;
        RECT 407.100 187.950 414.900 189.300 ;
        RECT 428.700 187.200 430.500 194.400 ;
        RECT 433.800 188.400 435.600 195.000 ;
        RECT 428.700 186.300 432.900 187.200 ;
        RECT 404.700 185.400 408.300 186.300 ;
        RECT 404.100 181.050 405.900 182.850 ;
        RECT 407.100 181.050 408.300 185.400 ;
        RECT 410.100 181.050 411.900 182.850 ;
        RECT 428.100 181.050 429.900 182.850 ;
        RECT 431.700 181.050 432.900 186.300 ;
        RECT 451.500 186.000 453.300 194.400 ;
        RECT 450.000 184.800 453.300 186.000 ;
        RECT 458.100 185.400 459.900 195.000 ;
        RECT 470.100 188.400 471.900 194.400 ;
        RECT 473.100 189.000 474.900 195.000 ;
        RECT 479.700 194.400 480.900 195.000 ;
        RECT 476.100 191.400 477.900 194.400 ;
        RECT 479.100 191.400 480.900 194.400 ;
        RECT 433.950 181.050 435.750 182.850 ;
        RECT 450.000 181.050 450.900 184.800 ;
        RECT 452.100 181.050 453.900 182.850 ;
        RECT 458.100 181.050 459.900 182.850 ;
        RECT 470.100 181.050 471.000 188.400 ;
        RECT 476.700 187.200 477.600 191.400 ;
        RECT 494.400 188.400 496.200 195.000 ;
        RECT 499.500 187.200 501.300 194.400 ;
        RECT 513.600 190.200 515.400 194.400 ;
        RECT 472.200 186.300 477.600 187.200 ;
        RECT 497.100 186.300 501.300 187.200 ;
        RECT 512.700 188.400 515.400 190.200 ;
        RECT 516.600 188.400 518.400 195.000 ;
        RECT 472.200 185.400 474.300 186.300 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 332.400 178.950 334.500 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 340.950 178.950 343.050 181.050 ;
        RECT 347.100 178.950 349.200 181.050 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 367.950 178.950 370.050 181.050 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 470.100 178.950 472.200 181.050 ;
        RECT 298.950 176.550 303.450 178.050 ;
        RECT 308.100 177.150 309.900 178.950 ;
        RECT 298.950 175.950 303.000 176.550 ;
        RECT 314.700 171.600 315.900 178.950 ;
        RECT 275.100 159.000 276.900 165.600 ;
        RECT 278.100 159.600 279.900 165.600 ;
        RECT 281.100 159.000 282.900 165.600 ;
        RECT 293.100 159.000 294.900 165.600 ;
        RECT 296.100 159.600 297.900 165.600 ;
        RECT 308.400 159.000 310.200 171.600 ;
        RECT 313.500 170.100 315.900 171.600 ;
        RECT 313.500 159.600 315.300 170.100 ;
        RECT 316.200 167.100 318.000 168.900 ;
        RECT 316.500 159.000 318.300 165.600 ;
        RECT 329.100 160.500 330.900 169.800 ;
        RECT 332.700 169.200 333.900 178.950 ;
        RECT 337.950 177.150 339.750 178.950 ;
        RECT 347.100 177.150 348.900 178.950 ;
        RECT 365.400 171.600 366.300 178.950 ;
        RECT 370.950 177.150 372.750 178.950 ;
        RECT 332.100 161.400 333.900 169.200 ;
        RECT 335.100 169.200 342.900 170.100 ;
        RECT 335.100 160.500 336.900 169.200 ;
        RECT 329.100 159.600 336.900 160.500 ;
        RECT 338.100 160.500 339.900 168.300 ;
        RECT 341.100 161.400 342.900 169.200 ;
        RECT 344.100 169.500 351.900 170.400 ;
        RECT 344.100 160.500 345.900 169.500 ;
        RECT 338.100 159.600 345.900 160.500 ;
        RECT 347.100 159.000 348.900 168.600 ;
        RECT 350.100 159.600 351.900 169.500 ;
        RECT 365.100 159.600 366.900 171.600 ;
        RECT 368.100 170.700 375.900 171.600 ;
        RECT 368.100 159.600 369.900 170.700 ;
        RECT 371.100 159.000 372.900 169.800 ;
        RECT 374.100 159.600 375.900 170.700 ;
        RECT 389.700 165.600 390.900 178.950 ;
        RECT 392.100 177.150 393.900 178.950 ;
        RECT 407.100 171.600 408.300 178.950 ;
        RECT 413.100 177.150 414.900 178.950 ;
        RECT 407.100 170.100 409.500 171.600 ;
        RECT 405.000 167.100 406.800 168.900 ;
        RECT 389.100 159.600 390.900 165.600 ;
        RECT 392.100 159.000 393.900 165.600 ;
        RECT 404.700 159.000 406.500 165.600 ;
        RECT 407.700 159.600 409.500 170.100 ;
        RECT 412.800 159.000 414.600 171.600 ;
        RECT 431.700 165.600 432.900 178.950 ;
        RECT 433.950 174.450 436.050 175.050 ;
        RECT 442.950 174.450 445.050 175.050 ;
        RECT 433.950 173.550 445.050 174.450 ;
        RECT 433.950 172.950 436.050 173.550 ;
        RECT 442.950 172.950 445.050 173.550 ;
        RECT 450.000 166.800 450.900 178.950 ;
        RECT 455.100 177.150 456.900 178.950 ;
        RECT 460.950 177.450 463.050 178.050 ;
        RECT 466.950 177.450 469.050 178.050 ;
        RECT 460.950 176.550 469.050 177.450 ;
        RECT 460.950 175.950 463.050 176.550 ;
        RECT 466.950 175.950 469.050 176.550 ;
        RECT 451.950 174.450 454.050 175.050 ;
        RECT 466.950 174.450 469.050 174.900 ;
        RECT 451.950 173.550 469.050 174.450 ;
        RECT 451.950 172.950 454.050 173.550 ;
        RECT 466.950 172.800 469.050 173.550 ;
        RECT 471.000 171.600 472.200 178.950 ;
        RECT 473.400 174.900 474.300 185.400 ;
        RECT 478.800 181.050 480.600 182.850 ;
        RECT 494.250 181.050 496.050 182.850 ;
        RECT 497.100 181.050 498.300 186.300 ;
        RECT 500.100 181.050 501.900 182.850 ;
        RECT 512.700 181.050 513.600 188.400 ;
        RECT 514.500 186.600 516.300 187.500 ;
        RECT 521.100 186.600 522.900 194.400 ;
        RECT 514.500 185.700 522.900 186.600 ;
        RECT 536.700 187.200 538.500 194.400 ;
        RECT 541.800 188.400 543.600 195.000 ;
        RECT 557.100 188.400 558.900 194.400 ;
        RECT 560.100 189.300 561.900 195.000 ;
        RECT 564.300 189.000 566.100 194.400 ;
        RECT 568.800 189.300 570.600 195.000 ;
        RECT 557.100 187.500 558.600 188.400 ;
        RECT 536.700 186.300 540.900 187.200 ;
        RECT 475.500 178.950 477.600 181.050 ;
        RECT 478.800 178.950 480.900 181.050 ;
        RECT 493.950 178.950 496.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 512.100 178.950 514.200 181.050 ;
        RECT 515.400 178.950 517.500 181.050 ;
        RECT 475.200 177.150 477.000 178.950 ;
        RECT 473.100 174.300 474.900 174.900 ;
        RECT 473.100 173.100 480.900 174.300 ;
        RECT 479.700 171.600 480.900 173.100 ;
        RECT 471.000 170.100 473.400 171.600 ;
        RECT 450.000 165.900 456.600 166.800 ;
        RECT 450.000 165.600 450.900 165.900 ;
        RECT 428.100 159.000 429.900 165.600 ;
        RECT 431.100 159.600 432.900 165.600 ;
        RECT 434.100 159.000 435.900 165.600 ;
        RECT 449.100 159.600 450.900 165.600 ;
        RECT 455.100 165.600 456.600 165.900 ;
        RECT 452.100 159.000 453.900 165.000 ;
        RECT 455.100 159.600 456.900 165.600 ;
        RECT 458.100 159.000 459.900 165.600 ;
        RECT 471.600 159.600 473.400 170.100 ;
        RECT 474.600 159.000 476.400 171.600 ;
        RECT 479.100 159.600 480.900 171.600 ;
        RECT 497.100 165.600 498.300 178.950 ;
        RECT 512.700 171.600 513.600 178.950 ;
        RECT 516.000 177.150 517.800 178.950 ;
        RECT 494.100 159.000 495.900 165.600 ;
        RECT 497.100 159.600 498.900 165.600 ;
        RECT 500.100 159.000 501.900 165.600 ;
        RECT 512.100 159.600 513.900 171.600 ;
        RECT 515.100 159.000 516.900 171.000 ;
        RECT 519.000 165.600 519.900 185.700 ;
        RECT 520.950 181.050 522.750 182.850 ;
        RECT 536.100 181.050 537.900 182.850 ;
        RECT 539.700 181.050 540.900 186.300 ;
        RECT 557.100 186.000 561.600 187.500 ;
        RECT 559.500 185.400 561.600 186.000 ;
        RECT 565.200 186.900 566.100 189.000 ;
        RECT 572.100 188.400 573.900 194.400 ;
        RECT 569.400 187.500 573.900 188.400 ;
        RECT 562.500 183.900 564.300 185.700 ;
        RECT 565.200 184.800 568.200 186.900 ;
        RECT 569.400 185.100 571.500 187.500 ;
        RECT 589.500 186.000 591.300 194.400 ;
        RECT 588.000 184.800 591.300 186.000 ;
        RECT 596.100 185.400 597.900 195.000 ;
        RECT 608.100 186.600 609.900 194.400 ;
        RECT 612.600 188.400 614.400 195.000 ;
        RECT 615.600 190.200 617.400 194.400 ;
        RECT 615.600 188.400 618.300 190.200 ;
        RECT 614.700 186.600 616.500 187.500 ;
        RECT 608.100 185.700 616.500 186.600 ;
        RECT 561.900 183.000 564.000 183.900 ;
        RECT 541.950 181.050 543.750 182.850 ;
        RECT 557.400 181.800 564.000 183.000 ;
        RECT 557.400 181.200 559.200 181.800 ;
        RECT 520.800 178.950 522.900 181.050 ;
        RECT 535.950 178.950 538.050 181.050 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 557.100 178.950 559.200 181.200 ;
        RECT 539.700 165.600 540.900 178.950 ;
        RECT 561.900 178.800 564.000 180.900 ;
        RECT 561.900 177.000 563.700 178.800 ;
        RECT 565.200 178.050 566.100 184.800 ;
        RECT 567.000 180.900 569.100 183.000 ;
        RECT 588.000 181.050 588.900 184.800 ;
        RECT 590.100 181.050 591.900 182.850 ;
        RECT 596.100 181.050 597.900 182.850 ;
        RECT 608.250 181.050 610.050 182.850 ;
        RECT 567.000 179.100 568.800 180.900 ;
        RECT 571.800 178.950 573.900 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 608.100 178.950 610.200 181.050 ;
        RECT 565.200 176.700 568.200 178.050 ;
        RECT 571.800 177.150 573.600 178.950 ;
        RECT 566.100 175.950 568.200 176.700 ;
        RECT 563.400 173.700 565.200 175.500 ;
        RECT 559.800 172.800 565.200 173.700 ;
        RECT 559.800 171.900 561.900 172.800 ;
        RECT 557.100 170.700 561.900 171.900 ;
        RECT 566.700 171.600 567.900 175.950 ;
        RECT 564.600 170.700 567.900 171.600 ;
        RECT 568.800 171.600 570.900 172.500 ;
        RECT 518.100 159.600 519.900 165.600 ;
        RECT 521.100 159.000 522.900 165.600 ;
        RECT 536.100 159.000 537.900 165.600 ;
        RECT 539.100 159.600 540.900 165.600 ;
        RECT 542.100 159.000 543.900 165.600 ;
        RECT 557.100 159.600 558.900 170.700 ;
        RECT 560.100 159.000 561.900 169.500 ;
        RECT 564.600 159.600 566.400 170.700 ;
        RECT 568.800 170.400 573.900 171.600 ;
        RECT 568.800 159.000 570.900 169.500 ;
        RECT 572.100 159.600 573.900 170.400 ;
        RECT 588.000 166.800 588.900 178.950 ;
        RECT 593.100 177.150 594.900 178.950 ;
        RECT 588.000 165.900 594.600 166.800 ;
        RECT 588.000 165.600 588.900 165.900 ;
        RECT 587.100 159.600 588.900 165.600 ;
        RECT 593.100 165.600 594.600 165.900 ;
        RECT 611.100 165.600 612.000 185.700 ;
        RECT 617.400 181.050 618.300 188.400 ;
        RECT 632.700 187.200 634.500 194.400 ;
        RECT 637.800 188.400 639.600 195.000 ;
        RECT 650.700 188.400 652.500 195.000 ;
        RECT 655.200 188.400 657.000 194.400 ;
        RECT 659.700 188.400 661.500 195.000 ;
        RECT 677.100 191.400 678.900 195.000 ;
        RECT 680.100 191.400 681.900 194.400 ;
        RECT 683.100 191.400 684.900 195.000 ;
        RECT 632.700 186.300 636.900 187.200 ;
        RECT 632.100 181.050 633.900 182.850 ;
        RECT 635.700 181.050 636.900 186.300 ;
        RECT 637.950 181.050 639.750 182.850 ;
        RECT 650.250 181.050 652.050 182.850 ;
        RECT 656.100 181.050 657.300 188.400 ;
        RECT 658.950 186.450 661.050 187.050 ;
        RECT 667.950 186.450 670.050 187.050 ;
        RECT 658.950 185.550 670.050 186.450 ;
        RECT 658.950 184.950 661.050 185.550 ;
        RECT 667.950 184.950 670.050 185.550 ;
        RECT 662.100 181.050 663.900 182.850 ;
        RECT 680.700 181.050 681.600 191.400 ;
        RECT 698.100 188.400 699.900 194.400 ;
        RECT 698.700 186.300 699.900 188.400 ;
        RECT 701.100 189.300 702.900 194.400 ;
        RECT 704.100 190.200 705.900 195.000 ;
        RECT 707.100 189.300 708.900 194.400 ;
        RECT 719.100 191.400 720.900 195.000 ;
        RECT 722.100 191.400 723.900 194.400 ;
        RECT 725.100 191.400 726.900 195.000 ;
        RECT 701.100 187.950 708.900 189.300 ;
        RECT 698.700 185.400 702.300 186.300 ;
        RECT 698.100 181.050 699.900 182.850 ;
        RECT 701.100 181.050 702.300 185.400 ;
        RECT 704.100 181.050 705.900 182.850 ;
        RECT 722.700 181.050 723.600 191.400 ;
        RECT 740.400 188.400 742.200 195.000 ;
        RECT 745.500 187.200 747.300 194.400 ;
        RECT 761.400 188.400 763.200 195.000 ;
        RECT 766.500 187.200 768.300 194.400 ;
        RECT 743.100 186.300 747.300 187.200 ;
        RECT 764.100 186.300 768.300 187.200 ;
        RECT 740.250 181.050 742.050 182.850 ;
        RECT 743.100 181.050 744.300 186.300 ;
        RECT 746.100 181.050 747.900 182.850 ;
        RECT 761.250 181.050 763.050 182.850 ;
        RECT 764.100 181.050 765.300 186.300 ;
        RECT 784.500 186.000 786.300 194.400 ;
        RECT 783.000 184.800 786.300 186.000 ;
        RECT 791.100 185.400 792.900 195.000 ;
        RECT 806.100 191.400 807.900 195.000 ;
        RECT 809.100 191.400 810.900 194.400 ;
        RECT 767.100 181.050 768.900 182.850 ;
        RECT 783.000 181.050 783.900 184.800 ;
        RECT 801.000 183.450 805.050 184.050 ;
        RECT 785.100 181.050 786.900 182.850 ;
        RECT 791.100 181.050 792.900 182.850 ;
        RECT 800.550 181.950 805.050 183.450 ;
        RECT 613.500 178.950 615.600 181.050 ;
        RECT 616.800 178.950 618.900 181.050 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 718.950 178.950 721.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 613.200 177.150 615.000 178.950 ;
        RECT 617.400 171.600 618.300 178.950 ;
        RECT 590.100 159.000 591.900 165.000 ;
        RECT 593.100 159.600 594.900 165.600 ;
        RECT 596.100 159.000 597.900 165.600 ;
        RECT 608.100 159.000 609.900 165.600 ;
        RECT 611.100 159.600 612.900 165.600 ;
        RECT 614.100 159.000 615.900 171.000 ;
        RECT 617.100 159.600 618.900 171.600 ;
        RECT 635.700 165.600 636.900 178.950 ;
        RECT 653.250 177.150 655.050 178.950 ;
        RECT 656.100 173.400 657.000 178.950 ;
        RECT 659.100 177.150 660.900 178.950 ;
        RECT 677.100 177.150 678.900 178.950 ;
        RECT 656.100 172.500 660.900 173.400 ;
        RECT 650.100 170.400 657.900 171.300 ;
        RECT 632.100 159.000 633.900 165.600 ;
        RECT 635.100 159.600 636.900 165.600 ;
        RECT 638.100 159.000 639.900 165.600 ;
        RECT 650.100 159.600 651.900 170.400 ;
        RECT 653.100 159.000 654.900 169.500 ;
        RECT 656.100 160.500 657.900 170.400 ;
        RECT 659.100 161.400 660.900 172.500 ;
        RECT 680.700 171.600 681.600 178.950 ;
        RECT 682.950 177.150 684.750 178.950 ;
        RECT 701.100 171.600 702.300 178.950 ;
        RECT 707.100 177.150 708.900 178.950 ;
        RECT 719.100 177.150 720.900 178.950 ;
        RECT 703.950 174.450 706.050 175.050 ;
        RECT 715.950 174.450 718.050 175.050 ;
        RECT 703.950 173.550 718.050 174.450 ;
        RECT 703.950 172.950 706.050 173.550 ;
        RECT 715.950 172.950 718.050 173.550 ;
        RECT 722.700 171.600 723.600 178.950 ;
        RECT 724.950 177.150 726.750 178.950 ;
        RECT 662.100 160.500 663.900 171.600 ;
        RECT 656.100 159.600 663.900 160.500 ;
        RECT 678.000 170.400 681.600 171.600 ;
        RECT 678.000 159.600 679.800 170.400 ;
        RECT 683.100 159.000 684.900 171.600 ;
        RECT 701.100 170.100 703.500 171.600 ;
        RECT 699.000 167.100 700.800 168.900 ;
        RECT 698.700 159.000 700.500 165.600 ;
        RECT 701.700 159.600 703.500 170.100 ;
        RECT 706.800 159.000 708.600 171.600 ;
        RECT 720.000 170.400 723.600 171.600 ;
        RECT 720.000 159.600 721.800 170.400 ;
        RECT 725.100 159.000 726.900 171.600 ;
        RECT 743.100 165.600 744.300 178.950 ;
        RECT 764.100 165.600 765.300 178.950 ;
        RECT 783.000 166.800 783.900 178.950 ;
        RECT 788.100 177.150 789.900 178.950 ;
        RECT 800.550 177.450 801.450 181.950 ;
        RECT 809.100 181.050 810.300 191.400 ;
        RECT 824.100 189.300 825.900 194.400 ;
        RECT 827.100 190.200 828.900 195.000 ;
        RECT 830.100 189.300 831.900 194.400 ;
        RECT 824.100 187.950 831.900 189.300 ;
        RECT 833.100 188.400 834.900 194.400 ;
        RECT 848.100 188.400 849.900 194.400 ;
        RECT 833.100 186.300 834.300 188.400 ;
        RECT 830.700 185.400 834.300 186.300 ;
        RECT 848.700 186.300 849.900 188.400 ;
        RECT 851.100 189.300 852.900 194.400 ;
        RECT 854.100 190.200 855.900 195.000 ;
        RECT 857.100 189.300 858.900 194.400 ;
        RECT 851.100 187.950 858.900 189.300 ;
        RECT 869.100 188.400 870.900 194.400 ;
        RECT 869.700 186.300 870.900 188.400 ;
        RECT 872.100 189.300 873.900 194.400 ;
        RECT 875.100 190.200 876.900 195.000 ;
        RECT 878.100 189.300 879.900 194.400 ;
        RECT 890.700 191.400 892.500 195.000 ;
        RECT 893.700 189.600 895.500 194.400 ;
        RECT 872.100 187.950 879.900 189.300 ;
        RECT 890.400 188.400 895.500 189.600 ;
        RECT 898.200 188.400 900.000 195.000 ;
        RECT 911.100 189.300 912.900 194.400 ;
        RECT 914.100 190.200 915.900 195.000 ;
        RECT 917.100 189.300 918.900 194.400 ;
        RECT 848.700 185.400 852.300 186.300 ;
        RECT 869.700 185.400 873.300 186.300 ;
        RECT 827.100 181.050 828.900 182.850 ;
        RECT 830.700 181.050 831.900 185.400 ;
        RECT 835.950 183.450 840.000 184.050 ;
        RECT 833.100 181.050 834.900 182.850 ;
        RECT 835.950 181.950 840.450 183.450 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 800.550 176.550 804.450 177.450 ;
        RECT 806.100 177.150 807.900 178.950 ;
        RECT 790.950 174.450 793.050 174.750 ;
        RECT 799.950 174.450 802.050 175.050 ;
        RECT 790.950 173.550 802.050 174.450 ;
        RECT 790.950 172.650 793.050 173.550 ;
        RECT 799.950 172.950 802.050 173.550 ;
        RECT 784.950 171.450 787.050 172.050 ;
        RECT 803.550 171.450 804.450 176.550 ;
        RECT 784.950 170.550 804.450 171.450 ;
        RECT 784.950 169.950 787.050 170.550 ;
        RECT 783.000 165.900 789.600 166.800 ;
        RECT 783.000 165.600 783.900 165.900 ;
        RECT 740.100 159.000 741.900 165.600 ;
        RECT 743.100 159.600 744.900 165.600 ;
        RECT 746.100 159.000 747.900 165.600 ;
        RECT 761.100 159.000 762.900 165.600 ;
        RECT 764.100 159.600 765.900 165.600 ;
        RECT 767.100 159.000 768.900 165.600 ;
        RECT 782.100 159.600 783.900 165.600 ;
        RECT 788.100 165.600 789.600 165.900 ;
        RECT 809.100 165.600 810.300 178.950 ;
        RECT 824.100 177.150 825.900 178.950 ;
        RECT 830.700 171.600 831.900 178.950 ;
        RECT 839.550 178.050 840.450 181.950 ;
        RECT 848.100 181.050 849.900 182.850 ;
        RECT 851.100 181.050 852.300 185.400 ;
        RECT 864.000 183.450 868.050 184.050 ;
        RECT 854.100 181.050 855.900 182.850 ;
        RECT 863.550 181.950 868.050 183.450 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 856.950 178.950 859.050 181.050 ;
        RECT 835.950 176.550 840.450 178.050 ;
        RECT 835.950 175.950 840.000 176.550 ;
        RECT 785.100 159.000 786.900 165.000 ;
        RECT 788.100 159.600 789.900 165.600 ;
        RECT 791.100 159.000 792.900 165.600 ;
        RECT 806.100 159.000 807.900 165.600 ;
        RECT 809.100 159.600 810.900 165.600 ;
        RECT 824.400 159.000 826.200 171.600 ;
        RECT 829.500 170.100 831.900 171.600 ;
        RECT 851.100 171.600 852.300 178.950 ;
        RECT 857.100 177.150 858.900 178.950 ;
        RECT 863.550 177.450 864.450 181.950 ;
        RECT 869.100 181.050 870.900 182.850 ;
        RECT 872.100 181.050 873.300 185.400 ;
        RECT 885.000 183.450 889.050 184.050 ;
        RECT 875.100 181.050 876.900 182.850 ;
        RECT 884.550 181.950 889.050 183.450 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 860.550 176.550 864.450 177.450 ;
        RECT 853.950 174.450 856.050 175.050 ;
        RECT 860.550 174.450 861.450 176.550 ;
        RECT 853.950 173.550 861.450 174.450 ;
        RECT 853.950 172.950 856.050 173.550 ;
        RECT 872.100 171.600 873.300 178.950 ;
        RECT 878.100 177.150 879.900 178.950 ;
        RECT 884.550 178.050 885.450 181.950 ;
        RECT 890.400 181.050 891.300 188.400 ;
        RECT 911.100 187.950 918.900 189.300 ;
        RECT 920.100 188.400 921.900 194.400 ;
        RECT 920.100 186.300 921.300 188.400 ;
        RECT 917.700 185.400 921.300 186.300 ;
        RECT 892.950 181.050 894.750 182.850 ;
        RECT 899.100 181.050 900.900 182.850 ;
        RECT 914.100 181.050 915.900 182.850 ;
        RECT 917.700 181.050 918.900 185.400 ;
        RECT 920.100 181.050 921.900 182.850 ;
        RECT 889.950 178.950 892.050 181.050 ;
        RECT 892.950 178.950 895.050 181.050 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 913.950 178.950 916.050 181.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 884.550 176.550 889.050 178.050 ;
        RECT 885.000 175.950 889.050 176.550 ;
        RECT 890.400 171.600 891.300 178.950 ;
        RECT 895.950 177.150 897.750 178.950 ;
        RECT 911.100 177.150 912.900 178.950 ;
        RECT 917.700 171.600 918.900 178.950 ;
        RECT 851.100 170.100 853.500 171.600 ;
        RECT 829.500 159.600 831.300 170.100 ;
        RECT 832.200 167.100 834.000 168.900 ;
        RECT 849.000 167.100 850.800 168.900 ;
        RECT 832.500 159.000 834.300 165.600 ;
        RECT 848.700 159.000 850.500 165.600 ;
        RECT 851.700 159.600 853.500 170.100 ;
        RECT 856.800 159.000 858.600 171.600 ;
        RECT 872.100 170.100 874.500 171.600 ;
        RECT 870.000 167.100 871.800 168.900 ;
        RECT 869.700 159.000 871.500 165.600 ;
        RECT 872.700 159.600 874.500 170.100 ;
        RECT 877.800 159.000 879.600 171.600 ;
        RECT 890.100 159.600 891.900 171.600 ;
        RECT 893.100 170.700 900.900 171.600 ;
        RECT 893.100 159.600 894.900 170.700 ;
        RECT 896.100 159.000 897.900 169.800 ;
        RECT 899.100 159.600 900.900 170.700 ;
        RECT 911.400 159.000 913.200 171.600 ;
        RECT 916.500 170.100 918.900 171.600 ;
        RECT 916.500 159.600 918.300 170.100 ;
        RECT 919.200 167.100 921.000 168.900 ;
        RECT 919.500 159.000 921.300 165.600 ;
        RECT 14.400 143.400 16.200 156.000 ;
        RECT 19.500 144.900 21.300 155.400 ;
        RECT 22.500 149.400 24.300 156.000 ;
        RECT 35.100 149.400 36.900 156.000 ;
        RECT 38.100 149.400 39.900 155.400 ;
        RECT 41.100 149.400 42.900 156.000 ;
        RECT 53.700 149.400 55.500 156.000 ;
        RECT 22.200 146.100 24.000 147.900 ;
        RECT 19.500 143.400 21.900 144.900 ;
        RECT 14.100 136.050 15.900 137.850 ;
        RECT 20.700 136.050 21.900 143.400 ;
        RECT 38.700 136.050 39.900 149.400 ;
        RECT 54.000 146.100 55.800 147.900 ;
        RECT 56.700 144.900 58.500 155.400 ;
        RECT 56.100 143.400 58.500 144.900 ;
        RECT 61.800 143.400 63.600 156.000 ;
        RECT 74.400 143.400 76.200 156.000 ;
        RECT 79.500 144.900 81.300 155.400 ;
        RECT 82.500 149.400 84.300 156.000 ;
        RECT 98.100 149.400 99.900 156.000 ;
        RECT 101.100 149.400 102.900 155.400 ;
        RECT 104.100 150.000 105.900 156.000 ;
        RECT 101.400 149.100 102.900 149.400 ;
        RECT 107.100 149.400 108.900 155.400 ;
        RECT 107.100 149.100 108.000 149.400 ;
        RECT 101.400 148.200 108.000 149.100 ;
        RECT 82.200 146.100 84.000 147.900 ;
        RECT 79.500 143.400 81.900 144.900 ;
        RECT 43.950 138.450 48.000 139.050 ;
        RECT 43.950 136.950 48.450 138.450 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 17.100 132.150 18.900 133.950 ;
        RECT 20.700 129.600 21.900 133.950 ;
        RECT 23.100 132.150 24.900 133.950 ;
        RECT 35.100 132.150 36.900 133.950 ;
        RECT 20.700 128.700 24.300 129.600 ;
        RECT 38.700 128.700 39.900 133.950 ;
        RECT 40.950 132.150 42.750 133.950 ;
        RECT 47.550 133.050 48.450 136.950 ;
        RECT 56.100 136.050 57.300 143.400 ;
        RECT 64.950 138.450 69.000 139.050 ;
        RECT 62.100 136.050 63.900 137.850 ;
        RECT 64.950 136.950 69.450 138.450 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 47.550 131.550 52.050 133.050 ;
        RECT 53.100 132.150 54.900 133.950 ;
        RECT 48.000 130.950 52.050 131.550 ;
        RECT 56.100 129.600 57.300 133.950 ;
        RECT 59.100 132.150 60.900 133.950 ;
        RECT 68.550 133.050 69.450 136.950 ;
        RECT 74.100 136.050 75.900 137.850 ;
        RECT 80.700 136.050 81.900 143.400 ;
        RECT 101.100 136.050 102.900 137.850 ;
        RECT 107.100 136.050 108.000 148.200 ;
        RECT 122.100 143.400 123.900 155.400 ;
        RECT 125.100 144.300 126.900 155.400 ;
        RECT 128.100 145.200 129.900 156.000 ;
        RECT 131.100 144.300 132.900 155.400 ;
        RECT 125.100 143.400 132.900 144.300 ;
        RECT 143.100 143.400 144.900 155.400 ;
        RECT 146.100 144.300 147.900 155.400 ;
        RECT 149.100 145.200 150.900 156.000 ;
        RECT 152.100 144.300 153.900 155.400 ;
        RECT 146.100 143.400 153.900 144.300 ;
        RECT 167.100 144.600 168.900 155.400 ;
        RECT 170.100 145.500 171.900 156.000 ;
        RECT 167.100 143.400 171.900 144.600 ;
        RECT 109.950 138.450 114.000 139.050 ;
        RECT 109.950 136.950 114.450 138.450 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 64.950 131.550 69.450 133.050 ;
        RECT 77.100 132.150 78.900 133.950 ;
        RECT 64.950 130.950 69.000 131.550 ;
        RECT 14.100 125.700 21.900 127.050 ;
        RECT 14.100 120.600 15.900 125.700 ;
        RECT 17.100 120.000 18.900 124.800 ;
        RECT 20.100 120.600 21.900 125.700 ;
        RECT 23.100 126.600 24.300 128.700 ;
        RECT 35.700 127.800 39.900 128.700 ;
        RECT 53.700 128.700 57.300 129.600 ;
        RECT 80.700 129.600 81.900 133.950 ;
        RECT 83.100 132.150 84.900 133.950 ;
        RECT 98.100 132.150 99.900 133.950 ;
        RECT 104.100 132.150 105.900 133.950 ;
        RECT 107.100 130.200 108.000 133.950 ;
        RECT 113.550 132.450 114.450 136.950 ;
        RECT 122.400 136.050 123.300 143.400 ;
        RECT 127.950 136.050 129.750 137.850 ;
        RECT 143.400 136.050 144.300 143.400 ;
        RECT 169.800 142.500 171.900 143.400 ;
        RECT 174.600 143.400 176.400 155.400 ;
        RECT 179.100 145.500 180.900 156.000 ;
        RECT 182.100 144.300 183.900 155.400 ;
        RECT 194.700 149.400 196.500 156.000 ;
        RECT 195.000 146.100 196.800 147.900 ;
        RECT 197.700 144.900 199.500 155.400 ;
        RECT 179.400 143.400 183.900 144.300 ;
        RECT 197.100 143.400 199.500 144.900 ;
        RECT 202.800 143.400 204.600 156.000 ;
        RECT 215.100 149.400 216.900 156.000 ;
        RECT 218.100 149.400 219.900 155.400 ;
        RECT 233.100 149.400 234.900 155.400 ;
        RECT 236.100 150.000 237.900 156.000 ;
        RECT 174.600 142.050 175.800 143.400 ;
        RECT 174.300 141.000 175.800 142.050 ;
        RECT 179.400 141.300 181.500 143.400 ;
        RECT 174.300 139.050 175.200 141.000 ;
        RECT 148.950 136.050 150.750 137.850 ;
        RECT 167.400 136.050 169.200 137.850 ;
        RECT 173.100 136.950 175.200 139.050 ;
        RECT 176.100 139.500 178.200 139.800 ;
        RECT 176.100 137.700 180.000 139.500 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 167.100 133.950 169.200 136.050 ;
        RECT 173.700 136.800 175.200 136.950 ;
        RECT 173.700 135.900 176.100 136.800 ;
        RECT 118.950 132.450 121.050 133.050 ;
        RECT 113.550 131.550 121.050 132.450 ;
        RECT 118.950 130.950 121.050 131.550 ;
        RECT 80.700 128.700 84.300 129.600 ;
        RECT 23.100 120.600 24.900 126.600 ;
        RECT 35.700 120.600 37.500 127.800 ;
        RECT 53.700 126.600 54.900 128.700 ;
        RECT 40.800 120.000 42.600 126.600 ;
        RECT 53.100 120.600 54.900 126.600 ;
        RECT 56.100 125.700 63.900 127.050 ;
        RECT 56.100 120.600 57.900 125.700 ;
        RECT 59.100 120.000 60.900 124.800 ;
        RECT 62.100 120.600 63.900 125.700 ;
        RECT 74.100 125.700 81.900 127.050 ;
        RECT 74.100 120.600 75.900 125.700 ;
        RECT 77.100 120.000 78.900 124.800 ;
        RECT 80.100 120.600 81.900 125.700 ;
        RECT 83.100 126.600 84.300 128.700 ;
        RECT 83.100 120.600 84.900 126.600 ;
        RECT 98.100 120.000 99.900 129.600 ;
        RECT 104.700 129.000 108.000 130.200 ;
        RECT 104.700 120.600 106.500 129.000 ;
        RECT 122.400 126.600 123.300 133.950 ;
        RECT 124.950 132.150 126.750 133.950 ;
        RECT 131.100 132.150 132.900 133.950 ;
        RECT 143.400 126.600 144.300 133.950 ;
        RECT 145.950 132.150 147.750 133.950 ;
        RECT 152.100 132.150 153.900 133.950 ;
        RECT 171.900 133.200 173.700 135.000 ;
        RECT 171.900 131.100 174.000 133.200 ;
        RECT 174.900 130.200 176.100 135.900 ;
        RECT 177.000 136.050 178.800 136.500 ;
        RECT 197.100 136.050 198.300 143.400 ;
        RECT 203.100 136.050 204.900 137.850 ;
        RECT 215.100 136.050 216.900 137.850 ;
        RECT 218.100 136.050 219.300 149.400 ;
        RECT 234.000 149.100 234.900 149.400 ;
        RECT 239.100 149.400 240.900 155.400 ;
        RECT 242.100 149.400 243.900 156.000 ;
        RECT 257.100 149.400 258.900 155.400 ;
        RECT 260.100 149.400 261.900 156.000 ;
        RECT 239.100 149.100 240.600 149.400 ;
        RECT 234.000 148.200 240.600 149.100 ;
        RECT 234.000 136.050 234.900 148.200 ;
        RECT 239.100 136.050 240.900 137.850 ;
        RECT 257.700 136.050 258.900 149.400 ;
        RECT 272.100 144.600 273.900 155.400 ;
        RECT 275.100 145.500 276.900 156.000 ;
        RECT 278.100 154.500 285.900 155.400 ;
        RECT 278.100 144.600 279.900 154.500 ;
        RECT 272.100 143.700 279.900 144.600 ;
        RECT 281.100 142.500 282.900 153.600 ;
        RECT 284.100 143.400 285.900 154.500 ;
        RECT 296.100 144.300 297.900 155.400 ;
        RECT 299.100 145.200 300.900 156.000 ;
        RECT 302.100 144.300 303.900 155.400 ;
        RECT 296.100 143.400 303.900 144.300 ;
        RECT 305.100 143.400 306.900 155.400 ;
        RECT 320.100 143.400 321.900 156.000 ;
        RECT 325.200 144.600 327.000 155.400 ;
        RECT 341.700 149.400 343.500 156.000 ;
        RECT 342.000 146.100 343.800 147.900 ;
        RECT 344.700 144.900 346.500 155.400 ;
        RECT 323.400 143.400 327.000 144.600 ;
        RECT 344.100 143.400 346.500 144.900 ;
        RECT 349.800 143.400 351.600 156.000 ;
        RECT 362.100 149.400 363.900 156.000 ;
        RECT 365.100 149.400 366.900 155.400 ;
        RECT 377.100 149.400 378.900 156.000 ;
        RECT 380.100 149.400 381.900 155.400 ;
        RECT 383.100 149.400 384.900 156.000 ;
        RECT 398.100 149.400 399.900 156.000 ;
        RECT 401.100 149.400 402.900 155.400 ;
        RECT 404.100 149.400 405.900 156.000 ;
        RECT 278.100 141.600 282.900 142.500 ;
        RECT 260.100 136.050 261.900 137.850 ;
        RECT 275.250 136.050 277.050 137.850 ;
        RECT 278.100 136.050 279.000 141.600 ;
        RECT 281.100 136.050 282.900 137.850 ;
        RECT 299.250 136.050 301.050 137.850 ;
        RECT 305.700 136.050 306.600 143.400 ;
        RECT 320.250 136.050 322.050 137.850 ;
        RECT 323.400 136.050 324.300 143.400 ;
        RECT 326.100 136.050 327.900 137.850 ;
        RECT 344.100 136.050 345.300 143.400 ;
        RECT 350.100 136.050 351.900 137.850 ;
        RECT 362.100 136.050 363.900 137.850 ;
        RECT 365.100 136.050 366.300 149.400 ;
        RECT 380.100 136.050 381.300 149.400 ;
        RECT 401.100 136.050 402.300 149.400 ;
        RECT 419.100 143.400 420.900 155.400 ;
        RECT 422.100 144.300 423.900 155.400 ;
        RECT 425.100 145.200 426.900 156.000 ;
        RECT 428.100 144.300 429.900 155.400 ;
        RECT 444.600 144.900 446.400 155.400 ;
        RECT 422.100 143.400 429.900 144.300 ;
        RECT 444.000 143.400 446.400 144.900 ;
        RECT 447.600 143.400 449.400 156.000 ;
        RECT 452.100 143.400 453.900 155.400 ;
        RECT 467.100 143.400 468.900 155.400 ;
        RECT 470.100 144.300 471.900 155.400 ;
        RECT 473.100 145.200 474.900 156.000 ;
        RECT 476.100 144.300 477.900 155.400 ;
        RECT 470.100 143.400 477.900 144.300 ;
        RECT 488.100 144.300 489.900 155.400 ;
        RECT 491.100 145.500 492.900 156.000 ;
        RECT 488.100 143.400 492.600 144.300 ;
        RECT 495.600 143.400 497.400 155.400 ;
        RECT 500.100 145.500 501.900 156.000 ;
        RECT 503.100 144.600 504.900 155.400 ;
        RECT 419.400 136.050 420.300 143.400 ;
        RECT 427.950 141.450 430.050 142.050 ;
        RECT 439.950 141.450 442.050 142.050 ;
        RECT 427.950 140.550 442.050 141.450 ;
        RECT 427.950 139.950 430.050 140.550 ;
        RECT 439.950 139.950 442.050 140.550 ;
        RECT 424.950 136.050 426.750 137.850 ;
        RECT 444.000 136.050 445.200 143.400 ;
        RECT 452.700 141.900 453.900 143.400 ;
        RECT 446.100 140.700 453.900 141.900 ;
        RECT 446.100 140.100 447.900 140.700 ;
        RECT 177.000 134.700 183.900 136.050 ;
        RECT 181.800 133.950 183.900 134.700 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 232.950 133.950 235.050 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 325.950 133.950 328.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 343.950 133.950 346.050 136.050 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 397.950 133.950 400.050 136.050 ;
        RECT 400.950 133.950 403.050 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 424.950 133.950 427.050 136.050 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 443.100 133.950 445.200 136.050 ;
        RECT 169.800 127.500 171.900 128.700 ;
        RECT 173.100 128.100 176.100 130.200 ;
        RECT 177.000 131.400 178.800 133.200 ;
        RECT 181.800 132.150 183.600 133.950 ;
        RECT 194.100 132.150 195.900 133.950 ;
        RECT 177.000 129.300 179.100 131.400 ;
        RECT 197.100 129.600 198.300 133.950 ;
        RECT 200.100 132.150 201.900 133.950 ;
        RECT 177.000 128.400 183.300 129.300 ;
        RECT 167.100 126.600 171.900 127.500 ;
        RECT 174.900 126.600 176.100 128.100 ;
        RECT 182.100 126.600 183.300 128.400 ;
        RECT 194.700 128.700 198.300 129.600 ;
        RECT 194.700 126.600 195.900 128.700 ;
        RECT 122.400 125.400 127.500 126.600 ;
        RECT 122.700 120.000 124.500 123.600 ;
        RECT 125.700 120.600 127.500 125.400 ;
        RECT 130.200 120.000 132.000 126.600 ;
        RECT 143.400 125.400 148.500 126.600 ;
        RECT 143.700 120.000 145.500 123.600 ;
        RECT 146.700 120.600 148.500 125.400 ;
        RECT 151.200 120.000 153.000 126.600 ;
        RECT 167.100 120.600 168.900 126.600 ;
        RECT 170.100 120.000 171.900 125.700 ;
        RECT 174.600 120.600 176.400 126.600 ;
        RECT 179.100 120.000 180.900 125.700 ;
        RECT 182.100 120.600 183.900 126.600 ;
        RECT 194.100 120.600 195.900 126.600 ;
        RECT 197.100 125.700 204.900 127.050 ;
        RECT 197.100 120.600 198.900 125.700 ;
        RECT 200.100 120.000 201.900 124.800 ;
        RECT 203.100 120.600 204.900 125.700 ;
        RECT 218.100 123.600 219.300 133.950 ;
        RECT 234.000 130.200 234.900 133.950 ;
        RECT 236.100 132.150 237.900 133.950 ;
        RECT 242.100 132.150 243.900 133.950 ;
        RECT 234.000 129.000 237.300 130.200 ;
        RECT 215.100 120.000 216.900 123.600 ;
        RECT 218.100 120.600 219.900 123.600 ;
        RECT 235.500 120.600 237.300 129.000 ;
        RECT 242.100 120.000 243.900 129.600 ;
        RECT 257.700 123.600 258.900 133.950 ;
        RECT 272.250 132.150 274.050 133.950 ;
        RECT 278.100 126.600 279.300 133.950 ;
        RECT 284.100 132.150 285.900 133.950 ;
        RECT 296.100 132.150 297.900 133.950 ;
        RECT 302.250 132.150 304.050 133.950 ;
        RECT 305.700 126.600 306.600 133.950 ;
        RECT 257.100 120.600 258.900 123.600 ;
        RECT 260.100 120.000 261.900 123.600 ;
        RECT 272.700 120.000 274.500 126.600 ;
        RECT 277.200 120.600 279.000 126.600 ;
        RECT 281.700 120.000 283.500 126.600 ;
        RECT 297.000 120.000 298.800 126.600 ;
        RECT 301.500 125.400 306.600 126.600 ;
        RECT 301.500 120.600 303.300 125.400 ;
        RECT 323.400 123.600 324.300 133.950 ;
        RECT 341.100 132.150 342.900 133.950 ;
        RECT 344.100 129.600 345.300 133.950 ;
        RECT 347.100 132.150 348.900 133.950 ;
        RECT 341.700 128.700 345.300 129.600 ;
        RECT 341.700 126.600 342.900 128.700 ;
        RECT 304.500 120.000 306.300 123.600 ;
        RECT 320.100 120.000 321.900 123.600 ;
        RECT 323.100 120.600 324.900 123.600 ;
        RECT 326.100 120.000 327.900 123.600 ;
        RECT 341.100 120.600 342.900 126.600 ;
        RECT 344.100 125.700 351.900 127.050 ;
        RECT 344.100 120.600 345.900 125.700 ;
        RECT 347.100 120.000 348.900 124.800 ;
        RECT 350.100 120.600 351.900 125.700 ;
        RECT 365.100 123.600 366.300 133.950 ;
        RECT 377.250 132.150 379.050 133.950 ;
        RECT 380.100 128.700 381.300 133.950 ;
        RECT 383.100 132.150 384.900 133.950 ;
        RECT 398.250 132.150 400.050 133.950 ;
        RECT 401.100 128.700 402.300 133.950 ;
        RECT 404.100 132.150 405.900 133.950 ;
        RECT 380.100 127.800 384.300 128.700 ;
        RECT 401.100 127.800 405.300 128.700 ;
        RECT 362.100 120.000 363.900 123.600 ;
        RECT 365.100 120.600 366.900 123.600 ;
        RECT 377.400 120.000 379.200 126.600 ;
        RECT 382.500 120.600 384.300 127.800 ;
        RECT 398.400 120.000 400.200 126.600 ;
        RECT 403.500 120.600 405.300 127.800 ;
        RECT 419.400 126.600 420.300 133.950 ;
        RECT 421.950 132.150 423.750 133.950 ;
        RECT 428.100 132.150 429.900 133.950 ;
        RECT 443.100 126.600 444.000 133.950 ;
        RECT 446.400 129.600 447.300 140.100 ;
        RECT 448.200 136.050 450.000 137.850 ;
        RECT 467.400 136.050 468.300 143.400 ;
        RECT 490.500 141.300 492.600 143.400 ;
        RECT 496.200 142.050 497.400 143.400 ;
        RECT 500.100 143.400 504.900 144.600 ;
        RECT 515.400 143.400 517.200 156.000 ;
        RECT 520.500 144.900 522.300 155.400 ;
        RECT 523.500 149.400 525.300 156.000 ;
        RECT 523.200 146.100 525.000 147.900 ;
        RECT 520.500 143.400 522.900 144.900 ;
        RECT 500.100 142.500 502.200 143.400 ;
        RECT 496.200 141.000 497.700 142.050 ;
        RECT 493.800 139.500 495.900 139.800 ;
        RECT 472.950 136.050 474.750 137.850 ;
        RECT 492.000 137.700 495.900 139.500 ;
        RECT 496.800 139.050 497.700 141.000 ;
        RECT 496.800 136.950 498.900 139.050 ;
        RECT 496.800 136.800 498.300 136.950 ;
        RECT 493.200 136.050 495.000 136.500 ;
        RECT 448.500 133.950 450.600 136.050 ;
        RECT 451.800 133.950 453.900 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 488.100 134.700 495.000 136.050 ;
        RECT 495.900 135.900 498.300 136.800 ;
        RECT 502.800 136.050 504.600 137.850 ;
        RECT 515.100 136.050 516.900 137.850 ;
        RECT 521.700 136.050 522.900 143.400 ;
        RECT 536.100 144.300 537.900 155.400 ;
        RECT 539.100 145.500 540.900 156.000 ;
        RECT 543.600 144.300 545.400 155.400 ;
        RECT 547.800 145.500 549.900 156.000 ;
        RECT 551.100 144.600 552.900 155.400 ;
        RECT 536.100 143.100 540.900 144.300 ;
        RECT 543.600 143.400 546.900 144.300 ;
        RECT 538.800 142.200 540.900 143.100 ;
        RECT 538.800 141.300 544.200 142.200 ;
        RECT 542.400 139.500 544.200 141.300 ;
        RECT 545.700 139.050 546.900 143.400 ;
        RECT 547.800 143.400 552.900 144.600 ;
        RECT 563.100 143.400 564.900 155.400 ;
        RECT 566.100 144.300 567.900 155.400 ;
        RECT 569.100 145.200 570.900 156.000 ;
        RECT 572.100 144.300 573.900 155.400 ;
        RECT 584.100 149.400 585.900 156.000 ;
        RECT 587.100 149.400 588.900 155.400 ;
        RECT 590.100 149.400 591.900 156.000 ;
        RECT 602.100 149.400 603.900 156.000 ;
        RECT 605.100 149.400 606.900 155.400 ;
        RECT 608.100 150.000 609.900 156.000 ;
        RECT 566.100 143.400 573.900 144.300 ;
        RECT 547.800 142.500 549.900 143.400 ;
        RECT 545.100 138.300 547.200 139.050 ;
        RECT 540.900 136.200 542.700 138.000 ;
        RECT 544.200 136.950 547.200 138.300 ;
        RECT 488.100 133.950 490.200 134.700 ;
        RECT 451.800 132.150 453.600 133.950 ;
        RECT 445.200 128.700 447.300 129.600 ;
        RECT 445.200 127.800 450.600 128.700 ;
        RECT 419.400 125.400 424.500 126.600 ;
        RECT 419.700 120.000 421.500 123.600 ;
        RECT 422.700 120.600 424.500 125.400 ;
        RECT 427.200 120.000 429.000 126.600 ;
        RECT 443.100 120.600 444.900 126.600 ;
        RECT 446.100 120.000 447.900 126.000 ;
        RECT 449.700 123.600 450.600 127.800 ;
        RECT 467.400 126.600 468.300 133.950 ;
        RECT 469.950 132.150 471.750 133.950 ;
        RECT 476.100 132.150 477.900 133.950 ;
        RECT 488.400 132.150 490.200 133.950 ;
        RECT 493.200 131.400 495.000 133.200 ;
        RECT 492.900 129.300 495.000 131.400 ;
        RECT 488.700 128.400 495.000 129.300 ;
        RECT 495.900 130.200 497.100 135.900 ;
        RECT 498.300 133.200 500.100 135.000 ;
        RECT 502.800 133.950 504.900 136.050 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 498.000 131.100 500.100 133.200 ;
        RECT 518.100 132.150 519.900 133.950 ;
        RECT 488.700 126.600 489.900 128.400 ;
        RECT 495.900 128.100 498.900 130.200 ;
        RECT 521.700 129.600 522.900 133.950 ;
        RECT 524.100 132.150 525.900 133.950 ;
        RECT 536.100 133.800 538.200 136.050 ;
        RECT 540.900 134.100 543.000 136.200 ;
        RECT 536.400 133.200 538.200 133.800 ;
        RECT 536.400 132.000 543.000 133.200 ;
        RECT 540.900 131.100 543.000 132.000 ;
        RECT 521.700 128.700 525.300 129.600 ;
        RECT 538.500 129.000 540.600 129.600 ;
        RECT 541.500 129.300 543.300 131.100 ;
        RECT 544.200 130.200 545.100 136.950 ;
        RECT 550.800 136.050 552.600 137.850 ;
        RECT 563.400 136.050 564.300 143.400 ;
        RECT 568.950 136.050 570.750 137.850 ;
        RECT 587.100 136.050 588.300 149.400 ;
        RECT 605.400 149.100 606.900 149.400 ;
        RECT 611.100 149.400 612.900 155.400 ;
        RECT 611.100 149.100 612.000 149.400 ;
        RECT 605.400 148.200 612.000 149.100 ;
        RECT 605.100 136.050 606.900 137.850 ;
        RECT 611.100 136.050 612.000 148.200 ;
        RECT 623.100 143.400 624.900 155.400 ;
        RECT 626.100 144.300 627.900 155.400 ;
        RECT 629.100 145.200 630.900 156.000 ;
        RECT 632.100 144.300 633.900 155.400 ;
        RECT 647.100 149.400 648.900 155.400 ;
        RECT 650.100 150.000 651.900 156.000 ;
        RECT 626.100 143.400 633.900 144.300 ;
        RECT 648.000 149.100 648.900 149.400 ;
        RECT 653.100 149.400 654.900 155.400 ;
        RECT 656.100 149.400 657.900 156.000 ;
        RECT 653.100 149.100 654.600 149.400 ;
        RECT 648.000 148.200 654.600 149.100 ;
        RECT 623.400 136.050 624.300 143.400 ;
        RECT 625.950 141.450 628.050 142.050 ;
        RECT 634.950 141.450 637.050 142.050 ;
        RECT 625.950 140.550 637.050 141.450 ;
        RECT 625.950 139.950 628.050 140.550 ;
        RECT 634.950 139.950 637.050 140.550 ;
        RECT 628.950 136.050 630.750 137.850 ;
        RECT 648.000 136.050 648.900 148.200 ;
        RECT 671.100 143.400 672.900 156.000 ;
        RECT 676.200 144.600 678.000 155.400 ;
        RECT 689.100 149.400 690.900 156.000 ;
        RECT 692.100 149.400 693.900 155.400 ;
        RECT 695.100 149.400 696.900 156.000 ;
        RECT 707.100 149.400 708.900 156.000 ;
        RECT 710.100 149.400 711.900 155.400 ;
        RECT 713.100 149.400 714.900 156.000 ;
        RECT 674.400 143.400 678.000 144.600 ;
        RECT 653.100 136.050 654.900 137.850 ;
        RECT 671.250 136.050 673.050 137.850 ;
        RECT 674.400 136.050 675.300 143.400 ;
        RECT 684.000 138.450 688.050 139.050 ;
        RECT 677.100 136.050 678.900 137.850 ;
        RECT 683.550 136.950 688.050 138.450 ;
        RECT 546.000 134.100 547.800 135.900 ;
        RECT 546.000 132.000 548.100 134.100 ;
        RECT 550.800 133.950 552.900 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 631.950 133.950 634.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 655.950 133.950 658.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 495.900 126.600 497.100 128.100 ;
        RECT 500.100 127.500 502.200 128.700 ;
        RECT 500.100 126.600 504.900 127.500 ;
        RECT 467.400 125.400 472.500 126.600 ;
        RECT 449.100 120.600 450.900 123.600 ;
        RECT 452.100 120.600 453.900 123.600 ;
        RECT 452.700 120.000 453.900 120.600 ;
        RECT 467.700 120.000 469.500 123.600 ;
        RECT 470.700 120.600 472.500 125.400 ;
        RECT 475.200 120.000 477.000 126.600 ;
        RECT 488.100 120.600 489.900 126.600 ;
        RECT 491.100 120.000 492.900 125.700 ;
        RECT 495.600 120.600 497.400 126.600 ;
        RECT 500.100 120.000 501.900 125.700 ;
        RECT 503.100 120.600 504.900 126.600 ;
        RECT 515.100 125.700 522.900 127.050 ;
        RECT 515.100 120.600 516.900 125.700 ;
        RECT 518.100 120.000 519.900 124.800 ;
        RECT 521.100 120.600 522.900 125.700 ;
        RECT 524.100 126.600 525.300 128.700 ;
        RECT 536.100 127.500 540.600 129.000 ;
        RECT 544.200 128.100 547.200 130.200 ;
        RECT 536.100 126.600 537.600 127.500 ;
        RECT 524.100 120.600 525.900 126.600 ;
        RECT 536.100 120.600 537.900 126.600 ;
        RECT 544.200 126.000 545.100 128.100 ;
        RECT 548.400 127.500 550.500 129.900 ;
        RECT 548.400 126.600 552.900 127.500 ;
        RECT 539.100 120.000 540.900 125.700 ;
        RECT 543.300 120.600 545.100 126.000 ;
        RECT 547.800 120.000 549.600 125.700 ;
        RECT 551.100 120.600 552.900 126.600 ;
        RECT 563.400 126.600 564.300 133.950 ;
        RECT 565.950 132.150 567.750 133.950 ;
        RECT 572.100 132.150 573.900 133.950 ;
        RECT 584.250 132.150 586.050 133.950 ;
        RECT 587.100 128.700 588.300 133.950 ;
        RECT 590.100 132.150 591.900 133.950 ;
        RECT 602.100 132.150 603.900 133.950 ;
        RECT 608.100 132.150 609.900 133.950 ;
        RECT 611.100 130.200 612.000 133.950 ;
        RECT 587.100 127.800 591.300 128.700 ;
        RECT 563.400 125.400 568.500 126.600 ;
        RECT 563.700 120.000 565.500 123.600 ;
        RECT 566.700 120.600 568.500 125.400 ;
        RECT 571.200 120.000 573.000 126.600 ;
        RECT 584.400 120.000 586.200 126.600 ;
        RECT 589.500 120.600 591.300 127.800 ;
        RECT 602.100 120.000 603.900 129.600 ;
        RECT 608.700 129.000 612.000 130.200 ;
        RECT 608.700 120.600 610.500 129.000 ;
        RECT 623.400 126.600 624.300 133.950 ;
        RECT 625.950 132.150 627.750 133.950 ;
        RECT 632.100 132.150 633.900 133.950 ;
        RECT 648.000 130.200 648.900 133.950 ;
        RECT 650.100 132.150 651.900 133.950 ;
        RECT 656.100 132.150 657.900 133.950 ;
        RECT 648.000 129.000 651.300 130.200 ;
        RECT 623.400 125.400 628.500 126.600 ;
        RECT 623.700 120.000 625.500 123.600 ;
        RECT 626.700 120.600 628.500 125.400 ;
        RECT 631.200 120.000 633.000 126.600 ;
        RECT 649.500 120.600 651.300 129.000 ;
        RECT 656.100 120.000 657.900 129.600 ;
        RECT 674.400 123.600 675.300 133.950 ;
        RECT 683.550 133.050 684.450 136.950 ;
        RECT 692.700 136.050 693.900 149.400 ;
        RECT 710.700 136.050 711.900 149.400 ;
        RECT 728.100 143.400 729.900 155.400 ;
        RECT 731.100 144.300 732.900 155.400 ;
        RECT 734.100 145.200 735.900 156.000 ;
        RECT 737.100 144.300 738.900 155.400 ;
        RECT 752.100 149.400 753.900 156.000 ;
        RECT 755.100 149.400 756.900 155.400 ;
        RECT 758.100 150.000 759.900 156.000 ;
        RECT 755.400 149.100 756.900 149.400 ;
        RECT 761.100 149.400 762.900 155.400 ;
        RECT 761.100 149.100 762.000 149.400 ;
        RECT 755.400 148.200 762.000 149.100 ;
        RECT 731.100 143.400 738.900 144.300 ;
        RECT 712.950 141.450 715.050 142.200 ;
        RECT 721.950 141.450 724.050 142.050 ;
        RECT 712.950 140.550 724.050 141.450 ;
        RECT 712.950 140.100 715.050 140.550 ;
        RECT 721.950 139.950 724.050 140.550 ;
        RECT 728.400 136.050 729.300 143.400 ;
        RECT 736.950 141.450 739.050 142.050 ;
        RECT 751.950 141.450 754.050 142.200 ;
        RECT 757.950 141.450 760.050 142.050 ;
        RECT 736.950 140.550 760.050 141.450 ;
        RECT 736.950 139.950 739.050 140.550 ;
        RECT 751.950 140.100 754.050 140.550 ;
        RECT 757.950 139.950 760.050 140.550 ;
        RECT 733.950 136.050 735.750 137.850 ;
        RECT 755.100 136.050 756.900 137.850 ;
        RECT 761.100 136.050 762.000 148.200 ;
        RECT 773.100 144.300 774.900 155.400 ;
        RECT 776.100 145.200 777.900 156.000 ;
        RECT 779.100 144.300 780.900 155.400 ;
        RECT 773.100 143.400 780.900 144.300 ;
        RECT 782.100 143.400 783.900 155.400 ;
        RECT 794.100 149.400 795.900 155.400 ;
        RECT 797.100 150.000 798.900 156.000 ;
        RECT 795.000 149.100 795.900 149.400 ;
        RECT 800.100 149.400 801.900 155.400 ;
        RECT 803.100 149.400 804.900 156.000 ;
        RECT 815.100 149.400 816.900 156.000 ;
        RECT 818.100 149.400 819.900 155.400 ;
        RECT 821.100 150.000 822.900 156.000 ;
        RECT 800.100 149.100 801.600 149.400 ;
        RECT 795.000 148.200 801.600 149.100 ;
        RECT 818.400 149.100 819.900 149.400 ;
        RECT 824.100 149.400 825.900 155.400 ;
        RECT 824.100 149.100 825.000 149.400 ;
        RECT 818.400 148.200 825.000 149.100 ;
        RECT 766.950 141.450 769.050 142.050 ;
        RECT 775.950 141.450 778.050 142.050 ;
        RECT 766.950 140.550 778.050 141.450 ;
        RECT 766.950 139.950 769.050 140.550 ;
        RECT 775.950 139.950 778.050 140.550 ;
        RECT 776.250 136.050 778.050 137.850 ;
        RECT 782.700 136.050 783.600 143.400 ;
        RECT 795.000 136.050 795.900 148.200 ;
        RECT 796.950 141.450 799.050 142.050 ;
        RECT 808.950 141.450 811.050 141.900 ;
        RECT 814.950 141.450 817.050 142.200 ;
        RECT 796.950 140.550 817.050 141.450 ;
        RECT 796.950 139.950 799.050 140.550 ;
        RECT 808.950 139.800 811.050 140.550 ;
        RECT 814.950 140.100 817.050 140.550 ;
        RECT 800.100 136.050 801.900 137.850 ;
        RECT 818.100 136.050 819.900 137.850 ;
        RECT 824.100 136.050 825.000 148.200 ;
        RECT 836.100 143.400 837.900 155.400 ;
        RECT 839.100 144.300 840.900 155.400 ;
        RECT 842.100 145.200 843.900 156.000 ;
        RECT 845.100 144.300 846.900 155.400 ;
        RECT 860.100 149.400 861.900 155.400 ;
        RECT 863.100 150.000 864.900 156.000 ;
        RECT 839.100 143.400 846.900 144.300 ;
        RECT 861.000 149.100 861.900 149.400 ;
        RECT 866.100 149.400 867.900 155.400 ;
        RECT 869.100 149.400 870.900 156.000 ;
        RECT 881.100 149.400 882.900 155.400 ;
        RECT 884.100 150.000 885.900 156.000 ;
        RECT 866.100 149.100 867.600 149.400 ;
        RECT 861.000 148.200 867.600 149.100 ;
        RECT 882.000 149.100 882.900 149.400 ;
        RECT 887.100 149.400 888.900 155.400 ;
        RECT 890.100 149.400 891.900 156.000 ;
        RECT 887.100 149.100 888.600 149.400 ;
        RECT 882.000 148.200 888.600 149.100 ;
        RECT 826.950 138.450 831.000 139.050 ;
        RECT 826.950 136.950 831.450 138.450 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 709.950 133.950 712.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 760.950 133.950 763.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 781.950 133.950 784.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 679.950 131.550 684.450 133.050 ;
        RECT 689.100 132.150 690.900 133.950 ;
        RECT 679.950 130.950 684.000 131.550 ;
        RECT 692.700 128.700 693.900 133.950 ;
        RECT 694.950 132.150 696.750 133.950 ;
        RECT 707.100 132.150 708.900 133.950 ;
        RECT 710.700 128.700 711.900 133.950 ;
        RECT 712.950 132.150 714.750 133.950 ;
        RECT 689.700 127.800 693.900 128.700 ;
        RECT 707.700 127.800 711.900 128.700 ;
        RECT 671.100 120.000 672.900 123.600 ;
        RECT 674.100 120.600 675.900 123.600 ;
        RECT 677.100 120.000 678.900 123.600 ;
        RECT 689.700 120.600 691.500 127.800 ;
        RECT 694.800 120.000 696.600 126.600 ;
        RECT 707.700 120.600 709.500 127.800 ;
        RECT 728.400 126.600 729.300 133.950 ;
        RECT 730.950 132.150 732.750 133.950 ;
        RECT 737.100 132.150 738.900 133.950 ;
        RECT 742.950 132.450 745.050 133.050 ;
        RECT 742.950 132.000 750.450 132.450 ;
        RECT 752.100 132.150 753.900 133.950 ;
        RECT 758.100 132.150 759.900 133.950 ;
        RECT 742.950 131.550 751.050 132.000 ;
        RECT 742.950 130.950 745.050 131.550 ;
        RECT 748.950 127.950 751.050 131.550 ;
        RECT 761.100 130.200 762.000 133.950 ;
        RECT 773.100 132.150 774.900 133.950 ;
        RECT 779.250 132.150 781.050 133.950 ;
        RECT 712.800 120.000 714.600 126.600 ;
        RECT 728.400 125.400 733.500 126.600 ;
        RECT 728.700 120.000 730.500 123.600 ;
        RECT 731.700 120.600 733.500 125.400 ;
        RECT 736.200 120.000 738.000 126.600 ;
        RECT 752.100 120.000 753.900 129.600 ;
        RECT 758.700 129.000 762.000 130.200 ;
        RECT 758.700 120.600 760.500 129.000 ;
        RECT 782.700 126.600 783.600 133.950 ;
        RECT 795.000 130.200 795.900 133.950 ;
        RECT 797.100 132.150 798.900 133.950 ;
        RECT 803.100 132.150 804.900 133.950 ;
        RECT 815.100 132.150 816.900 133.950 ;
        RECT 821.100 132.150 822.900 133.950 ;
        RECT 824.100 130.200 825.000 133.950 ;
        RECT 830.550 133.050 831.450 136.950 ;
        RECT 836.400 136.050 837.300 143.400 ;
        RECT 841.950 136.050 843.750 137.850 ;
        RECT 861.000 136.050 861.900 148.200 ;
        RECT 871.950 138.450 876.000 139.050 ;
        RECT 866.100 136.050 867.900 137.850 ;
        RECT 871.950 136.950 876.450 138.450 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 844.950 133.950 847.050 136.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 868.950 133.950 871.050 136.050 ;
        RECT 830.550 131.550 835.050 133.050 ;
        RECT 831.000 130.950 835.050 131.550 ;
        RECT 795.000 129.000 798.300 130.200 ;
        RECT 774.000 120.000 775.800 126.600 ;
        RECT 778.500 125.400 783.600 126.600 ;
        RECT 778.500 120.600 780.300 125.400 ;
        RECT 781.500 120.000 783.300 123.600 ;
        RECT 796.500 120.600 798.300 129.000 ;
        RECT 803.100 120.000 804.900 129.600 ;
        RECT 815.100 120.000 816.900 129.600 ;
        RECT 821.700 129.000 825.000 130.200 ;
        RECT 821.700 120.600 823.500 129.000 ;
        RECT 836.400 126.600 837.300 133.950 ;
        RECT 838.950 132.150 840.750 133.950 ;
        RECT 845.100 132.150 846.900 133.950 ;
        RECT 861.000 130.200 861.900 133.950 ;
        RECT 863.100 132.150 864.900 133.950 ;
        RECT 869.100 132.150 870.900 133.950 ;
        RECT 875.550 133.050 876.450 136.950 ;
        RECT 882.000 136.050 882.900 148.200 ;
        RECT 902.100 143.400 903.900 155.400 ;
        RECT 905.100 144.300 906.900 155.400 ;
        RECT 908.100 145.200 909.900 156.000 ;
        RECT 911.100 144.300 912.900 155.400 ;
        RECT 905.100 143.400 912.900 144.300 ;
        RECT 887.100 136.050 888.900 137.850 ;
        RECT 902.400 136.050 903.300 143.400 ;
        RECT 907.950 136.050 909.750 137.850 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 901.950 133.950 904.050 136.050 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 875.550 131.550 880.050 133.050 ;
        RECT 876.000 130.950 880.050 131.550 ;
        RECT 882.000 130.200 882.900 133.950 ;
        RECT 884.100 132.150 885.900 133.950 ;
        RECT 890.100 132.150 891.900 133.950 ;
        RECT 861.000 129.000 864.300 130.200 ;
        RECT 836.400 125.400 841.500 126.600 ;
        RECT 836.700 120.000 838.500 123.600 ;
        RECT 839.700 120.600 841.500 125.400 ;
        RECT 844.200 120.000 846.000 126.600 ;
        RECT 862.500 120.600 864.300 129.000 ;
        RECT 869.100 120.000 870.900 129.600 ;
        RECT 882.000 129.000 885.300 130.200 ;
        RECT 883.500 120.600 885.300 129.000 ;
        RECT 890.100 120.000 891.900 129.600 ;
        RECT 902.400 126.600 903.300 133.950 ;
        RECT 904.950 132.150 906.750 133.950 ;
        RECT 911.100 132.150 912.900 133.950 ;
        RECT 907.950 129.450 910.050 130.050 ;
        RECT 922.950 129.450 925.050 130.050 ;
        RECT 907.950 128.550 925.050 129.450 ;
        RECT 907.950 127.950 910.050 128.550 ;
        RECT 922.950 127.950 925.050 128.550 ;
        RECT 902.400 125.400 907.500 126.600 ;
        RECT 902.700 120.000 904.500 123.600 ;
        RECT 905.700 120.600 907.500 125.400 ;
        RECT 910.200 120.000 912.000 126.600 ;
        RECT 11.100 113.400 12.900 116.400 ;
        RECT 11.100 109.500 12.300 113.400 ;
        RECT 14.100 110.400 15.900 117.000 ;
        RECT 17.100 110.400 18.900 116.400 ;
        RECT 29.100 110.400 30.900 116.400 ;
        RECT 32.100 111.300 33.900 117.000 ;
        RECT 36.600 110.400 38.400 116.400 ;
        RECT 41.100 111.300 42.900 117.000 ;
        RECT 44.100 110.400 45.900 116.400 ;
        RECT 59.100 113.400 60.900 116.400 ;
        RECT 62.100 113.400 63.900 117.000 ;
        RECT 74.100 113.400 75.900 117.000 ;
        RECT 77.100 113.400 78.900 116.400 ;
        RECT 80.100 113.400 81.900 117.000 ;
        RECT 11.100 108.600 16.800 109.500 ;
        RECT 15.000 107.700 16.800 108.600 ;
        RECT 11.400 100.950 13.500 103.050 ;
        RECT 11.400 99.150 13.200 100.950 ;
        RECT 15.000 96.300 15.900 107.700 ;
        RECT 17.700 103.050 18.900 110.400 ;
        RECT 29.700 108.600 30.900 110.400 ;
        RECT 36.900 108.900 38.100 110.400 ;
        RECT 41.100 109.500 45.900 110.400 ;
        RECT 29.700 107.700 36.000 108.600 ;
        RECT 33.900 105.600 36.000 107.700 ;
        RECT 29.400 103.050 31.200 104.850 ;
        RECT 34.200 103.800 36.000 105.600 ;
        RECT 36.900 106.800 39.900 108.900 ;
        RECT 41.100 108.300 43.200 109.500 ;
        RECT 16.800 100.950 18.900 103.050 ;
        RECT 29.100 102.300 31.200 103.050 ;
        RECT 29.100 100.950 36.000 102.300 ;
        RECT 15.000 95.400 16.800 96.300 ;
        RECT 11.100 94.500 16.800 95.400 ;
        RECT 11.100 87.600 12.300 94.500 ;
        RECT 17.700 93.600 18.900 100.950 ;
        RECT 34.200 100.500 36.000 100.950 ;
        RECT 36.900 101.100 38.100 106.800 ;
        RECT 39.000 103.800 41.100 105.900 ;
        RECT 39.300 102.000 41.100 103.800 ;
        RECT 59.700 103.050 60.900 113.400 ;
        RECT 77.400 103.050 78.300 113.400 ;
        RECT 95.100 110.400 96.900 116.400 ;
        RECT 95.700 108.300 96.900 110.400 ;
        RECT 98.100 111.300 99.900 116.400 ;
        RECT 101.100 112.200 102.900 117.000 ;
        RECT 104.100 111.300 105.900 116.400 ;
        RECT 98.100 109.950 105.900 111.300 ;
        RECT 119.400 110.400 121.200 117.000 ;
        RECT 124.500 109.200 126.300 116.400 ;
        RECT 122.100 108.300 126.300 109.200 ;
        RECT 95.700 107.400 99.300 108.300 ;
        RECT 95.100 103.050 96.900 104.850 ;
        RECT 98.100 103.050 99.300 107.400 ;
        RECT 101.100 103.050 102.900 104.850 ;
        RECT 119.250 103.050 121.050 104.850 ;
        RECT 122.100 103.050 123.300 108.300 ;
        RECT 140.100 107.400 141.900 117.000 ;
        RECT 146.700 108.000 148.500 116.400 ;
        RECT 161.700 110.400 163.500 117.000 ;
        RECT 166.200 110.400 168.000 116.400 ;
        RECT 170.700 110.400 172.500 117.000 ;
        RECT 185.100 113.400 186.900 117.000 ;
        RECT 188.100 113.400 189.900 116.400 ;
        RECT 146.700 106.800 150.000 108.000 ;
        RECT 125.100 103.050 126.900 104.850 ;
        RECT 140.100 103.050 141.900 104.850 ;
        RECT 146.100 103.050 147.900 104.850 ;
        RECT 149.100 103.050 150.000 106.800 ;
        RECT 161.250 103.050 163.050 104.850 ;
        RECT 167.100 103.050 168.300 110.400 ;
        RECT 173.100 103.050 174.900 104.850 ;
        RECT 188.100 103.050 189.300 113.400 ;
        RECT 205.500 108.000 207.300 116.400 ;
        RECT 204.000 106.800 207.300 108.000 ;
        RECT 212.100 107.400 213.900 117.000 ;
        RECT 224.700 109.200 226.500 116.400 ;
        RECT 229.800 110.400 231.600 117.000 ;
        RECT 245.100 111.300 246.900 116.400 ;
        RECT 248.100 112.200 249.900 117.000 ;
        RECT 251.100 111.300 252.900 116.400 ;
        RECT 245.100 109.950 252.900 111.300 ;
        RECT 254.100 110.400 255.900 116.400 ;
        RECT 266.100 113.400 267.900 116.400 ;
        RECT 269.100 113.400 270.900 117.000 ;
        RECT 224.700 108.300 228.900 109.200 ;
        RECT 254.100 108.300 255.300 110.400 ;
        RECT 198.000 105.450 202.050 106.050 ;
        RECT 197.550 103.950 202.050 105.450 ;
        RECT 36.900 100.200 39.300 101.100 ;
        RECT 37.800 100.050 39.300 100.200 ;
        RECT 43.800 100.950 45.900 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 76.950 100.950 79.050 103.050 ;
        RECT 79.950 100.950 82.050 103.050 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 121.950 100.950 124.050 103.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 33.000 97.500 36.900 99.300 ;
        RECT 34.800 97.200 36.900 97.500 ;
        RECT 37.800 97.950 39.900 100.050 ;
        RECT 43.800 99.150 45.600 100.950 ;
        RECT 37.800 96.000 38.700 97.950 ;
        RECT 31.500 93.600 33.600 95.700 ;
        RECT 37.200 94.950 38.700 96.000 ;
        RECT 37.200 93.600 38.400 94.950 ;
        RECT 11.100 81.600 12.900 87.600 ;
        RECT 14.100 81.000 15.900 91.800 ;
        RECT 17.100 81.600 18.900 93.600 ;
        RECT 29.100 92.700 33.600 93.600 ;
        RECT 29.100 81.600 30.900 92.700 ;
        RECT 32.100 81.000 33.900 91.500 ;
        RECT 36.600 81.600 38.400 93.600 ;
        RECT 41.100 93.600 43.200 94.500 ;
        RECT 41.100 92.400 45.900 93.600 ;
        RECT 41.100 81.000 42.900 91.500 ;
        RECT 44.100 81.600 45.900 92.400 ;
        RECT 59.700 87.600 60.900 100.950 ;
        RECT 62.100 99.150 63.900 100.950 ;
        RECT 74.250 99.150 76.050 100.950 ;
        RECT 77.400 93.600 78.300 100.950 ;
        RECT 80.100 99.150 81.900 100.950 ;
        RECT 98.100 93.600 99.300 100.950 ;
        RECT 104.100 99.150 105.900 100.950 ;
        RECT 59.100 81.600 60.900 87.600 ;
        RECT 62.100 81.000 63.900 87.600 ;
        RECT 74.100 81.000 75.900 93.600 ;
        RECT 77.400 92.400 81.000 93.600 ;
        RECT 79.200 81.600 81.000 92.400 ;
        RECT 98.100 92.100 100.500 93.600 ;
        RECT 96.000 89.100 97.800 90.900 ;
        RECT 95.700 81.000 97.500 87.600 ;
        RECT 98.700 81.600 100.500 92.100 ;
        RECT 103.800 81.000 105.600 93.600 ;
        RECT 122.100 87.600 123.300 100.950 ;
        RECT 143.100 99.150 144.900 100.950 ;
        RECT 124.950 96.450 127.050 97.050 ;
        RECT 145.950 96.450 148.050 97.050 ;
        RECT 124.950 95.550 148.050 96.450 ;
        RECT 124.950 94.950 127.050 95.550 ;
        RECT 145.950 94.950 148.050 95.550 ;
        RECT 149.100 88.800 150.000 100.950 ;
        RECT 164.250 99.150 166.050 100.950 ;
        RECT 167.100 95.400 168.000 100.950 ;
        RECT 170.100 99.150 171.900 100.950 ;
        RECT 185.100 99.150 186.900 100.950 ;
        RECT 167.100 94.500 171.900 95.400 ;
        RECT 143.400 87.900 150.000 88.800 ;
        RECT 143.400 87.600 144.900 87.900 ;
        RECT 119.100 81.000 120.900 87.600 ;
        RECT 122.100 81.600 123.900 87.600 ;
        RECT 125.100 81.000 126.900 87.600 ;
        RECT 140.100 81.000 141.900 87.600 ;
        RECT 143.100 81.600 144.900 87.600 ;
        RECT 149.100 87.600 150.000 87.900 ;
        RECT 161.100 92.400 168.900 93.300 ;
        RECT 146.100 81.000 147.900 87.000 ;
        RECT 149.100 81.600 150.900 87.600 ;
        RECT 161.100 81.600 162.900 92.400 ;
        RECT 164.100 81.000 165.900 91.500 ;
        RECT 167.100 82.500 168.900 92.400 ;
        RECT 170.100 83.400 171.900 94.500 ;
        RECT 173.100 82.500 174.900 93.600 ;
        RECT 188.100 87.600 189.300 100.950 ;
        RECT 197.550 100.050 198.450 103.950 ;
        RECT 204.000 103.050 204.900 106.800 ;
        RECT 206.100 103.050 207.900 104.850 ;
        RECT 212.100 103.050 213.900 104.850 ;
        RECT 224.100 103.050 225.900 104.850 ;
        RECT 227.700 103.050 228.900 108.300 ;
        RECT 251.700 107.400 255.300 108.300 ;
        RECT 229.950 103.050 231.750 104.850 ;
        RECT 248.100 103.050 249.900 104.850 ;
        RECT 251.700 103.050 252.900 107.400 ;
        RECT 254.100 103.050 255.900 104.850 ;
        RECT 266.700 103.050 267.900 113.400 ;
        RECT 281.400 110.400 283.200 117.000 ;
        RECT 286.500 109.200 288.300 116.400 ;
        RECT 302.100 110.400 303.900 116.400 ;
        RECT 284.100 108.300 288.300 109.200 ;
        RECT 302.700 108.300 303.900 110.400 ;
        RECT 305.100 111.300 306.900 116.400 ;
        RECT 308.100 112.200 309.900 117.000 ;
        RECT 311.100 111.300 312.900 116.400 ;
        RECT 305.100 109.950 312.900 111.300 ;
        RECT 326.700 109.200 328.500 116.400 ;
        RECT 331.800 110.400 333.600 117.000 ;
        RECT 344.100 113.400 345.900 117.000 ;
        RECT 347.100 113.400 348.900 116.400 ;
        RECT 362.100 113.400 363.900 116.400 ;
        RECT 365.100 113.400 366.900 117.000 ;
        RECT 326.700 108.300 330.900 109.200 ;
        RECT 281.250 103.050 283.050 104.850 ;
        RECT 284.100 103.050 285.300 108.300 ;
        RECT 302.700 107.400 306.300 108.300 ;
        RECT 297.000 105.450 301.050 106.050 ;
        RECT 287.100 103.050 288.900 104.850 ;
        RECT 296.550 103.950 301.050 105.450 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 197.550 98.550 202.050 100.050 ;
        RECT 198.000 97.950 202.050 98.550 ;
        RECT 204.000 88.800 204.900 100.950 ;
        RECT 209.100 99.150 210.900 100.950 ;
        RECT 205.950 96.450 208.050 97.050 ;
        RECT 217.950 96.450 220.050 97.050 ;
        RECT 205.950 95.550 220.050 96.450 ;
        RECT 205.950 94.950 208.050 95.550 ;
        RECT 217.950 94.950 220.050 95.550 ;
        RECT 204.000 87.900 210.600 88.800 ;
        RECT 204.000 87.600 204.900 87.900 ;
        RECT 167.100 81.600 174.900 82.500 ;
        RECT 185.100 81.000 186.900 87.600 ;
        RECT 188.100 81.600 189.900 87.600 ;
        RECT 203.100 81.600 204.900 87.600 ;
        RECT 209.100 87.600 210.600 87.900 ;
        RECT 227.700 87.600 228.900 100.950 ;
        RECT 245.100 99.150 246.900 100.950 ;
        RECT 251.700 93.600 252.900 100.950 ;
        RECT 206.100 81.000 207.900 87.000 ;
        RECT 209.100 81.600 210.900 87.600 ;
        RECT 212.100 81.000 213.900 87.600 ;
        RECT 224.100 81.000 225.900 87.600 ;
        RECT 227.100 81.600 228.900 87.600 ;
        RECT 230.100 81.000 231.900 87.600 ;
        RECT 245.400 81.000 247.200 93.600 ;
        RECT 250.500 92.100 252.900 93.600 ;
        RECT 250.500 81.600 252.300 92.100 ;
        RECT 253.200 89.100 255.000 90.900 ;
        RECT 266.700 87.600 267.900 100.950 ;
        RECT 269.100 99.150 270.900 100.950 ;
        RECT 284.100 87.600 285.300 100.950 ;
        RECT 296.550 100.050 297.450 103.950 ;
        RECT 302.100 103.050 303.900 104.850 ;
        RECT 305.100 103.050 306.300 107.400 ;
        RECT 308.100 103.050 309.900 104.850 ;
        RECT 326.100 103.050 327.900 104.850 ;
        RECT 329.700 103.050 330.900 108.300 ;
        RECT 331.950 103.050 333.750 104.850 ;
        RECT 347.100 103.050 348.300 113.400 ;
        RECT 362.700 103.050 363.900 113.400 ;
        RECT 377.700 109.200 379.500 116.400 ;
        RECT 382.800 110.400 384.600 117.000 ;
        RECT 399.600 112.200 401.400 116.400 ;
        RECT 398.700 110.400 401.400 112.200 ;
        RECT 402.600 110.400 404.400 117.000 ;
        RECT 364.950 108.450 367.050 109.050 ;
        RECT 370.950 108.450 373.050 109.050 ;
        RECT 364.950 107.550 373.050 108.450 ;
        RECT 377.700 108.300 381.900 109.200 ;
        RECT 364.950 106.950 367.050 107.550 ;
        RECT 370.950 106.950 373.050 107.550 ;
        RECT 377.100 103.050 378.900 104.850 ;
        RECT 380.700 103.050 381.900 108.300 ;
        RECT 382.950 103.050 384.750 104.850 ;
        RECT 398.700 103.050 399.600 110.400 ;
        RECT 400.500 108.600 402.300 109.500 ;
        RECT 407.100 108.600 408.900 116.400 ;
        RECT 421.500 110.400 423.300 117.000 ;
        RECT 426.000 110.400 427.800 116.400 ;
        RECT 430.500 110.400 432.300 117.000 ;
        RECT 400.500 107.700 408.900 108.600 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 328.950 100.950 331.050 103.050 ;
        RECT 331.950 100.950 334.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 398.100 100.950 400.200 103.050 ;
        RECT 401.400 100.950 403.500 103.050 ;
        RECT 296.550 98.550 301.050 100.050 ;
        RECT 297.000 97.950 301.050 98.550 ;
        RECT 292.950 96.450 295.050 97.050 ;
        RECT 301.950 96.450 304.050 97.050 ;
        RECT 292.950 95.550 304.050 96.450 ;
        RECT 292.950 94.950 295.050 95.550 ;
        RECT 301.950 94.950 304.050 95.550 ;
        RECT 286.950 93.450 289.050 94.050 ;
        RECT 298.950 93.450 301.050 94.050 ;
        RECT 286.950 92.550 301.050 93.450 ;
        RECT 286.950 91.950 289.050 92.550 ;
        RECT 298.950 91.950 301.050 92.550 ;
        RECT 305.100 93.600 306.300 100.950 ;
        RECT 311.100 99.150 312.900 100.950 ;
        RECT 305.100 92.100 307.500 93.600 ;
        RECT 303.000 89.100 304.800 90.900 ;
        RECT 253.500 81.000 255.300 87.600 ;
        RECT 266.100 81.600 267.900 87.600 ;
        RECT 269.100 81.000 270.900 87.600 ;
        RECT 281.100 81.000 282.900 87.600 ;
        RECT 284.100 81.600 285.900 87.600 ;
        RECT 287.100 81.000 288.900 87.600 ;
        RECT 302.700 81.000 304.500 87.600 ;
        RECT 305.700 81.600 307.500 92.100 ;
        RECT 310.800 81.000 312.600 93.600 ;
        RECT 329.700 87.600 330.900 100.950 ;
        RECT 344.100 99.150 345.900 100.950 ;
        RECT 347.100 87.600 348.300 100.950 ;
        RECT 362.700 87.600 363.900 100.950 ;
        RECT 365.100 99.150 366.900 100.950 ;
        RECT 380.700 87.600 381.900 100.950 ;
        RECT 398.700 93.600 399.600 100.950 ;
        RECT 402.000 99.150 403.800 100.950 ;
        RECT 326.100 81.000 327.900 87.600 ;
        RECT 329.100 81.600 330.900 87.600 ;
        RECT 332.100 81.000 333.900 87.600 ;
        RECT 344.100 81.000 345.900 87.600 ;
        RECT 347.100 81.600 348.900 87.600 ;
        RECT 362.100 81.600 363.900 87.600 ;
        RECT 365.100 81.000 366.900 87.600 ;
        RECT 377.100 81.000 378.900 87.600 ;
        RECT 380.100 81.600 381.900 87.600 ;
        RECT 383.100 81.000 384.900 87.600 ;
        RECT 398.100 81.600 399.900 93.600 ;
        RECT 401.100 81.000 402.900 93.000 ;
        RECT 405.000 87.600 405.900 107.700 ;
        RECT 406.950 103.050 408.750 104.850 ;
        RECT 419.100 103.050 420.900 104.850 ;
        RECT 425.700 103.050 426.900 110.400 ;
        RECT 445.500 108.000 447.300 116.400 ;
        RECT 444.000 106.800 447.300 108.000 ;
        RECT 452.100 107.400 453.900 117.000 ;
        RECT 467.700 113.400 469.500 117.000 ;
        RECT 470.700 111.600 472.500 116.400 ;
        RECT 467.400 110.400 472.500 111.600 ;
        RECT 475.200 110.400 477.000 117.000 ;
        RECT 488.400 110.400 490.200 117.000 ;
        RECT 430.950 103.050 432.750 104.850 ;
        RECT 444.000 103.050 444.900 106.800 ;
        RECT 446.100 103.050 447.900 104.850 ;
        RECT 452.100 103.050 453.900 104.850 ;
        RECT 467.400 103.050 468.300 110.400 ;
        RECT 493.500 109.200 495.300 116.400 ;
        RECT 509.100 113.400 510.900 117.000 ;
        RECT 512.100 113.400 513.900 116.400 ;
        RECT 515.100 113.400 516.900 117.000 ;
        RECT 491.100 108.300 495.300 109.200 ;
        RECT 469.950 103.050 471.750 104.850 ;
        RECT 476.100 103.050 477.900 104.850 ;
        RECT 488.250 103.050 490.050 104.850 ;
        RECT 491.100 103.050 492.300 108.300 ;
        RECT 494.100 103.050 495.900 104.850 ;
        RECT 512.700 103.050 513.600 113.400 ;
        RECT 530.400 110.400 532.200 117.000 ;
        RECT 535.500 109.200 537.300 116.400 ;
        RECT 551.100 110.400 552.900 116.400 ;
        RECT 533.100 108.300 537.300 109.200 ;
        RECT 551.700 108.300 552.900 110.400 ;
        RECT 554.100 111.300 555.900 116.400 ;
        RECT 557.100 112.200 558.900 117.000 ;
        RECT 560.100 111.300 561.900 116.400 ;
        RECT 554.100 109.950 561.900 111.300 ;
        RECT 575.100 111.300 576.900 116.400 ;
        RECT 578.100 112.200 579.900 117.000 ;
        RECT 581.100 111.300 582.900 116.400 ;
        RECT 575.100 109.950 582.900 111.300 ;
        RECT 584.100 110.400 585.900 116.400 ;
        RECT 596.400 110.400 598.200 117.000 ;
        RECT 584.100 108.300 585.300 110.400 ;
        RECT 601.500 109.200 603.300 116.400 ;
        RECT 617.100 113.400 618.900 117.000 ;
        RECT 620.100 113.400 621.900 116.400 ;
        RECT 623.100 113.400 624.900 117.000 ;
        RECT 530.250 103.050 532.050 104.850 ;
        RECT 533.100 103.050 534.300 108.300 ;
        RECT 551.700 107.400 555.300 108.300 ;
        RECT 536.100 103.050 537.900 104.850 ;
        RECT 551.100 103.050 552.900 104.850 ;
        RECT 554.100 103.050 555.300 107.400 ;
        RECT 581.700 107.400 585.300 108.300 ;
        RECT 599.100 108.300 603.300 109.200 ;
        RECT 557.100 103.050 558.900 104.850 ;
        RECT 578.100 103.050 579.900 104.850 ;
        RECT 581.700 103.050 582.900 107.400 ;
        RECT 584.100 103.050 585.900 104.850 ;
        RECT 596.250 103.050 598.050 104.850 ;
        RECT 599.100 103.050 600.300 108.300 ;
        RECT 602.100 103.050 603.900 104.850 ;
        RECT 620.700 103.050 621.600 113.400 ;
        RECT 639.000 110.400 640.800 117.000 ;
        RECT 643.500 111.600 645.300 116.400 ;
        RECT 646.500 113.400 648.300 117.000 ;
        RECT 643.500 110.400 648.600 111.600 ;
        RECT 659.100 110.400 660.900 116.400 ;
        RECT 625.950 105.450 628.050 106.050 ;
        RECT 625.950 104.550 633.450 105.450 ;
        RECT 625.950 103.950 628.050 104.550 ;
        RECT 406.800 100.950 408.900 103.050 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 448.950 100.950 451.050 103.050 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 422.100 99.150 423.900 100.950 ;
        RECT 426.000 95.400 426.900 100.950 ;
        RECT 427.950 99.150 429.750 100.950 ;
        RECT 422.100 94.500 426.900 95.400 ;
        RECT 404.100 81.600 405.900 87.600 ;
        RECT 407.100 81.000 408.900 87.600 ;
        RECT 419.100 82.500 420.900 93.600 ;
        RECT 422.100 83.400 423.900 94.500 ;
        RECT 425.100 92.400 432.900 93.300 ;
        RECT 425.100 82.500 426.900 92.400 ;
        RECT 419.100 81.600 426.900 82.500 ;
        RECT 428.100 81.000 429.900 91.500 ;
        RECT 431.100 81.600 432.900 92.400 ;
        RECT 444.000 88.800 444.900 100.950 ;
        RECT 449.100 99.150 450.900 100.950 ;
        RECT 467.400 93.600 468.300 100.950 ;
        RECT 472.950 99.150 474.750 100.950 ;
        RECT 444.000 87.900 450.600 88.800 ;
        RECT 444.000 87.600 444.900 87.900 ;
        RECT 443.100 81.600 444.900 87.600 ;
        RECT 449.100 87.600 450.600 87.900 ;
        RECT 446.100 81.000 447.900 87.000 ;
        RECT 449.100 81.600 450.900 87.600 ;
        RECT 452.100 81.000 453.900 87.600 ;
        RECT 467.100 81.600 468.900 93.600 ;
        RECT 470.100 92.700 477.900 93.600 ;
        RECT 470.100 81.600 471.900 92.700 ;
        RECT 473.100 81.000 474.900 91.800 ;
        RECT 476.100 81.600 477.900 92.700 ;
        RECT 491.100 87.600 492.300 100.950 ;
        RECT 509.100 99.150 510.900 100.950 ;
        RECT 512.700 93.600 513.600 100.950 ;
        RECT 514.950 99.150 516.750 100.950 ;
        RECT 510.000 92.400 513.600 93.600 ;
        RECT 488.100 81.000 489.900 87.600 ;
        RECT 491.100 81.600 492.900 87.600 ;
        RECT 494.100 81.000 495.900 87.600 ;
        RECT 510.000 81.600 511.800 92.400 ;
        RECT 515.100 81.000 516.900 93.600 ;
        RECT 533.100 87.600 534.300 100.950 ;
        RECT 554.100 93.600 555.300 100.950 ;
        RECT 560.100 99.150 561.900 100.950 ;
        RECT 575.100 99.150 576.900 100.950 ;
        RECT 556.950 96.450 559.050 97.050 ;
        RECT 568.950 96.450 571.050 97.050 ;
        RECT 556.950 95.550 571.050 96.450 ;
        RECT 556.950 94.950 559.050 95.550 ;
        RECT 568.950 94.950 571.050 95.550 ;
        RECT 581.700 93.600 582.900 100.950 ;
        RECT 554.100 92.100 556.500 93.600 ;
        RECT 552.000 89.100 553.800 90.900 ;
        RECT 530.100 81.000 531.900 87.600 ;
        RECT 533.100 81.600 534.900 87.600 ;
        RECT 536.100 81.000 537.900 87.600 ;
        RECT 551.700 81.000 553.500 87.600 ;
        RECT 554.700 81.600 556.500 92.100 ;
        RECT 559.800 81.000 561.600 93.600 ;
        RECT 575.400 81.000 577.200 93.600 ;
        RECT 580.500 92.100 582.900 93.600 ;
        RECT 580.500 81.600 582.300 92.100 ;
        RECT 583.200 89.100 585.000 90.900 ;
        RECT 599.100 87.600 600.300 100.950 ;
        RECT 617.100 99.150 618.900 100.950 ;
        RECT 620.700 93.600 621.600 100.950 ;
        RECT 622.950 99.150 624.750 100.950 ;
        RECT 632.550 100.050 633.450 104.550 ;
        RECT 638.100 103.050 639.900 104.850 ;
        RECT 644.250 103.050 646.050 104.850 ;
        RECT 647.700 103.050 648.600 110.400 ;
        RECT 659.700 108.300 660.900 110.400 ;
        RECT 662.100 111.300 663.900 116.400 ;
        RECT 665.100 112.200 666.900 117.000 ;
        RECT 668.100 111.300 669.900 116.400 ;
        RECT 662.100 109.950 669.900 111.300 ;
        RECT 659.700 107.400 663.300 108.300 ;
        RECT 685.500 108.000 687.300 116.400 ;
        RECT 659.100 103.050 660.900 104.850 ;
        RECT 662.100 103.050 663.300 107.400 ;
        RECT 684.000 106.800 687.300 108.000 ;
        RECT 692.100 107.400 693.900 117.000 ;
        RECT 706.500 110.400 708.300 117.000 ;
        RECT 711.000 110.400 712.800 116.400 ;
        RECT 715.500 110.400 717.300 117.000 ;
        RECT 731.100 113.400 732.900 117.000 ;
        RECT 734.100 113.400 735.900 116.400 ;
        RECT 746.700 113.400 748.500 117.000 ;
        RECT 665.100 103.050 666.900 104.850 ;
        RECT 684.000 103.050 684.900 106.800 ;
        RECT 686.100 103.050 687.900 104.850 ;
        RECT 692.100 103.050 693.900 104.850 ;
        RECT 704.100 103.050 705.900 104.850 ;
        RECT 710.700 103.050 711.900 110.400 ;
        RECT 715.950 103.050 717.750 104.850 ;
        RECT 734.100 103.050 735.300 113.400 ;
        RECT 749.700 111.600 751.500 116.400 ;
        RECT 746.400 110.400 751.500 111.600 ;
        RECT 754.200 110.400 756.000 117.000 ;
        RECT 746.400 103.050 747.300 110.400 ;
        RECT 767.100 107.400 768.900 117.000 ;
        RECT 773.700 108.000 775.500 116.400 ;
        RECT 789.000 110.400 790.800 117.000 ;
        RECT 793.500 111.600 795.300 116.400 ;
        RECT 796.500 113.400 798.300 117.000 ;
        RECT 793.500 110.400 798.600 111.600 ;
        RECT 773.700 106.800 777.000 108.000 ;
        RECT 748.950 103.050 750.750 104.850 ;
        RECT 755.100 103.050 756.900 104.850 ;
        RECT 767.100 103.050 768.900 104.850 ;
        RECT 773.100 103.050 774.900 104.850 ;
        RECT 776.100 103.050 777.000 106.800 ;
        RECT 788.100 103.050 789.900 104.850 ;
        RECT 794.250 103.050 796.050 104.850 ;
        RECT 797.700 103.050 798.600 110.400 ;
        RECT 809.100 111.300 810.900 116.400 ;
        RECT 812.100 112.200 813.900 117.000 ;
        RECT 815.100 111.300 816.900 116.400 ;
        RECT 809.100 109.950 816.900 111.300 ;
        RECT 818.100 110.400 819.900 116.400 ;
        RECT 831.000 110.400 832.800 117.000 ;
        RECT 835.500 111.600 837.300 116.400 ;
        RECT 838.500 113.400 840.300 117.000 ;
        RECT 835.500 110.400 840.600 111.600 ;
        RECT 818.100 108.300 819.300 110.400 ;
        RECT 815.700 107.400 819.300 108.300 ;
        RECT 812.100 103.050 813.900 104.850 ;
        RECT 815.700 103.050 816.900 107.400 ;
        RECT 818.100 103.050 819.900 104.850 ;
        RECT 830.100 103.050 831.900 104.850 ;
        RECT 836.250 103.050 838.050 104.850 ;
        RECT 839.700 103.050 840.600 110.400 ;
        RECT 854.100 107.400 855.900 117.000 ;
        RECT 860.700 108.000 862.500 116.400 ;
        RECT 878.100 111.300 879.900 116.400 ;
        RECT 881.100 112.200 882.900 117.000 ;
        RECT 884.100 111.300 885.900 116.400 ;
        RECT 878.100 109.950 885.900 111.300 ;
        RECT 887.100 110.400 888.900 116.400 ;
        RECT 902.100 111.300 903.900 116.400 ;
        RECT 905.100 112.200 906.900 117.000 ;
        RECT 908.100 111.300 909.900 116.400 ;
        RECT 887.100 108.300 888.300 110.400 ;
        RECT 902.100 109.950 909.900 111.300 ;
        RECT 911.100 110.400 912.900 116.400 ;
        RECT 911.100 108.300 912.300 110.400 ;
        RECT 860.700 106.800 864.000 108.000 ;
        RECT 854.100 103.050 855.900 104.850 ;
        RECT 860.100 103.050 861.900 104.850 ;
        RECT 863.100 103.050 864.000 106.800 ;
        RECT 884.700 107.400 888.300 108.300 ;
        RECT 908.700 107.400 912.300 108.300 ;
        RECT 881.100 103.050 882.900 104.850 ;
        RECT 884.700 103.050 885.900 107.400 ;
        RECT 887.100 103.050 888.900 104.850 ;
        RECT 905.100 103.050 906.900 104.850 ;
        RECT 908.700 103.050 909.900 107.400 ;
        RECT 911.100 103.050 912.900 104.850 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 745.950 100.950 748.050 103.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 751.950 100.950 754.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 814.950 100.950 817.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 880.950 100.950 883.050 103.050 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 901.950 100.950 904.050 103.050 ;
        RECT 904.950 100.950 907.050 103.050 ;
        RECT 907.950 100.950 910.050 103.050 ;
        RECT 910.950 100.950 913.050 103.050 ;
        RECT 632.550 98.550 637.050 100.050 ;
        RECT 641.250 99.150 643.050 100.950 ;
        RECT 633.000 97.950 637.050 98.550 ;
        RECT 647.700 93.600 648.600 100.950 ;
        RECT 662.100 93.600 663.300 100.950 ;
        RECT 668.100 99.150 669.900 100.950 ;
        RECT 618.000 92.400 621.600 93.600 ;
        RECT 583.500 81.000 585.300 87.600 ;
        RECT 596.100 81.000 597.900 87.600 ;
        RECT 599.100 81.600 600.900 87.600 ;
        RECT 602.100 81.000 603.900 87.600 ;
        RECT 618.000 81.600 619.800 92.400 ;
        RECT 623.100 81.000 624.900 93.600 ;
        RECT 638.100 92.700 645.900 93.600 ;
        RECT 638.100 81.600 639.900 92.700 ;
        RECT 641.100 81.000 642.900 91.800 ;
        RECT 644.100 81.600 645.900 92.700 ;
        RECT 647.100 81.600 648.900 93.600 ;
        RECT 662.100 92.100 664.500 93.600 ;
        RECT 660.000 89.100 661.800 90.900 ;
        RECT 659.700 81.000 661.500 87.600 ;
        RECT 662.700 81.600 664.500 92.100 ;
        RECT 667.800 81.000 669.600 93.600 ;
        RECT 684.000 88.800 684.900 100.950 ;
        RECT 689.100 99.150 690.900 100.950 ;
        RECT 707.100 99.150 708.900 100.950 ;
        RECT 711.000 95.400 711.900 100.950 ;
        RECT 712.950 99.150 714.750 100.950 ;
        RECT 731.100 99.150 732.900 100.950 ;
        RECT 707.100 94.500 711.900 95.400 ;
        RECT 684.000 87.900 690.600 88.800 ;
        RECT 684.000 87.600 684.900 87.900 ;
        RECT 683.100 81.600 684.900 87.600 ;
        RECT 689.100 87.600 690.600 87.900 ;
        RECT 686.100 81.000 687.900 87.000 ;
        RECT 689.100 81.600 690.900 87.600 ;
        RECT 692.100 81.000 693.900 87.600 ;
        RECT 704.100 82.500 705.900 93.600 ;
        RECT 707.100 83.400 708.900 94.500 ;
        RECT 710.100 92.400 717.900 93.300 ;
        RECT 710.100 82.500 711.900 92.400 ;
        RECT 704.100 81.600 711.900 82.500 ;
        RECT 713.100 81.000 714.900 91.500 ;
        RECT 716.100 81.600 717.900 92.400 ;
        RECT 734.100 87.600 735.300 100.950 ;
        RECT 746.400 93.600 747.300 100.950 ;
        RECT 751.950 99.150 753.750 100.950 ;
        RECT 770.100 99.150 771.900 100.950 ;
        RECT 731.100 81.000 732.900 87.600 ;
        RECT 734.100 81.600 735.900 87.600 ;
        RECT 746.100 81.600 747.900 93.600 ;
        RECT 749.100 92.700 756.900 93.600 ;
        RECT 749.100 81.600 750.900 92.700 ;
        RECT 752.100 81.000 753.900 91.800 ;
        RECT 755.100 81.600 756.900 92.700 ;
        RECT 776.100 88.800 777.000 100.950 ;
        RECT 791.250 99.150 793.050 100.950 ;
        RECT 797.700 93.600 798.600 100.950 ;
        RECT 809.100 99.150 810.900 100.950 ;
        RECT 815.700 93.600 816.900 100.950 ;
        RECT 833.250 99.150 835.050 100.950 ;
        RECT 839.700 93.600 840.600 100.950 ;
        RECT 857.100 99.150 858.900 100.950 ;
        RECT 770.400 87.900 777.000 88.800 ;
        RECT 770.400 87.600 771.900 87.900 ;
        RECT 767.100 81.000 768.900 87.600 ;
        RECT 770.100 81.600 771.900 87.600 ;
        RECT 776.100 87.600 777.000 87.900 ;
        RECT 788.100 92.700 795.900 93.600 ;
        RECT 773.100 81.000 774.900 87.000 ;
        RECT 776.100 81.600 777.900 87.600 ;
        RECT 788.100 81.600 789.900 92.700 ;
        RECT 791.100 81.000 792.900 91.800 ;
        RECT 794.100 81.600 795.900 92.700 ;
        RECT 797.100 81.600 798.900 93.600 ;
        RECT 809.400 81.000 811.200 93.600 ;
        RECT 814.500 92.100 816.900 93.600 ;
        RECT 830.100 92.700 837.900 93.600 ;
        RECT 814.500 81.600 816.300 92.100 ;
        RECT 817.200 89.100 819.000 90.900 ;
        RECT 817.500 81.000 819.300 87.600 ;
        RECT 830.100 81.600 831.900 92.700 ;
        RECT 833.100 81.000 834.900 91.800 ;
        RECT 836.100 81.600 837.900 92.700 ;
        RECT 839.100 81.600 840.900 93.600 ;
        RECT 863.100 88.800 864.000 100.950 ;
        RECT 878.100 99.150 879.900 100.950 ;
        RECT 884.700 93.600 885.900 100.950 ;
        RECT 889.950 99.450 892.050 100.050 ;
        RECT 895.950 99.450 898.050 100.050 ;
        RECT 889.950 98.550 898.050 99.450 ;
        RECT 902.100 99.150 903.900 100.950 ;
        RECT 889.950 97.950 892.050 98.550 ;
        RECT 895.950 97.950 898.050 98.550 ;
        RECT 908.700 93.600 909.900 100.950 ;
        RECT 857.400 87.900 864.000 88.800 ;
        RECT 857.400 87.600 858.900 87.900 ;
        RECT 854.100 81.000 855.900 87.600 ;
        RECT 857.100 81.600 858.900 87.600 ;
        RECT 863.100 87.600 864.000 87.900 ;
        RECT 860.100 81.000 861.900 87.000 ;
        RECT 863.100 81.600 864.900 87.600 ;
        RECT 878.400 81.000 880.200 93.600 ;
        RECT 883.500 92.100 885.900 93.600 ;
        RECT 883.500 81.600 885.300 92.100 ;
        RECT 886.200 89.100 888.000 90.900 ;
        RECT 886.500 81.000 888.300 87.600 ;
        RECT 902.400 81.000 904.200 93.600 ;
        RECT 907.500 92.100 909.900 93.600 ;
        RECT 907.500 81.600 909.300 92.100 ;
        RECT 910.200 89.100 912.000 90.900 ;
        RECT 910.500 81.000 912.300 87.600 ;
        RECT 14.100 71.400 15.900 77.400 ;
        RECT 17.100 71.400 18.900 78.000 ;
        RECT 14.700 58.050 15.900 71.400 ;
        RECT 29.100 65.400 30.900 77.400 ;
        RECT 32.100 66.300 33.900 77.400 ;
        RECT 35.100 67.200 36.900 78.000 ;
        RECT 38.100 66.300 39.900 77.400 ;
        RECT 50.700 71.400 52.500 78.000 ;
        RECT 51.000 68.100 52.800 69.900 ;
        RECT 53.700 66.900 55.500 77.400 ;
        RECT 32.100 65.400 39.900 66.300 ;
        RECT 53.100 65.400 55.500 66.900 ;
        RECT 58.800 65.400 60.600 78.000 ;
        RECT 75.000 66.600 76.800 77.400 ;
        RECT 75.000 65.400 78.600 66.600 ;
        RECT 80.100 65.400 81.900 78.000 ;
        RECT 92.100 71.400 93.900 77.400 ;
        RECT 95.100 72.000 96.900 78.000 ;
        RECT 93.000 71.100 93.900 71.400 ;
        RECT 98.100 71.400 99.900 77.400 ;
        RECT 101.100 71.400 102.900 78.000 ;
        RECT 116.100 71.400 117.900 78.000 ;
        RECT 119.100 71.400 120.900 77.400 ;
        RECT 122.100 71.400 123.900 78.000 ;
        RECT 134.100 71.400 135.900 77.400 ;
        RECT 137.100 72.000 138.900 78.000 ;
        RECT 98.100 71.100 99.600 71.400 ;
        RECT 93.000 70.200 99.600 71.100 ;
        RECT 85.950 67.950 88.050 70.050 ;
        RECT 17.100 58.050 18.900 59.850 ;
        RECT 29.400 58.050 30.300 65.400 ;
        RECT 31.950 63.450 34.050 64.200 ;
        RECT 43.950 63.450 46.050 64.050 ;
        RECT 49.950 63.450 52.050 64.050 ;
        RECT 31.950 62.550 42.450 63.450 ;
        RECT 31.950 62.100 34.050 62.550 ;
        RECT 41.550 60.450 42.450 62.550 ;
        RECT 43.950 62.550 52.050 63.450 ;
        RECT 43.950 61.950 46.050 62.550 ;
        RECT 49.950 61.950 52.050 62.550 ;
        RECT 46.950 60.450 49.050 60.900 ;
        RECT 34.950 58.050 36.750 59.850 ;
        RECT 41.550 59.550 49.050 60.450 ;
        RECT 46.950 58.800 49.050 59.550 ;
        RECT 53.100 58.050 54.300 65.400 ;
        RECT 55.950 63.450 58.050 64.050 ;
        RECT 55.950 62.550 63.450 63.450 ;
        RECT 55.950 61.950 58.050 62.550 ;
        RECT 62.550 60.450 63.450 62.550 ;
        RECT 59.100 58.050 60.900 59.850 ;
        RECT 62.550 59.550 66.450 60.450 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 28.950 55.950 31.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 49.950 55.950 52.050 58.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 14.700 45.600 15.900 55.950 ;
        RECT 29.400 48.600 30.300 55.950 ;
        RECT 31.950 54.150 33.750 55.950 ;
        RECT 38.100 54.150 39.900 55.950 ;
        RECT 50.100 54.150 51.900 55.950 ;
        RECT 53.100 51.600 54.300 55.950 ;
        RECT 56.100 54.150 57.900 55.950 ;
        RECT 65.550 55.050 66.450 59.550 ;
        RECT 74.100 58.050 75.900 59.850 ;
        RECT 77.700 58.050 78.600 65.400 ;
        RECT 79.950 58.050 81.750 59.850 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 61.950 53.550 66.450 55.050 ;
        RECT 61.950 52.950 66.000 53.550 ;
        RECT 50.700 50.700 54.300 51.600 ;
        RECT 50.700 48.600 51.900 50.700 ;
        RECT 29.400 47.400 34.500 48.600 ;
        RECT 14.100 42.600 15.900 45.600 ;
        RECT 17.100 42.000 18.900 45.600 ;
        RECT 29.700 42.000 31.500 45.600 ;
        RECT 32.700 42.600 34.500 47.400 ;
        RECT 37.200 42.000 39.000 48.600 ;
        RECT 50.100 42.600 51.900 48.600 ;
        RECT 53.100 47.700 60.900 49.050 ;
        RECT 53.100 42.600 54.900 47.700 ;
        RECT 56.100 42.000 57.900 46.800 ;
        RECT 59.100 42.600 60.900 47.700 ;
        RECT 77.700 45.600 78.600 55.950 ;
        RECT 86.550 55.050 87.450 67.950 ;
        RECT 93.000 58.050 93.900 70.200 ;
        RECT 106.950 63.450 109.050 64.050 ;
        RECT 115.950 63.450 118.050 64.200 ;
        RECT 106.950 62.550 118.050 63.450 ;
        RECT 106.950 61.950 109.050 62.550 ;
        RECT 115.950 62.100 118.050 62.550 ;
        RECT 98.100 58.050 99.900 59.850 ;
        RECT 119.700 58.050 120.900 71.400 ;
        RECT 135.000 71.100 135.900 71.400 ;
        RECT 140.100 71.400 141.900 77.400 ;
        RECT 143.100 71.400 144.900 78.000 ;
        RECT 158.100 71.400 159.900 78.000 ;
        RECT 161.100 71.400 162.900 77.400 ;
        RECT 164.100 71.400 165.900 78.000 ;
        RECT 176.100 71.400 177.900 77.400 ;
        RECT 179.100 71.400 180.900 78.000 ;
        RECT 194.100 71.400 195.900 77.400 ;
        RECT 197.100 72.000 198.900 78.000 ;
        RECT 140.100 71.100 141.600 71.400 ;
        RECT 135.000 70.200 141.600 71.100 ;
        RECT 135.000 58.050 135.900 70.200 ;
        RECT 140.100 58.050 141.900 59.850 ;
        RECT 161.100 58.050 162.300 71.400 ;
        RECT 176.700 58.050 177.900 71.400 ;
        RECT 195.000 71.100 195.900 71.400 ;
        RECT 200.100 71.400 201.900 77.400 ;
        RECT 203.100 71.400 204.900 78.000 ;
        RECT 200.100 71.100 201.600 71.400 ;
        RECT 195.000 70.200 201.600 71.100 ;
        RECT 179.100 58.050 180.900 59.850 ;
        RECT 195.000 58.050 195.900 70.200 ;
        RECT 218.100 66.300 219.900 77.400 ;
        RECT 221.100 67.200 222.900 78.000 ;
        RECT 224.100 66.300 225.900 77.400 ;
        RECT 218.100 65.400 225.900 66.300 ;
        RECT 227.100 65.400 228.900 77.400 ;
        RECT 239.400 65.400 241.200 78.000 ;
        RECT 244.500 66.900 246.300 77.400 ;
        RECT 247.500 71.400 249.300 78.000 ;
        RECT 263.100 71.400 264.900 77.400 ;
        RECT 266.100 72.000 267.900 78.000 ;
        RECT 264.000 71.100 264.900 71.400 ;
        RECT 269.100 71.400 270.900 77.400 ;
        RECT 272.100 71.400 273.900 78.000 ;
        RECT 287.100 71.400 288.900 78.000 ;
        RECT 290.100 71.400 291.900 77.400 ;
        RECT 293.100 71.400 294.900 78.000 ;
        RECT 308.100 71.400 309.900 78.000 ;
        RECT 311.100 71.400 312.900 77.400 ;
        RECT 314.100 71.400 315.900 78.000 ;
        RECT 269.100 71.100 270.600 71.400 ;
        RECT 264.000 70.200 270.600 71.100 ;
        RECT 247.200 68.100 249.000 69.900 ;
        RECT 244.500 65.400 246.900 66.900 ;
        RECT 196.950 63.450 199.050 64.050 ;
        RECT 217.950 63.450 220.050 64.050 ;
        RECT 196.950 62.550 220.050 63.450 ;
        RECT 196.950 61.950 199.050 62.550 ;
        RECT 217.950 61.950 220.050 62.550 ;
        RECT 200.100 58.050 201.900 59.850 ;
        RECT 221.250 58.050 223.050 59.850 ;
        RECT 227.700 58.050 228.600 65.400 ;
        RECT 239.100 58.050 240.900 59.850 ;
        RECT 245.700 58.050 246.900 65.400 ;
        RECT 264.000 58.050 264.900 70.200 ;
        RECT 269.100 58.050 270.900 59.850 ;
        RECT 290.700 58.050 291.900 71.400 ;
        RECT 311.100 58.050 312.300 71.400 ;
        RECT 329.100 65.400 330.900 77.400 ;
        RECT 332.100 66.300 333.900 77.400 ;
        RECT 335.100 67.200 336.900 78.000 ;
        RECT 338.100 66.300 339.900 77.400 ;
        RECT 353.100 71.400 354.900 77.400 ;
        RECT 356.100 72.000 357.900 78.000 ;
        RECT 332.100 65.400 339.900 66.300 ;
        RECT 354.000 71.100 354.900 71.400 ;
        RECT 359.100 71.400 360.900 77.400 ;
        RECT 362.100 71.400 363.900 78.000 ;
        RECT 359.100 71.100 360.600 71.400 ;
        RECT 354.000 70.200 360.600 71.100 ;
        RECT 316.950 60.450 321.000 61.050 ;
        RECT 316.950 58.950 321.450 60.450 ;
        RECT 91.950 55.950 94.050 58.050 ;
        RECT 94.950 55.950 97.050 58.050 ;
        RECT 97.950 55.950 100.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 115.950 55.950 118.050 58.050 ;
        RECT 118.950 55.950 121.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 220.950 55.950 223.050 58.050 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 86.550 53.550 91.050 55.050 ;
        RECT 87.000 52.950 91.050 53.550 ;
        RECT 93.000 52.200 93.900 55.950 ;
        RECT 95.100 54.150 96.900 55.950 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 116.100 54.150 117.900 55.950 ;
        RECT 93.000 51.000 96.300 52.200 ;
        RECT 74.100 42.000 75.900 45.600 ;
        RECT 77.100 42.600 78.900 45.600 ;
        RECT 80.100 42.000 81.900 45.600 ;
        RECT 94.500 42.600 96.300 51.000 ;
        RECT 101.100 42.000 102.900 51.600 ;
        RECT 119.700 50.700 120.900 55.950 ;
        RECT 121.950 54.150 123.750 55.950 ;
        RECT 135.000 52.200 135.900 55.950 ;
        RECT 137.100 54.150 138.900 55.950 ;
        RECT 143.100 54.150 144.900 55.950 ;
        RECT 158.250 54.150 160.050 55.950 ;
        RECT 135.000 51.000 138.300 52.200 ;
        RECT 116.700 49.800 120.900 50.700 ;
        RECT 116.700 42.600 118.500 49.800 ;
        RECT 121.800 42.000 123.600 48.600 ;
        RECT 136.500 42.600 138.300 51.000 ;
        RECT 143.100 42.000 144.900 51.600 ;
        RECT 161.100 50.700 162.300 55.950 ;
        RECT 164.100 54.150 165.900 55.950 ;
        RECT 161.100 49.800 165.300 50.700 ;
        RECT 158.400 42.000 160.200 48.600 ;
        RECT 163.500 42.600 165.300 49.800 ;
        RECT 176.700 45.600 177.900 55.950 ;
        RECT 195.000 52.200 195.900 55.950 ;
        RECT 197.100 54.150 198.900 55.950 ;
        RECT 203.100 54.150 204.900 55.950 ;
        RECT 218.100 54.150 219.900 55.950 ;
        RECT 224.250 54.150 226.050 55.950 ;
        RECT 195.000 51.000 198.300 52.200 ;
        RECT 176.100 42.600 177.900 45.600 ;
        RECT 179.100 42.000 180.900 45.600 ;
        RECT 196.500 42.600 198.300 51.000 ;
        RECT 203.100 42.000 204.900 51.600 ;
        RECT 208.950 51.450 211.050 52.050 ;
        RECT 223.950 51.450 226.050 52.050 ;
        RECT 208.950 50.550 226.050 51.450 ;
        RECT 208.950 49.950 211.050 50.550 ;
        RECT 223.950 49.950 226.050 50.550 ;
        RECT 227.700 48.600 228.600 55.950 ;
        RECT 242.100 54.150 243.900 55.950 ;
        RECT 245.700 51.600 246.900 55.950 ;
        RECT 248.100 54.150 249.900 55.950 ;
        RECT 264.000 52.200 264.900 55.950 ;
        RECT 266.100 54.150 267.900 55.950 ;
        RECT 272.100 54.150 273.900 55.950 ;
        RECT 287.100 54.150 288.900 55.950 ;
        RECT 245.700 50.700 249.300 51.600 ;
        RECT 264.000 51.000 267.300 52.200 ;
        RECT 219.000 42.000 220.800 48.600 ;
        RECT 223.500 47.400 228.600 48.600 ;
        RECT 229.950 48.450 232.050 49.050 ;
        RECT 235.950 48.450 238.050 49.050 ;
        RECT 229.950 47.550 238.050 48.450 ;
        RECT 223.500 42.600 225.300 47.400 ;
        RECT 229.950 46.950 232.050 47.550 ;
        RECT 235.950 46.950 238.050 47.550 ;
        RECT 239.100 47.700 246.900 49.050 ;
        RECT 226.500 42.000 228.300 45.600 ;
        RECT 239.100 42.600 240.900 47.700 ;
        RECT 242.100 42.000 243.900 46.800 ;
        RECT 245.100 42.600 246.900 47.700 ;
        RECT 248.100 48.600 249.300 50.700 ;
        RECT 248.100 42.600 249.900 48.600 ;
        RECT 265.500 42.600 267.300 51.000 ;
        RECT 272.100 42.000 273.900 51.600 ;
        RECT 290.700 50.700 291.900 55.950 ;
        RECT 292.950 54.150 294.750 55.950 ;
        RECT 308.250 54.150 310.050 55.950 ;
        RECT 287.700 49.800 291.900 50.700 ;
        RECT 311.100 50.700 312.300 55.950 ;
        RECT 314.100 54.150 315.900 55.950 ;
        RECT 320.550 51.900 321.450 58.950 ;
        RECT 329.400 58.050 330.300 65.400 ;
        RECT 334.950 58.050 336.750 59.850 ;
        RECT 354.000 58.050 354.900 70.200 ;
        RECT 374.100 65.400 375.900 77.400 ;
        RECT 377.100 66.300 378.900 77.400 ;
        RECT 380.100 67.200 381.900 78.000 ;
        RECT 383.100 66.300 384.900 77.400 ;
        RECT 398.100 71.400 399.900 77.400 ;
        RECT 401.100 72.000 402.900 78.000 ;
        RECT 377.100 65.400 384.900 66.300 ;
        RECT 399.000 71.100 399.900 71.400 ;
        RECT 404.100 71.400 405.900 77.400 ;
        RECT 407.100 71.400 408.900 78.000 ;
        RECT 419.100 71.400 420.900 78.000 ;
        RECT 422.100 71.400 423.900 77.400 ;
        RECT 425.100 72.000 426.900 78.000 ;
        RECT 404.100 71.100 405.600 71.400 ;
        RECT 399.000 70.200 405.600 71.100 ;
        RECT 422.400 71.100 423.900 71.400 ;
        RECT 428.100 71.400 429.900 77.400 ;
        RECT 440.700 71.400 442.500 78.000 ;
        RECT 428.100 71.100 429.000 71.400 ;
        RECT 422.400 70.200 429.000 71.100 ;
        RECT 361.950 63.450 364.050 64.050 ;
        RECT 370.950 63.450 373.050 64.050 ;
        RECT 361.950 62.550 373.050 63.450 ;
        RECT 361.950 61.950 364.050 62.550 ;
        RECT 370.950 61.950 373.050 62.550 ;
        RECT 359.100 58.050 360.900 59.850 ;
        RECT 374.400 58.050 375.300 65.400 ;
        RECT 379.950 58.050 381.750 59.850 ;
        RECT 399.000 58.050 399.900 70.200 ;
        RECT 414.000 60.450 418.050 61.050 ;
        RECT 404.100 58.050 405.900 59.850 ;
        RECT 413.550 58.950 418.050 60.450 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 400.950 55.950 403.050 58.050 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 311.100 49.800 315.300 50.700 ;
        RECT 319.950 49.800 322.050 51.900 ;
        RECT 287.700 42.600 289.500 49.800 ;
        RECT 292.800 42.000 294.600 48.600 ;
        RECT 308.400 42.000 310.200 48.600 ;
        RECT 313.500 42.600 315.300 49.800 ;
        RECT 329.400 48.600 330.300 55.950 ;
        RECT 331.950 54.150 333.750 55.950 ;
        RECT 338.100 54.150 339.900 55.950 ;
        RECT 354.000 52.200 354.900 55.950 ;
        RECT 356.100 54.150 357.900 55.950 ;
        RECT 362.100 54.150 363.900 55.950 ;
        RECT 354.000 51.000 357.300 52.200 ;
        RECT 329.400 47.400 334.500 48.600 ;
        RECT 329.700 42.000 331.500 45.600 ;
        RECT 332.700 42.600 334.500 47.400 ;
        RECT 337.200 42.000 339.000 48.600 ;
        RECT 355.500 42.600 357.300 51.000 ;
        RECT 362.100 42.000 363.900 51.600 ;
        RECT 374.400 48.600 375.300 55.950 ;
        RECT 376.950 54.150 378.750 55.950 ;
        RECT 383.100 54.150 384.900 55.950 ;
        RECT 399.000 52.200 399.900 55.950 ;
        RECT 401.100 54.150 402.900 55.950 ;
        RECT 407.100 54.150 408.900 55.950 ;
        RECT 413.550 55.050 414.450 58.950 ;
        RECT 422.100 58.050 423.900 59.850 ;
        RECT 428.100 58.050 429.000 70.200 ;
        RECT 441.000 68.100 442.800 69.900 ;
        RECT 443.700 66.900 445.500 77.400 ;
        RECT 443.100 65.400 445.500 66.900 ;
        RECT 448.800 65.400 450.600 78.000 ;
        RECT 461.400 65.400 463.200 78.000 ;
        RECT 466.500 66.900 468.300 77.400 ;
        RECT 469.500 71.400 471.300 78.000 ;
        RECT 485.100 71.400 486.900 77.400 ;
        RECT 488.100 72.000 489.900 78.000 ;
        RECT 486.000 71.100 486.900 71.400 ;
        RECT 491.100 71.400 492.900 77.400 ;
        RECT 494.100 71.400 495.900 78.000 ;
        RECT 509.100 71.400 510.900 77.400 ;
        RECT 512.100 71.400 513.900 78.000 ;
        RECT 491.100 71.100 492.600 71.400 ;
        RECT 486.000 70.200 492.600 71.100 ;
        RECT 469.200 68.100 471.000 69.900 ;
        RECT 466.500 65.400 468.900 66.900 ;
        RECT 443.100 58.050 444.300 65.400 ;
        RECT 445.950 63.450 448.050 64.050 ;
        RECT 463.950 63.450 466.050 64.050 ;
        RECT 445.950 62.550 466.050 63.450 ;
        RECT 445.950 61.950 448.050 62.550 ;
        RECT 463.950 61.950 466.050 62.550 ;
        RECT 449.100 58.050 450.900 59.850 ;
        RECT 461.100 58.050 462.900 59.850 ;
        RECT 467.700 58.050 468.900 65.400 ;
        RECT 486.000 58.050 486.900 70.200 ;
        RECT 491.100 58.050 492.900 59.850 ;
        RECT 509.700 58.050 510.900 71.400 ;
        RECT 524.100 65.400 525.900 77.400 ;
        RECT 527.100 66.300 528.900 77.400 ;
        RECT 530.100 67.200 531.900 78.000 ;
        RECT 533.100 66.300 534.900 77.400 ;
        RECT 527.100 65.400 534.900 66.300 ;
        RECT 548.100 66.300 549.900 77.400 ;
        RECT 551.100 67.200 552.900 78.000 ;
        RECT 554.100 66.300 555.900 77.400 ;
        RECT 548.100 65.400 555.900 66.300 ;
        RECT 557.100 65.400 558.900 77.400 ;
        RECT 572.100 71.400 573.900 78.000 ;
        RECT 575.100 71.400 576.900 77.400 ;
        RECT 578.100 72.000 579.900 78.000 ;
        RECT 575.400 71.100 576.900 71.400 ;
        RECT 581.100 71.400 582.900 77.400 ;
        RECT 581.100 71.100 582.000 71.400 ;
        RECT 575.400 70.200 582.000 71.100 ;
        RECT 512.100 58.050 513.900 59.850 ;
        RECT 524.400 58.050 525.300 65.400 ;
        RECT 529.950 58.050 531.750 59.850 ;
        RECT 551.250 58.050 553.050 59.850 ;
        RECT 557.700 58.050 558.600 65.400 ;
        RECT 575.100 58.050 576.900 59.850 ;
        RECT 581.100 58.050 582.000 70.200 ;
        RECT 593.100 65.400 594.900 77.400 ;
        RECT 596.100 66.300 597.900 77.400 ;
        RECT 599.100 67.200 600.900 78.000 ;
        RECT 602.100 66.300 603.900 77.400 ;
        RECT 614.100 71.400 615.900 78.000 ;
        RECT 617.100 71.400 618.900 77.400 ;
        RECT 620.100 72.000 621.900 78.000 ;
        RECT 617.400 71.100 618.900 71.400 ;
        RECT 623.100 71.400 624.900 77.400 ;
        RECT 635.100 71.400 636.900 78.000 ;
        RECT 638.100 71.400 639.900 77.400 ;
        RECT 641.100 72.000 642.900 78.000 ;
        RECT 623.100 71.100 624.000 71.400 ;
        RECT 617.400 70.200 624.000 71.100 ;
        RECT 638.400 71.100 639.900 71.400 ;
        RECT 644.100 71.400 645.900 77.400 ;
        RECT 656.700 71.400 658.500 78.000 ;
        RECT 644.100 71.100 645.000 71.400 ;
        RECT 638.400 70.200 645.000 71.100 ;
        RECT 596.100 65.400 603.900 66.300 ;
        RECT 593.400 58.050 594.300 65.400 ;
        RECT 598.950 58.050 600.750 59.850 ;
        RECT 617.100 58.050 618.900 59.850 ;
        RECT 623.100 58.050 624.000 70.200 ;
        RECT 638.100 58.050 639.900 59.850 ;
        RECT 644.100 58.050 645.000 70.200 ;
        RECT 657.000 68.100 658.800 69.900 ;
        RECT 659.700 66.900 661.500 77.400 ;
        RECT 659.100 65.400 661.500 66.900 ;
        RECT 664.800 65.400 666.600 78.000 ;
        RECT 680.400 65.400 682.200 78.000 ;
        RECT 685.500 66.900 687.300 77.400 ;
        RECT 688.500 71.400 690.300 78.000 ;
        RECT 688.200 68.100 690.000 69.900 ;
        RECT 685.500 65.400 687.900 66.900 ;
        RECT 704.100 65.400 705.900 78.000 ;
        RECT 709.200 66.600 711.000 77.400 ;
        RECT 722.100 71.400 723.900 78.000 ;
        RECT 725.100 71.400 726.900 77.400 ;
        RECT 707.400 65.400 711.000 66.600 ;
        RECT 659.100 58.050 660.300 65.400 ;
        RECT 665.100 58.050 666.900 59.850 ;
        RECT 680.100 58.050 681.900 59.850 ;
        RECT 686.700 58.050 687.900 65.400 ;
        RECT 704.250 58.050 706.050 59.850 ;
        RECT 707.400 58.050 708.300 65.400 ;
        RECT 710.100 58.050 711.900 59.850 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 448.950 55.950 451.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 580.950 55.950 583.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 722.100 55.950 724.200 58.050 ;
        RECT 409.950 53.550 414.450 55.050 ;
        RECT 419.100 54.150 420.900 55.950 ;
        RECT 425.100 54.150 426.900 55.950 ;
        RECT 409.950 52.950 414.000 53.550 ;
        RECT 428.100 52.200 429.000 55.950 ;
        RECT 440.100 54.150 441.900 55.950 ;
        RECT 399.000 51.000 402.300 52.200 ;
        RECT 374.400 47.400 379.500 48.600 ;
        RECT 374.700 42.000 376.500 45.600 ;
        RECT 377.700 42.600 379.500 47.400 ;
        RECT 382.200 42.000 384.000 48.600 ;
        RECT 385.950 45.450 388.050 46.050 ;
        RECT 394.950 45.450 397.050 46.050 ;
        RECT 385.950 44.550 397.050 45.450 ;
        RECT 385.950 43.950 388.050 44.550 ;
        RECT 394.950 43.950 397.050 44.550 ;
        RECT 400.500 42.600 402.300 51.000 ;
        RECT 407.100 42.000 408.900 51.600 ;
        RECT 419.100 42.000 420.900 51.600 ;
        RECT 425.700 51.000 429.000 52.200 ;
        RECT 443.100 51.600 444.300 55.950 ;
        RECT 446.100 54.150 447.900 55.950 ;
        RECT 464.100 54.150 465.900 55.950 ;
        RECT 425.700 42.600 427.500 51.000 ;
        RECT 440.700 50.700 444.300 51.600 ;
        RECT 467.700 51.600 468.900 55.950 ;
        RECT 470.100 54.150 471.900 55.950 ;
        RECT 486.000 52.200 486.900 55.950 ;
        RECT 488.100 54.150 489.900 55.950 ;
        RECT 494.100 54.150 495.900 55.950 ;
        RECT 467.700 50.700 471.300 51.600 ;
        RECT 486.000 51.000 489.300 52.200 ;
        RECT 440.700 48.600 441.900 50.700 ;
        RECT 440.100 42.600 441.900 48.600 ;
        RECT 443.100 47.700 450.900 49.050 ;
        RECT 443.100 42.600 444.900 47.700 ;
        RECT 446.100 42.000 447.900 46.800 ;
        RECT 449.100 42.600 450.900 47.700 ;
        RECT 461.100 47.700 468.900 49.050 ;
        RECT 461.100 42.600 462.900 47.700 ;
        RECT 464.100 42.000 465.900 46.800 ;
        RECT 467.100 42.600 468.900 47.700 ;
        RECT 470.100 48.600 471.300 50.700 ;
        RECT 470.100 42.600 471.900 48.600 ;
        RECT 487.500 42.600 489.300 51.000 ;
        RECT 494.100 42.000 495.900 51.600 ;
        RECT 509.700 45.600 510.900 55.950 ;
        RECT 524.400 48.600 525.300 55.950 ;
        RECT 526.950 54.150 528.750 55.950 ;
        RECT 533.100 54.150 534.900 55.950 ;
        RECT 548.100 54.150 549.900 55.950 ;
        RECT 554.250 54.150 556.050 55.950 ;
        RECT 529.950 51.450 532.050 52.050 ;
        RECT 550.950 51.450 553.050 52.050 ;
        RECT 529.950 50.550 553.050 51.450 ;
        RECT 529.950 49.950 532.050 50.550 ;
        RECT 550.950 49.950 553.050 50.550 ;
        RECT 557.700 48.600 558.600 55.950 ;
        RECT 572.100 54.150 573.900 55.950 ;
        RECT 578.100 54.150 579.900 55.950 ;
        RECT 581.100 52.200 582.000 55.950 ;
        RECT 524.400 47.400 529.500 48.600 ;
        RECT 509.100 42.600 510.900 45.600 ;
        RECT 512.100 42.000 513.900 45.600 ;
        RECT 524.700 42.000 526.500 45.600 ;
        RECT 527.700 42.600 529.500 47.400 ;
        RECT 532.200 42.000 534.000 48.600 ;
        RECT 549.000 42.000 550.800 48.600 ;
        RECT 553.500 47.400 558.600 48.600 ;
        RECT 553.500 42.600 555.300 47.400 ;
        RECT 556.500 42.000 558.300 45.600 ;
        RECT 572.100 42.000 573.900 51.600 ;
        RECT 578.700 51.000 582.000 52.200 ;
        RECT 578.700 42.600 580.500 51.000 ;
        RECT 593.400 48.600 594.300 55.950 ;
        RECT 595.950 54.150 597.750 55.950 ;
        RECT 602.100 54.150 603.900 55.950 ;
        RECT 614.100 54.150 615.900 55.950 ;
        RECT 620.100 54.150 621.900 55.950 ;
        RECT 623.100 52.200 624.000 55.950 ;
        RECT 635.100 54.150 636.900 55.950 ;
        RECT 641.100 54.150 642.900 55.950 ;
        RECT 644.100 52.200 645.000 55.950 ;
        RECT 656.100 54.150 657.900 55.950 ;
        RECT 595.950 51.450 598.050 52.050 ;
        RECT 610.950 51.450 613.050 52.050 ;
        RECT 595.950 50.550 613.050 51.450 ;
        RECT 595.950 49.950 598.050 50.550 ;
        RECT 610.950 49.950 613.050 50.550 ;
        RECT 593.400 47.400 598.500 48.600 ;
        RECT 593.700 42.000 595.500 45.600 ;
        RECT 596.700 42.600 598.500 47.400 ;
        RECT 601.200 42.000 603.000 48.600 ;
        RECT 614.100 42.000 615.900 51.600 ;
        RECT 620.700 51.000 624.000 52.200 ;
        RECT 620.700 42.600 622.500 51.000 ;
        RECT 635.100 42.000 636.900 51.600 ;
        RECT 641.700 51.000 645.000 52.200 ;
        RECT 659.100 51.600 660.300 55.950 ;
        RECT 662.100 54.150 663.900 55.950 ;
        RECT 683.100 54.150 684.900 55.950 ;
        RECT 641.700 42.600 643.500 51.000 ;
        RECT 656.700 50.700 660.300 51.600 ;
        RECT 686.700 51.600 687.900 55.950 ;
        RECT 689.100 54.150 690.900 55.950 ;
        RECT 686.700 50.700 690.300 51.600 ;
        RECT 656.700 48.600 657.900 50.700 ;
        RECT 656.100 42.600 657.900 48.600 ;
        RECT 659.100 47.700 666.900 49.050 ;
        RECT 659.100 42.600 660.900 47.700 ;
        RECT 662.100 42.000 663.900 46.800 ;
        RECT 665.100 42.600 666.900 47.700 ;
        RECT 680.100 47.700 687.900 49.050 ;
        RECT 680.100 42.600 681.900 47.700 ;
        RECT 683.100 42.000 684.900 46.800 ;
        RECT 686.100 42.600 687.900 47.700 ;
        RECT 689.100 48.600 690.300 50.700 ;
        RECT 689.100 42.600 690.900 48.600 ;
        RECT 707.400 45.600 708.300 55.950 ;
        RECT 722.250 54.150 724.050 55.950 ;
        RECT 709.950 51.450 712.050 52.050 ;
        RECT 715.950 51.450 718.050 52.050 ;
        RECT 709.950 50.550 718.050 51.450 ;
        RECT 725.100 51.300 726.000 71.400 ;
        RECT 728.100 66.000 729.900 78.000 ;
        RECT 731.100 65.400 732.900 77.400 ;
        RECT 743.400 65.400 745.200 78.000 ;
        RECT 748.500 66.900 750.300 77.400 ;
        RECT 751.500 71.400 753.300 78.000 ;
        RECT 764.100 71.400 765.900 78.000 ;
        RECT 767.100 71.400 768.900 77.400 ;
        RECT 751.200 68.100 753.000 69.900 ;
        RECT 748.500 65.400 750.900 66.900 ;
        RECT 727.200 58.050 729.000 59.850 ;
        RECT 731.400 58.050 732.300 65.400 ;
        RECT 743.100 58.050 744.900 59.850 ;
        RECT 749.700 58.050 750.900 65.400 ;
        RECT 764.100 58.050 765.900 59.850 ;
        RECT 767.100 58.050 768.300 71.400 ;
        RECT 782.400 65.400 784.200 78.000 ;
        RECT 787.500 66.900 789.300 77.400 ;
        RECT 790.500 71.400 792.300 78.000 ;
        RECT 790.200 68.100 792.000 69.900 ;
        RECT 787.500 65.400 789.900 66.900 ;
        RECT 806.400 65.400 808.200 78.000 ;
        RECT 811.500 66.900 813.300 77.400 ;
        RECT 814.500 71.400 816.300 78.000 ;
        RECT 814.200 68.100 816.000 69.900 ;
        RECT 830.100 67.500 831.900 77.400 ;
        RECT 833.100 68.400 834.900 78.000 ;
        RECT 836.100 76.500 843.900 77.400 ;
        RECT 836.100 67.500 837.900 76.500 ;
        RECT 811.500 65.400 813.900 66.900 ;
        RECT 830.100 66.600 837.900 67.500 ;
        RECT 839.100 67.800 840.900 75.600 ;
        RECT 842.100 68.700 843.900 76.500 ;
        RECT 845.100 76.500 852.900 77.400 ;
        RECT 845.100 67.800 846.900 76.500 ;
        RECT 839.100 66.900 846.900 67.800 ;
        RECT 848.100 67.800 849.900 75.600 ;
        RECT 782.100 58.050 783.900 59.850 ;
        RECT 788.700 58.050 789.900 65.400 ;
        RECT 806.100 58.050 807.900 59.850 ;
        RECT 812.700 58.050 813.900 65.400 ;
        RECT 814.950 63.450 817.050 64.050 ;
        RECT 823.950 63.450 826.050 64.050 ;
        RECT 814.950 62.550 826.050 63.450 ;
        RECT 814.950 61.950 817.050 62.550 ;
        RECT 823.950 61.950 826.050 62.550 ;
        RECT 833.100 58.050 834.900 59.850 ;
        RECT 842.250 58.050 844.050 59.850 ;
        RECT 848.100 58.050 849.300 67.800 ;
        RECT 851.100 67.200 852.900 76.500 ;
        RECT 863.100 66.300 864.900 77.400 ;
        RECT 866.100 67.200 867.900 78.000 ;
        RECT 869.100 66.300 870.900 77.400 ;
        RECT 863.100 65.400 870.900 66.300 ;
        RECT 872.100 65.400 873.900 77.400 ;
        RECT 874.950 75.450 877.050 76.050 ;
        RECT 883.950 75.450 886.050 76.050 ;
        RECT 874.950 74.550 886.050 75.450 ;
        RECT 874.950 73.950 877.050 74.550 ;
        RECT 883.950 73.950 886.050 74.550 ;
        RECT 887.400 65.400 889.200 78.000 ;
        RECT 892.500 66.900 894.300 77.400 ;
        RECT 895.500 71.400 897.300 78.000 ;
        RECT 908.100 71.400 909.900 78.000 ;
        RECT 911.100 71.400 912.900 77.400 ;
        RECT 914.100 72.000 915.900 78.000 ;
        RECT 911.400 71.100 912.900 71.400 ;
        RECT 917.100 71.400 918.900 77.400 ;
        RECT 917.100 71.100 918.000 71.400 ;
        RECT 911.400 70.200 918.000 71.100 ;
        RECT 895.200 68.100 897.000 69.900 ;
        RECT 892.500 65.400 894.900 66.900 ;
        RECT 868.950 63.450 871.050 64.200 ;
        RECT 854.550 62.550 871.050 63.450 ;
        RECT 727.500 55.950 729.600 58.050 ;
        RECT 730.800 55.950 732.900 58.050 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 745.950 55.950 748.050 58.050 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 811.950 55.950 814.050 58.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 832.800 55.950 834.900 58.050 ;
        RECT 838.950 55.950 841.050 58.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 847.500 55.950 849.600 58.050 ;
        RECT 709.950 49.950 712.050 50.550 ;
        RECT 715.950 49.950 718.050 50.550 ;
        RECT 722.100 50.400 730.500 51.300 ;
        RECT 704.100 42.000 705.900 45.600 ;
        RECT 707.100 42.600 708.900 45.600 ;
        RECT 710.100 42.000 711.900 45.600 ;
        RECT 722.100 42.600 723.900 50.400 ;
        RECT 728.700 49.500 730.500 50.400 ;
        RECT 731.400 48.600 732.300 55.950 ;
        RECT 746.100 54.150 747.900 55.950 ;
        RECT 749.700 51.600 750.900 55.950 ;
        RECT 752.100 54.150 753.900 55.950 ;
        RECT 749.700 50.700 753.300 51.600 ;
        RECT 726.600 42.000 728.400 48.600 ;
        RECT 729.600 46.800 732.300 48.600 ;
        RECT 743.100 47.700 750.900 49.050 ;
        RECT 729.600 42.600 731.400 46.800 ;
        RECT 743.100 42.600 744.900 47.700 ;
        RECT 746.100 42.000 747.900 46.800 ;
        RECT 749.100 42.600 750.900 47.700 ;
        RECT 752.100 48.600 753.300 50.700 ;
        RECT 752.100 42.600 753.900 48.600 ;
        RECT 767.100 45.600 768.300 55.950 ;
        RECT 785.100 54.150 786.900 55.950 ;
        RECT 788.700 51.600 789.900 55.950 ;
        RECT 791.100 54.150 792.900 55.950 ;
        RECT 809.100 54.150 810.900 55.950 ;
        RECT 812.700 51.600 813.900 55.950 ;
        RECT 815.100 54.150 816.900 55.950 ;
        RECT 838.950 54.150 840.750 55.950 ;
        RECT 788.700 50.700 792.300 51.600 ;
        RECT 812.700 50.700 816.300 51.600 ;
        RECT 782.100 47.700 789.900 49.050 ;
        RECT 764.100 42.000 765.900 45.600 ;
        RECT 767.100 42.600 768.900 45.600 ;
        RECT 782.100 42.600 783.900 47.700 ;
        RECT 785.100 42.000 786.900 46.800 ;
        RECT 788.100 42.600 789.900 47.700 ;
        RECT 791.100 48.600 792.300 50.700 ;
        RECT 791.100 42.600 792.900 48.600 ;
        RECT 806.100 47.700 813.900 49.050 ;
        RECT 806.100 42.600 807.900 47.700 ;
        RECT 809.100 42.000 810.900 46.800 ;
        RECT 812.100 42.600 813.900 47.700 ;
        RECT 815.100 48.600 816.300 50.700 ;
        RECT 820.950 51.450 823.050 52.050 ;
        RECT 832.950 51.450 835.050 52.050 ;
        RECT 820.950 50.550 835.050 51.450 ;
        RECT 820.950 49.950 823.050 50.550 ;
        RECT 832.950 49.950 835.050 50.550 ;
        RECT 815.100 42.600 816.900 48.600 ;
        RECT 848.100 47.400 849.300 55.950 ;
        RECT 854.550 51.900 855.450 62.550 ;
        RECT 868.950 62.100 871.050 62.550 ;
        RECT 866.250 58.050 868.050 59.850 ;
        RECT 872.700 58.050 873.600 65.400 ;
        RECT 887.100 58.050 888.900 59.850 ;
        RECT 893.700 58.050 894.900 65.400 ;
        RECT 898.950 60.450 903.000 61.050 ;
        RECT 898.950 58.950 903.450 60.450 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 886.950 55.950 889.050 58.050 ;
        RECT 889.950 55.950 892.050 58.050 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 863.100 54.150 864.900 55.950 ;
        RECT 869.250 54.150 871.050 55.950 ;
        RECT 853.950 49.800 856.050 51.900 ;
        RECT 872.700 48.600 873.600 55.950 ;
        RECT 890.100 54.150 891.900 55.950 ;
        RECT 893.700 51.600 894.900 55.950 ;
        RECT 896.100 54.150 897.900 55.950 ;
        RECT 902.550 55.050 903.450 58.950 ;
        RECT 911.100 58.050 912.900 59.850 ;
        RECT 917.100 58.050 918.000 70.200 ;
        RECT 907.950 55.950 910.050 58.050 ;
        RECT 910.950 55.950 913.050 58.050 ;
        RECT 913.950 55.950 916.050 58.050 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 902.550 53.550 907.050 55.050 ;
        RECT 908.100 54.150 909.900 55.950 ;
        RECT 914.100 54.150 915.900 55.950 ;
        RECT 903.000 52.950 907.050 53.550 ;
        RECT 917.100 52.200 918.000 55.950 ;
        RECT 893.700 50.700 897.300 51.600 ;
        RECT 836.700 46.500 849.300 47.400 ;
        RECT 836.700 45.600 837.600 46.500 ;
        RECT 843.900 45.600 844.800 46.500 ;
        RECT 832.800 42.000 834.900 45.600 ;
        RECT 836.100 42.600 837.900 45.600 ;
        RECT 839.100 42.000 840.900 45.600 ;
        RECT 842.100 42.600 844.800 45.600 ;
        RECT 864.000 42.000 865.800 48.600 ;
        RECT 868.500 47.400 873.600 48.600 ;
        RECT 887.100 47.700 894.900 49.050 ;
        RECT 868.500 42.600 870.300 47.400 ;
        RECT 871.500 42.000 873.300 45.600 ;
        RECT 887.100 42.600 888.900 47.700 ;
        RECT 890.100 42.000 891.900 46.800 ;
        RECT 893.100 42.600 894.900 47.700 ;
        RECT 896.100 48.600 897.300 50.700 ;
        RECT 896.100 42.600 897.900 48.600 ;
        RECT 908.100 42.000 909.900 51.600 ;
        RECT 914.700 51.000 918.000 52.200 ;
        RECT 914.700 42.600 916.500 51.000 ;
        RECT 14.100 35.400 15.900 38.400 ;
        RECT 14.100 31.500 15.300 35.400 ;
        RECT 17.100 32.400 18.900 39.000 ;
        RECT 20.100 32.400 21.900 38.400 ;
        RECT 14.100 30.600 19.800 31.500 ;
        RECT 18.000 29.700 19.800 30.600 ;
        RECT 14.400 22.950 16.500 25.050 ;
        RECT 14.400 21.150 16.200 22.950 ;
        RECT 18.000 18.300 18.900 29.700 ;
        RECT 20.700 25.050 21.900 32.400 ;
        RECT 19.800 22.950 21.900 25.050 ;
        RECT 18.000 17.400 19.800 18.300 ;
        RECT 14.100 16.500 19.800 17.400 ;
        RECT 14.100 9.600 15.300 16.500 ;
        RECT 20.700 15.600 21.900 22.950 ;
        RECT 14.100 3.600 15.900 9.600 ;
        RECT 17.100 3.000 18.900 13.800 ;
        RECT 20.100 3.600 21.900 15.600 ;
        RECT 32.100 32.400 33.900 38.400 ;
        RECT 35.100 32.400 36.900 39.000 ;
        RECT 38.100 35.400 39.900 38.400 ;
        RECT 32.100 25.050 33.300 32.400 ;
        RECT 38.700 31.500 39.900 35.400 ;
        RECT 34.200 30.600 39.900 31.500 ;
        RECT 50.100 32.400 51.900 38.400 ;
        RECT 53.100 32.400 54.900 39.000 ;
        RECT 56.100 35.400 57.900 38.400 ;
        RECT 71.100 35.400 72.900 38.400 ;
        RECT 74.100 35.400 75.900 39.000 ;
        RECT 89.100 35.400 90.900 38.400 ;
        RECT 34.200 29.700 36.000 30.600 ;
        RECT 32.100 22.950 34.200 25.050 ;
        RECT 32.100 15.600 33.300 22.950 ;
        RECT 35.100 18.300 36.000 29.700 ;
        RECT 50.100 25.050 51.300 32.400 ;
        RECT 56.700 31.500 57.900 35.400 ;
        RECT 52.200 30.600 57.900 31.500 ;
        RECT 52.200 29.700 54.000 30.600 ;
        RECT 37.500 22.950 39.600 25.050 ;
        RECT 37.800 21.150 39.600 22.950 ;
        RECT 50.100 22.950 52.200 25.050 ;
        RECT 34.200 17.400 36.000 18.300 ;
        RECT 34.200 16.500 39.900 17.400 ;
        RECT 32.100 3.600 33.900 15.600 ;
        RECT 35.100 3.000 36.900 13.800 ;
        RECT 38.700 9.600 39.900 16.500 ;
        RECT 38.100 3.600 39.900 9.600 ;
        RECT 50.100 15.600 51.300 22.950 ;
        RECT 53.100 18.300 54.000 29.700 ;
        RECT 71.700 25.050 72.900 35.400 ;
        RECT 89.100 31.500 90.300 35.400 ;
        RECT 92.100 32.400 93.900 39.000 ;
        RECT 95.100 32.400 96.900 38.400 ;
        RECT 107.400 32.400 109.200 39.000 ;
        RECT 89.100 30.600 94.800 31.500 ;
        RECT 93.000 29.700 94.800 30.600 ;
        RECT 55.500 22.950 57.600 25.050 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 89.400 22.950 91.500 25.050 ;
        RECT 55.800 21.150 57.600 22.950 ;
        RECT 52.200 17.400 54.000 18.300 ;
        RECT 52.200 16.500 57.900 17.400 ;
        RECT 50.100 3.600 51.900 15.600 ;
        RECT 53.100 3.000 54.900 13.800 ;
        RECT 56.700 9.600 57.900 16.500 ;
        RECT 71.700 9.600 72.900 22.950 ;
        RECT 74.100 21.150 75.900 22.950 ;
        RECT 89.400 21.150 91.200 22.950 ;
        RECT 93.000 18.300 93.900 29.700 ;
        RECT 95.700 25.050 96.900 32.400 ;
        RECT 112.500 31.200 114.300 38.400 ;
        RECT 110.100 30.300 114.300 31.200 ;
        RECT 107.250 25.050 109.050 26.850 ;
        RECT 110.100 25.050 111.300 30.300 ;
        RECT 127.500 30.000 129.300 38.400 ;
        RECT 126.000 28.800 129.300 30.000 ;
        RECT 134.100 29.400 135.900 39.000 ;
        RECT 149.100 32.400 150.900 38.400 ;
        RECT 152.100 33.000 153.900 39.000 ;
        RECT 158.700 38.400 159.900 39.000 ;
        RECT 155.100 35.400 156.900 38.400 ;
        RECT 158.100 35.400 159.900 38.400 ;
        RECT 113.100 25.050 114.900 26.850 ;
        RECT 126.000 25.050 126.900 28.800 ;
        RECT 128.100 25.050 129.900 26.850 ;
        RECT 134.100 25.050 135.900 26.850 ;
        RECT 149.100 25.050 150.000 32.400 ;
        RECT 155.700 31.200 156.600 35.400 ;
        RECT 151.200 30.300 156.600 31.200 ;
        RECT 151.200 29.400 153.300 30.300 ;
        RECT 173.100 29.400 174.900 39.000 ;
        RECT 179.700 30.000 181.500 38.400 ;
        RECT 194.100 35.400 195.900 38.400 ;
        RECT 197.100 35.400 198.900 39.000 ;
        RECT 94.800 22.950 96.900 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 149.100 22.950 151.200 25.050 ;
        RECT 93.000 17.400 94.800 18.300 ;
        RECT 89.100 16.500 94.800 17.400 ;
        RECT 89.100 9.600 90.300 16.500 ;
        RECT 95.700 15.600 96.900 22.950 ;
        RECT 56.100 3.600 57.900 9.600 ;
        RECT 71.100 3.600 72.900 9.600 ;
        RECT 74.100 3.000 75.900 9.600 ;
        RECT 89.100 3.600 90.900 9.600 ;
        RECT 92.100 3.000 93.900 13.800 ;
        RECT 95.100 3.600 96.900 15.600 ;
        RECT 110.100 9.600 111.300 22.950 ;
        RECT 126.000 10.800 126.900 22.950 ;
        RECT 131.100 21.150 132.900 22.950 ;
        RECT 133.950 18.450 136.050 19.050 ;
        RECT 145.950 18.450 148.050 19.050 ;
        RECT 133.950 17.550 148.050 18.450 ;
        RECT 133.950 16.950 136.050 17.550 ;
        RECT 145.950 16.950 148.050 17.550 ;
        RECT 150.000 15.600 151.200 22.950 ;
        RECT 152.400 18.900 153.300 29.400 ;
        RECT 179.700 28.800 183.000 30.000 ;
        RECT 157.800 25.050 159.600 26.850 ;
        RECT 173.100 25.050 174.900 26.850 ;
        RECT 179.100 25.050 180.900 26.850 ;
        RECT 182.100 25.050 183.000 28.800 ;
        RECT 194.700 25.050 195.900 35.400 ;
        RECT 209.100 29.400 210.900 39.000 ;
        RECT 215.700 30.000 217.500 38.400 ;
        RECT 223.950 36.450 226.050 37.050 ;
        RECT 229.950 36.450 232.050 37.050 ;
        RECT 223.950 35.550 232.050 36.450 ;
        RECT 223.950 34.950 226.050 35.550 ;
        RECT 229.950 34.950 232.050 35.550 ;
        RECT 233.100 33.300 234.900 38.400 ;
        RECT 236.100 34.200 237.900 39.000 ;
        RECT 239.100 33.300 240.900 38.400 ;
        RECT 233.100 31.950 240.900 33.300 ;
        RECT 242.100 32.400 243.900 38.400 ;
        RECT 242.100 30.300 243.300 32.400 ;
        RECT 215.700 28.800 219.000 30.000 ;
        RECT 209.100 25.050 210.900 26.850 ;
        RECT 215.100 25.050 216.900 26.850 ;
        RECT 218.100 25.050 219.000 28.800 ;
        RECT 239.700 29.400 243.300 30.300 ;
        RECT 254.100 29.400 255.900 39.000 ;
        RECT 260.700 30.000 262.500 38.400 ;
        RECT 275.100 35.400 276.900 38.400 ;
        RECT 278.100 35.400 279.900 39.000 ;
        RECT 236.100 25.050 237.900 26.850 ;
        RECT 239.700 25.050 240.900 29.400 ;
        RECT 260.700 28.800 264.000 30.000 ;
        RECT 242.100 25.050 243.900 26.850 ;
        RECT 254.100 25.050 255.900 26.850 ;
        RECT 260.100 25.050 261.900 26.850 ;
        RECT 263.100 25.050 264.000 28.800 ;
        RECT 275.700 25.050 276.900 35.400 ;
        RECT 290.400 32.400 292.200 39.000 ;
        RECT 295.500 31.200 297.300 38.400 ;
        RECT 293.100 30.300 297.300 31.200 ;
        RECT 290.250 25.050 292.050 26.850 ;
        RECT 293.100 25.050 294.300 30.300 ;
        RECT 308.100 29.400 309.900 39.000 ;
        RECT 314.700 30.000 316.500 38.400 ;
        RECT 334.500 30.000 336.300 38.400 ;
        RECT 314.700 28.800 318.000 30.000 ;
        RECT 296.100 25.050 297.900 26.850 ;
        RECT 308.100 25.050 309.900 26.850 ;
        RECT 314.100 25.050 315.900 26.850 ;
        RECT 317.100 25.050 318.000 28.800 ;
        RECT 333.000 28.800 336.300 30.000 ;
        RECT 341.100 29.400 342.900 39.000 ;
        RECT 356.100 32.400 357.900 38.400 ;
        RECT 356.700 30.300 357.900 32.400 ;
        RECT 359.100 33.300 360.900 38.400 ;
        RECT 362.100 34.200 363.900 39.000 ;
        RECT 365.100 33.300 366.900 38.400 ;
        RECT 359.100 31.950 366.900 33.300 ;
        RECT 380.100 32.400 381.900 38.400 ;
        RECT 380.700 30.300 381.900 32.400 ;
        RECT 383.100 33.300 384.900 38.400 ;
        RECT 386.100 34.200 387.900 39.000 ;
        RECT 389.100 33.300 390.900 38.400 ;
        RECT 383.100 31.950 390.900 33.300 ;
        RECT 401.100 33.300 402.900 38.400 ;
        RECT 404.100 34.200 405.900 39.000 ;
        RECT 407.100 33.300 408.900 38.400 ;
        RECT 401.100 31.950 408.900 33.300 ;
        RECT 410.100 32.400 411.900 38.400 ;
        RECT 425.100 35.400 426.900 38.400 ;
        RECT 428.100 35.400 429.900 39.000 ;
        RECT 410.100 30.300 411.300 32.400 ;
        RECT 356.700 29.400 360.300 30.300 ;
        RECT 380.700 29.400 384.300 30.300 ;
        RECT 328.950 27.450 331.050 28.050 ;
        RECT 323.550 26.550 331.050 27.450 ;
        RECT 154.500 22.950 156.600 25.050 ;
        RECT 157.800 22.950 159.900 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 181.950 22.950 184.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 307.950 22.950 310.050 25.050 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 154.200 21.150 156.000 22.950 ;
        RECT 176.100 21.150 177.900 22.950 ;
        RECT 152.100 18.300 153.900 18.900 ;
        RECT 152.100 17.100 159.900 18.300 ;
        RECT 158.700 15.600 159.900 17.100 ;
        RECT 150.000 14.100 152.400 15.600 ;
        RECT 126.000 9.900 132.600 10.800 ;
        RECT 126.000 9.600 126.900 9.900 ;
        RECT 107.100 3.000 108.900 9.600 ;
        RECT 110.100 3.600 111.900 9.600 ;
        RECT 113.100 3.000 114.900 9.600 ;
        RECT 125.100 3.600 126.900 9.600 ;
        RECT 131.100 9.600 132.600 9.900 ;
        RECT 128.100 3.000 129.900 9.000 ;
        RECT 131.100 3.600 132.900 9.600 ;
        RECT 134.100 3.000 135.900 9.600 ;
        RECT 150.600 3.600 152.400 14.100 ;
        RECT 153.600 3.000 155.400 15.600 ;
        RECT 158.100 3.600 159.900 15.600 ;
        RECT 182.100 10.800 183.000 22.950 ;
        RECT 176.400 9.900 183.000 10.800 ;
        RECT 176.400 9.600 177.900 9.900 ;
        RECT 173.100 3.000 174.900 9.600 ;
        RECT 176.100 3.600 177.900 9.600 ;
        RECT 182.100 9.600 183.000 9.900 ;
        RECT 194.700 9.600 195.900 22.950 ;
        RECT 197.100 21.150 198.900 22.950 ;
        RECT 212.100 21.150 213.900 22.950 ;
        RECT 218.100 10.800 219.000 22.950 ;
        RECT 233.100 21.150 234.900 22.950 ;
        RECT 239.700 15.600 240.900 22.950 ;
        RECT 257.100 21.150 258.900 22.950 ;
        RECT 244.950 18.450 247.050 19.050 ;
        RECT 259.950 18.450 262.050 19.050 ;
        RECT 244.950 17.550 262.050 18.450 ;
        RECT 244.950 16.950 247.050 17.550 ;
        RECT 259.950 16.950 262.050 17.550 ;
        RECT 212.400 9.900 219.000 10.800 ;
        RECT 212.400 9.600 213.900 9.900 ;
        RECT 179.100 3.000 180.900 9.000 ;
        RECT 182.100 3.600 183.900 9.600 ;
        RECT 194.100 3.600 195.900 9.600 ;
        RECT 197.100 3.000 198.900 9.600 ;
        RECT 209.100 3.000 210.900 9.600 ;
        RECT 212.100 3.600 213.900 9.600 ;
        RECT 218.100 9.600 219.000 9.900 ;
        RECT 215.100 3.000 216.900 9.000 ;
        RECT 218.100 3.600 219.900 9.600 ;
        RECT 233.400 3.000 235.200 15.600 ;
        RECT 238.500 14.100 240.900 15.600 ;
        RECT 238.500 3.600 240.300 14.100 ;
        RECT 241.200 11.100 243.000 12.900 ;
        RECT 263.100 10.800 264.000 22.950 ;
        RECT 257.400 9.900 264.000 10.800 ;
        RECT 257.400 9.600 258.900 9.900 ;
        RECT 241.500 3.000 243.300 9.600 ;
        RECT 254.100 3.000 255.900 9.600 ;
        RECT 257.100 3.600 258.900 9.600 ;
        RECT 263.100 9.600 264.000 9.900 ;
        RECT 275.700 9.600 276.900 22.950 ;
        RECT 278.100 21.150 279.900 22.950 ;
        RECT 283.950 15.450 286.050 16.050 ;
        RECT 289.950 15.450 292.050 16.050 ;
        RECT 283.950 14.550 292.050 15.450 ;
        RECT 283.950 13.950 286.050 14.550 ;
        RECT 289.950 13.950 292.050 14.550 ;
        RECT 293.100 9.600 294.300 22.950 ;
        RECT 311.100 21.150 312.900 22.950 ;
        RECT 317.100 10.800 318.000 22.950 ;
        RECT 323.550 21.450 324.450 26.550 ;
        RECT 328.950 25.950 331.050 26.550 ;
        RECT 333.000 25.050 333.900 28.800 ;
        RECT 335.100 25.050 336.900 26.850 ;
        RECT 341.100 25.050 342.900 26.850 ;
        RECT 356.100 25.050 357.900 26.850 ;
        RECT 359.100 25.050 360.300 29.400 ;
        RECT 362.100 25.050 363.900 26.850 ;
        RECT 380.100 25.050 381.900 26.850 ;
        RECT 383.100 25.050 384.300 29.400 ;
        RECT 407.700 29.400 411.300 30.300 ;
        RECT 386.100 25.050 387.900 26.850 ;
        RECT 404.100 25.050 405.900 26.850 ;
        RECT 407.700 25.050 408.900 29.400 ;
        RECT 410.100 25.050 411.900 26.850 ;
        RECT 425.700 25.050 426.900 35.400 ;
        RECT 427.950 30.450 430.050 31.050 ;
        RECT 433.950 30.450 436.050 31.050 ;
        RECT 427.950 29.550 436.050 30.450 ;
        RECT 427.950 28.950 430.050 29.550 ;
        RECT 433.950 28.950 436.050 29.550 ;
        RECT 440.100 29.400 441.900 39.000 ;
        RECT 446.700 30.000 448.500 38.400 ;
        RECT 463.500 30.000 465.300 38.400 ;
        RECT 446.700 28.800 450.000 30.000 ;
        RECT 440.100 25.050 441.900 26.850 ;
        RECT 446.100 25.050 447.900 26.850 ;
        RECT 449.100 25.050 450.000 28.800 ;
        RECT 462.000 28.800 465.300 30.000 ;
        RECT 470.100 29.400 471.900 39.000 ;
        RECT 482.700 31.200 484.500 38.400 ;
        RECT 487.800 32.400 489.600 39.000 ;
        RECT 482.700 30.300 486.900 31.200 ;
        RECT 462.000 25.050 462.900 28.800 ;
        RECT 464.100 25.050 465.900 26.850 ;
        RECT 470.100 25.050 471.900 26.850 ;
        RECT 482.100 25.050 483.900 26.850 ;
        RECT 485.700 25.050 486.900 30.300 ;
        RECT 505.500 30.000 507.300 38.400 ;
        RECT 504.000 28.800 507.300 30.000 ;
        RECT 512.100 29.400 513.900 39.000 ;
        RECT 527.700 35.400 529.500 39.000 ;
        RECT 530.700 33.600 532.500 38.400 ;
        RECT 527.400 32.400 532.500 33.600 ;
        RECT 535.200 32.400 537.000 39.000 ;
        RECT 487.950 25.050 489.750 26.850 ;
        RECT 504.000 25.050 504.900 28.800 ;
        RECT 506.100 25.050 507.900 26.850 ;
        RECT 512.100 25.050 513.900 26.850 ;
        RECT 527.400 25.050 528.300 32.400 ;
        RECT 550.500 30.000 552.300 38.400 ;
        RECT 549.000 28.800 552.300 30.000 ;
        RECT 557.100 29.400 558.900 39.000 ;
        RECT 572.100 32.400 573.900 38.400 ;
        RECT 572.700 30.300 573.900 32.400 ;
        RECT 575.100 33.300 576.900 38.400 ;
        RECT 578.100 34.200 579.900 39.000 ;
        RECT 581.100 33.300 582.900 38.400 ;
        RECT 575.100 31.950 582.900 33.300 ;
        RECT 572.700 29.400 576.300 30.300 ;
        RECT 598.500 30.000 600.300 38.400 ;
        RECT 529.950 25.050 531.750 26.850 ;
        RECT 536.100 25.050 537.900 26.850 ;
        RECT 549.000 25.050 549.900 28.800 ;
        RECT 551.100 25.050 552.900 26.850 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 572.100 25.050 573.900 26.850 ;
        RECT 575.100 25.050 576.300 29.400 ;
        RECT 597.000 28.800 600.300 30.000 ;
        RECT 605.100 29.400 606.900 39.000 ;
        RECT 619.500 30.000 621.300 38.400 ;
        RECT 618.000 28.800 621.300 30.000 ;
        RECT 626.100 29.400 627.900 39.000 ;
        RECT 638.100 35.400 639.900 39.000 ;
        RECT 641.100 35.400 642.900 38.400 ;
        RECT 578.100 25.050 579.900 26.850 ;
        RECT 597.000 25.050 597.900 28.800 ;
        RECT 599.100 25.050 600.900 26.850 ;
        RECT 605.100 25.050 606.900 26.850 ;
        RECT 618.000 25.050 618.900 28.800 ;
        RECT 620.100 25.050 621.900 26.850 ;
        RECT 626.100 25.050 627.900 26.850 ;
        RECT 641.100 25.050 642.300 35.400 ;
        RECT 656.100 29.400 657.900 39.000 ;
        RECT 662.700 30.000 664.500 38.400 ;
        RECT 662.700 28.800 666.000 30.000 ;
        RECT 677.100 29.400 678.900 39.000 ;
        RECT 683.700 30.000 685.500 38.400 ;
        RECT 701.100 33.300 702.900 38.400 ;
        RECT 704.100 34.200 705.900 39.000 ;
        RECT 707.100 33.300 708.900 38.400 ;
        RECT 701.100 31.950 708.900 33.300 ;
        RECT 710.100 32.400 711.900 38.400 ;
        RECT 725.400 32.400 727.200 39.000 ;
        RECT 743.100 38.400 744.300 39.000 ;
        RECT 710.100 30.300 711.300 32.400 ;
        RECT 730.500 31.200 732.300 38.400 ;
        RECT 743.100 35.400 744.900 38.400 ;
        RECT 746.100 35.400 747.900 38.400 ;
        RECT 683.700 28.800 687.000 30.000 ;
        RECT 656.100 25.050 657.900 26.850 ;
        RECT 662.100 25.050 663.900 26.850 ;
        RECT 665.100 25.050 666.000 28.800 ;
        RECT 677.100 25.050 678.900 26.850 ;
        RECT 683.100 25.050 684.900 26.850 ;
        RECT 686.100 25.050 687.000 28.800 ;
        RECT 707.700 29.400 711.300 30.300 ;
        RECT 728.100 30.300 732.300 31.200 ;
        RECT 746.400 31.200 747.300 35.400 ;
        RECT 749.100 33.000 750.900 39.000 ;
        RECT 752.100 32.400 753.900 38.400 ;
        RECT 746.400 30.300 751.800 31.200 ;
        RECT 704.100 25.050 705.900 26.850 ;
        RECT 707.700 25.050 708.900 29.400 ;
        RECT 710.100 25.050 711.900 26.850 ;
        RECT 725.250 25.050 727.050 26.850 ;
        RECT 728.100 25.050 729.300 30.300 ;
        RECT 749.700 29.400 751.800 30.300 ;
        RECT 731.100 25.050 732.900 26.850 ;
        RECT 743.400 25.050 745.200 26.850 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 382.950 22.950 385.050 25.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 445.950 22.950 448.050 25.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 469.950 22.950 472.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 724.950 22.950 727.050 25.050 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 743.100 22.950 745.200 25.050 ;
        RECT 746.400 22.950 748.500 25.050 ;
        RECT 320.550 21.000 324.450 21.450 ;
        RECT 319.950 20.550 324.450 21.000 ;
        RECT 319.950 16.950 322.050 20.550 ;
        RECT 311.400 9.900 318.000 10.800 ;
        RECT 311.400 9.600 312.900 9.900 ;
        RECT 260.100 3.000 261.900 9.000 ;
        RECT 263.100 3.600 264.900 9.600 ;
        RECT 275.100 3.600 276.900 9.600 ;
        RECT 278.100 3.000 279.900 9.600 ;
        RECT 290.100 3.000 291.900 9.600 ;
        RECT 293.100 3.600 294.900 9.600 ;
        RECT 296.100 3.000 297.900 9.600 ;
        RECT 308.100 3.000 309.900 9.600 ;
        RECT 311.100 3.600 312.900 9.600 ;
        RECT 317.100 9.600 318.000 9.900 ;
        RECT 333.000 10.800 333.900 22.950 ;
        RECT 338.100 21.150 339.900 22.950 ;
        RECT 343.950 21.450 346.050 22.050 ;
        RECT 349.950 21.450 352.050 22.050 ;
        RECT 343.950 20.550 352.050 21.450 ;
        RECT 343.950 19.950 346.050 20.550 ;
        RECT 349.950 19.950 352.050 20.550 ;
        RECT 359.100 15.600 360.300 22.950 ;
        RECT 365.100 21.150 366.900 22.950 ;
        RECT 383.100 15.600 384.300 22.950 ;
        RECT 389.100 21.150 390.900 22.950 ;
        RECT 401.100 21.150 402.900 22.950 ;
        RECT 407.700 15.600 408.900 22.950 ;
        RECT 359.100 14.100 361.500 15.600 ;
        RECT 357.000 11.100 358.800 12.900 ;
        RECT 333.000 9.900 339.600 10.800 ;
        RECT 333.000 9.600 333.900 9.900 ;
        RECT 314.100 3.000 315.900 9.000 ;
        RECT 317.100 3.600 318.900 9.600 ;
        RECT 332.100 3.600 333.900 9.600 ;
        RECT 338.100 9.600 339.600 9.900 ;
        RECT 335.100 3.000 336.900 9.000 ;
        RECT 338.100 3.600 339.900 9.600 ;
        RECT 341.100 3.000 342.900 9.600 ;
        RECT 356.700 3.000 358.500 9.600 ;
        RECT 359.700 3.600 361.500 14.100 ;
        RECT 364.800 3.000 366.600 15.600 ;
        RECT 383.100 14.100 385.500 15.600 ;
        RECT 381.000 11.100 382.800 12.900 ;
        RECT 380.700 3.000 382.500 9.600 ;
        RECT 383.700 3.600 385.500 14.100 ;
        RECT 388.800 3.000 390.600 15.600 ;
        RECT 401.400 3.000 403.200 15.600 ;
        RECT 406.500 14.100 408.900 15.600 ;
        RECT 406.500 3.600 408.300 14.100 ;
        RECT 409.200 11.100 411.000 12.900 ;
        RECT 425.700 9.600 426.900 22.950 ;
        RECT 428.100 21.150 429.900 22.950 ;
        RECT 443.100 21.150 444.900 22.950 ;
        RECT 433.950 18.450 436.050 19.050 ;
        RECT 445.950 18.450 448.050 19.050 ;
        RECT 433.950 17.550 448.050 18.450 ;
        RECT 433.950 16.950 436.050 17.550 ;
        RECT 445.950 16.950 448.050 17.550 ;
        RECT 449.100 10.800 450.000 22.950 ;
        RECT 443.400 9.900 450.000 10.800 ;
        RECT 443.400 9.600 444.900 9.900 ;
        RECT 409.500 3.000 411.300 9.600 ;
        RECT 425.100 3.600 426.900 9.600 ;
        RECT 428.100 3.000 429.900 9.600 ;
        RECT 440.100 3.000 441.900 9.600 ;
        RECT 443.100 3.600 444.900 9.600 ;
        RECT 449.100 9.600 450.000 9.900 ;
        RECT 462.000 10.800 462.900 22.950 ;
        RECT 467.100 21.150 468.900 22.950 ;
        RECT 462.000 9.900 468.600 10.800 ;
        RECT 462.000 9.600 462.900 9.900 ;
        RECT 446.100 3.000 447.900 9.000 ;
        RECT 449.100 3.600 450.900 9.600 ;
        RECT 461.100 3.600 462.900 9.600 ;
        RECT 467.100 9.600 468.600 9.900 ;
        RECT 485.700 9.600 486.900 22.950 ;
        RECT 490.950 21.450 493.050 22.050 ;
        RECT 496.950 21.450 499.050 22.050 ;
        RECT 490.950 20.550 499.050 21.450 ;
        RECT 490.950 19.950 493.050 20.550 ;
        RECT 496.950 19.950 499.050 20.550 ;
        RECT 504.000 10.800 504.900 22.950 ;
        RECT 509.100 21.150 510.900 22.950 ;
        RECT 527.400 15.600 528.300 22.950 ;
        RECT 532.950 21.150 534.750 22.950 ;
        RECT 529.950 18.450 532.050 19.050 ;
        RECT 538.950 18.450 541.050 19.050 ;
        RECT 529.950 17.550 541.050 18.450 ;
        RECT 529.950 16.950 532.050 17.550 ;
        RECT 538.950 16.950 541.050 17.550 ;
        RECT 504.000 9.900 510.600 10.800 ;
        RECT 504.000 9.600 504.900 9.900 ;
        RECT 464.100 3.000 465.900 9.000 ;
        RECT 467.100 3.600 468.900 9.600 ;
        RECT 470.100 3.000 471.900 9.600 ;
        RECT 482.100 3.000 483.900 9.600 ;
        RECT 485.100 3.600 486.900 9.600 ;
        RECT 488.100 3.000 489.900 9.600 ;
        RECT 503.100 3.600 504.900 9.600 ;
        RECT 509.100 9.600 510.600 9.900 ;
        RECT 506.100 3.000 507.900 9.000 ;
        RECT 509.100 3.600 510.900 9.600 ;
        RECT 512.100 3.000 513.900 9.600 ;
        RECT 527.100 3.600 528.900 15.600 ;
        RECT 530.100 14.700 537.900 15.600 ;
        RECT 530.100 3.600 531.900 14.700 ;
        RECT 533.100 3.000 534.900 13.800 ;
        RECT 536.100 3.600 537.900 14.700 ;
        RECT 549.000 10.800 549.900 22.950 ;
        RECT 554.100 21.150 555.900 22.950 ;
        RECT 550.950 18.450 553.050 19.050 ;
        RECT 565.950 18.450 568.050 19.050 ;
        RECT 550.950 17.550 568.050 18.450 ;
        RECT 550.950 16.950 553.050 17.550 ;
        RECT 565.950 16.950 568.050 17.550 ;
        RECT 575.100 15.600 576.300 22.950 ;
        RECT 581.100 21.150 582.900 22.950 ;
        RECT 586.950 21.450 589.050 22.050 ;
        RECT 592.950 21.450 595.050 22.050 ;
        RECT 586.950 20.550 595.050 21.450 ;
        RECT 586.950 19.950 589.050 20.550 ;
        RECT 592.950 19.950 595.050 20.550 ;
        RECT 575.100 14.100 577.500 15.600 ;
        RECT 573.000 11.100 574.800 12.900 ;
        RECT 549.000 9.900 555.600 10.800 ;
        RECT 549.000 9.600 549.900 9.900 ;
        RECT 548.100 3.600 549.900 9.600 ;
        RECT 554.100 9.600 555.600 9.900 ;
        RECT 551.100 3.000 552.900 9.000 ;
        RECT 554.100 3.600 555.900 9.600 ;
        RECT 557.100 3.000 558.900 9.600 ;
        RECT 572.700 3.000 574.500 9.600 ;
        RECT 575.700 3.600 577.500 14.100 ;
        RECT 580.800 3.000 582.600 15.600 ;
        RECT 597.000 10.800 597.900 22.950 ;
        RECT 602.100 21.150 603.900 22.950 ;
        RECT 601.950 15.450 604.050 16.050 ;
        RECT 607.950 15.450 610.050 16.050 ;
        RECT 601.950 14.550 610.050 15.450 ;
        RECT 601.950 13.950 604.050 14.550 ;
        RECT 607.950 13.950 610.050 14.550 ;
        RECT 618.000 10.800 618.900 22.950 ;
        RECT 623.100 21.150 624.900 22.950 ;
        RECT 638.100 21.150 639.900 22.950 ;
        RECT 597.000 9.900 603.600 10.800 ;
        RECT 597.000 9.600 597.900 9.900 ;
        RECT 596.100 3.600 597.900 9.600 ;
        RECT 602.100 9.600 603.600 9.900 ;
        RECT 618.000 9.900 624.600 10.800 ;
        RECT 618.000 9.600 618.900 9.900 ;
        RECT 599.100 3.000 600.900 9.000 ;
        RECT 602.100 3.600 603.900 9.600 ;
        RECT 605.100 3.000 606.900 9.600 ;
        RECT 617.100 3.600 618.900 9.600 ;
        RECT 623.100 9.600 624.600 9.900 ;
        RECT 641.100 9.600 642.300 22.950 ;
        RECT 659.100 21.150 660.900 22.950 ;
        RECT 665.100 10.800 666.000 22.950 ;
        RECT 680.100 21.150 681.900 22.950 ;
        RECT 686.100 10.800 687.000 22.950 ;
        RECT 701.100 21.150 702.900 22.950 ;
        RECT 707.700 15.600 708.900 22.950 ;
        RECT 659.400 9.900 666.000 10.800 ;
        RECT 659.400 9.600 660.900 9.900 ;
        RECT 620.100 3.000 621.900 9.000 ;
        RECT 623.100 3.600 624.900 9.600 ;
        RECT 626.100 3.000 627.900 9.600 ;
        RECT 638.100 3.000 639.900 9.600 ;
        RECT 641.100 3.600 642.900 9.600 ;
        RECT 656.100 3.000 657.900 9.600 ;
        RECT 659.100 3.600 660.900 9.600 ;
        RECT 665.100 9.600 666.000 9.900 ;
        RECT 680.400 9.900 687.000 10.800 ;
        RECT 680.400 9.600 681.900 9.900 ;
        RECT 662.100 3.000 663.900 9.000 ;
        RECT 665.100 3.600 666.900 9.600 ;
        RECT 677.100 3.000 678.900 9.600 ;
        RECT 680.100 3.600 681.900 9.600 ;
        RECT 686.100 9.600 687.000 9.900 ;
        RECT 683.100 3.000 684.900 9.000 ;
        RECT 686.100 3.600 687.900 9.600 ;
        RECT 701.400 3.000 703.200 15.600 ;
        RECT 706.500 14.100 708.900 15.600 ;
        RECT 706.500 3.600 708.300 14.100 ;
        RECT 709.200 11.100 711.000 12.900 ;
        RECT 728.100 9.600 729.300 22.950 ;
        RECT 747.000 21.150 748.800 22.950 ;
        RECT 749.700 18.900 750.600 29.400 ;
        RECT 753.000 25.050 753.900 32.400 ;
        RECT 767.100 29.400 768.900 39.000 ;
        RECT 773.700 30.000 775.500 38.400 ;
        RECT 791.700 31.200 793.500 38.400 ;
        RECT 796.800 32.400 798.600 39.000 ;
        RECT 791.700 30.300 795.900 31.200 ;
        RECT 773.700 28.800 777.000 30.000 ;
        RECT 767.100 25.050 768.900 26.850 ;
        RECT 773.100 25.050 774.900 26.850 ;
        RECT 776.100 25.050 777.000 28.800 ;
        RECT 791.100 25.050 792.900 26.850 ;
        RECT 794.700 25.050 795.900 30.300 ;
        RECT 809.100 30.600 810.900 38.400 ;
        RECT 813.600 32.400 815.400 39.000 ;
        RECT 816.600 34.200 818.400 38.400 ;
        RECT 816.600 32.400 819.300 34.200 ;
        RECT 833.700 32.400 835.500 39.000 ;
        RECT 838.200 32.400 840.000 38.400 ;
        RECT 842.700 32.400 844.500 39.000 ;
        RECT 815.700 30.600 817.500 31.500 ;
        RECT 809.100 29.700 817.500 30.600 ;
        RECT 796.950 25.050 798.750 26.850 ;
        RECT 809.250 25.050 811.050 26.850 ;
        RECT 751.800 22.950 753.900 25.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 809.100 22.950 811.200 25.050 ;
        RECT 749.100 18.300 750.900 18.900 ;
        RECT 743.100 17.100 750.900 18.300 ;
        RECT 743.100 15.600 744.300 17.100 ;
        RECT 751.800 15.600 753.000 22.950 ;
        RECT 770.100 21.150 771.900 22.950 ;
        RECT 754.950 18.450 757.050 19.050 ;
        RECT 772.950 18.450 775.050 19.050 ;
        RECT 754.950 17.550 775.050 18.450 ;
        RECT 754.950 16.950 757.050 17.550 ;
        RECT 772.950 16.950 775.050 17.550 ;
        RECT 709.500 3.000 711.300 9.600 ;
        RECT 725.100 3.000 726.900 9.600 ;
        RECT 728.100 3.600 729.900 9.600 ;
        RECT 731.100 3.000 732.900 9.600 ;
        RECT 743.100 3.600 744.900 15.600 ;
        RECT 747.600 3.000 749.400 15.600 ;
        RECT 750.600 14.100 753.000 15.600 ;
        RECT 750.600 3.600 752.400 14.100 ;
        RECT 776.100 10.800 777.000 22.950 ;
        RECT 770.400 9.900 777.000 10.800 ;
        RECT 770.400 9.600 771.900 9.900 ;
        RECT 767.100 3.000 768.900 9.600 ;
        RECT 770.100 3.600 771.900 9.600 ;
        RECT 776.100 9.600 777.000 9.900 ;
        RECT 794.700 9.600 795.900 22.950 ;
        RECT 812.100 9.600 813.000 29.700 ;
        RECT 818.400 25.050 819.300 32.400 ;
        RECT 833.250 25.050 835.050 26.850 ;
        RECT 839.100 25.050 840.300 32.400 ;
        RECT 857.100 29.400 858.900 39.000 ;
        RECT 863.700 30.000 865.500 38.400 ;
        RECT 863.700 28.800 867.000 30.000 ;
        RECT 881.100 29.400 882.900 39.000 ;
        RECT 887.700 30.000 889.500 38.400 ;
        RECT 903.600 34.200 905.400 38.400 ;
        RECT 902.700 32.400 905.400 34.200 ;
        RECT 906.600 32.400 908.400 39.000 ;
        RECT 887.700 28.800 891.000 30.000 ;
        RECT 845.100 25.050 846.900 26.850 ;
        RECT 857.100 25.050 858.900 26.850 ;
        RECT 863.100 25.050 864.900 26.850 ;
        RECT 866.100 25.050 867.000 28.800 ;
        RECT 881.100 25.050 882.900 26.850 ;
        RECT 887.100 25.050 888.900 26.850 ;
        RECT 890.100 25.050 891.000 28.800 ;
        RECT 902.700 25.050 903.600 32.400 ;
        RECT 904.500 30.600 906.300 31.500 ;
        RECT 911.100 30.600 912.900 38.400 ;
        RECT 904.500 29.700 912.900 30.600 ;
        RECT 814.500 22.950 816.600 25.050 ;
        RECT 817.800 22.950 819.900 25.050 ;
        RECT 832.950 22.950 835.050 25.050 ;
        RECT 835.950 22.950 838.050 25.050 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 856.950 22.950 859.050 25.050 ;
        RECT 859.950 22.950 862.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 880.950 22.950 883.050 25.050 ;
        RECT 883.950 22.950 886.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 902.100 22.950 904.200 25.050 ;
        RECT 905.400 22.950 907.500 25.050 ;
        RECT 814.200 21.150 816.000 22.950 ;
        RECT 818.400 15.600 819.300 22.950 ;
        RECT 836.250 21.150 838.050 22.950 ;
        RECT 839.100 17.400 840.000 22.950 ;
        RECT 842.100 21.150 843.900 22.950 ;
        RECT 860.100 21.150 861.900 22.950 ;
        RECT 839.100 16.500 843.900 17.400 ;
        RECT 773.100 3.000 774.900 9.000 ;
        RECT 776.100 3.600 777.900 9.600 ;
        RECT 791.100 3.000 792.900 9.600 ;
        RECT 794.100 3.600 795.900 9.600 ;
        RECT 797.100 3.000 798.900 9.600 ;
        RECT 809.100 3.000 810.900 9.600 ;
        RECT 812.100 3.600 813.900 9.600 ;
        RECT 815.100 3.000 816.900 15.000 ;
        RECT 818.100 3.600 819.900 15.600 ;
        RECT 833.100 14.400 840.900 15.300 ;
        RECT 833.100 3.600 834.900 14.400 ;
        RECT 836.100 3.000 837.900 13.500 ;
        RECT 839.100 4.500 840.900 14.400 ;
        RECT 842.100 5.400 843.900 16.500 ;
        RECT 845.100 4.500 846.900 15.600 ;
        RECT 866.100 10.800 867.000 22.950 ;
        RECT 884.100 21.150 885.900 22.950 ;
        RECT 890.100 10.800 891.000 22.950 ;
        RECT 902.700 15.600 903.600 22.950 ;
        RECT 906.000 21.150 907.800 22.950 ;
        RECT 860.400 9.900 867.000 10.800 ;
        RECT 860.400 9.600 861.900 9.900 ;
        RECT 839.100 3.600 846.900 4.500 ;
        RECT 857.100 3.000 858.900 9.600 ;
        RECT 860.100 3.600 861.900 9.600 ;
        RECT 866.100 9.600 867.000 9.900 ;
        RECT 884.400 9.900 891.000 10.800 ;
        RECT 884.400 9.600 885.900 9.900 ;
        RECT 863.100 3.000 864.900 9.000 ;
        RECT 866.100 3.600 867.900 9.600 ;
        RECT 881.100 3.000 882.900 9.600 ;
        RECT 884.100 3.600 885.900 9.600 ;
        RECT 890.100 9.600 891.000 9.900 ;
        RECT 887.100 3.000 888.900 9.000 ;
        RECT 890.100 3.600 891.900 9.600 ;
        RECT 902.100 3.600 903.900 15.600 ;
        RECT 905.100 3.000 906.900 15.000 ;
        RECT 909.000 9.600 909.900 29.700 ;
        RECT 910.950 25.050 912.750 26.850 ;
        RECT 910.800 22.950 912.900 25.050 ;
        RECT 908.100 3.600 909.900 9.600 ;
        RECT 911.100 3.000 912.900 9.600 ;
      LAYER metal2 ;
        RECT 367.950 934.950 370.050 937.050 ;
        RECT 577.950 934.950 580.050 937.050 ;
        RECT 91.950 931.950 94.050 934.050 ;
        RECT 133.950 931.950 136.050 934.050 ;
        RECT 61.950 928.950 64.050 931.050 ;
        RECT 16.950 917.100 19.050 919.200 ;
        RECT 22.950 917.100 25.050 919.200 ;
        RECT 34.950 917.100 37.050 922.050 ;
        RECT 46.950 919.950 49.050 922.050 ;
        RECT 40.950 917.100 43.050 919.200 ;
        RECT 17.400 916.350 18.600 917.100 ;
        RECT 23.400 916.350 24.600 917.100 ;
        RECT 35.400 916.350 36.600 917.100 ;
        RECT 41.400 916.350 42.600 917.100 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 19.950 913.950 22.050 916.050 ;
        RECT 22.950 913.950 25.050 916.050 ;
        RECT 34.950 913.950 37.050 916.050 ;
        RECT 37.950 913.950 40.050 916.050 ;
        RECT 40.950 913.950 43.050 916.050 ;
        RECT 14.400 911.400 15.600 913.650 ;
        RECT 20.400 912.000 21.600 913.650 ;
        RECT 14.400 892.050 15.450 911.400 ;
        RECT 19.950 907.950 22.050 912.000 ;
        RECT 38.400 911.400 39.600 913.650 ;
        RECT 38.400 892.050 39.450 911.400 ;
        RECT 43.950 907.950 46.050 913.050 ;
        RECT 47.400 901.050 48.450 919.950 ;
        RECT 49.950 918.600 54.000 919.050 ;
        RECT 49.950 916.950 54.600 918.600 ;
        RECT 53.400 916.350 54.600 916.950 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 55.950 913.950 58.050 916.050 ;
        RECT 49.950 910.950 52.050 913.050 ;
        RECT 56.400 912.000 57.600 913.650 ;
        RECT 50.400 907.050 51.450 910.950 ;
        RECT 55.950 907.950 58.050 912.000 ;
        RECT 62.400 910.050 63.450 928.950 ;
        RECT 73.950 922.950 76.050 925.050 ;
        RECT 85.950 922.950 88.050 925.050 ;
        RECT 67.950 917.100 70.050 919.200 ;
        RECT 74.400 918.600 75.450 922.950 ;
        RECT 86.400 918.600 87.450 922.950 ;
        RECT 92.400 918.600 93.450 931.950 ;
        RECT 124.950 928.950 127.050 931.050 ;
        RECT 100.950 922.950 103.050 925.050 ;
        RECT 68.400 916.350 69.600 917.100 ;
        RECT 74.400 916.350 75.600 918.600 ;
        RECT 86.400 916.350 87.600 918.600 ;
        RECT 92.400 916.350 93.600 918.600 ;
        RECT 97.950 917.100 100.050 919.200 ;
        RECT 67.950 913.950 70.050 916.050 ;
        RECT 70.950 913.950 73.050 916.050 ;
        RECT 73.950 913.950 76.050 916.050 ;
        RECT 85.950 913.950 88.050 916.050 ;
        RECT 88.950 913.950 91.050 916.050 ;
        RECT 91.950 913.950 94.050 916.050 ;
        RECT 71.400 911.400 72.600 913.650 ;
        RECT 61.950 907.950 64.050 910.050 ;
        RECT 49.950 904.950 52.050 907.050 ;
        RECT 46.950 898.950 49.050 901.050 ;
        RECT 46.950 892.950 49.050 895.050 ;
        RECT 1.950 889.950 4.050 892.050 ;
        RECT 13.950 889.950 16.050 892.050 ;
        RECT 25.950 889.950 28.050 892.050 ;
        RECT 37.950 889.950 40.050 892.050 ;
        RECT 2.400 879.900 3.450 889.950 ;
        RECT 4.950 883.950 7.050 886.050 ;
        RECT 13.950 884.100 16.050 886.200 ;
        RECT 1.950 877.800 4.050 879.900 ;
        RECT 2.400 834.900 3.450 877.800 ;
        RECT 5.400 850.050 6.450 883.950 ;
        RECT 14.400 883.350 15.600 884.100 ;
        RECT 22.950 883.950 25.050 886.050 ;
        RECT 10.950 880.950 13.050 883.050 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 11.400 879.900 12.600 880.650 ;
        RECT 17.400 879.900 18.600 880.650 ;
        RECT 23.400 879.900 24.450 883.950 ;
        RECT 10.950 877.800 13.050 879.900 ;
        RECT 16.950 877.800 19.050 879.900 ;
        RECT 22.950 877.800 25.050 879.900 ;
        RECT 4.950 847.950 7.050 850.050 ;
        RECT 17.400 844.200 18.450 877.800 ;
        RECT 26.400 846.450 27.450 889.950 ;
        RECT 31.950 884.100 34.050 886.200 ;
        RECT 37.950 884.100 40.050 886.200 ;
        RECT 32.400 883.350 33.600 884.100 ;
        RECT 38.400 883.350 39.600 884.100 ;
        RECT 31.950 880.950 34.050 883.050 ;
        RECT 34.950 880.950 37.050 883.050 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 35.400 879.900 36.600 880.650 ;
        RECT 34.950 877.800 37.050 879.900 ;
        RECT 41.400 878.400 42.600 880.650 ;
        RECT 47.400 879.900 48.450 892.950 ;
        RECT 56.400 892.050 57.450 907.950 ;
        RECT 71.400 907.050 72.450 911.400 ;
        RECT 76.950 910.950 79.050 913.050 ;
        RECT 89.400 911.400 90.600 913.650 ;
        RECT 70.950 904.950 73.050 907.050 ;
        RECT 77.400 906.450 78.450 910.950 ;
        RECT 77.400 905.400 81.450 906.450 ;
        RECT 55.950 889.950 58.050 892.050 ;
        RECT 80.400 886.200 81.450 905.400 ;
        RECT 89.400 895.050 90.450 911.400 ;
        RECT 98.400 903.450 99.450 917.100 ;
        RECT 101.400 912.450 102.450 922.950 ;
        RECT 109.950 917.100 112.050 919.200 ;
        RECT 115.950 918.000 118.050 922.050 ;
        RECT 121.950 919.950 124.050 922.050 ;
        RECT 110.400 916.350 111.600 917.100 ;
        RECT 116.400 916.350 117.600 918.000 ;
        RECT 106.950 913.950 109.050 916.050 ;
        RECT 109.950 913.950 112.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 101.400 911.400 105.450 912.450 ;
        RECT 95.400 902.400 99.450 903.450 ;
        RECT 88.950 892.950 91.050 895.050 ;
        RECT 95.400 889.050 96.450 902.400 ;
        RECT 97.950 898.950 100.050 901.050 ;
        RECT 88.950 886.950 91.050 889.050 ;
        RECT 94.950 886.950 97.050 889.050 ;
        RECT 55.950 884.100 58.050 886.200 ;
        RECT 56.400 883.350 57.600 884.100 ;
        RECT 64.950 883.800 67.050 885.900 ;
        RECT 73.950 884.100 76.050 886.200 ;
        RECT 79.950 884.100 82.050 886.200 ;
        RECT 52.950 880.950 55.050 883.050 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 53.400 879.900 54.600 880.650 ;
        RECT 59.400 879.900 60.600 880.650 ;
        RECT 65.400 879.900 66.450 883.800 ;
        RECT 74.400 883.350 75.600 884.100 ;
        RECT 80.400 883.350 81.600 884.100 ;
        RECT 73.950 880.950 76.050 883.050 ;
        RECT 76.950 880.950 79.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 41.400 874.050 42.450 878.400 ;
        RECT 46.950 877.800 49.050 879.900 ;
        RECT 52.950 877.800 55.050 879.900 ;
        RECT 58.950 877.800 61.050 879.900 ;
        RECT 64.950 877.800 67.050 879.900 ;
        RECT 77.400 879.000 78.600 880.650 ;
        RECT 55.950 874.950 58.050 877.050 ;
        RECT 40.950 871.950 43.050 874.050 ;
        RECT 56.400 847.050 57.450 874.950 ;
        RECT 59.400 874.050 60.450 877.800 ;
        RECT 76.950 874.950 79.050 879.000 ;
        RECT 83.400 878.400 84.600 880.650 ;
        RECT 58.950 871.950 61.050 874.050 ;
        RECT 83.400 862.050 84.450 878.400 ;
        RECT 89.400 876.450 90.450 886.950 ;
        RECT 98.400 885.600 99.450 898.950 ;
        RECT 98.400 883.350 99.600 885.600 ;
        RECT 94.950 880.950 97.050 883.050 ;
        RECT 97.950 880.950 100.050 883.050 ;
        RECT 95.400 879.900 96.600 880.650 ;
        RECT 94.950 877.800 97.050 879.900 ;
        RECT 91.950 876.450 94.050 877.050 ;
        RECT 89.400 875.400 94.050 876.450 ;
        RECT 91.950 874.950 94.050 875.400 ;
        RECT 82.950 859.950 85.050 862.050 ;
        RECT 73.950 856.950 76.050 859.050 ;
        RECT 58.950 847.950 61.050 850.050 ;
        RECT 23.400 845.400 27.450 846.450 ;
        RECT 10.950 840.000 13.050 844.050 ;
        RECT 16.950 842.100 19.050 844.200 ;
        RECT 23.400 841.050 24.450 845.400 ;
        RECT 55.950 844.950 58.050 847.050 ;
        RECT 25.950 841.950 28.050 844.050 ;
        RECT 11.400 838.350 12.600 840.000 ;
        RECT 16.950 838.950 19.050 841.050 ;
        RECT 22.950 838.950 25.050 841.050 ;
        RECT 17.400 838.350 18.600 838.950 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 16.950 835.950 19.050 838.050 ;
        RECT 19.950 835.950 22.050 838.050 ;
        RECT 14.400 834.900 15.600 835.650 ;
        RECT 1.950 832.800 4.050 834.900 ;
        RECT 13.950 832.800 16.050 834.900 ;
        RECT 20.400 833.400 21.600 835.650 ;
        RECT 16.950 829.950 19.050 832.050 ;
        RECT 7.950 817.950 10.050 820.050 ;
        RECT 8.400 799.050 9.450 817.950 ;
        RECT 17.400 808.200 18.450 829.950 ;
        RECT 20.400 829.050 21.450 833.400 ;
        RECT 22.950 832.950 25.050 835.050 ;
        RECT 19.950 826.950 22.050 829.050 ;
        RECT 23.400 811.200 24.450 832.950 ;
        RECT 26.400 829.050 27.450 841.950 ;
        RECT 34.950 840.000 37.050 844.050 ;
        RECT 35.400 838.350 36.600 840.000 ;
        RECT 40.950 839.100 43.050 841.200 ;
        RECT 46.950 839.100 49.050 841.200 ;
        RECT 59.400 840.600 60.450 847.950 ;
        RECT 74.400 841.050 75.450 856.950 ;
        RECT 79.950 844.950 82.050 847.050 ;
        RECT 66.000 840.600 70.050 841.050 ;
        RECT 41.400 838.350 42.600 839.100 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 37.950 835.950 40.050 838.050 ;
        RECT 40.950 835.950 43.050 838.050 ;
        RECT 38.400 834.900 39.600 835.650 ;
        RECT 28.950 832.800 31.050 834.900 ;
        RECT 37.950 832.800 40.050 834.900 ;
        RECT 25.950 826.950 28.050 829.050 ;
        RECT 22.950 809.100 25.050 811.200 ;
        RECT 16.950 806.100 19.050 808.200 ;
        RECT 17.400 805.350 18.600 806.100 ;
        RECT 22.950 805.950 25.050 808.050 ;
        RECT 23.400 805.350 24.600 805.950 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 16.950 802.950 19.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 10.950 799.950 13.050 802.050 ;
        RECT 14.400 801.000 15.600 802.650 ;
        RECT 20.400 801.900 21.600 802.650 ;
        RECT 7.950 796.950 10.050 799.050 ;
        RECT 7.950 790.950 10.050 793.050 ;
        RECT 8.400 754.050 9.450 790.950 ;
        RECT 11.400 763.050 12.450 799.950 ;
        RECT 13.950 796.950 16.050 801.000 ;
        RECT 19.950 799.800 22.050 801.900 ;
        RECT 29.400 793.050 30.450 832.800 ;
        RECT 47.400 823.050 48.450 839.100 ;
        RECT 59.400 838.350 60.600 840.600 ;
        RECT 65.400 838.950 70.050 840.600 ;
        RECT 73.950 838.950 76.050 841.050 ;
        RECT 80.400 840.600 81.450 844.950 ;
        RECT 65.400 838.350 66.600 838.950 ;
        RECT 80.400 838.350 81.600 840.600 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 61.950 835.950 64.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 76.950 835.950 79.050 838.050 ;
        RECT 79.950 835.950 82.050 838.050 ;
        RECT 82.950 835.950 85.050 838.050 ;
        RECT 85.950 835.950 88.050 838.050 ;
        RECT 56.400 833.400 57.600 835.650 ;
        RECT 62.400 833.400 63.600 835.650 ;
        RECT 49.950 829.950 52.050 832.050 ;
        RECT 46.950 820.950 49.050 823.050 ;
        RECT 31.950 811.950 34.050 814.050 ;
        RECT 28.950 790.950 31.050 793.050 ;
        RECT 13.950 775.950 16.050 778.050 ;
        RECT 25.950 775.950 28.050 778.050 ;
        RECT 10.950 760.950 13.050 763.050 ;
        RECT 14.400 762.600 15.450 775.950 ;
        RECT 14.400 760.350 15.600 762.600 ;
        RECT 19.950 761.100 22.050 763.200 ;
        RECT 20.400 760.350 21.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 17.400 755.400 18.600 757.650 ;
        RECT 7.950 751.950 10.050 754.050 ;
        RECT 17.400 729.600 18.450 755.400 ;
        RECT 22.950 754.950 25.050 757.050 ;
        RECT 19.950 751.950 22.050 754.050 ;
        RECT 20.400 730.050 21.450 751.950 ;
        RECT 17.400 727.350 18.600 729.600 ;
        RECT 19.950 727.950 22.050 730.050 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 14.400 722.400 15.600 724.650 ;
        RECT 10.950 718.950 13.050 721.050 ;
        RECT 7.950 691.950 10.050 694.050 ;
        RECT 1.950 688.950 4.050 691.050 ;
        RECT 2.400 532.050 3.450 688.950 ;
        RECT 8.400 652.200 9.450 691.950 ;
        RECT 11.400 679.050 12.450 718.950 ;
        RECT 14.400 694.050 15.450 722.400 ;
        RECT 23.400 721.050 24.450 754.950 ;
        RECT 26.400 748.050 27.450 775.950 ;
        RECT 32.400 765.450 33.450 811.950 ;
        RECT 40.950 806.100 43.050 808.200 ;
        RECT 41.400 805.350 42.600 806.100 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 38.400 801.900 39.600 802.650 ;
        RECT 50.400 801.900 51.450 829.950 ;
        RECT 56.400 828.450 57.450 833.400 ;
        RECT 62.400 829.050 63.450 833.400 ;
        RECT 73.950 832.950 76.050 835.050 ;
        RECT 77.400 833.400 78.600 835.650 ;
        RECT 83.400 834.000 84.600 835.650 ;
        RECT 70.950 829.950 73.050 832.050 ;
        RECT 56.400 827.400 60.450 828.450 ;
        RECT 55.950 823.950 58.050 826.050 ;
        RECT 56.400 811.050 57.450 823.950 ;
        RECT 59.400 823.050 60.450 827.400 ;
        RECT 61.950 826.950 64.050 829.050 ;
        RECT 58.950 820.950 61.050 823.050 ;
        RECT 71.400 820.050 72.450 829.950 ;
        RECT 74.400 828.450 75.450 832.950 ;
        RECT 77.400 831.450 78.450 833.400 ;
        RECT 82.950 832.050 85.050 834.000 ;
        RECT 92.400 832.050 93.450 874.950 ;
        RECT 104.400 859.050 105.450 911.400 ;
        RECT 107.400 911.400 108.600 913.650 ;
        RECT 113.400 912.000 114.600 913.650 ;
        RECT 107.400 898.050 108.450 911.400 ;
        RECT 112.950 907.950 115.050 912.000 ;
        RECT 115.950 907.950 118.050 910.050 ;
        RECT 116.400 901.050 117.450 907.950 ;
        RECT 115.950 898.950 118.050 901.050 ;
        RECT 106.950 895.950 109.050 898.050 ;
        RECT 109.950 885.000 112.050 889.050 ;
        RECT 116.400 885.600 117.450 898.950 ;
        RECT 122.400 898.050 123.450 919.950 ;
        RECT 125.400 904.050 126.450 928.950 ;
        RECT 134.400 919.200 135.450 931.950 ;
        RECT 160.950 928.950 163.050 931.050 ;
        RECT 181.950 928.950 184.050 931.050 ;
        RECT 361.950 928.950 364.050 931.050 ;
        RECT 133.950 917.100 136.050 919.200 ;
        RECT 139.950 917.100 142.050 919.200 ;
        RECT 154.950 917.100 157.050 919.200 ;
        RECT 161.400 918.600 162.450 928.950 ;
        RECT 182.400 925.050 183.450 928.950 ;
        RECT 328.950 925.950 331.050 928.050 ;
        RECT 181.950 922.950 184.050 925.050 ;
        RECT 134.400 916.350 135.600 917.100 ;
        RECT 140.400 916.350 141.600 917.100 ;
        RECT 155.400 916.350 156.600 917.100 ;
        RECT 161.400 916.350 162.600 918.600 ;
        RECT 169.950 917.100 172.050 919.200 ;
        RECT 175.950 917.100 178.050 919.200 ;
        RECT 182.400 918.600 183.450 922.950 ;
        RECT 199.500 921.300 201.600 923.400 ;
        RECT 209.100 922.500 211.200 924.600 ;
        RECT 214.950 922.950 217.050 925.050 ;
        RECT 229.950 922.950 232.050 925.050 ;
        RECT 322.950 922.950 325.050 925.050 ;
        RECT 130.950 913.950 133.050 916.050 ;
        RECT 133.950 913.950 136.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 154.950 913.950 157.050 916.050 ;
        RECT 157.950 913.950 160.050 916.050 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 131.400 911.400 132.600 913.650 ;
        RECT 137.400 911.400 138.600 913.650 ;
        RECT 158.400 912.900 159.600 913.650 ;
        RECT 164.400 912.900 165.600 913.650 ;
        RECT 124.950 901.950 127.050 904.050 ;
        RECT 131.400 898.050 132.450 911.400 ;
        RECT 121.950 895.950 124.050 898.050 ;
        RECT 130.950 895.950 133.050 898.050 ;
        RECT 110.400 883.350 111.600 885.000 ;
        RECT 116.400 883.350 117.600 885.600 ;
        RECT 118.950 883.950 121.050 889.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 112.950 880.950 115.050 883.050 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 113.400 879.900 114.600 880.650 ;
        RECT 112.950 877.800 115.050 879.900 ;
        RECT 118.950 877.950 121.050 880.050 ;
        RECT 106.950 871.950 109.050 874.050 ;
        RECT 103.950 856.950 106.050 859.050 ;
        RECT 107.400 841.200 108.450 871.950 ;
        RECT 112.950 859.950 115.050 862.050 ;
        RECT 94.950 839.100 97.050 841.200 ;
        RECT 100.950 839.100 103.050 841.200 ;
        RECT 106.950 839.100 109.050 841.200 ;
        RECT 95.400 834.450 96.450 839.100 ;
        RECT 101.400 838.350 102.600 839.100 ;
        RECT 107.400 838.350 108.600 839.100 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 103.950 835.950 106.050 838.050 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 95.400 833.400 99.450 834.450 ;
        RECT 77.400 831.000 81.450 831.450 ;
        RECT 82.800 831.000 85.050 832.050 ;
        RECT 77.400 830.400 82.050 831.000 ;
        RECT 74.400 827.400 78.450 828.450 ;
        RECT 70.950 817.950 73.050 820.050 ;
        RECT 64.950 811.950 67.050 814.050 ;
        RECT 55.950 808.950 58.050 811.050 ;
        RECT 58.950 806.100 61.050 808.200 ;
        RECT 65.400 808.050 66.450 811.950 ;
        RECT 59.400 805.350 60.600 806.100 ;
        RECT 64.950 805.950 67.050 808.050 ;
        RECT 77.400 807.600 78.450 827.400 ;
        RECT 79.950 826.950 82.050 830.400 ;
        RECT 82.800 829.950 84.900 831.000 ;
        RECT 91.950 829.950 94.050 832.050 ;
        RECT 98.400 829.050 99.450 833.400 ;
        RECT 104.400 833.400 105.600 835.650 ;
        RECT 104.400 832.050 105.450 833.400 ;
        RECT 109.950 832.950 112.050 835.050 ;
        RECT 100.950 830.400 105.450 832.050 ;
        RECT 100.950 829.950 105.000 830.400 ;
        RECT 106.950 829.950 109.050 832.050 ;
        RECT 97.950 826.950 100.050 829.050 ;
        RECT 107.400 817.050 108.450 829.950 ;
        RECT 106.950 814.950 109.050 817.050 ;
        RECT 77.400 805.350 78.600 807.600 ;
        RECT 82.950 807.000 85.050 811.050 ;
        RECT 83.400 805.350 84.600 807.000 ;
        RECT 97.950 806.100 100.050 808.200 ;
        RECT 98.400 805.350 99.600 806.100 ;
        RECT 55.950 802.950 58.050 805.050 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 76.950 802.950 79.050 805.050 ;
        RECT 79.950 802.950 82.050 805.050 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 94.950 802.950 97.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 37.950 799.800 40.050 801.900 ;
        RECT 49.800 799.800 51.900 801.900 ;
        RECT 56.400 801.000 57.600 802.650 ;
        RECT 62.400 801.900 63.600 802.650 ;
        RECT 32.400 764.400 36.450 765.450 ;
        RECT 35.400 763.200 36.450 764.400 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 40.950 761.100 43.050 763.200 ;
        RECT 46.950 761.100 49.050 763.200 ;
        RECT 35.400 760.350 36.600 761.100 ;
        RECT 41.400 760.350 42.600 761.100 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 28.950 754.950 31.050 757.050 ;
        RECT 32.400 755.400 33.600 757.650 ;
        RECT 38.400 755.400 39.600 757.650 ;
        RECT 47.400 757.050 48.450 761.100 ;
        RECT 25.950 745.950 28.050 748.050 ;
        RECT 29.400 736.050 30.450 754.950 ;
        RECT 32.400 736.050 33.450 755.400 ;
        RECT 38.400 748.050 39.450 755.400 ;
        RECT 46.950 754.950 49.050 757.050 ;
        RECT 50.400 753.450 51.450 799.800 ;
        RECT 55.950 796.950 58.050 801.000 ;
        RECT 61.950 799.800 64.050 801.900 ;
        RECT 74.400 800.400 75.600 802.650 ;
        RECT 80.400 801.900 81.600 802.650 ;
        RECT 74.400 793.050 75.450 800.400 ;
        RECT 79.950 799.800 82.050 801.900 ;
        RECT 91.950 799.950 94.050 802.050 ;
        RECT 95.400 800.400 96.600 802.650 ;
        RECT 101.400 801.900 102.600 802.650 ;
        RECT 73.950 790.950 76.050 793.050 ;
        RECT 73.950 781.950 76.050 784.050 ;
        RECT 55.500 765.300 57.600 767.400 ;
        RECT 65.100 766.500 67.200 768.600 ;
        RECT 52.950 761.100 55.050 763.200 ;
        RECT 53.400 760.350 54.600 761.100 ;
        RECT 53.100 757.950 55.200 760.050 ;
        RECT 56.400 756.300 57.300 765.300 ;
        RECT 58.800 761.700 60.900 763.800 ;
        RECT 62.400 763.350 63.600 765.600 ;
        RECT 60.000 759.300 60.900 761.700 ;
        RECT 61.800 760.950 63.900 763.050 ;
        RECT 65.700 759.300 66.900 766.500 ;
        RECT 60.000 758.100 66.900 759.300 ;
        RECT 63.000 756.300 65.100 757.200 ;
        RECT 56.400 755.100 65.100 756.300 ;
        RECT 47.400 752.400 51.450 753.450 ;
        RECT 57.900 753.300 60.000 755.100 ;
        RECT 37.950 745.950 40.050 748.050 ;
        RECT 47.400 736.050 48.450 752.400 ;
        RECT 61.800 752.100 63.900 754.200 ;
        RECT 66.000 752.700 66.900 758.100 ;
        RECT 67.800 757.950 69.900 760.050 ;
        RECT 68.400 756.900 69.600 757.650 ;
        RECT 67.950 754.800 70.050 756.900 ;
        RECT 49.950 750.450 54.000 751.050 ;
        RECT 49.950 750.000 54.450 750.450 ;
        RECT 49.950 748.950 55.050 750.000 ;
        RECT 52.950 745.950 55.050 748.950 ;
        RECT 62.400 749.550 63.600 751.800 ;
        RECT 65.100 750.600 67.200 752.700 ;
        RECT 62.400 736.050 63.450 749.550 ;
        RECT 70.950 736.950 73.050 739.050 ;
        RECT 28.950 733.950 31.050 736.050 ;
        RECT 31.950 733.950 34.050 736.050 ;
        RECT 46.950 733.950 49.050 736.050 ;
        RECT 61.950 733.950 64.050 736.050 ;
        RECT 31.950 728.100 34.050 730.200 ;
        RECT 47.400 729.600 48.450 733.950 ;
        RECT 32.400 727.350 33.600 728.100 ;
        RECT 47.400 727.350 48.600 729.600 ;
        RECT 52.950 728.100 55.050 730.200 ;
        RECT 58.950 728.100 61.050 730.200 ;
        RECT 71.400 729.600 72.450 736.950 ;
        RECT 53.400 727.350 54.600 728.100 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 46.950 724.950 49.050 727.050 ;
        RECT 49.950 724.950 52.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 29.400 722.400 30.600 724.650 ;
        RECT 50.400 722.400 51.600 724.650 ;
        RECT 22.950 718.950 25.050 721.050 ;
        RECT 13.950 691.950 16.050 694.050 ;
        RECT 22.950 688.950 25.050 691.050 ;
        RECT 23.400 684.600 24.450 688.950 ;
        RECT 23.400 682.350 24.600 684.600 ;
        RECT 14.100 679.950 16.200 682.050 ;
        RECT 17.400 679.950 19.500 682.050 ;
        RECT 22.800 679.950 24.900 682.050 ;
        RECT 10.950 676.950 13.050 679.050 ;
        RECT 17.400 678.900 18.600 679.650 ;
        RECT 16.950 676.800 19.050 678.900 ;
        RECT 7.950 650.100 10.050 652.200 ;
        RECT 13.950 650.100 16.050 652.200 ;
        RECT 19.950 650.100 22.050 652.200 ;
        RECT 25.950 650.100 28.050 652.200 ;
        RECT 14.400 649.350 15.600 650.100 ;
        RECT 20.400 649.350 21.600 650.100 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 17.400 644.400 18.600 646.650 ;
        RECT 7.950 610.950 10.050 613.050 ;
        RECT 8.400 535.050 9.450 610.950 ;
        RECT 17.400 609.450 18.450 644.400 ;
        RECT 26.400 643.050 27.450 650.100 ;
        RECT 25.950 640.950 28.050 643.050 ;
        RECT 29.400 613.050 30.450 722.400 ;
        RECT 46.800 683.100 48.900 685.200 ;
        RECT 50.400 685.050 51.450 722.400 ;
        RECT 59.400 712.050 60.450 728.100 ;
        RECT 71.400 727.350 72.600 729.600 ;
        RECT 74.400 729.450 75.450 781.950 ;
        RECT 80.400 775.050 81.450 799.800 ;
        RECT 92.400 778.050 93.450 799.950 ;
        RECT 95.400 796.050 96.450 800.400 ;
        RECT 100.950 799.800 103.050 801.900 ;
        RECT 103.950 799.950 106.050 802.050 ;
        RECT 107.400 801.900 108.450 814.950 ;
        RECT 110.400 811.050 111.450 832.950 ;
        RECT 113.400 832.050 114.450 859.950 ;
        RECT 115.950 844.950 118.050 847.050 ;
        RECT 112.950 829.950 115.050 832.050 ;
        RECT 116.400 828.450 117.450 844.950 ;
        RECT 119.400 841.050 120.450 877.950 ;
        RECT 122.400 862.050 123.450 895.950 ;
        RECT 137.400 889.050 138.450 911.400 ;
        RECT 157.950 910.800 160.050 912.900 ;
        RECT 163.950 910.800 166.050 912.900 ;
        RECT 170.400 910.050 171.450 917.100 ;
        RECT 176.400 916.350 177.600 917.100 ;
        RECT 182.400 916.350 183.600 918.600 ;
        RECT 190.950 916.950 193.050 919.050 ;
        RECT 197.400 918.450 198.600 918.600 ;
        RECT 194.400 917.400 198.600 918.450 ;
        RECT 175.950 913.950 178.050 916.050 ;
        RECT 178.950 913.950 181.050 916.050 ;
        RECT 181.950 913.950 184.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 172.950 910.800 175.050 912.900 ;
        RECT 179.400 912.000 180.600 913.650 ;
        RECT 185.400 912.900 186.600 913.650 ;
        RECT 169.950 907.950 172.050 910.050 ;
        RECT 157.950 901.950 160.050 904.050 ;
        RECT 158.400 891.450 159.450 901.950 ;
        RECT 124.950 886.950 127.050 889.050 ;
        RECT 136.950 886.950 139.050 889.050 ;
        RECT 154.800 888.300 156.900 890.400 ;
        RECT 158.400 889.200 159.600 891.450 ;
        RECT 125.400 879.900 126.450 886.950 ;
        RECT 133.950 884.100 136.050 886.200 ;
        RECT 139.950 884.100 142.050 886.200 ;
        RECT 152.400 885.450 153.600 885.600 ;
        RECT 149.400 884.400 153.600 885.450 ;
        RECT 134.400 883.350 135.600 884.100 ;
        RECT 140.400 883.350 141.600 884.100 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 124.950 877.800 127.050 879.900 ;
        RECT 131.400 878.400 132.600 880.650 ;
        RECT 137.400 879.900 138.600 880.650 ;
        RECT 131.400 874.050 132.450 878.400 ;
        RECT 136.950 877.800 139.050 879.900 ;
        RECT 142.950 877.950 145.050 880.050 ;
        RECT 130.950 871.950 133.050 874.050 ;
        RECT 121.950 859.950 124.050 862.050 ;
        RECT 133.950 856.950 136.050 859.050 ;
        RECT 118.950 838.950 121.050 841.050 ;
        RECT 124.950 839.100 127.050 841.200 ;
        RECT 134.400 841.050 135.450 856.950 ;
        RECT 143.400 847.050 144.450 877.950 ;
        RECT 149.400 870.450 150.450 884.400 ;
        RECT 152.400 883.350 153.600 884.400 ;
        RECT 152.100 880.950 154.200 883.050 ;
        RECT 155.100 882.900 156.000 888.300 ;
        RECT 158.100 886.800 160.200 888.900 ;
        RECT 162.000 885.900 164.100 887.700 ;
        RECT 156.900 884.700 165.600 885.900 ;
        RECT 156.900 883.800 159.000 884.700 ;
        RECT 155.100 881.700 162.000 882.900 ;
        RECT 155.100 874.500 156.300 881.700 ;
        RECT 158.100 877.950 160.200 880.050 ;
        RECT 161.100 879.300 162.000 881.700 ;
        RECT 158.400 875.400 159.600 877.650 ;
        RECT 161.100 877.200 163.200 879.300 ;
        RECT 164.700 875.700 165.600 884.700 ;
        RECT 169.950 883.950 172.050 886.050 ;
        RECT 166.800 880.950 168.900 883.050 ;
        RECT 167.400 879.450 168.600 880.650 ;
        RECT 170.400 879.450 171.450 883.950 ;
        RECT 167.400 878.400 171.450 879.450 ;
        RECT 154.800 872.400 156.900 874.500 ;
        RECT 164.400 873.600 166.500 875.700 ;
        RECT 149.400 869.400 153.450 870.450 ;
        RECT 142.950 844.950 145.050 847.050 ;
        RECT 148.950 844.950 151.050 847.050 ;
        RECT 149.400 841.200 150.450 844.950 ;
        RECT 125.400 838.350 126.600 839.100 ;
        RECT 130.950 838.950 133.050 841.050 ;
        RECT 133.950 838.950 136.050 841.050 ;
        RECT 136.950 839.100 139.050 841.200 ;
        RECT 142.950 839.100 145.050 841.200 ;
        RECT 148.950 839.100 151.050 841.200 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 124.950 835.950 127.050 838.050 ;
        RECT 118.950 834.450 121.050 835.050 ;
        RECT 122.400 834.450 123.600 835.650 ;
        RECT 118.950 833.400 123.600 834.450 ;
        RECT 118.950 832.950 121.050 833.400 ;
        RECT 127.950 832.950 130.050 835.050 ;
        RECT 113.400 827.400 117.450 828.450 ;
        RECT 109.950 808.950 112.050 811.050 ;
        RECT 113.400 807.450 114.450 827.400 ;
        RECT 119.400 811.050 120.450 832.950 ;
        RECT 124.950 822.450 127.050 823.050 ;
        RECT 128.400 822.450 129.450 832.950 ;
        RECT 131.400 829.050 132.450 838.950 ;
        RECT 137.400 838.350 138.600 839.100 ;
        RECT 143.400 838.350 144.600 839.100 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 142.950 835.950 145.050 838.050 ;
        RECT 145.950 835.950 148.050 838.050 ;
        RECT 133.950 832.950 136.050 835.050 ;
        RECT 140.400 833.400 141.600 835.650 ;
        RECT 146.400 833.400 147.600 835.650 ;
        RECT 134.400 829.050 135.450 832.950 ;
        RECT 136.950 829.950 139.050 832.050 ;
        RECT 130.800 826.950 132.900 829.050 ;
        RECT 133.950 826.950 136.050 829.050 ;
        RECT 130.950 823.800 133.050 825.900 ;
        RECT 124.950 821.400 129.450 822.450 ;
        RECT 124.950 820.950 127.050 821.400 ;
        RECT 118.950 808.950 121.050 811.050 ;
        RECT 110.400 806.400 114.450 807.450 ;
        RECT 119.400 807.600 120.450 808.950 ;
        RECT 125.400 807.600 126.450 820.950 ;
        RECT 104.400 796.050 105.450 799.950 ;
        RECT 106.950 799.800 109.050 801.900 ;
        RECT 94.950 793.950 97.050 796.050 ;
        RECT 103.950 793.950 106.050 796.050 ;
        RECT 91.950 775.950 94.050 778.050 ;
        RECT 79.950 772.950 82.050 775.050 ;
        RECT 85.950 772.950 88.050 775.050 ;
        RECT 79.950 766.950 82.050 769.050 ;
        RECT 80.400 762.600 81.450 766.950 ;
        RECT 86.400 762.600 87.450 772.950 ;
        RECT 97.950 766.950 100.050 769.050 ;
        RECT 80.400 760.350 81.600 762.600 ;
        RECT 86.400 760.350 87.600 762.600 ;
        RECT 91.950 761.100 94.050 763.200 ;
        RECT 92.400 760.350 93.600 761.100 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 91.950 757.950 94.050 760.050 ;
        RECT 83.400 756.900 84.600 757.650 ;
        RECT 82.950 754.800 85.050 756.900 ;
        RECT 89.400 756.000 90.600 757.650 ;
        RECT 83.400 753.450 84.450 754.800 ;
        RECT 80.400 752.400 84.450 753.450 ;
        RECT 80.400 730.050 81.450 752.400 ;
        RECT 88.950 751.950 91.050 756.000 ;
        RECT 94.950 754.950 97.050 757.050 ;
        RECT 95.400 742.050 96.450 754.950 ;
        RECT 98.400 751.050 99.450 766.950 ;
        RECT 100.950 760.950 103.050 763.050 ;
        RECT 101.400 754.050 102.450 760.950 ;
        RECT 100.950 751.950 103.050 754.050 ;
        RECT 97.950 748.950 100.050 751.050 ;
        RECT 97.950 742.950 100.050 745.050 ;
        RECT 94.950 739.950 97.050 742.050 ;
        RECT 82.950 736.950 85.050 739.050 ;
        RECT 83.400 733.050 84.450 736.950 ;
        RECT 85.950 733.950 88.050 736.050 ;
        RECT 82.950 730.950 85.050 733.050 ;
        RECT 74.400 728.400 78.450 729.450 ;
        RECT 67.950 724.950 70.050 727.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 68.400 723.900 69.600 724.650 ;
        RECT 67.950 721.800 70.050 723.900 ;
        RECT 58.950 709.950 61.050 712.050 ;
        RECT 77.400 694.050 78.450 728.400 ;
        RECT 79.950 727.950 82.050 730.050 ;
        RECT 86.400 729.600 87.450 733.950 ;
        RECT 98.400 730.050 99.450 742.950 ;
        RECT 86.400 727.350 87.600 729.600 ;
        RECT 97.950 727.950 100.050 730.050 ;
        RECT 104.400 729.600 105.450 793.950 ;
        RECT 107.400 793.050 108.450 799.800 ;
        RECT 106.950 790.950 109.050 793.050 ;
        RECT 110.400 766.050 111.450 806.400 ;
        RECT 119.400 805.350 120.600 807.600 ;
        RECT 125.400 805.350 126.600 807.600 ;
        RECT 115.950 802.950 118.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 116.400 801.900 117.600 802.650 ;
        RECT 122.400 801.900 123.600 802.650 ;
        RECT 115.950 799.800 118.050 801.900 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 112.950 784.950 115.050 787.050 ;
        RECT 113.400 766.050 114.450 784.950 ;
        RECT 131.400 784.050 132.450 823.800 ;
        RECT 137.400 811.050 138.450 829.950 ;
        RECT 140.400 817.050 141.450 833.400 ;
        RECT 146.400 829.050 147.450 833.400 ;
        RECT 152.400 829.050 153.450 869.400 ;
        RECT 173.400 865.050 174.450 910.800 ;
        RECT 178.950 907.950 181.050 912.000 ;
        RECT 184.950 910.800 187.050 912.900 ;
        RECT 187.950 910.950 190.050 913.050 ;
        RECT 191.400 912.900 192.450 916.950 ;
        RECT 188.400 892.050 189.450 910.950 ;
        RECT 190.950 910.800 193.050 912.900 ;
        RECT 194.400 904.050 195.450 917.400 ;
        RECT 197.400 916.350 198.600 917.400 ;
        RECT 197.100 913.950 199.200 916.050 ;
        RECT 200.400 912.300 201.300 921.300 ;
        RECT 202.800 917.700 204.900 919.800 ;
        RECT 206.400 919.350 207.600 921.600 ;
        RECT 204.000 915.300 204.900 917.700 ;
        RECT 205.800 916.950 207.900 919.050 ;
        RECT 209.700 915.300 210.900 922.500 ;
        RECT 204.000 914.100 210.900 915.300 ;
        RECT 207.000 912.300 209.100 913.200 ;
        RECT 200.400 911.100 209.100 912.300 ;
        RECT 201.900 909.300 204.000 911.100 ;
        RECT 205.800 908.100 207.900 910.200 ;
        RECT 210.000 908.700 210.900 914.100 ;
        RECT 211.800 913.950 213.900 916.050 ;
        RECT 212.400 912.900 213.600 913.650 ;
        RECT 211.950 910.800 214.050 912.900 ;
        RECT 206.400 905.550 207.600 907.800 ;
        RECT 209.100 906.600 211.200 908.700 ;
        RECT 193.950 901.950 196.050 904.050 ;
        RECT 206.400 895.050 207.450 905.550 ;
        RECT 199.950 892.950 202.050 895.050 ;
        RECT 205.950 892.950 208.050 895.050 ;
        RECT 175.950 889.950 178.050 892.050 ;
        RECT 187.950 889.950 190.050 892.050 ;
        RECT 172.950 862.950 175.050 865.050 ;
        RECT 176.400 859.050 177.450 889.950 ;
        RECT 181.950 884.100 184.050 886.200 ;
        RECT 188.400 885.600 189.450 889.950 ;
        RECT 182.400 883.350 183.600 884.100 ;
        RECT 188.400 883.350 189.600 885.600 ;
        RECT 196.950 883.950 199.050 886.050 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 187.950 880.950 190.050 883.050 ;
        RECT 190.950 880.950 193.050 883.050 ;
        RECT 185.400 879.900 186.600 880.650 ;
        RECT 184.950 877.800 187.050 879.900 ;
        RECT 191.400 878.400 192.600 880.650 ;
        RECT 197.400 879.900 198.450 883.950 ;
        RECT 191.400 865.050 192.450 878.400 ;
        RECT 196.950 877.800 199.050 879.900 ;
        RECT 193.950 865.950 196.050 868.050 ;
        RECT 190.950 862.950 193.050 865.050 ;
        RECT 175.950 856.950 178.050 859.050 ;
        RECT 154.950 853.950 157.050 856.050 ;
        RECT 155.400 832.050 156.450 853.950 ;
        RECT 160.500 843.300 162.600 845.400 ;
        RECT 170.100 844.500 172.200 846.600 ;
        RECT 157.950 839.100 160.050 841.200 ;
        RECT 158.400 838.350 159.600 839.100 ;
        RECT 158.100 835.950 160.200 838.050 ;
        RECT 161.400 834.300 162.300 843.300 ;
        RECT 163.800 839.700 165.900 841.800 ;
        RECT 167.400 841.350 168.600 843.600 ;
        RECT 165.000 837.300 165.900 839.700 ;
        RECT 166.800 838.950 168.900 841.050 ;
        RECT 170.700 837.300 171.900 844.500 ;
        RECT 191.400 840.450 192.600 840.600 ;
        RECT 194.400 840.450 195.450 865.950 ;
        RECT 196.950 859.950 199.050 862.050 ;
        RECT 191.400 839.400 195.450 840.450 ;
        RECT 191.400 838.350 192.600 839.400 ;
        RECT 197.400 838.050 198.450 859.950 ;
        RECT 165.000 836.100 171.900 837.300 ;
        RECT 168.000 834.300 170.100 835.200 ;
        RECT 161.400 833.100 170.100 834.300 ;
        RECT 154.950 829.950 157.050 832.050 ;
        RECT 162.900 831.300 165.000 833.100 ;
        RECT 166.800 830.100 168.900 832.200 ;
        RECT 171.000 830.700 171.900 836.100 ;
        RECT 172.800 835.950 174.900 838.050 ;
        RECT 173.400 834.450 174.600 835.650 ;
        RECT 175.950 834.450 178.050 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 187.950 835.950 190.050 838.050 ;
        RECT 190.950 835.950 193.050 838.050 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 173.400 834.000 178.050 834.450 ;
        RECT 173.400 833.400 177.450 834.000 ;
        RECT 188.400 833.400 189.600 835.650 ;
        RECT 145.950 826.950 148.050 829.050 ;
        RECT 151.950 826.950 154.050 829.050 ;
        RECT 167.400 827.550 168.600 829.800 ;
        RECT 170.100 828.600 172.200 830.700 ;
        RECT 175.950 829.950 178.050 832.050 ;
        RECT 188.400 831.450 189.450 833.400 ;
        RECT 193.950 832.950 196.050 835.050 ;
        RECT 185.400 830.400 189.450 831.450 ;
        RECT 139.950 814.950 142.050 817.050 ;
        RECT 139.950 811.800 142.050 813.900 ;
        RECT 136.950 808.950 139.050 811.050 ;
        RECT 140.400 807.600 141.450 811.800 ;
        RECT 140.400 805.350 141.600 807.600 ;
        RECT 136.950 802.950 139.050 805.050 ;
        RECT 139.950 802.950 142.050 805.050 ;
        RECT 137.400 801.900 138.600 802.650 ;
        RECT 136.950 799.800 139.050 801.900 ;
        RECT 146.400 787.050 147.450 826.950 ;
        RECT 167.400 820.050 168.450 827.550 ;
        RECT 169.950 820.950 172.050 823.050 ;
        RECT 166.950 817.950 169.050 820.050 ;
        RECT 148.950 806.100 151.050 808.200 ;
        RECT 157.950 806.100 160.050 808.200 ;
        RECT 163.950 806.100 166.050 808.200 ;
        RECT 145.950 784.950 148.050 787.050 ;
        RECT 130.950 781.950 133.050 784.050 ;
        RECT 149.400 781.050 150.450 806.100 ;
        RECT 158.400 805.350 159.600 806.100 ;
        RECT 164.400 805.350 165.600 806.100 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 160.950 802.950 163.050 805.050 ;
        RECT 163.950 802.950 166.050 805.050 ;
        RECT 155.400 801.900 156.600 802.650 ;
        RECT 161.400 801.900 162.600 802.650 ;
        RECT 154.950 799.800 157.050 801.900 ;
        RECT 160.950 799.800 163.050 801.900 ;
        RECT 170.400 781.050 171.450 820.950 ;
        RECT 176.400 807.450 177.450 829.950 ;
        RECT 185.400 808.200 186.450 830.400 ;
        RECT 187.950 826.950 190.050 829.050 ;
        RECT 173.400 806.400 177.450 807.450 ;
        RECT 173.400 801.900 174.450 806.400 ;
        RECT 184.950 806.100 187.050 808.200 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 181.950 802.950 184.050 805.050 ;
        RECT 172.950 799.800 175.050 801.900 ;
        RECT 182.400 800.400 183.600 802.650 ;
        RECT 188.400 802.050 189.450 826.950 ;
        RECT 194.400 814.050 195.450 832.950 ;
        RECT 193.950 811.950 196.050 814.050 ;
        RECT 196.950 807.000 199.050 811.050 ;
        RECT 200.400 807.450 201.450 892.950 ;
        RECT 211.950 889.950 214.050 892.050 ;
        RECT 205.950 884.100 208.050 889.050 ;
        RECT 212.400 885.600 213.450 889.950 ;
        RECT 215.400 889.050 216.450 922.950 ;
        RECT 230.400 919.200 231.450 922.950 ;
        RECT 229.950 917.100 232.050 919.200 ;
        RECT 238.950 917.100 241.050 919.200 ;
        RECT 247.950 917.100 250.050 919.200 ;
        RECT 254.400 918.450 255.600 918.600 ;
        RECT 254.400 917.400 261.450 918.450 ;
        RECT 230.400 916.350 231.600 917.100 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 232.950 913.950 235.050 916.050 ;
        RECT 227.400 911.400 228.600 913.650 ;
        RECT 233.400 912.000 234.600 913.650 ;
        RECT 239.400 912.900 240.450 917.100 ;
        RECT 248.400 916.350 249.600 917.100 ;
        RECT 254.400 916.350 255.600 917.400 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 251.400 912.900 252.600 913.650 ;
        RECT 227.400 895.050 228.450 911.400 ;
        RECT 232.950 907.950 235.050 912.000 ;
        RECT 238.950 910.800 241.050 912.900 ;
        RECT 250.950 910.800 253.050 912.900 ;
        RECT 239.400 901.050 240.450 910.800 ;
        RECT 241.950 907.950 244.050 910.050 ;
        RECT 238.950 898.950 241.050 901.050 ;
        RECT 226.950 892.950 229.050 895.050 ;
        RECT 235.950 892.950 238.050 895.050 ;
        RECT 214.950 886.950 217.050 889.050 ;
        RECT 236.400 886.200 237.450 892.950 ;
        RECT 206.400 883.350 207.600 884.100 ;
        RECT 212.400 883.350 213.600 885.600 ;
        RECT 229.950 884.100 232.050 886.200 ;
        RECT 235.950 884.100 238.050 886.200 ;
        RECT 230.400 883.350 231.600 884.100 ;
        RECT 236.400 883.350 237.600 884.100 ;
        RECT 205.950 880.950 208.050 883.050 ;
        RECT 208.950 880.950 211.050 883.050 ;
        RECT 211.950 880.950 214.050 883.050 ;
        RECT 214.950 880.950 217.050 883.050 ;
        RECT 226.950 880.950 229.050 883.050 ;
        RECT 229.950 880.950 232.050 883.050 ;
        RECT 232.950 880.950 235.050 883.050 ;
        RECT 235.950 880.950 238.050 883.050 ;
        RECT 209.400 879.900 210.600 880.650 ;
        RECT 215.400 879.900 216.600 880.650 ;
        RECT 208.950 877.800 211.050 879.900 ;
        RECT 214.950 877.800 217.050 879.900 ;
        RECT 227.400 878.400 228.600 880.650 ;
        RECT 233.400 878.400 234.600 880.650 ;
        RECT 202.950 844.950 205.050 847.050 ;
        RECT 203.400 841.050 204.450 844.950 ;
        RECT 202.950 838.950 205.050 841.050 ;
        RECT 208.950 839.100 211.050 841.200 ;
        RECT 215.400 840.600 216.450 877.800 ;
        RECT 227.400 859.050 228.450 878.400 ;
        RECT 233.400 874.050 234.450 878.400 ;
        RECT 232.950 871.950 235.050 874.050 ;
        RECT 242.400 859.050 243.450 907.950 ;
        RECT 260.400 904.050 261.450 917.400 ;
        RECT 262.950 917.100 265.050 919.200 ;
        RECT 268.950 917.100 271.050 919.200 ;
        RECT 274.950 917.100 277.050 919.200 ;
        RECT 292.950 917.100 295.050 919.200 ;
        RECT 263.400 913.050 264.450 917.100 ;
        RECT 269.400 916.350 270.600 917.100 ;
        RECT 275.400 916.350 276.600 917.100 ;
        RECT 293.400 916.350 294.600 917.100 ;
        RECT 298.950 916.950 301.050 919.050 ;
        RECT 307.950 918.000 310.050 922.050 ;
        RECT 313.950 918.000 316.050 922.050 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 277.950 913.950 280.050 916.050 ;
        RECT 289.950 913.950 292.050 916.050 ;
        RECT 292.950 913.950 295.050 916.050 ;
        RECT 262.950 910.950 265.050 913.050 ;
        RECT 272.400 911.400 273.600 913.650 ;
        RECT 278.400 911.400 279.600 913.650 ;
        RECT 290.400 911.400 291.600 913.650 ;
        RECT 295.800 912.000 297.900 913.050 ;
        RECT 299.400 912.900 300.450 916.950 ;
        RECT 308.400 916.350 309.600 918.000 ;
        RECT 314.400 916.350 315.600 918.000 ;
        RECT 304.950 913.950 307.050 916.050 ;
        RECT 307.950 913.950 310.050 916.050 ;
        RECT 310.950 913.950 313.050 916.050 ;
        RECT 313.950 913.950 316.050 916.050 ;
        RECT 305.400 913.050 306.600 913.650 ;
        RECT 259.950 901.950 262.050 904.050 ;
        RECT 272.400 895.050 273.450 911.400 ;
        RECT 271.950 894.450 274.050 895.050 ;
        RECT 271.950 893.400 276.450 894.450 ;
        RECT 271.950 892.950 274.050 893.400 ;
        RECT 256.950 889.950 259.050 892.050 ;
        RECT 244.950 884.100 247.050 886.200 ;
        RECT 245.400 879.450 246.450 884.100 ;
        RECT 248.100 880.950 250.200 883.050 ;
        RECT 253.500 880.950 255.600 883.050 ;
        RECT 248.400 879.900 249.600 880.650 ;
        RECT 247.950 879.450 250.050 879.900 ;
        RECT 245.400 878.400 250.050 879.450 ;
        RECT 247.950 877.800 250.050 878.400 ;
        RECT 257.400 874.050 258.450 889.950 ;
        RECT 266.400 880.950 268.500 883.050 ;
        RECT 271.800 880.950 273.900 883.050 ;
        RECT 259.950 877.950 262.050 880.050 ;
        RECT 272.400 878.400 273.600 880.650 ;
        RECT 256.950 871.950 259.050 874.050 ;
        RECT 226.950 856.950 229.050 859.050 ;
        RECT 241.950 856.950 244.050 859.050 ;
        RECT 223.950 847.950 226.050 850.050 ;
        RECT 209.400 838.350 210.600 839.100 ;
        RECT 215.400 838.350 216.600 840.600 ;
        RECT 220.950 839.100 223.050 841.200 ;
        RECT 224.400 841.050 225.450 847.950 ;
        RECT 205.950 835.950 208.050 838.050 ;
        RECT 208.950 835.950 211.050 838.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 214.950 835.950 217.050 838.050 ;
        RECT 206.400 834.900 207.600 835.650 ;
        RECT 205.950 832.800 208.050 834.900 ;
        RECT 212.400 833.400 213.600 835.650 ;
        RECT 221.400 835.050 222.450 839.100 ;
        RECT 223.950 838.950 226.050 841.050 ;
        RECT 227.400 840.600 228.450 856.950 ;
        RECT 232.950 847.950 235.050 850.050 ;
        RECT 233.400 840.600 234.450 847.950 ;
        RECT 227.400 838.350 228.600 840.600 ;
        RECT 233.400 838.350 234.600 840.600 ;
        RECT 226.950 835.950 229.050 838.050 ;
        RECT 229.950 835.950 232.050 838.050 ;
        RECT 232.950 835.950 235.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 212.400 832.050 213.450 833.400 ;
        RECT 220.950 832.950 223.050 835.050 ;
        RECT 230.400 834.900 231.600 835.650 ;
        RECT 229.950 832.800 232.050 834.900 ;
        RECT 236.400 834.000 237.600 835.650 ;
        RECT 211.950 829.950 214.050 832.050 ;
        RECT 235.950 829.950 238.050 834.000 ;
        RECT 205.950 814.950 208.050 817.050 ;
        RECT 206.400 808.050 207.450 814.950 ;
        RECT 212.400 811.200 213.450 829.950 ;
        RECT 232.950 826.950 235.050 829.050 ;
        RECT 217.950 811.950 220.050 814.050 ;
        RECT 223.950 811.950 226.050 814.050 ;
        RECT 211.950 809.100 214.050 811.200 ;
        RECT 197.400 805.350 198.600 807.000 ;
        RECT 200.400 806.400 204.450 807.450 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 182.400 796.050 183.450 800.400 ;
        RECT 187.950 799.950 190.050 802.050 ;
        RECT 194.400 801.900 195.600 802.650 ;
        RECT 203.400 801.900 204.450 806.400 ;
        RECT 205.950 805.950 208.050 808.050 ;
        RECT 211.950 805.950 214.050 808.050 ;
        RECT 218.400 807.600 219.450 811.950 ;
        RECT 212.400 805.350 213.600 805.950 ;
        RECT 218.400 805.350 219.600 807.600 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 217.950 802.950 220.050 805.050 ;
        RECT 193.950 799.800 196.050 801.900 ;
        RECT 202.950 799.800 205.050 801.900 ;
        RECT 205.950 799.950 208.050 802.050 ;
        RECT 209.400 801.900 210.600 802.650 ;
        RECT 181.950 793.950 184.050 796.050 ;
        RECT 194.400 790.050 195.450 799.800 ;
        RECT 193.950 787.950 196.050 790.050 ;
        RECT 148.950 778.950 151.050 781.050 ;
        RECT 160.950 778.950 163.050 781.050 ;
        RECT 169.950 778.950 172.050 781.050 ;
        RECT 154.950 772.950 157.050 775.050 ;
        RECT 124.950 766.950 127.050 769.050 ;
        RECT 142.950 766.950 145.050 772.050 ;
        RECT 148.950 766.950 154.050 769.050 ;
        RECT 109.800 763.950 111.900 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 106.950 761.100 109.050 763.200 ;
        RECT 116.400 762.450 117.600 762.600 ;
        RECT 116.400 761.400 120.450 762.450 ;
        RECT 107.400 760.350 108.600 761.100 ;
        RECT 116.400 760.350 117.600 761.400 ;
        RECT 107.100 757.950 109.200 760.050 ;
        RECT 112.500 757.950 114.600 760.050 ;
        RECT 115.800 757.950 117.900 760.050 ;
        RECT 113.400 756.900 114.600 757.650 ;
        RECT 112.950 754.800 115.050 756.900 ;
        RECT 109.800 751.950 111.900 754.050 ;
        RECT 110.400 745.050 111.450 751.950 ;
        RECT 115.950 748.950 118.050 754.050 ;
        RECT 119.400 748.050 120.450 761.400 ;
        RECT 125.400 751.050 126.450 766.950 ;
        RECT 130.950 761.100 133.050 763.200 ;
        RECT 136.950 761.100 139.050 763.200 ;
        RECT 155.400 762.600 156.450 772.950 ;
        RECT 161.400 766.050 162.450 778.950 ;
        RECT 193.950 772.950 196.050 775.050 ;
        RECT 181.950 769.950 184.050 772.050 ;
        RECT 131.400 760.350 132.600 761.100 ;
        RECT 137.400 760.350 138.600 761.100 ;
        RECT 155.400 760.350 156.600 762.600 ;
        RECT 160.950 762.000 163.050 766.050 ;
        RECT 166.950 763.950 169.050 766.050 ;
        RECT 161.400 760.350 162.600 762.000 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 133.950 757.950 136.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 154.950 757.950 157.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 127.950 754.950 130.050 757.050 ;
        RECT 134.400 755.400 135.600 757.650 ;
        RECT 140.400 755.400 141.600 757.650 ;
        RECT 121.950 748.950 124.050 751.050 ;
        RECT 124.950 748.950 127.050 751.050 ;
        RECT 115.800 745.800 117.900 747.900 ;
        RECT 118.950 745.950 121.050 748.050 ;
        RECT 109.950 742.950 112.050 745.050 ;
        RECT 116.400 736.050 117.450 745.800 ;
        RECT 122.400 736.050 123.450 748.950 ;
        RECT 128.400 744.450 129.450 754.950 ;
        RECT 130.950 744.450 133.050 745.050 ;
        RECT 128.400 743.400 133.050 744.450 ;
        RECT 130.950 742.950 133.050 743.400 ;
        RECT 115.950 733.950 118.050 736.050 ;
        RECT 121.950 733.950 124.050 736.050 ;
        RECT 104.400 727.350 105.600 729.600 ;
        RECT 109.950 728.100 112.050 733.050 ;
        RECT 110.400 727.350 111.600 728.100 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 83.400 723.900 84.600 724.650 ;
        RECT 82.950 721.800 85.050 723.900 ;
        RECT 91.950 721.800 94.050 723.900 ;
        RECT 97.950 721.950 100.050 724.050 ;
        RECT 101.400 723.900 102.600 724.650 ;
        RECT 76.950 691.950 79.050 694.050 ;
        RECT 47.400 682.350 48.600 683.100 ;
        RECT 49.950 682.950 52.050 685.050 ;
        RECT 55.950 682.950 58.050 688.050 ;
        RECT 61.950 684.000 64.050 688.050 ;
        RECT 73.950 685.950 79.050 688.050 ;
        RECT 75.000 684.900 78.000 685.050 ;
        RECT 73.950 684.600 78.000 684.900 ;
        RECT 62.400 682.350 63.600 684.000 ;
        RECT 73.950 682.950 78.600 684.600 ;
        RECT 85.950 684.000 88.050 688.050 ;
        RECT 73.950 682.800 76.050 682.950 ;
        RECT 77.400 682.350 78.600 682.950 ;
        RECT 86.400 682.350 87.600 684.000 ;
        RECT 88.950 682.950 91.050 685.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 40.950 679.950 43.050 682.050 ;
        RECT 43.950 679.950 46.050 682.050 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 77.100 679.950 79.200 682.050 ;
        RECT 82.500 679.950 84.600 682.050 ;
        RECT 85.800 679.950 87.900 682.050 ;
        RECT 44.400 677.400 45.600 679.650 ;
        RECT 65.400 679.050 66.600 679.650 ;
        RECT 44.400 661.050 45.450 677.400 ;
        RECT 55.950 676.950 58.050 679.050 ;
        RECT 65.400 677.400 70.050 679.050 ;
        RECT 66.000 676.950 70.050 677.400 ;
        RECT 56.400 664.050 57.450 676.950 ;
        RECT 71.400 673.050 72.450 679.950 ;
        RECT 83.400 678.900 84.600 679.650 ;
        RECT 89.400 678.900 90.450 682.950 ;
        RECT 82.950 676.800 85.050 678.900 ;
        RECT 88.950 676.800 91.050 678.900 ;
        RECT 92.400 673.050 93.450 721.800 ;
        RECT 98.400 712.050 99.450 721.950 ;
        RECT 100.950 721.800 103.050 723.900 ;
        RECT 107.400 723.000 108.600 724.650 ;
        RECT 106.950 718.950 109.050 723.000 ;
        RECT 112.950 718.950 115.050 723.900 ;
        RECT 116.400 721.050 117.450 733.950 ;
        RECT 124.950 728.100 127.050 730.200 ;
        RECT 131.400 729.600 132.450 742.950 ;
        RECT 134.400 730.050 135.450 755.400 ;
        RECT 140.400 754.050 141.450 755.400 ;
        RECT 142.950 754.950 145.050 757.050 ;
        RECT 152.400 755.400 153.600 757.650 ;
        RECT 158.400 756.900 159.600 757.650 ;
        RECT 136.950 752.400 141.450 754.050 ;
        RECT 136.950 751.950 141.000 752.400 ;
        RECT 136.950 748.800 139.050 750.900 ;
        RECT 137.400 742.050 138.450 748.800 ;
        RECT 143.400 748.050 144.450 754.950 ;
        RECT 142.950 747.450 145.050 748.050 ;
        RECT 140.400 746.400 145.050 747.450 ;
        RECT 136.950 739.950 139.050 742.050 ;
        RECT 125.400 727.350 126.600 728.100 ;
        RECT 131.400 727.350 132.600 729.600 ;
        RECT 133.950 727.950 136.050 730.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 118.950 721.950 121.050 724.050 ;
        RECT 122.400 723.000 123.600 724.650 ;
        RECT 128.400 723.000 129.600 724.650 ;
        RECT 115.950 718.950 118.050 721.050 ;
        RECT 97.950 709.950 100.050 712.050 ;
        RECT 109.950 709.950 112.050 712.050 ;
        RECT 94.950 691.950 97.050 694.050 ;
        RECT 95.400 678.900 96.450 691.950 ;
        RECT 103.950 683.100 106.050 685.200 ;
        RECT 110.400 685.050 111.450 709.950 ;
        RECT 112.950 691.950 115.050 694.050 ;
        RECT 104.400 682.350 105.600 683.100 ;
        RECT 109.950 682.950 112.050 685.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 101.400 678.900 102.600 679.650 ;
        RECT 107.400 678.900 108.600 679.650 ;
        RECT 113.400 679.050 114.450 691.950 ;
        RECT 119.400 685.200 120.450 721.950 ;
        RECT 121.950 718.950 124.050 723.000 ;
        RECT 127.950 718.950 130.050 723.000 ;
        RECT 140.400 721.050 141.450 746.400 ;
        RECT 142.950 745.950 145.050 746.400 ;
        RECT 152.400 742.050 153.450 755.400 ;
        RECT 157.950 754.800 160.050 756.900 ;
        RECT 151.950 739.950 154.050 742.050 ;
        RECT 145.800 732.300 147.900 734.400 ;
        RECT 148.950 733.950 151.050 736.050 ;
        RECT 149.400 733.200 150.600 733.950 ;
        RECT 158.400 733.050 159.450 754.800 ;
        RECT 167.400 736.050 168.450 763.950 ;
        RECT 169.950 760.950 172.050 763.050 ;
        RECT 175.950 761.100 178.050 763.200 ;
        RECT 182.400 763.050 183.450 769.950 ;
        RECT 184.950 766.950 187.050 769.050 ;
        RECT 170.400 756.900 171.450 760.950 ;
        RECT 176.400 760.350 177.600 761.100 ;
        RECT 181.950 760.950 184.050 763.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 179.400 756.900 180.600 757.650 ;
        RECT 185.400 756.900 186.450 766.950 ;
        RECT 194.400 762.600 195.450 772.950 ;
        RECT 194.400 760.350 195.600 762.600 ;
        RECT 199.950 760.950 202.050 766.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 196.950 757.950 199.050 760.050 ;
        RECT 197.400 756.900 198.600 757.650 ;
        RECT 169.950 754.800 172.050 756.900 ;
        RECT 178.950 754.800 181.050 756.900 ;
        RECT 184.950 754.800 187.050 756.900 ;
        RECT 196.950 754.800 199.050 756.900 ;
        RECT 197.400 751.050 198.450 754.800 ;
        RECT 196.950 748.950 199.050 751.050 ;
        RECT 160.950 733.950 163.050 736.050 ;
        RECT 166.950 733.950 169.050 736.050 ;
        RECT 175.950 733.950 178.050 736.050 ;
        RECT 142.950 728.100 145.050 730.200 ;
        RECT 143.400 727.350 144.600 728.100 ;
        RECT 143.100 724.950 145.200 727.050 ;
        RECT 146.100 726.900 147.000 732.300 ;
        RECT 149.100 730.800 151.200 732.900 ;
        RECT 153.000 729.900 155.100 731.700 ;
        RECT 157.950 730.950 160.050 733.050 ;
        RECT 147.900 728.700 156.600 729.900 ;
        RECT 147.900 727.800 150.000 728.700 ;
        RECT 146.100 725.700 153.000 726.900 ;
        RECT 139.950 718.950 142.050 721.050 ;
        RECT 146.100 718.500 147.300 725.700 ;
        RECT 149.100 721.950 151.200 724.050 ;
        RECT 152.100 723.300 153.000 725.700 ;
        RECT 149.400 719.400 150.600 721.650 ;
        RECT 152.100 721.200 154.200 723.300 ;
        RECT 155.700 719.700 156.600 728.700 ;
        RECT 157.800 724.950 159.900 727.050 ;
        RECT 158.400 723.450 159.600 724.650 ;
        RECT 161.400 723.450 162.450 733.950 ;
        RECT 176.400 729.600 177.450 733.950 ;
        RECT 203.400 730.200 204.450 799.800 ;
        RECT 206.400 787.050 207.450 799.950 ;
        RECT 208.950 799.800 211.050 801.900 ;
        RECT 215.400 800.400 216.600 802.650 ;
        RECT 215.400 796.050 216.450 800.400 ;
        RECT 224.400 799.050 225.450 811.950 ;
        RECT 233.400 811.050 234.450 826.950 ;
        RECT 238.950 820.950 241.050 823.050 ;
        RECT 239.400 814.050 240.450 820.950 ;
        RECT 238.950 811.950 241.050 814.050 ;
        RECT 242.400 811.050 243.450 856.950 ;
        RECT 247.950 853.950 250.050 856.050 ;
        RECT 248.400 841.200 249.450 853.950 ;
        RECT 247.950 839.100 250.050 841.200 ;
        RECT 253.950 839.100 256.050 841.200 ;
        RECT 248.400 838.350 249.600 839.100 ;
        RECT 254.400 838.350 255.600 839.100 ;
        RECT 247.950 835.950 250.050 838.050 ;
        RECT 250.950 835.950 253.050 838.050 ;
        RECT 253.950 835.950 256.050 838.050 ;
        RECT 251.400 833.400 252.600 835.650 ;
        RECT 251.400 826.050 252.450 833.400 ;
        RECT 260.400 832.050 261.450 877.950 ;
        RECT 262.950 874.950 265.050 877.050 ;
        RECT 263.400 859.050 264.450 874.950 ;
        RECT 262.950 856.950 265.050 859.050 ;
        RECT 262.950 847.950 265.050 850.050 ;
        RECT 259.950 829.950 262.050 832.050 ;
        RECT 263.400 829.050 264.450 847.950 ;
        RECT 272.400 846.450 273.450 878.400 ;
        RECT 275.400 850.050 276.450 893.400 ;
        RECT 278.400 868.050 279.450 911.400 ;
        RECT 290.400 907.050 291.450 911.400 ;
        RECT 295.800 910.950 298.050 912.000 ;
        RECT 295.950 907.950 298.050 910.950 ;
        RECT 298.950 910.800 301.050 912.900 ;
        RECT 301.950 911.400 306.600 913.050 ;
        RECT 311.400 912.900 312.600 913.650 ;
        RECT 301.950 910.950 306.000 911.400 ;
        RECT 310.950 910.800 313.050 912.900 ;
        RECT 289.950 904.950 292.050 907.050 ;
        RECT 283.950 901.950 286.050 904.050 ;
        RECT 284.400 886.050 285.450 901.950 ;
        RECT 290.400 901.050 291.450 904.950 ;
        RECT 289.950 898.950 292.050 901.050 ;
        RECT 299.400 889.050 300.450 910.800 ;
        RECT 319.950 904.950 322.050 907.050 ;
        RECT 283.950 883.950 286.050 886.050 ;
        RECT 289.950 885.000 292.050 889.050 ;
        RECT 295.950 885.000 298.050 889.050 ;
        RECT 298.950 886.950 301.050 889.050 ;
        RECT 301.950 886.950 304.050 892.050 ;
        RECT 290.400 883.350 291.600 885.000 ;
        RECT 296.400 883.350 297.600 885.000 ;
        RECT 307.950 884.100 310.050 886.200 ;
        RECT 313.950 884.100 316.050 886.200 ;
        RECT 320.400 885.600 321.450 904.950 ;
        RECT 323.400 892.050 324.450 922.950 ;
        RECT 329.400 922.050 330.450 925.950 ;
        RECT 328.950 919.950 331.050 922.050 ;
        RECT 329.400 918.600 330.450 919.950 ;
        RECT 329.400 916.350 330.600 918.600 ;
        RECT 334.950 917.100 337.050 919.200 ;
        RECT 340.950 917.100 343.050 919.200 ;
        RECT 346.950 918.000 349.050 922.050 ;
        RECT 335.400 916.350 336.600 917.100 ;
        RECT 328.950 913.950 331.050 916.050 ;
        RECT 331.950 913.950 334.050 916.050 ;
        RECT 334.950 913.950 337.050 916.050 ;
        RECT 332.400 911.400 333.600 913.650 ;
        RECT 341.400 913.050 342.450 917.100 ;
        RECT 347.400 916.350 348.600 918.000 ;
        RECT 352.950 917.100 355.050 919.200 ;
        RECT 353.400 916.350 354.600 917.100 ;
        RECT 346.950 913.950 349.050 916.050 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 355.950 913.950 358.050 916.050 ;
        RECT 332.400 898.050 333.450 911.400 ;
        RECT 340.950 910.950 343.050 913.050 ;
        RECT 350.400 911.400 351.600 913.650 ;
        RECT 356.400 911.400 357.600 913.650 ;
        RECT 350.400 904.050 351.450 911.400 ;
        RECT 356.400 907.050 357.450 911.400 ;
        RECT 362.400 907.050 363.450 928.950 ;
        RECT 368.400 919.200 369.450 934.950 ;
        RECT 412.950 928.950 415.050 931.050 ;
        RECT 463.950 928.950 466.050 931.050 ;
        RECT 502.950 928.950 505.050 931.050 ;
        RECT 514.950 928.950 517.050 931.050 ;
        RECT 367.950 917.100 370.050 919.200 ;
        RECT 373.950 917.100 376.050 919.200 ;
        RECT 379.950 917.100 382.050 919.200 ;
        RECT 385.950 918.000 388.050 922.050 ;
        RECT 391.950 918.000 394.050 922.050 ;
        RECT 400.950 919.950 403.050 922.050 ;
        RECT 368.400 916.350 369.600 917.100 ;
        RECT 374.400 916.350 375.600 917.100 ;
        RECT 367.950 913.950 370.050 916.050 ;
        RECT 370.950 913.950 373.050 916.050 ;
        RECT 373.950 913.950 376.050 916.050 ;
        RECT 371.400 912.900 372.600 913.650 ;
        RECT 380.400 913.050 381.450 917.100 ;
        RECT 386.400 916.350 387.600 918.000 ;
        RECT 392.400 916.350 393.600 918.000 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 388.950 913.950 391.050 916.050 ;
        RECT 391.950 913.950 394.050 916.050 ;
        RECT 394.950 913.950 397.050 916.050 ;
        RECT 370.950 910.800 373.050 912.900 ;
        RECT 379.950 910.950 382.050 913.050 ;
        RECT 389.400 912.900 390.600 913.650 ;
        RECT 388.950 910.800 391.050 912.900 ;
        RECT 395.400 911.400 396.600 913.650 ;
        RECT 401.400 913.050 402.450 919.950 ;
        RECT 413.400 918.600 414.450 928.950 ;
        RECT 418.950 925.950 424.050 928.050 ;
        RECT 424.950 922.950 427.050 928.050 ;
        RECT 421.950 919.950 424.050 922.050 ;
        RECT 413.400 916.350 414.600 918.600 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 412.950 913.950 415.050 916.050 ;
        RECT 415.950 913.950 418.050 916.050 ;
        RECT 395.400 907.050 396.450 911.400 ;
        RECT 400.950 910.950 403.050 913.050 ;
        RECT 410.400 912.900 411.600 913.650 ;
        RECT 409.950 910.800 412.050 912.900 ;
        RECT 416.400 911.400 417.600 913.650 ;
        RECT 422.400 913.050 423.450 919.950 ;
        RECT 424.950 917.100 427.050 919.200 ;
        RECT 430.950 917.100 433.050 919.200 ;
        RECT 436.950 917.100 439.050 919.200 ;
        RECT 445.950 917.100 448.050 919.200 ;
        RECT 448.950 918.600 453.000 919.050 ;
        RECT 410.400 909.450 411.450 910.800 ;
        RECT 410.400 908.400 414.450 909.450 ;
        RECT 355.950 904.950 358.050 907.050 ;
        RECT 361.950 904.950 364.050 907.050 ;
        RECT 394.950 904.950 397.050 907.050 ;
        RECT 349.950 901.950 352.050 904.050 ;
        RECT 331.950 895.950 334.050 898.050 ;
        RECT 400.950 895.950 403.050 898.050 ;
        RECT 409.950 895.950 412.050 898.050 ;
        RECT 401.400 892.050 402.450 895.950 ;
        RECT 322.950 889.950 325.050 892.050 ;
        RECT 346.950 891.450 349.050 892.050 ;
        RECT 338.400 890.400 349.050 891.450 ;
        RECT 338.400 889.050 339.450 890.400 ;
        RECT 346.950 889.950 349.050 890.400 ;
        RECT 355.950 891.450 360.000 892.050 ;
        RECT 355.950 891.000 360.450 891.450 ;
        RECT 355.950 889.950 361.050 891.000 ;
        RECT 400.950 889.950 403.050 892.050 ;
        RECT 334.950 887.400 339.450 889.050 ;
        RECT 340.950 888.450 345.000 889.050 ;
        RECT 334.950 886.950 339.000 887.400 ;
        RECT 340.950 886.950 345.450 888.450 ;
        RECT 358.950 886.950 361.050 889.950 ;
        RECT 286.950 880.950 289.050 883.050 ;
        RECT 289.950 880.950 292.050 883.050 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 287.400 879.900 288.600 880.650 ;
        RECT 286.950 877.800 289.050 879.900 ;
        RECT 293.400 878.400 294.600 880.650 ;
        RECT 299.400 878.400 300.600 880.650 ;
        RECT 277.950 865.950 280.050 868.050 ;
        RECT 274.950 847.950 277.050 850.050 ;
        RECT 272.400 846.000 276.450 846.450 ;
        RECT 272.400 845.400 277.050 846.000 ;
        RECT 274.950 841.950 277.050 845.400 ;
        RECT 271.950 839.100 274.050 841.200 ;
        RECT 278.400 841.050 279.450 865.950 ;
        RECT 293.400 853.050 294.450 878.400 ;
        RECT 299.400 871.050 300.450 878.400 ;
        RECT 308.400 871.050 309.450 884.100 ;
        RECT 314.400 883.350 315.600 884.100 ;
        RECT 320.400 883.350 321.600 885.600 ;
        RECT 328.950 883.950 331.050 886.050 ;
        RECT 337.950 884.100 340.050 886.200 ;
        RECT 344.400 885.600 345.450 886.950 ;
        RECT 313.950 880.950 316.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 322.950 880.950 325.050 883.050 ;
        RECT 317.400 879.900 318.600 880.650 ;
        RECT 316.950 877.800 319.050 879.900 ;
        RECT 323.400 879.000 324.600 880.650 ;
        RECT 322.950 874.950 325.050 879.000 ;
        RECT 329.400 877.050 330.450 883.950 ;
        RECT 338.400 883.350 339.600 884.100 ;
        RECT 344.400 883.350 345.600 885.600 ;
        RECT 349.950 884.100 352.050 886.200 ;
        RECT 355.950 884.100 358.050 886.200 ;
        RECT 376.950 885.000 379.050 889.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 343.950 880.950 346.050 883.050 ;
        RECT 335.400 878.400 336.600 880.650 ;
        RECT 341.400 879.900 342.600 880.650 ;
        RECT 350.400 880.050 351.450 884.100 ;
        RECT 356.400 883.350 357.600 884.100 ;
        RECT 377.400 883.350 378.600 885.000 ;
        RECT 382.950 884.100 385.050 886.200 ;
        RECT 383.400 883.350 384.600 884.100 ;
        RECT 388.950 883.950 391.050 886.050 ;
        RECT 394.950 884.100 397.050 886.200 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 358.950 880.950 361.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 382.950 880.950 385.050 883.050 ;
        RECT 328.950 874.950 331.050 877.050 ;
        RECT 335.400 871.050 336.450 878.400 ;
        RECT 340.950 877.800 343.050 879.900 ;
        RECT 349.950 877.950 352.050 880.050 ;
        RECT 359.400 879.900 360.600 880.650 ;
        RECT 374.400 879.900 375.600 880.650 ;
        RECT 358.950 877.800 361.050 879.900 ;
        RECT 373.950 877.800 376.050 879.900 ;
        RECT 380.400 879.000 381.600 880.650 ;
        RECT 298.950 868.950 301.050 871.050 ;
        RECT 307.950 868.950 310.050 871.050 ;
        RECT 334.950 868.950 337.050 871.050 ;
        RECT 337.950 865.950 340.050 868.050 ;
        RECT 334.950 853.950 337.050 856.050 ;
        RECT 292.950 850.950 295.050 853.050 ;
        RECT 313.950 850.950 316.050 853.050 ;
        RECT 289.800 844.200 291.900 846.300 ;
        RECT 298.800 844.500 300.900 846.600 ;
        RECT 310.950 844.950 313.050 847.050 ;
        RECT 283.950 841.950 286.050 844.050 ;
        RECT 272.400 838.350 273.600 839.100 ;
        RECT 277.950 838.950 280.050 841.050 ;
        RECT 268.950 835.950 271.050 838.050 ;
        RECT 271.950 835.950 274.050 838.050 ;
        RECT 274.950 835.950 277.050 838.050 ;
        RECT 269.400 834.900 270.600 835.650 ;
        RECT 268.950 832.800 271.050 834.900 ;
        RECT 275.400 833.400 276.600 835.650 ;
        RECT 262.950 826.950 265.050 829.050 ;
        RECT 275.400 826.050 276.450 833.400 ;
        RECT 250.950 823.950 253.050 826.050 ;
        RECT 274.950 823.950 277.050 826.050 ;
        RECT 268.950 817.950 271.050 820.050 ;
        RECT 280.950 817.950 283.050 820.050 ;
        RECT 250.950 811.950 253.050 814.050 ;
        RECT 262.950 811.950 265.050 814.050 ;
        RECT 232.950 808.950 235.050 811.050 ;
        RECT 241.950 808.950 244.050 811.050 ;
        RECT 247.950 808.950 250.050 811.050 ;
        RECT 233.400 807.450 234.600 807.600 ;
        RECT 227.400 806.400 234.600 807.450 ;
        RECT 223.950 796.950 226.050 799.050 ;
        RECT 214.950 793.950 217.050 796.050 ;
        RECT 205.950 784.950 208.050 787.050 ;
        RECT 217.950 784.950 220.050 787.050 ;
        RECT 214.950 772.950 217.050 775.050 ;
        RECT 208.950 761.100 211.050 763.200 ;
        RECT 215.400 762.600 216.450 772.950 ;
        RECT 218.400 772.050 219.450 784.950 ;
        RECT 227.400 775.050 228.450 806.400 ;
        RECT 233.400 805.350 234.600 806.400 ;
        RECT 238.950 806.100 241.050 808.200 ;
        RECT 239.400 805.350 240.600 806.100 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 238.950 802.950 241.050 805.050 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 236.400 801.900 237.600 802.650 ;
        RECT 242.400 801.900 243.600 802.650 ;
        RECT 235.950 799.800 238.050 801.900 ;
        RECT 241.950 799.800 244.050 801.900 ;
        RECT 248.400 799.050 249.450 808.950 ;
        RECT 251.400 799.050 252.450 811.950 ;
        RECT 256.950 806.100 259.050 808.200 ;
        RECT 263.400 807.600 264.450 811.950 ;
        RECT 269.400 807.600 270.450 817.950 ;
        RECT 277.950 814.950 280.050 817.050 ;
        RECT 278.400 808.050 279.450 814.950 ;
        RECT 281.400 813.450 282.450 817.950 ;
        RECT 284.400 817.050 285.450 841.950 ;
        RECT 286.950 839.100 289.050 841.200 ;
        RECT 287.400 838.350 288.600 839.100 ;
        RECT 287.100 835.950 289.200 838.050 ;
        RECT 290.100 831.600 291.000 844.200 ;
        RECT 296.400 841.350 297.600 843.600 ;
        RECT 296.100 838.950 298.200 841.050 ;
        RECT 291.900 837.900 294.000 838.200 ;
        RECT 300.000 837.900 300.900 844.500 ;
        RECT 291.900 837.000 300.900 837.900 ;
        RECT 291.900 836.100 294.000 837.000 ;
        RECT 297.000 835.200 299.100 836.100 ;
        RECT 291.900 834.000 299.100 835.200 ;
        RECT 291.900 833.100 294.000 834.000 ;
        RECT 289.500 829.500 291.600 831.600 ;
        RECT 292.950 828.450 295.050 832.050 ;
        RECT 296.100 830.100 298.200 832.200 ;
        RECT 300.000 831.900 300.900 837.000 ;
        RECT 301.800 835.950 303.900 838.050 ;
        RECT 302.400 834.450 303.600 835.650 ;
        RECT 304.950 834.450 307.050 834.900 ;
        RECT 302.400 833.400 307.050 834.450 ;
        RECT 304.950 832.800 307.050 833.400 ;
        RECT 299.400 829.800 301.500 831.900 ;
        RECT 296.400 828.450 297.600 829.800 ;
        RECT 292.950 828.000 297.600 828.450 ;
        RECT 293.400 827.550 297.600 828.000 ;
        RECT 293.400 827.400 297.450 827.550 ;
        RECT 286.950 823.950 289.050 826.050 ;
        RECT 292.800 823.950 294.900 826.050 ;
        RECT 295.950 823.950 298.050 826.050 ;
        RECT 287.400 820.050 288.450 823.950 ;
        RECT 286.950 817.950 289.050 820.050 ;
        RECT 283.950 814.950 286.050 817.050 ;
        RECT 281.400 812.400 285.450 813.450 ;
        RECT 257.400 805.350 258.600 806.100 ;
        RECT 263.400 805.350 264.600 807.600 ;
        RECT 269.400 805.350 270.600 807.600 ;
        RECT 277.950 805.950 280.050 808.050 ;
        RECT 284.400 807.600 285.450 812.400 ;
        RECT 284.400 805.350 285.600 807.600 ;
        RECT 289.950 806.100 292.050 808.200 ;
        RECT 293.400 808.050 294.450 823.950 ;
        RECT 296.400 820.050 297.450 823.950 ;
        RECT 298.950 820.950 301.050 823.050 ;
        RECT 295.950 817.950 298.050 820.050 ;
        RECT 290.400 805.350 291.600 806.100 ;
        RECT 292.950 805.950 295.050 808.050 ;
        RECT 295.950 806.100 298.050 808.200 ;
        RECT 256.950 802.950 259.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 280.950 802.950 283.050 805.050 ;
        RECT 283.950 802.950 286.050 805.050 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 253.950 799.950 256.050 802.050 ;
        RECT 260.400 800.400 261.600 802.650 ;
        RECT 266.400 800.400 267.600 802.650 ;
        RECT 281.400 800.400 282.600 802.650 ;
        RECT 287.400 801.900 288.600 802.650 ;
        RECT 241.950 796.650 244.050 798.750 ;
        RECT 247.950 796.950 250.050 799.050 ;
        RECT 250.950 796.950 253.050 799.050 ;
        RECT 229.950 793.950 232.050 796.050 ;
        RECT 230.400 781.050 231.450 793.950 ;
        RECT 229.950 778.950 232.050 781.050 ;
        RECT 226.950 772.950 229.050 775.050 ;
        RECT 217.950 769.950 220.050 772.050 ;
        RECT 209.400 760.350 210.600 761.100 ;
        RECT 215.400 760.350 216.600 762.600 ;
        RECT 223.950 761.100 226.050 763.200 ;
        RECT 229.950 761.100 232.050 763.200 ;
        RECT 235.950 762.000 238.050 766.050 ;
        RECT 242.400 762.450 243.450 796.650 ;
        RECT 254.400 796.050 255.450 799.950 ;
        RECT 247.950 793.800 250.050 795.900 ;
        RECT 253.950 793.950 256.050 796.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 217.950 757.950 220.050 760.050 ;
        RECT 205.950 751.950 208.050 757.050 ;
        RECT 212.400 756.000 213.600 757.650 ;
        RECT 218.400 756.900 219.600 757.650 ;
        RECT 211.950 751.950 214.050 756.000 ;
        RECT 217.950 754.800 220.050 756.900 ;
        RECT 224.400 751.050 225.450 761.100 ;
        RECT 230.400 760.350 231.600 761.100 ;
        RECT 236.400 760.350 237.600 762.000 ;
        RECT 242.400 761.400 246.450 762.450 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 233.400 756.900 234.600 757.650 ;
        RECT 239.400 756.900 240.600 757.650 ;
        RECT 232.950 754.800 235.050 756.900 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 223.950 748.950 226.050 751.050 ;
        RECT 245.400 750.450 246.450 761.400 ;
        RECT 242.400 749.400 246.450 750.450 ;
        RECT 205.950 745.950 208.050 748.050 ;
        RECT 176.400 727.350 177.600 729.600 ;
        RECT 193.950 728.100 196.050 730.200 ;
        RECT 202.950 728.100 205.050 730.200 ;
        RECT 206.400 729.600 207.450 745.950 ;
        RECT 211.950 736.950 214.050 739.050 ;
        RECT 212.400 733.050 213.450 736.950 ;
        RECT 223.950 733.950 226.050 736.050 ;
        RECT 211.950 730.950 214.050 733.050 ;
        RECT 212.400 729.600 213.450 730.950 ;
        RECT 194.400 727.350 195.600 728.100 ;
        RECT 206.400 727.350 207.600 729.600 ;
        RECT 212.400 727.350 213.600 729.600 ;
        RECT 220.950 727.950 223.050 730.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 205.950 724.950 208.050 727.050 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 158.400 722.400 162.450 723.450 ;
        RECT 173.400 722.400 174.600 724.650 ;
        RECT 191.400 723.000 192.600 724.650 ;
        RECT 209.400 723.900 210.600 724.650 ;
        RECT 145.800 716.400 147.900 718.500 ;
        RECT 155.400 717.600 157.500 719.700 ;
        RECT 169.950 718.950 172.050 721.050 ;
        RECT 139.950 691.950 142.050 694.050 ;
        RECT 118.950 683.100 121.050 685.200 ;
        RECT 124.950 683.100 127.050 685.200 ;
        RECT 140.400 684.600 141.450 691.950 ;
        RECT 145.950 688.950 148.050 691.050 ;
        RECT 146.400 684.600 147.450 688.950 ;
        RECT 170.400 685.050 171.450 718.950 ;
        RECT 173.400 706.050 174.450 722.400 ;
        RECT 190.950 718.950 193.050 723.000 ;
        RECT 208.950 721.800 211.050 723.900 ;
        RECT 215.400 722.400 216.600 724.650 ;
        RECT 221.400 723.900 222.450 727.950 ;
        RECT 208.950 718.650 211.050 720.750 ;
        RECT 175.950 706.950 178.050 709.050 ;
        RECT 172.950 703.950 175.050 706.050 ;
        RECT 176.400 691.050 177.450 706.950 ;
        RECT 202.950 691.950 205.050 694.050 ;
        RECT 175.950 688.950 178.050 691.050 ;
        RECT 119.400 682.350 120.600 683.100 ;
        RECT 125.400 682.350 126.600 683.100 ;
        RECT 140.400 682.350 141.600 684.600 ;
        RECT 146.400 682.350 147.600 684.600 ;
        RECT 154.950 682.950 157.050 685.050 ;
        RECT 163.950 682.950 166.050 685.050 ;
        RECT 169.950 682.950 172.050 685.050 ;
        RECT 181.950 683.100 184.050 685.200 ;
        RECT 187.950 684.000 190.050 688.050 ;
        RECT 193.950 685.950 196.050 688.050 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 121.950 679.950 124.050 682.050 ;
        RECT 124.950 679.950 127.050 682.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 145.950 679.950 148.050 682.050 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 94.950 676.800 97.050 678.900 ;
        RECT 100.950 676.800 103.050 678.900 ;
        RECT 106.950 676.800 109.050 678.900 ;
        RECT 112.950 676.950 115.050 679.050 ;
        RECT 122.400 678.900 123.600 679.650 ;
        RECT 121.950 676.800 124.050 678.900 ;
        RECT 143.400 677.400 144.600 679.650 ;
        RECT 149.400 678.900 150.600 679.650 ;
        RECT 148.950 678.450 151.050 678.900 ;
        RECT 148.950 678.000 153.450 678.450 ;
        RECT 148.950 677.400 154.050 678.000 ;
        RECT 112.950 673.800 115.050 675.900 ;
        RECT 70.950 670.950 73.050 673.050 ;
        RECT 85.950 670.950 88.050 673.050 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 103.950 670.950 106.050 673.050 ;
        RECT 55.950 661.950 58.050 664.050 ;
        RECT 43.950 658.950 46.050 661.050 ;
        RECT 49.950 658.950 52.050 661.050 ;
        RECT 50.400 651.600 51.450 658.950 ;
        RECT 86.400 652.200 87.450 670.950 ;
        RECT 50.400 649.350 51.600 651.600 ;
        RECT 55.950 650.100 58.050 652.200 ;
        RECT 56.400 649.350 57.600 650.100 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 85.950 650.100 88.050 652.200 ;
        RECT 104.400 651.600 105.450 670.950 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 38.400 644.400 39.600 646.650 ;
        RECT 53.400 644.400 54.600 646.650 ;
        RECT 59.400 645.000 60.600 646.650 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 28.950 610.950 31.050 613.050 ;
        RECT 14.400 608.400 18.450 609.450 ;
        RECT 14.400 592.050 15.450 608.400 ;
        RECT 31.950 607.950 34.050 610.050 ;
        RECT 22.950 605.100 25.050 607.200 ;
        RECT 28.950 605.100 31.050 607.200 ;
        RECT 23.400 604.350 24.600 605.100 ;
        RECT 17.100 601.950 19.200 604.050 ;
        RECT 23.100 601.950 25.200 604.050 ;
        RECT 29.400 601.050 30.450 605.100 ;
        RECT 19.950 598.950 22.050 601.050 ;
        RECT 25.950 598.950 28.050 601.050 ;
        RECT 28.950 598.950 31.050 601.050 ;
        RECT 13.950 589.950 16.050 592.050 ;
        RECT 16.950 572.100 19.050 574.200 ;
        RECT 17.400 571.350 18.600 572.100 ;
        RECT 11.100 568.950 13.200 571.050 ;
        RECT 16.500 568.950 18.600 571.050 ;
        RECT 20.400 550.050 21.450 598.950 ;
        RECT 26.400 573.450 27.450 598.950 ;
        RECT 28.950 582.450 31.050 583.050 ;
        RECT 32.400 582.450 33.450 607.950 ;
        RECT 35.400 607.050 36.450 628.950 ;
        RECT 38.400 619.050 39.450 644.400 ;
        RECT 53.400 637.050 54.450 644.400 ;
        RECT 58.950 640.950 61.050 645.000 ;
        RECT 52.950 634.950 55.050 637.050 ;
        RECT 58.950 634.950 61.050 637.050 ;
        RECT 37.950 616.950 40.050 619.050 ;
        RECT 55.950 616.950 58.050 619.050 ;
        RECT 34.950 604.950 37.050 607.050 ;
        RECT 40.950 606.000 43.050 610.050 ;
        RECT 41.400 604.350 42.600 606.000 ;
        RECT 46.950 605.100 49.050 607.200 ;
        RECT 52.950 605.100 55.050 607.200 ;
        RECT 47.400 604.350 48.600 605.100 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 46.950 601.950 49.050 604.050 ;
        RECT 28.950 581.400 33.450 582.450 ;
        RECT 38.400 599.400 39.600 601.650 ;
        RECT 44.400 599.400 45.600 601.650 ;
        RECT 28.950 580.950 31.050 581.400 ;
        RECT 23.400 572.400 27.450 573.450 ;
        RECT 29.400 573.600 30.450 580.950 ;
        RECT 38.400 576.450 39.450 599.400 ;
        RECT 44.400 592.050 45.450 599.400 ;
        RECT 53.400 595.050 54.450 605.100 ;
        RECT 52.950 592.950 55.050 595.050 ;
        RECT 56.400 592.050 57.450 616.950 ;
        RECT 59.400 607.050 60.450 634.950 ;
        RECT 65.400 625.050 66.450 649.950 ;
        RECT 86.400 649.350 87.600 650.100 ;
        RECT 104.400 649.350 105.600 651.600 ;
        RECT 70.950 646.950 73.050 649.050 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 88.950 646.950 91.050 649.050 ;
        RECT 91.950 646.950 94.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 71.400 645.900 72.600 646.650 ;
        RECT 70.950 643.800 73.050 645.900 ;
        RECT 89.400 644.400 90.600 646.650 ;
        RECT 64.950 622.950 67.050 625.050 ;
        RECT 89.400 619.050 90.450 644.400 ;
        RECT 97.950 643.950 100.050 646.050 ;
        RECT 107.400 644.400 108.600 646.650 ;
        RECT 94.950 640.950 97.050 643.050 ;
        RECT 88.950 616.950 91.050 619.050 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 64.950 605.100 67.050 607.200 ;
        RECT 85.950 605.100 88.050 607.200 ;
        RECT 65.400 604.350 66.600 605.100 ;
        RECT 86.400 604.350 87.600 605.100 ;
        RECT 95.400 604.050 96.450 640.950 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 85.950 601.950 88.050 604.050 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 94.950 601.950 97.050 604.050 ;
        RECT 62.400 600.900 63.600 601.650 ;
        RECT 61.950 598.800 64.050 600.900 ;
        RECT 83.400 599.400 84.600 601.650 ;
        RECT 89.400 599.400 90.600 601.650 ;
        RECT 43.950 589.950 46.050 592.050 ;
        RECT 55.950 589.950 58.050 592.050 ;
        RECT 62.400 589.050 63.450 598.800 ;
        RECT 64.950 592.950 67.050 595.050 ;
        RECT 61.950 586.950 64.050 589.050 ;
        RECT 65.400 586.050 66.450 592.950 ;
        RECT 79.950 589.950 82.050 592.050 ;
        RECT 64.950 583.950 67.050 586.050 ;
        RECT 58.950 580.950 61.050 583.050 ;
        RECT 59.400 577.050 60.450 580.950 ;
        RECT 38.400 576.000 42.450 576.450 ;
        RECT 38.400 575.400 43.050 576.000 ;
        RECT 23.400 565.050 24.450 572.400 ;
        RECT 29.400 571.350 30.600 573.600 ;
        RECT 34.950 572.100 37.050 574.200 ;
        RECT 35.400 571.350 36.600 572.100 ;
        RECT 40.950 571.950 43.050 575.400 ;
        RECT 58.950 574.950 61.050 577.050 ;
        RECT 64.950 574.950 67.050 577.050 ;
        RECT 43.950 571.950 46.050 574.050 ;
        RECT 52.950 572.100 55.050 574.200 ;
        RECT 61.950 572.100 64.050 574.200 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 25.950 565.950 28.050 568.050 ;
        RECT 32.400 567.000 33.600 568.650 ;
        RECT 22.950 562.950 25.050 565.050 ;
        RECT 26.400 556.050 27.450 565.950 ;
        RECT 31.950 562.950 34.050 567.000 ;
        RECT 38.400 566.400 39.600 568.650 ;
        RECT 38.400 562.050 39.450 566.400 ;
        RECT 37.950 559.950 40.050 562.050 ;
        RECT 25.950 553.950 28.050 556.050 ;
        RECT 13.950 547.950 16.050 550.050 ;
        RECT 19.950 547.950 22.050 550.050 ;
        RECT 14.400 544.050 15.450 547.950 ;
        RECT 44.400 547.050 45.450 571.950 ;
        RECT 53.400 571.350 54.600 572.100 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 46.950 565.950 49.050 568.050 ;
        RECT 50.400 567.000 51.600 568.650 ;
        RECT 56.400 567.000 57.600 568.650 ;
        RECT 47.400 547.050 48.450 565.950 ;
        RECT 49.950 562.950 52.050 567.000 ;
        RECT 55.950 562.950 58.050 567.000 ;
        RECT 28.950 544.950 31.050 547.050 ;
        RECT 43.800 544.950 45.900 547.050 ;
        RECT 46.950 544.950 49.050 547.050 ;
        RECT 58.950 544.950 61.050 547.050 ;
        RECT 13.950 541.950 16.050 544.050 ;
        RECT 7.950 532.950 10.050 535.050 ;
        RECT 1.800 529.950 3.900 532.050 ;
        RECT 4.950 530.100 7.050 532.200 ;
        RECT 5.400 529.350 6.600 530.100 ;
        RECT 4.800 526.950 6.900 529.050 ;
        RECT 10.800 526.950 12.900 529.050 ;
        RECT 1.950 523.950 4.050 526.050 ;
        RECT 7.950 523.950 10.050 526.050 ;
        RECT 2.400 418.200 3.450 523.950 ;
        RECT 4.950 493.950 7.050 496.050 ;
        RECT 5.400 453.450 6.450 493.950 ;
        RECT 8.400 487.050 9.450 523.950 ;
        RECT 14.400 511.050 15.450 541.950 ;
        RECT 17.400 540.300 20.400 542.400 ;
        RECT 21.300 540.300 23.400 542.400 ;
        RECT 17.400 521.400 18.900 540.300 ;
        RECT 21.300 534.300 22.500 540.300 ;
        RECT 20.400 532.200 22.500 534.300 ;
        RECT 17.400 519.300 19.500 521.400 ;
        RECT 18.300 515.700 19.500 519.300 ;
        RECT 21.300 515.700 22.500 532.200 ;
        RECT 23.700 537.300 25.800 539.400 ;
        RECT 23.700 515.700 24.900 537.300 ;
        RECT 29.400 525.600 30.450 544.950 ;
        RECT 40.200 540.300 42.300 542.400 ;
        RECT 32.400 535.800 34.500 537.900 ;
        RECT 37.800 537.300 39.900 539.400 ;
        RECT 32.400 529.200 33.300 535.800 ;
        RECT 38.100 530.100 39.300 537.300 ;
        RECT 40.800 535.500 42.300 540.300 ;
        RECT 43.200 537.300 45.300 542.400 ;
        RECT 40.800 533.400 42.900 535.500 ;
        RECT 32.400 527.100 34.500 529.200 ;
        RECT 37.800 528.000 39.900 530.100 ;
        RECT 29.400 523.350 30.600 525.600 ;
        RECT 28.800 520.950 30.900 523.050 ;
        RECT 32.400 516.600 33.300 527.100 ;
        RECT 35.100 520.500 37.200 522.600 ;
        RECT 17.700 513.600 19.800 515.700 ;
        RECT 20.700 513.600 22.800 515.700 ;
        RECT 23.700 513.600 25.800 515.700 ;
        RECT 31.800 514.500 33.900 516.600 ;
        RECT 38.100 515.700 39.300 528.000 ;
        RECT 40.800 515.700 42.300 533.400 ;
        RECT 44.100 515.700 45.300 537.300 ;
        RECT 37.200 513.600 39.300 515.700 ;
        RECT 40.200 513.600 42.300 515.700 ;
        RECT 43.200 513.600 45.300 515.700 ;
        RECT 46.200 540.300 48.300 542.400 ;
        RECT 46.200 535.500 47.700 540.300 ;
        RECT 46.200 533.400 48.300 535.500 ;
        RECT 46.200 515.700 47.700 533.400 ;
        RECT 49.950 529.950 52.050 532.050 ;
        RECT 46.200 513.600 48.300 515.700 ;
        RECT 13.950 508.950 16.050 511.050 ;
        RECT 19.950 508.950 22.050 511.050 ;
        RECT 28.950 508.950 31.050 511.050 ;
        RECT 10.950 502.950 13.050 505.050 ;
        RECT 7.950 484.950 10.050 487.050 ;
        RECT 11.400 460.050 12.450 502.950 ;
        RECT 20.400 496.200 21.450 508.950 ;
        RECT 19.950 494.100 22.050 496.200 ;
        RECT 20.400 493.350 21.600 494.100 ;
        RECT 29.400 493.050 30.450 508.950 ;
        RECT 50.400 508.050 51.450 529.950 ;
        RECT 55.800 526.950 57.900 529.050 ;
        RECT 56.400 525.000 57.600 526.650 ;
        RECT 55.950 520.950 58.050 525.000 ;
        RECT 59.400 511.050 60.450 544.950 ;
        RECT 62.400 532.050 63.450 572.100 ;
        RECT 65.400 547.050 66.450 574.950 ;
        RECT 73.950 573.000 76.050 577.050 ;
        RECT 80.400 574.200 81.450 589.950 ;
        RECT 83.400 577.050 84.450 599.400 ;
        RECT 89.400 592.050 90.450 599.400 ;
        RECT 91.950 598.950 94.050 601.050 ;
        RECT 88.950 589.950 91.050 592.050 ;
        RECT 82.950 574.950 85.050 577.050 ;
        RECT 88.950 574.950 91.050 577.050 ;
        RECT 74.400 571.350 75.600 573.000 ;
        RECT 79.950 572.100 82.050 574.200 ;
        RECT 80.400 571.350 81.600 572.100 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 71.400 567.900 72.600 568.650 ;
        RECT 70.950 565.800 73.050 567.900 ;
        RECT 77.400 566.400 78.600 568.650 ;
        RECT 83.400 566.400 84.600 568.650 ;
        RECT 67.950 553.950 70.050 556.050 ;
        RECT 64.950 544.950 67.050 547.050 ;
        RECT 61.950 529.950 64.050 532.050 ;
        RECT 68.400 529.050 69.450 553.950 ;
        RECT 71.400 553.050 72.450 565.800 ;
        RECT 77.400 565.050 78.450 566.400 ;
        RECT 73.950 563.550 78.450 565.050 ;
        RECT 73.950 562.950 78.000 563.550 ;
        RECT 73.950 559.800 76.050 561.900 ;
        RECT 70.950 550.950 73.050 553.050 ;
        RECT 74.400 549.450 75.450 559.800 ;
        RECT 71.400 548.400 75.450 549.450 ;
        RECT 64.800 526.950 66.900 529.050 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 65.400 525.450 66.600 526.650 ;
        RECT 67.950 525.450 70.050 529.050 ;
        RECT 65.400 525.000 70.050 525.450 ;
        RECT 65.400 524.400 69.450 525.000 ;
        RECT 62.400 517.050 63.450 523.950 ;
        RECT 71.400 523.050 72.450 548.400 ;
        RECT 83.400 538.050 84.450 566.400 ;
        RECT 85.950 565.950 88.050 568.050 ;
        RECT 86.400 559.050 87.450 565.950 ;
        RECT 89.400 565.050 90.450 574.950 ;
        RECT 92.400 574.050 93.450 598.950 ;
        RECT 98.400 598.050 99.450 643.950 ;
        RECT 107.400 622.050 108.450 644.400 ;
        RECT 113.400 637.050 114.450 673.800 ;
        RECT 143.400 667.050 144.450 677.400 ;
        RECT 148.950 676.800 151.050 677.400 ;
        RECT 151.950 673.950 154.050 677.400 ;
        RECT 115.950 664.950 118.050 667.050 ;
        RECT 142.800 664.950 144.900 667.050 ;
        RECT 145.950 664.950 148.050 667.050 ;
        RECT 151.950 664.950 154.050 667.050 ;
        RECT 112.950 634.950 115.050 637.050 ;
        RECT 106.950 619.950 109.050 622.050 ;
        RECT 116.400 616.050 117.450 664.950 ;
        RECT 121.950 661.950 124.050 664.050 ;
        RECT 122.400 651.600 123.450 661.950 ;
        RECT 133.950 658.950 136.050 661.050 ;
        RECT 122.400 649.350 123.600 651.600 ;
        RECT 127.950 650.100 130.050 652.200 ;
        RECT 128.400 649.350 129.600 650.100 ;
        RECT 121.950 646.950 124.050 649.050 ;
        RECT 124.950 646.950 127.050 649.050 ;
        RECT 127.950 646.950 130.050 649.050 ;
        RECT 125.400 645.900 126.600 646.650 ;
        RECT 134.400 646.050 135.450 658.950 ;
        RECT 142.950 651.450 145.050 652.200 ;
        RECT 146.400 651.450 147.450 664.950 ;
        RECT 142.950 650.400 147.450 651.450 ;
        RECT 142.950 650.100 145.050 650.400 ;
        RECT 143.400 649.350 144.600 650.100 ;
        RECT 148.950 649.950 151.050 652.050 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 142.950 646.950 145.050 649.050 ;
        RECT 124.950 643.800 127.050 645.900 ;
        RECT 133.950 643.950 136.050 646.050 ;
        RECT 140.400 645.900 141.600 646.650 ;
        RECT 149.400 645.900 150.450 649.950 ;
        RECT 139.950 640.950 142.050 645.900 ;
        RECT 148.950 643.800 151.050 645.900 ;
        RECT 139.950 634.950 142.050 637.050 ;
        RECT 124.950 622.950 127.050 625.050 ;
        RECT 106.950 613.950 109.050 616.050 ;
        RECT 115.950 613.950 118.050 616.050 ;
        RECT 121.950 613.950 124.050 616.050 ;
        RECT 107.400 606.600 108.450 613.950 ;
        RECT 115.950 610.800 118.050 612.900 ;
        RECT 107.400 604.350 108.600 606.600 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 106.950 601.950 109.050 604.050 ;
        RECT 109.950 601.950 112.050 604.050 ;
        RECT 110.400 600.000 111.600 601.650 ;
        RECT 97.950 595.950 100.050 598.050 ;
        RECT 103.950 595.950 106.050 598.050 ;
        RECT 109.950 595.950 112.050 600.000 ;
        RECT 104.400 577.050 105.450 595.950 ;
        RECT 116.400 595.050 117.450 610.800 ;
        RECT 109.950 589.950 112.050 594.900 ;
        RECT 115.950 592.950 118.050 595.050 ;
        RECT 122.400 592.050 123.450 613.950 ;
        RECT 125.400 606.600 126.450 622.950 ;
        RECT 125.400 604.350 126.600 606.600 ;
        RECT 134.400 606.450 135.600 606.600 ;
        RECT 134.400 605.400 138.450 606.450 ;
        RECT 134.400 604.350 135.600 605.400 ;
        RECT 125.100 601.950 127.200 604.050 ;
        RECT 128.400 601.950 130.500 604.050 ;
        RECT 133.800 601.950 135.900 604.050 ;
        RECT 128.400 599.400 129.600 601.650 ;
        RECT 128.400 595.050 129.450 599.400 ;
        RECT 127.950 592.950 130.050 595.050 ;
        RECT 121.950 589.950 124.050 592.050 ;
        RECT 106.950 586.950 109.050 589.050 ;
        RECT 107.400 583.050 108.450 586.950 ;
        RECT 137.400 586.050 138.450 605.400 ;
        RECT 140.400 598.050 141.450 634.950 ;
        RECT 142.950 619.950 145.050 622.050 ;
        RECT 143.400 607.050 144.450 619.950 ;
        RECT 145.950 610.950 148.050 613.050 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 146.400 606.600 147.450 610.950 ;
        RECT 146.400 604.350 147.600 606.600 ;
        RECT 152.400 606.450 153.450 664.950 ;
        RECT 155.400 658.050 156.450 682.950 ;
        RECT 164.400 682.350 165.600 682.950 ;
        RECT 182.400 682.350 183.600 683.100 ;
        RECT 188.400 682.350 189.600 684.000 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 679.950 169.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 167.400 678.900 168.600 679.650 ;
        RECT 179.400 678.900 180.600 679.650 ;
        RECT 166.950 676.800 169.050 678.900 ;
        RECT 178.950 676.800 181.050 678.900 ;
        RECT 185.400 677.400 186.600 679.650 ;
        RECT 185.400 661.050 186.450 677.400 ;
        RECT 194.400 676.050 195.450 685.950 ;
        RECT 203.400 685.200 204.450 691.950 ;
        RECT 196.950 683.100 199.050 685.200 ;
        RECT 202.950 683.100 205.050 685.200 ;
        RECT 209.400 684.600 210.450 718.650 ;
        RECT 215.400 715.050 216.450 722.400 ;
        RECT 220.950 721.800 223.050 723.900 ;
        RECT 224.400 721.050 225.450 733.950 ;
        RECT 232.950 728.100 235.050 730.200 ;
        RECT 238.950 728.100 241.050 730.200 ;
        RECT 242.400 730.050 243.450 749.400 ;
        RECT 248.400 736.050 249.450 793.800 ;
        RECT 260.400 787.050 261.450 800.400 ;
        RECT 266.400 787.050 267.450 800.400 ;
        RECT 281.400 799.050 282.450 800.400 ;
        RECT 286.950 799.800 289.050 801.900 ;
        RECT 292.950 799.950 295.050 802.050 ;
        RECT 268.950 796.950 274.050 799.050 ;
        RECT 280.950 796.950 283.050 799.050 ;
        RECT 283.950 796.950 286.050 799.050 ;
        RECT 281.400 793.050 282.450 796.950 ;
        RECT 280.950 790.950 283.050 793.050 ;
        RECT 259.950 784.950 262.050 787.050 ;
        RECT 265.950 784.950 268.050 787.050 ;
        RECT 250.800 781.950 252.900 784.050 ;
        RECT 253.950 781.950 256.050 784.050 ;
        RECT 251.400 763.050 252.450 781.950 ;
        RECT 254.400 772.050 255.450 781.950 ;
        RECT 253.950 769.950 256.050 772.050 ;
        RECT 262.950 766.950 265.050 769.050 ;
        RECT 250.950 760.950 253.050 763.050 ;
        RECT 256.950 761.100 259.050 766.050 ;
        RECT 263.400 762.600 264.450 766.950 ;
        RECT 257.400 760.350 258.600 761.100 ;
        RECT 263.400 760.350 264.600 762.600 ;
        RECT 271.950 761.100 274.050 766.050 ;
        RECT 284.400 763.200 285.450 796.950 ;
        RECT 293.400 790.050 294.450 799.950 ;
        RECT 292.950 787.950 295.050 790.050 ;
        RECT 292.950 781.950 295.050 784.050 ;
        RECT 277.950 761.100 280.050 763.200 ;
        RECT 283.950 761.100 286.050 763.200 ;
        RECT 278.400 760.350 279.600 761.100 ;
        RECT 284.400 760.350 285.600 761.100 ;
        RECT 289.950 760.950 292.050 763.050 ;
        RECT 253.950 757.950 256.050 760.050 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 283.950 757.950 286.050 760.050 ;
        RECT 254.400 756.900 255.600 757.650 ;
        RECT 253.950 754.800 256.050 756.900 ;
        RECT 260.400 755.400 261.600 757.650 ;
        RECT 260.400 751.050 261.450 755.400 ;
        RECT 271.950 754.950 274.050 757.050 ;
        RECT 275.400 756.900 276.600 757.650 ;
        RECT 256.950 749.400 261.450 751.050 ;
        RECT 256.950 748.950 261.000 749.400 ;
        RECT 259.950 745.950 262.050 748.050 ;
        RECT 247.950 733.950 250.050 736.050 ;
        RECT 233.400 727.350 234.600 728.100 ;
        RECT 239.400 727.350 240.600 728.100 ;
        RECT 241.950 727.950 244.050 730.050 ;
        RECT 244.950 727.950 247.050 730.050 ;
        RECT 253.950 729.000 256.050 733.050 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 230.400 723.000 231.600 724.650 ;
        RECT 236.400 723.900 237.600 724.650 ;
        RECT 223.950 718.950 226.050 721.050 ;
        RECT 229.950 718.950 232.050 723.000 ;
        RECT 235.950 721.800 238.050 723.900 ;
        RECT 241.950 718.950 244.050 724.050 ;
        RECT 245.400 715.050 246.450 727.950 ;
        RECT 254.400 727.350 255.600 729.000 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 251.400 723.900 252.600 724.650 ;
        RECT 250.950 721.800 253.050 723.900 ;
        RECT 214.950 712.950 217.050 715.050 ;
        RECT 244.950 712.950 247.050 715.050 ;
        RECT 211.950 703.950 214.050 706.050 ;
        RECT 212.400 688.050 213.450 703.950 ;
        RECT 227.400 696.300 230.400 698.400 ;
        RECT 231.300 696.300 233.400 698.400 ;
        RECT 250.200 696.300 252.300 698.400 ;
        RECT 211.800 685.950 213.900 688.050 ;
        RECT 214.950 686.100 217.050 688.200 ;
        RECT 215.400 685.350 216.600 686.100 ;
        RECT 193.950 673.950 196.050 676.050 ;
        RECT 178.950 658.950 181.050 661.050 ;
        RECT 184.950 658.950 187.050 661.050 ;
        RECT 154.950 655.950 157.050 658.050 ;
        RECT 163.950 655.950 166.050 658.050 ;
        RECT 157.950 650.100 160.050 652.200 ;
        RECT 164.400 651.600 165.450 655.950 ;
        RECT 179.400 651.600 180.450 658.950 ;
        RECT 158.400 649.350 159.600 650.100 ;
        RECT 164.400 649.350 165.600 651.600 ;
        RECT 179.400 649.350 180.600 651.600 ;
        RECT 184.950 650.100 187.050 652.200 ;
        RECT 185.400 649.350 186.600 650.100 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 160.950 646.950 163.050 649.050 ;
        RECT 163.950 646.950 166.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 187.950 646.950 190.050 649.050 ;
        RECT 161.400 645.900 162.600 646.650 ;
        RECT 160.950 643.800 163.050 645.900 ;
        RECT 172.950 643.950 175.050 646.050 ;
        RECT 176.400 644.400 177.600 646.650 ;
        RECT 182.400 644.400 183.600 646.650 ;
        RECT 188.400 645.000 189.600 646.650 ;
        RECT 173.400 624.450 174.450 643.950 ;
        RECT 176.400 628.050 177.450 644.400 ;
        RECT 182.400 631.050 183.450 644.400 ;
        RECT 187.950 640.950 190.050 645.000 ;
        RECT 197.400 634.050 198.450 683.100 ;
        RECT 203.400 682.350 204.600 683.100 ;
        RECT 209.400 682.350 210.600 684.600 ;
        RECT 214.800 682.950 216.900 685.050 ;
        RECT 220.800 682.950 222.900 685.050 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 199.950 676.800 202.050 678.900 ;
        RECT 206.400 678.000 207.600 679.650 ;
        RECT 200.400 652.200 201.450 676.800 ;
        RECT 205.950 673.950 208.050 678.000 ;
        RECT 211.950 676.950 214.050 679.050 ;
        RECT 208.950 655.950 211.050 658.050 ;
        RECT 199.950 650.100 202.050 652.200 ;
        RECT 200.400 649.350 201.600 650.100 ;
        RECT 200.400 646.950 202.500 649.050 ;
        RECT 205.500 646.950 207.600 649.050 ;
        RECT 199.950 637.950 202.050 643.050 ;
        RECT 209.400 640.050 210.450 655.950 ;
        RECT 212.400 652.200 213.450 676.950 ;
        RECT 218.400 664.050 219.450 679.950 ;
        RECT 227.400 677.400 228.900 696.300 ;
        RECT 231.300 690.300 232.500 696.300 ;
        RECT 230.400 688.200 232.500 690.300 ;
        RECT 227.400 675.300 229.500 677.400 ;
        RECT 223.950 670.950 226.050 673.050 ;
        RECT 228.300 671.700 229.500 675.300 ;
        RECT 231.300 671.700 232.500 688.200 ;
        RECT 233.700 693.300 235.800 695.400 ;
        RECT 233.700 671.700 234.900 693.300 ;
        RECT 238.950 691.950 241.050 694.050 ;
        RECT 239.400 685.200 240.450 691.950 ;
        RECT 242.400 691.800 244.500 693.900 ;
        RECT 247.800 693.300 249.900 695.400 ;
        RECT 242.400 685.200 243.300 691.800 ;
        RECT 248.100 686.100 249.300 693.300 ;
        RECT 250.800 691.500 252.300 696.300 ;
        RECT 253.200 693.300 255.300 698.400 ;
        RECT 250.800 689.400 252.900 691.500 ;
        RECT 238.950 683.100 241.050 685.200 ;
        RECT 242.400 683.100 244.500 685.200 ;
        RECT 247.800 684.000 249.900 686.100 ;
        RECT 238.950 679.950 241.050 682.050 ;
        RECT 239.400 679.350 240.600 679.950 ;
        RECT 238.800 676.950 240.900 679.050 ;
        RECT 242.400 672.600 243.300 683.100 ;
        RECT 245.100 676.500 247.200 678.600 ;
        RECT 217.950 661.950 220.050 664.050 ;
        RECT 214.950 658.950 217.050 661.050 ;
        RECT 211.950 650.100 214.050 652.200 ;
        RECT 208.950 637.950 211.050 640.050 ;
        RECT 196.950 631.950 199.050 634.050 ;
        RECT 181.950 628.950 184.050 631.050 ;
        RECT 175.950 625.950 178.050 628.050 ;
        RECT 173.400 623.400 177.450 624.450 ;
        RECT 163.950 613.950 166.050 616.050 ;
        RECT 172.950 613.950 175.050 616.050 ;
        RECT 164.400 606.600 165.450 613.950 ;
        RECT 173.400 610.050 174.450 613.950 ;
        RECT 172.950 607.950 175.050 610.050 ;
        RECT 152.400 605.400 156.450 606.450 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 148.950 601.950 151.050 604.050 ;
        RECT 142.950 598.950 145.050 601.050 ;
        RECT 149.400 600.450 150.600 601.650 ;
        RECT 149.400 600.000 153.450 600.450 ;
        RECT 149.400 599.400 154.050 600.000 ;
        RECT 139.950 595.950 142.050 598.050 ;
        RECT 143.400 586.050 144.450 598.950 ;
        RECT 145.950 595.950 148.050 598.050 ;
        RECT 151.950 595.950 154.050 599.400 ;
        RECT 124.950 583.950 127.050 586.050 ;
        RECT 136.950 583.950 139.050 586.050 ;
        RECT 142.950 583.950 145.050 586.050 ;
        RECT 106.950 580.950 109.050 583.050 ;
        RECT 121.950 580.950 124.050 583.050 ;
        RECT 103.950 574.950 106.050 577.050 ;
        RECT 122.400 576.450 123.450 580.950 ;
        RECT 125.400 580.050 126.450 583.950 ;
        RECT 124.950 577.950 127.050 580.050 ;
        RECT 127.950 577.950 130.050 580.050 ;
        RECT 142.950 577.950 145.050 580.050 ;
        RECT 122.400 575.400 126.450 576.450 ;
        RECT 91.950 571.950 94.050 574.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 95.400 567.900 96.600 568.650 ;
        RECT 94.950 565.800 97.050 567.900 ;
        RECT 88.950 562.950 91.050 565.050 ;
        RECT 100.950 562.950 103.050 568.050 ;
        RECT 94.950 559.950 97.050 562.050 ;
        RECT 86.400 557.400 91.050 559.050 ;
        RECT 87.000 556.950 91.050 557.400 ;
        RECT 88.950 550.950 91.050 553.050 ;
        RECT 89.400 541.050 90.450 550.950 ;
        RECT 91.950 544.950 94.050 547.050 ;
        RECT 88.950 538.950 91.050 541.050 ;
        RECT 82.950 535.950 85.050 538.050 ;
        RECT 79.950 527.100 82.050 529.200 ;
        RECT 85.950 527.100 88.050 529.200 ;
        RECT 92.400 529.050 93.450 544.950 ;
        RECT 80.400 526.350 81.600 527.100 ;
        RECT 86.400 526.350 87.600 527.100 ;
        RECT 91.950 526.950 94.050 529.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 85.950 523.950 88.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 64.950 520.950 67.050 523.050 ;
        RECT 70.950 520.950 73.050 523.050 ;
        RECT 83.400 522.900 84.600 523.650 ;
        RECT 89.400 522.900 90.600 523.650 ;
        RECT 61.950 514.950 64.050 517.050 ;
        RECT 65.400 511.050 66.450 520.950 ;
        RECT 82.950 520.800 85.050 522.900 ;
        RECT 88.950 520.800 91.050 522.900 ;
        RECT 95.400 522.450 96.450 559.950 ;
        RECT 97.950 553.950 100.050 556.050 ;
        RECT 98.400 544.050 99.450 553.950 ;
        RECT 100.950 550.950 103.050 553.050 ;
        RECT 97.950 541.950 100.050 544.050 ;
        RECT 101.400 532.050 102.450 550.950 ;
        RECT 104.400 532.050 105.450 574.950 ;
        RECT 106.950 573.600 111.000 574.050 ;
        RECT 106.950 571.950 111.600 573.600 ;
        RECT 115.950 572.100 118.050 574.200 ;
        RECT 110.400 571.350 111.600 571.950 ;
        RECT 116.400 571.350 117.600 572.100 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 113.400 567.900 114.600 568.650 ;
        RECT 112.950 565.800 115.050 567.900 ;
        RECT 119.400 567.450 120.600 568.650 ;
        RECT 119.400 566.400 123.450 567.450 ;
        RECT 113.400 562.050 114.450 565.800 ;
        RECT 112.950 559.950 115.050 562.050 ;
        RECT 112.950 556.800 115.050 558.900 ;
        RECT 118.950 556.950 121.050 559.050 ;
        RECT 106.950 547.950 109.050 550.050 ;
        RECT 107.400 538.050 108.450 547.950 ;
        RECT 113.400 547.050 114.450 556.800 ;
        RECT 112.950 544.950 115.050 547.050 ;
        RECT 119.400 540.450 120.450 556.950 ;
        RECT 122.400 555.450 123.450 566.400 ;
        RECT 125.400 559.050 126.450 575.400 ;
        RECT 128.400 574.050 129.450 577.950 ;
        RECT 127.950 571.950 130.050 574.050 ;
        RECT 133.950 572.100 136.050 574.200 ;
        RECT 139.950 572.100 142.050 574.200 ;
        RECT 143.400 574.050 144.450 577.950 ;
        RECT 134.400 571.350 135.600 572.100 ;
        RECT 140.400 571.350 141.600 572.100 ;
        RECT 142.950 571.950 145.050 574.050 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 131.400 566.400 132.600 568.650 ;
        RECT 137.400 567.900 138.600 568.650 ;
        RECT 128.400 562.050 129.450 565.950 ;
        RECT 127.950 559.950 130.050 562.050 ;
        RECT 124.950 556.950 127.050 559.050 ;
        RECT 122.400 554.400 126.450 555.450 ;
        RECT 119.400 539.400 123.450 540.450 ;
        RECT 106.950 535.950 109.050 538.050 ;
        RECT 118.950 535.950 121.050 538.050 ;
        RECT 100.950 529.950 103.050 532.050 ;
        RECT 103.950 529.950 106.050 532.050 ;
        RECT 97.950 528.450 100.050 529.050 ;
        RECT 104.400 528.450 105.600 528.600 ;
        RECT 97.950 527.400 105.600 528.450 ;
        RECT 97.950 526.950 100.050 527.400 ;
        RECT 92.400 521.400 96.450 522.450 ;
        RECT 70.950 514.950 73.050 517.050 ;
        RECT 58.950 508.950 61.050 511.050 ;
        RECT 64.950 508.950 67.050 511.050 ;
        RECT 49.950 505.950 52.050 508.050 ;
        RECT 38.700 501.300 40.800 503.400 ;
        RECT 41.700 501.300 43.800 503.400 ;
        RECT 44.700 501.300 46.800 503.400 ;
        RECT 39.300 497.700 40.500 501.300 ;
        RECT 38.400 495.600 40.500 497.700 ;
        RECT 14.100 490.950 16.200 493.050 ;
        RECT 19.500 490.950 21.600 493.050 ;
        RECT 28.950 490.950 31.050 493.050 ;
        RECT 32.400 492.450 33.600 492.600 ;
        RECT 32.400 491.400 36.450 492.450 ;
        RECT 14.400 489.000 15.600 490.650 ;
        RECT 32.400 490.350 33.600 491.400 ;
        RECT 13.950 484.950 16.050 489.000 ;
        RECT 25.800 487.950 27.900 490.050 ;
        RECT 31.800 487.950 33.900 490.050 ;
        RECT 35.400 487.050 36.450 491.400 ;
        RECT 34.950 484.950 37.050 487.050 ;
        RECT 38.400 476.700 39.900 495.600 ;
        RECT 42.300 484.800 43.500 501.300 ;
        RECT 41.400 482.700 43.500 484.800 ;
        RECT 42.300 476.700 43.500 482.700 ;
        RECT 44.700 479.700 45.900 501.300 ;
        RECT 52.800 500.400 54.900 502.500 ;
        RECT 58.200 501.300 60.300 503.400 ;
        RECT 61.200 501.300 63.300 503.400 ;
        RECT 64.200 501.300 66.300 503.400 ;
        RECT 49.800 493.950 51.900 496.050 ;
        RECT 46.800 490.950 48.900 493.050 ;
        RECT 50.400 492.900 51.600 493.650 ;
        RECT 47.400 483.450 48.450 490.950 ;
        RECT 49.950 490.800 52.050 492.900 ;
        RECT 53.400 489.900 54.300 500.400 ;
        RECT 56.100 494.400 58.200 496.500 ;
        RECT 53.400 487.800 55.500 489.900 ;
        RECT 59.100 489.000 60.300 501.300 ;
        RECT 47.400 482.400 51.450 483.450 ;
        RECT 44.700 477.600 46.800 479.700 ;
        RECT 38.400 474.600 41.400 476.700 ;
        RECT 42.300 474.600 44.400 476.700 ;
        RECT 50.400 469.050 51.450 482.400 ;
        RECT 53.400 481.200 54.300 487.800 ;
        RECT 58.800 486.900 60.900 489.000 ;
        RECT 53.400 479.100 55.500 481.200 ;
        RECT 59.100 479.700 60.300 486.900 ;
        RECT 61.800 483.600 63.300 501.300 ;
        RECT 61.800 481.500 63.900 483.600 ;
        RECT 58.800 477.600 60.900 479.700 ;
        RECT 61.800 476.700 63.300 481.500 ;
        RECT 65.100 479.700 66.300 501.300 ;
        RECT 61.200 474.600 63.300 476.700 ;
        RECT 64.200 474.600 66.300 479.700 ;
        RECT 67.200 501.300 69.300 503.400 ;
        RECT 67.200 483.600 68.700 501.300 ;
        RECT 71.400 496.050 72.450 514.950 ;
        RECT 89.400 511.050 90.450 520.800 ;
        RECT 76.950 508.950 79.050 511.050 ;
        RECT 88.950 508.950 91.050 511.050 ;
        RECT 70.950 493.950 73.050 496.050 ;
        RECT 77.400 492.600 78.450 508.950 ;
        RECT 89.400 496.200 90.450 508.950 ;
        RECT 88.950 494.100 91.050 496.200 ;
        RECT 77.400 492.450 78.600 492.600 ;
        RECT 86.400 492.450 87.600 492.600 ;
        RECT 89.400 492.450 90.450 494.100 ;
        RECT 77.400 491.400 81.450 492.450 ;
        RECT 77.400 490.350 78.600 491.400 ;
        RECT 76.800 487.950 78.900 490.050 ;
        RECT 67.200 481.500 69.300 483.600 ;
        RECT 67.200 476.700 68.700 481.500 ;
        RECT 80.400 478.050 81.450 491.400 ;
        RECT 86.400 491.400 90.450 492.450 ;
        RECT 86.400 490.350 87.600 491.400 ;
        RECT 85.800 487.950 87.900 490.050 ;
        RECT 82.950 484.950 85.050 487.050 ;
        RECT 67.200 474.600 69.300 476.700 ;
        RECT 73.950 475.950 76.050 478.050 ;
        RECT 79.950 475.950 82.050 478.050 ;
        RECT 74.400 469.050 75.450 475.950 ;
        RECT 37.950 466.950 40.050 469.050 ;
        RECT 49.950 466.950 52.050 469.050 ;
        RECT 73.950 466.950 76.050 469.050 ;
        RECT 10.950 457.950 13.050 460.050 ;
        RECT 28.950 457.950 31.050 460.050 ;
        RECT 5.400 452.400 9.450 453.450 ;
        RECT 4.950 449.100 7.050 451.200 ;
        RECT 5.400 436.050 6.450 449.100 ;
        RECT 4.950 433.950 7.050 436.050 ;
        RECT 8.400 427.050 9.450 452.400 ;
        RECT 13.950 449.100 16.050 451.200 ;
        RECT 14.400 448.350 15.600 449.100 ;
        RECT 23.100 448.950 25.200 451.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 23.400 447.000 24.600 448.650 ;
        RECT 17.400 444.900 18.600 445.650 ;
        RECT 16.950 442.800 19.050 444.900 ;
        RECT 22.950 442.800 25.050 447.000 ;
        RECT 7.950 424.950 10.050 427.050 ;
        RECT 7.950 418.950 10.050 421.050 ;
        RECT 1.950 416.100 4.050 418.200 ;
        RECT 8.400 295.050 9.450 418.950 ;
        RECT 17.400 417.600 18.450 442.800 ;
        RECT 17.400 415.350 18.600 417.600 ;
        RECT 11.100 412.950 13.200 415.050 ;
        RECT 16.500 412.950 18.600 415.050 ;
        RECT 29.400 391.050 30.450 457.950 ;
        RECT 32.100 448.950 34.200 451.050 ;
        RECT 32.400 446.400 33.600 448.650 ;
        RECT 32.400 433.050 33.450 446.400 ;
        RECT 31.950 430.950 34.050 433.050 ;
        RECT 38.400 421.050 39.450 466.950 ;
        RECT 41.700 462.300 43.800 464.400 ;
        RECT 42.300 457.500 43.800 462.300 ;
        RECT 41.700 455.400 43.800 457.500 ;
        RECT 42.300 437.700 43.800 455.400 ;
        RECT 41.700 435.600 43.800 437.700 ;
        RECT 44.700 459.300 46.800 464.400 ;
        RECT 47.700 462.300 49.800 464.400 ;
        RECT 66.600 462.300 68.700 464.400 ;
        RECT 69.600 462.300 72.600 464.400 ;
        RECT 44.700 437.700 45.900 459.300 ;
        RECT 47.700 457.500 49.200 462.300 ;
        RECT 50.100 459.300 52.200 461.400 ;
        RECT 47.100 455.400 49.200 457.500 ;
        RECT 47.700 437.700 49.200 455.400 ;
        RECT 50.700 452.100 51.900 459.300 ;
        RECT 55.500 457.800 57.600 459.900 ;
        RECT 64.200 459.300 66.300 461.400 ;
        RECT 50.100 450.000 52.200 452.100 ;
        RECT 56.700 451.200 57.600 457.800 ;
        RECT 50.700 437.700 51.900 450.000 ;
        RECT 55.500 449.100 57.600 451.200 ;
        RECT 52.800 442.500 54.900 444.600 ;
        RECT 56.700 438.600 57.600 449.100 ;
        RECT 58.950 446.100 61.050 448.200 ;
        RECT 59.400 445.350 60.600 446.100 ;
        RECT 59.100 442.950 61.200 445.050 ;
        RECT 44.700 435.600 46.800 437.700 ;
        RECT 47.700 435.600 49.800 437.700 ;
        RECT 50.700 435.600 52.800 437.700 ;
        RECT 56.100 436.500 58.200 438.600 ;
        RECT 65.100 437.700 66.300 459.300 ;
        RECT 67.500 456.300 68.700 462.300 ;
        RECT 67.500 454.200 69.600 456.300 ;
        RECT 67.500 437.700 68.700 454.200 ;
        RECT 71.100 443.400 72.600 462.300 ;
        RECT 70.500 441.300 72.600 443.400 ;
        RECT 70.500 437.700 71.700 441.300 ;
        RECT 64.200 435.600 66.300 437.700 ;
        RECT 67.200 435.600 69.300 437.700 ;
        RECT 70.200 435.600 72.300 437.700 ;
        RECT 74.400 433.050 75.450 466.950 ;
        RECT 83.400 453.600 84.450 484.950 ;
        RECT 83.400 451.350 84.600 453.600 ;
        RECT 77.100 448.950 79.200 451.050 ;
        RECT 83.100 448.950 85.200 451.050 ;
        RECT 43.950 430.950 46.050 433.050 ;
        RECT 73.950 430.950 76.050 433.050 ;
        RECT 37.950 418.950 40.050 421.050 ;
        RECT 38.400 417.450 39.600 417.600 ;
        RECT 38.400 416.400 42.450 417.450 ;
        RECT 38.400 415.350 39.600 416.400 ;
        RECT 32.100 412.950 34.200 415.050 ;
        RECT 37.500 412.950 39.600 415.050 ;
        RECT 41.400 397.050 42.450 416.400 ;
        RECT 40.950 394.950 43.050 397.050 ;
        RECT 28.950 388.950 31.050 391.050 ;
        RECT 40.950 385.950 43.050 388.050 ;
        RECT 34.950 372.000 37.050 376.050 ;
        RECT 35.400 370.350 36.600 372.000 ;
        RECT 16.800 367.950 18.900 370.050 ;
        RECT 34.800 367.950 36.900 370.050 ;
        RECT 22.950 361.950 25.050 364.050 ;
        RECT 16.800 334.950 18.900 337.050 ;
        RECT 19.950 298.950 22.050 301.050 ;
        RECT 7.950 292.950 10.050 295.050 ;
        RECT 13.950 293.100 16.050 295.200 ;
        RECT 14.400 292.350 15.600 293.100 ;
        RECT 10.950 289.950 13.050 292.050 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 7.950 286.950 10.050 289.050 ;
        RECT 11.400 287.400 12.600 289.650 ;
        RECT 4.950 264.450 7.050 265.050 ;
        RECT 2.400 263.400 7.050 264.450 ;
        RECT 2.400 106.200 3.450 263.400 ;
        RECT 4.950 262.950 7.050 263.400 ;
        RECT 5.400 258.600 6.450 262.950 ;
        RECT 5.400 256.350 6.600 258.600 ;
        RECT 8.400 258.450 9.450 286.950 ;
        RECT 11.400 265.050 12.450 287.400 ;
        RECT 13.950 271.950 16.050 274.050 ;
        RECT 10.950 262.950 13.050 265.050 ;
        RECT 14.400 258.600 15.450 271.950 ;
        RECT 20.400 258.900 21.450 298.950 ;
        RECT 23.400 288.900 24.450 361.950 ;
        RECT 28.950 352.950 31.050 355.050 ;
        RECT 29.400 298.050 30.450 352.950 ;
        RECT 37.950 337.950 40.050 340.050 ;
        RECT 34.800 334.950 36.900 337.050 ;
        RECT 35.400 333.450 36.600 334.650 ;
        RECT 38.400 333.450 39.450 337.950 ;
        RECT 35.400 332.400 39.450 333.450 ;
        RECT 38.400 304.050 39.450 332.400 ;
        RECT 41.400 325.050 42.450 385.950 ;
        RECT 44.400 376.050 45.450 430.950 ;
        RECT 70.950 424.950 73.050 427.050 ;
        RECT 88.950 424.950 91.050 427.050 ;
        RECT 52.950 416.100 55.050 418.200 ;
        RECT 58.950 416.100 61.050 418.200 ;
        RECT 71.400 417.600 72.450 424.950 ;
        RECT 79.950 421.950 82.050 424.050 ;
        RECT 53.400 415.350 54.600 416.100 ;
        RECT 59.400 415.350 60.600 416.100 ;
        RECT 71.400 415.350 72.600 417.600 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 55.950 412.950 58.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 71.400 412.950 73.500 415.050 ;
        RECT 76.800 412.950 78.900 415.050 ;
        RECT 50.400 410.400 51.600 412.650 ;
        RECT 56.400 410.400 57.600 412.650 ;
        RECT 50.400 403.050 51.450 410.400 ;
        RECT 49.950 400.950 52.050 403.050 ;
        RECT 56.400 388.050 57.450 410.400 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 77.400 410.400 78.600 412.650 ;
        RECT 55.950 385.950 58.050 388.050 ;
        RECT 43.950 373.950 46.050 376.050 ;
        RECT 62.400 375.450 63.450 409.950 ;
        RECT 77.400 406.050 78.450 410.400 ;
        RECT 76.950 403.950 79.050 406.050 ;
        RECT 80.400 403.050 81.450 421.950 ;
        RECT 89.400 417.600 90.450 424.950 ;
        RECT 92.400 424.050 93.450 521.400 ;
        RECT 94.950 517.950 97.050 520.050 ;
        RECT 95.400 505.050 96.450 517.950 ;
        RECT 98.400 517.050 99.450 526.950 ;
        RECT 104.400 526.350 105.600 527.400 ;
        RECT 109.950 527.100 112.050 529.200 ;
        RECT 110.400 526.350 111.600 527.100 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 107.400 521.400 108.600 523.650 ;
        RECT 113.400 521.400 114.600 523.650 ;
        RECT 97.950 514.950 100.050 517.050 ;
        RECT 101.400 513.450 102.450 520.950 ;
        RECT 98.400 512.400 102.450 513.450 ;
        RECT 94.950 502.950 97.050 505.050 ;
        RECT 98.400 481.050 99.450 512.400 ;
        RECT 107.400 505.050 108.450 521.400 ;
        RECT 109.950 514.950 112.050 517.050 ;
        RECT 106.950 502.950 109.050 505.050 ;
        RECT 103.950 494.100 106.050 496.200 ;
        RECT 110.400 495.600 111.450 514.950 ;
        RECT 113.400 499.050 114.450 521.400 ;
        RECT 115.950 520.950 118.050 523.050 ;
        RECT 112.950 496.950 115.050 499.050 ;
        RECT 116.400 496.050 117.450 520.950 ;
        RECT 119.400 520.050 120.450 535.950 ;
        RECT 122.400 523.050 123.450 539.400 ;
        RECT 125.400 529.050 126.450 554.400 ;
        RECT 131.400 547.050 132.450 566.400 ;
        RECT 136.950 565.800 139.050 567.900 ;
        RECT 142.950 565.800 145.050 567.900 ;
        RECT 139.950 559.950 142.050 562.050 ;
        RECT 136.950 553.950 139.050 556.050 ;
        RECT 130.950 544.950 133.050 547.050 ;
        RECT 137.400 544.050 138.450 553.950 ;
        RECT 136.950 541.950 139.050 544.050 ;
        RECT 127.950 538.950 130.050 541.050 ;
        RECT 128.400 535.050 129.450 538.950 ;
        RECT 127.950 532.950 130.050 535.050 ;
        RECT 124.950 526.950 127.050 529.050 ;
        RECT 127.950 528.000 130.050 531.900 ;
        RECT 128.400 526.350 129.600 528.000 ;
        RECT 133.950 527.100 136.050 529.200 ;
        RECT 140.400 529.050 141.450 559.950 ;
        RECT 143.400 550.050 144.450 565.800 ;
        RECT 142.950 547.950 145.050 550.050 ;
        RECT 146.400 538.050 147.450 595.950 ;
        RECT 148.950 594.900 153.000 595.050 ;
        RECT 148.950 592.950 154.050 594.900 ;
        RECT 151.950 592.800 154.050 592.950 ;
        RECT 155.400 583.050 156.450 605.400 ;
        RECT 164.400 604.350 165.600 606.600 ;
        RECT 169.950 605.100 172.050 607.200 ;
        RECT 176.400 607.050 177.450 623.400 ;
        RECT 178.950 616.950 181.050 619.050 ;
        RECT 202.950 616.950 205.050 619.050 ;
        RECT 170.400 604.350 171.600 605.100 ;
        RECT 175.950 604.950 178.050 607.050 ;
        RECT 160.950 601.950 163.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 161.400 600.000 162.600 601.650 ;
        RECT 160.950 595.950 163.050 600.000 ;
        RECT 167.400 599.400 168.600 601.650 ;
        RECT 173.400 600.900 174.600 601.650 ;
        RECT 179.400 601.050 180.450 616.950 ;
        RECT 187.950 610.950 190.050 613.050 ;
        RECT 181.950 607.950 184.050 610.050 ;
        RECT 167.400 597.450 168.450 599.400 ;
        RECT 172.950 598.800 175.050 600.900 ;
        RECT 178.800 598.950 180.900 601.050 ;
        RECT 182.400 600.900 183.450 607.950 ;
        RECT 184.950 604.950 187.050 610.050 ;
        RECT 188.400 606.600 189.450 610.950 ;
        RECT 188.400 604.350 189.600 606.600 ;
        RECT 193.950 605.100 196.050 607.200 ;
        RECT 199.950 605.100 202.050 607.200 ;
        RECT 203.400 607.050 204.450 616.950 ;
        RECT 215.400 613.050 216.450 658.950 ;
        RECT 224.400 655.050 225.450 670.950 ;
        RECT 227.700 669.600 229.800 671.700 ;
        RECT 230.700 669.600 232.800 671.700 ;
        RECT 233.700 669.600 235.800 671.700 ;
        RECT 241.800 670.500 243.900 672.600 ;
        RECT 248.100 671.700 249.300 684.000 ;
        RECT 250.800 671.700 252.300 689.400 ;
        RECT 254.100 671.700 255.300 693.300 ;
        RECT 247.200 669.600 249.300 671.700 ;
        RECT 250.200 669.600 252.300 671.700 ;
        RECT 253.200 669.600 255.300 671.700 ;
        RECT 256.200 696.300 258.300 698.400 ;
        RECT 256.200 691.500 257.700 696.300 ;
        RECT 256.200 689.400 258.300 691.500 ;
        RECT 256.200 671.700 257.700 689.400 ;
        RECT 256.200 669.600 258.300 671.700 ;
        RECT 260.400 667.050 261.450 745.950 ;
        RECT 268.950 742.950 271.050 745.050 ;
        RECT 265.950 739.950 268.050 742.050 ;
        RECT 266.400 733.050 267.450 739.950 ;
        RECT 269.400 736.050 270.450 742.950 ;
        RECT 268.950 733.950 271.050 736.050 ;
        RECT 265.950 730.950 268.050 733.050 ;
        RECT 272.400 729.600 273.450 754.950 ;
        RECT 274.950 754.800 277.050 756.900 ;
        RECT 281.400 755.400 282.600 757.650 ;
        RECT 290.400 757.050 291.450 760.950 ;
        RECT 277.950 751.950 280.050 754.050 ;
        RECT 278.400 730.200 279.450 751.950 ;
        RECT 281.400 733.050 282.450 755.400 ;
        RECT 289.950 754.950 292.050 757.050 ;
        RECT 293.400 756.900 294.450 781.950 ;
        RECT 292.950 754.800 295.050 756.900 ;
        RECT 289.950 751.800 292.050 753.900 ;
        RECT 286.950 745.950 289.050 748.050 ;
        RECT 280.950 730.950 283.050 733.050 ;
        RECT 272.400 727.350 273.600 729.600 ;
        RECT 277.950 728.100 280.050 730.200 ;
        RECT 278.400 727.350 279.600 728.100 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 265.950 721.800 268.050 723.900 ;
        RECT 269.400 723.000 270.600 724.650 ;
        RECT 266.400 706.050 267.450 721.800 ;
        RECT 268.950 718.950 271.050 723.000 ;
        RECT 275.400 722.400 276.600 724.650 ;
        RECT 275.400 718.050 276.450 722.400 ;
        RECT 274.950 715.950 277.050 718.050 ;
        RECT 287.400 717.450 288.450 745.950 ;
        RECT 290.400 723.450 291.450 751.800 ;
        RECT 293.400 748.050 294.450 754.800 ;
        RECT 296.400 748.050 297.450 806.100 ;
        RECT 299.400 796.050 300.450 820.950 ;
        RECT 305.400 817.050 306.450 832.800 ;
        RECT 304.950 814.950 307.050 817.050 ;
        RECT 301.950 805.950 304.050 811.050 ;
        RECT 305.400 807.600 306.450 814.950 ;
        RECT 311.400 807.600 312.450 844.950 ;
        RECT 314.400 841.200 315.450 850.950 ;
        RECT 319.500 843.300 321.600 845.400 ;
        RECT 329.100 844.500 331.200 846.600 ;
        RECT 313.950 840.450 316.050 841.200 ;
        RECT 317.400 840.450 318.600 840.600 ;
        RECT 313.950 839.400 318.600 840.450 ;
        RECT 313.950 839.100 316.050 839.400 ;
        RECT 314.400 811.050 315.450 839.100 ;
        RECT 317.400 838.350 318.600 839.400 ;
        RECT 317.100 835.950 319.200 838.050 ;
        RECT 320.400 834.300 321.300 843.300 ;
        RECT 322.800 839.700 324.900 841.800 ;
        RECT 326.400 841.350 327.600 843.600 ;
        RECT 324.000 837.300 324.900 839.700 ;
        RECT 325.800 838.950 327.900 841.050 ;
        RECT 329.700 837.300 330.900 844.500 ;
        RECT 324.000 836.100 330.900 837.300 ;
        RECT 327.000 834.300 329.100 835.200 ;
        RECT 320.400 833.100 329.100 834.300 ;
        RECT 321.900 831.300 324.000 833.100 ;
        RECT 325.800 830.100 327.900 832.200 ;
        RECT 330.000 830.700 330.900 836.100 ;
        RECT 331.800 835.950 333.900 838.050 ;
        RECT 332.400 834.900 333.600 835.650 ;
        RECT 331.950 832.800 334.050 834.900 ;
        RECT 335.400 832.050 336.450 853.950 ;
        RECT 326.400 827.550 327.600 829.800 ;
        RECT 329.100 828.600 331.200 830.700 ;
        RECT 334.950 829.950 337.050 832.050 ;
        RECT 326.400 814.050 327.450 827.550 ;
        RECT 338.400 826.050 339.450 865.950 ;
        RECT 341.400 838.050 342.450 877.800 ;
        RECT 367.950 874.950 370.050 877.050 ;
        RECT 379.950 874.950 382.050 879.000 ;
        RECT 349.950 871.950 352.050 874.050 ;
        RECT 350.400 847.050 351.450 871.950 ;
        RECT 349.950 844.950 352.050 847.050 ;
        RECT 346.950 840.000 349.050 844.050 ;
        RECT 347.400 838.350 348.600 840.000 ;
        RECT 352.950 839.100 355.050 841.200 ;
        RECT 361.950 839.100 364.050 841.200 ;
        RECT 368.400 840.600 369.450 874.950 ;
        RECT 376.950 856.950 379.050 859.050 ;
        RECT 377.400 849.450 378.450 856.950 ;
        RECT 374.400 848.400 378.450 849.450 ;
        RECT 374.400 840.600 375.450 848.400 ;
        RECT 382.950 844.950 385.050 847.050 ;
        RECT 353.400 838.350 354.600 839.100 ;
        RECT 340.950 835.950 343.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 352.950 835.950 355.050 838.050 ;
        RECT 355.950 835.950 358.050 838.050 ;
        RECT 350.400 834.000 351.600 835.650 ;
        RECT 356.400 834.900 357.600 835.650 ;
        RECT 362.400 835.050 363.450 839.100 ;
        RECT 368.400 838.350 369.600 840.600 ;
        RECT 374.400 838.350 375.600 840.600 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 376.950 835.950 379.050 838.050 ;
        RECT 349.950 829.950 352.050 834.000 ;
        RECT 355.950 832.800 358.050 834.900 ;
        RECT 361.950 832.950 364.050 835.050 ;
        RECT 371.400 834.900 372.600 835.650 ;
        RECT 377.400 834.900 378.600 835.650 ;
        RECT 370.950 832.800 373.050 834.900 ;
        RECT 376.950 832.800 379.050 834.900 ;
        RECT 337.950 823.950 340.050 826.050 ;
        RECT 325.950 811.950 328.050 814.050 ;
        RECT 313.950 808.950 316.050 811.050 ;
        RECT 305.400 805.350 306.600 807.600 ;
        RECT 311.400 805.350 312.600 807.600 ;
        RECT 328.950 806.100 331.050 808.200 ;
        RECT 329.400 805.350 330.600 806.100 ;
        RECT 304.950 802.950 307.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 313.950 802.950 316.050 805.050 ;
        RECT 325.950 802.950 328.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 308.400 801.000 309.600 802.650 ;
        RECT 307.950 796.950 310.050 801.000 ;
        RECT 314.400 800.400 315.600 802.650 ;
        RECT 326.400 801.900 327.600 802.650 ;
        RECT 332.400 801.900 333.600 802.650 ;
        RECT 298.950 793.950 301.050 796.050 ;
        RECT 314.400 793.050 315.450 800.400 ;
        RECT 325.950 799.800 328.050 801.900 ;
        RECT 331.950 799.800 334.050 801.900 ;
        RECT 310.800 790.950 312.900 793.050 ;
        RECT 313.950 790.950 316.050 793.050 ;
        RECT 304.950 787.950 307.050 790.050 ;
        RECT 298.950 772.950 301.050 775.050 ;
        RECT 299.400 766.050 300.450 772.950 ;
        RECT 305.400 766.050 306.450 787.950 ;
        RECT 307.950 778.950 310.050 781.050 ;
        RECT 298.950 763.950 301.050 766.050 ;
        RECT 304.950 763.950 307.050 766.050 ;
        RECT 299.400 762.600 300.450 763.950 ;
        RECT 308.400 762.600 309.450 778.950 ;
        RECT 311.400 766.050 312.450 790.950 ;
        RECT 316.950 787.050 319.050 790.050 ;
        RECT 313.950 786.000 319.050 787.050 ;
        RECT 313.950 785.400 318.450 786.000 ;
        RECT 313.950 784.950 318.000 785.400 ;
        RECT 326.400 781.050 327.450 799.800 ;
        RECT 328.950 793.950 331.050 796.050 ;
        RECT 329.400 781.050 330.450 793.950 ;
        RECT 325.800 778.950 327.900 781.050 ;
        RECT 328.950 778.950 331.050 781.050 ;
        RECT 316.950 777.450 319.050 778.050 ;
        RECT 316.950 777.000 324.450 777.450 ;
        RECT 316.950 776.400 325.050 777.000 ;
        RECT 316.950 775.950 319.050 776.400 ;
        RECT 322.950 772.950 325.050 776.400 ;
        RECT 313.950 766.950 316.050 769.050 ;
        RECT 322.950 766.950 325.050 769.050 ;
        RECT 310.950 763.950 313.050 766.050 ;
        RECT 299.400 760.350 300.600 762.600 ;
        RECT 308.400 760.350 309.600 762.600 ;
        RECT 310.950 760.800 313.050 762.900 ;
        RECT 299.100 757.950 301.200 760.050 ;
        RECT 304.500 757.950 306.600 760.050 ;
        RECT 307.800 757.950 309.900 760.050 ;
        RECT 305.400 756.900 306.600 757.650 ;
        RECT 304.950 754.800 307.050 756.900 ;
        RECT 304.950 748.950 307.050 751.050 ;
        RECT 292.950 745.950 295.050 748.050 ;
        RECT 295.950 745.950 298.050 748.050 ;
        RECT 305.400 730.200 306.450 748.950 ;
        RECT 311.400 742.050 312.450 760.800 ;
        RECT 314.400 757.050 315.450 766.950 ;
        RECT 323.400 762.600 324.450 766.950 ;
        RECT 323.400 760.350 324.600 762.600 ;
        RECT 328.950 761.100 331.050 763.200 ;
        RECT 334.950 761.100 337.050 763.200 ;
        RECT 329.400 760.350 330.600 761.100 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 325.950 757.950 328.050 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 313.950 754.950 316.050 757.050 ;
        RECT 316.950 754.950 319.050 757.050 ;
        RECT 320.400 755.400 321.600 757.650 ;
        RECT 326.400 756.900 327.600 757.650 ;
        RECT 310.800 739.950 312.900 742.050 ;
        RECT 313.950 739.950 316.050 742.050 ;
        RECT 298.950 728.100 301.050 730.200 ;
        RECT 304.950 728.100 307.050 730.200 ;
        RECT 314.400 729.600 315.450 739.950 ;
        RECT 317.400 733.050 318.450 754.950 ;
        RECT 316.950 730.950 319.050 733.050 ;
        RECT 320.400 729.600 321.450 755.400 ;
        RECT 325.950 754.800 328.050 756.900 ;
        RECT 331.950 751.950 334.050 757.050 ;
        RECT 328.950 739.950 331.050 742.050 ;
        RECT 299.400 727.350 300.600 728.100 ;
        RECT 293.100 724.950 295.200 727.050 ;
        RECT 298.500 724.950 300.600 727.050 ;
        RECT 301.800 724.950 303.900 727.050 ;
        RECT 293.400 723.450 294.600 724.650 ;
        RECT 290.400 722.400 294.600 723.450 ;
        RECT 302.400 722.400 303.600 724.650 ;
        RECT 284.400 716.400 288.450 717.450 ;
        RECT 277.950 712.950 280.050 715.050 ;
        RECT 268.950 706.950 271.050 709.050 ;
        RECT 265.950 703.950 268.050 706.050 ;
        RECT 269.400 703.050 270.450 706.950 ;
        RECT 268.950 700.950 271.050 703.050 ;
        RECT 268.950 694.950 271.050 697.050 ;
        RECT 265.800 682.950 267.900 685.050 ;
        RECT 262.950 679.950 265.050 682.050 ;
        RECT 266.400 680.400 267.600 682.650 ;
        RECT 244.950 664.950 247.050 667.050 ;
        RECT 253.950 664.950 256.050 667.050 ;
        RECT 259.950 664.950 262.050 667.050 ;
        RECT 232.800 661.950 234.900 664.050 ;
        RECT 235.950 661.950 238.050 664.050 ;
        RECT 223.950 652.950 226.050 655.050 ;
        RECT 229.950 652.950 232.050 655.050 ;
        RECT 220.950 646.950 223.050 649.050 ;
        RECT 223.950 646.950 226.050 649.050 ;
        RECT 224.400 645.450 225.600 646.650 ;
        RECT 224.400 644.400 228.450 645.450 ;
        RECT 217.950 625.950 220.050 628.050 ;
        RECT 223.950 625.950 226.050 628.050 ;
        RECT 205.950 610.950 208.050 613.050 ;
        RECT 214.950 610.950 217.050 613.050 ;
        RECT 194.400 604.350 195.600 605.100 ;
        RECT 200.400 604.350 201.600 605.100 ;
        RECT 202.950 604.950 205.050 607.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 181.950 598.800 184.050 600.900 ;
        RECT 184.950 598.950 187.050 601.050 ;
        RECT 191.400 600.900 192.600 601.650 ;
        RECT 164.400 596.400 168.450 597.450 ;
        RECT 157.950 594.450 160.050 595.050 ;
        RECT 164.400 594.450 165.450 596.400 ;
        RECT 178.950 595.800 181.050 597.900 ;
        RECT 157.950 593.400 165.450 594.450 ;
        RECT 157.950 592.950 160.050 593.400 ;
        RECT 166.950 592.950 169.050 595.050 ;
        RECT 163.950 589.950 166.050 592.050 ;
        RECT 155.400 581.400 160.050 583.050 ;
        RECT 156.000 580.950 160.050 581.400 ;
        RECT 154.950 579.450 157.050 580.050 ;
        RECT 149.400 578.400 157.050 579.450 ;
        RECT 149.400 574.050 150.450 578.400 ;
        RECT 154.950 577.950 157.050 578.400 ;
        RECT 148.950 571.950 151.050 574.050 ;
        RECT 151.950 573.000 154.050 577.050 ;
        RECT 152.400 571.350 153.600 573.000 ;
        RECT 157.950 572.100 160.050 574.200 ;
        RECT 164.400 574.050 165.450 589.950 ;
        RECT 158.400 571.350 159.600 572.100 ;
        RECT 163.950 571.950 166.050 574.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 148.950 565.950 151.050 568.050 ;
        RECT 155.400 566.400 156.600 568.650 ;
        RECT 161.400 567.000 162.600 568.650 ;
        RECT 149.400 553.050 150.450 565.950 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 148.950 550.950 151.050 553.050 ;
        RECT 152.400 547.050 153.450 562.950 ;
        RECT 155.400 559.050 156.450 566.400 ;
        RECT 160.950 562.950 163.050 567.000 ;
        RECT 163.950 565.950 166.050 568.050 ;
        RECT 154.950 556.950 157.050 559.050 ;
        RECT 151.950 544.950 154.050 547.050 ;
        RECT 164.400 543.450 165.450 565.950 ;
        RECT 167.400 562.050 168.450 592.950 ;
        RECT 179.400 592.050 180.450 595.800 ;
        RECT 172.950 589.950 175.050 592.050 ;
        RECT 178.950 589.950 181.050 592.050 ;
        RECT 169.950 580.950 172.050 583.050 ;
        RECT 170.400 565.050 171.450 580.950 ;
        RECT 173.400 568.050 174.450 589.950 ;
        RECT 178.950 577.950 181.050 580.050 ;
        RECT 179.400 573.600 180.450 577.950 ;
        RECT 185.400 576.450 186.450 598.950 ;
        RECT 190.950 598.800 193.050 600.900 ;
        RECT 197.400 600.000 198.600 601.650 ;
        RECT 196.950 595.950 199.050 600.000 ;
        RECT 206.400 589.050 207.450 610.950 ;
        RECT 211.950 605.100 214.050 607.200 ;
        RECT 218.400 607.050 219.450 625.950 ;
        RECT 220.950 610.950 223.050 613.050 ;
        RECT 212.400 604.350 213.600 605.100 ;
        RECT 217.950 604.950 220.050 607.050 ;
        RECT 211.950 601.950 214.050 604.050 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 215.400 600.900 216.600 601.650 ;
        RECT 214.950 598.800 217.050 600.900 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 190.950 586.950 193.050 589.050 ;
        RECT 205.950 586.950 208.050 589.050 ;
        RECT 185.400 575.400 189.450 576.450 ;
        RECT 179.400 571.350 180.600 573.600 ;
        RECT 176.100 568.950 178.200 571.050 ;
        RECT 179.400 568.950 181.500 571.050 ;
        RECT 184.800 568.950 186.900 571.050 ;
        RECT 172.950 565.950 175.050 568.050 ;
        RECT 176.400 566.400 177.600 568.650 ;
        RECT 185.400 567.450 186.600 568.650 ;
        RECT 188.400 567.450 189.450 575.400 ;
        RECT 185.400 566.400 189.450 567.450 ;
        RECT 176.400 565.050 177.450 566.400 ;
        RECT 169.950 562.950 172.050 565.050 ;
        RECT 174.000 564.900 177.450 565.050 ;
        RECT 172.950 563.400 177.450 564.900 ;
        RECT 172.950 562.950 177.000 563.400 ;
        RECT 166.950 559.950 169.050 562.050 ;
        RECT 170.400 550.050 171.450 562.950 ;
        RECT 172.950 562.800 175.050 562.950 ;
        RECT 181.950 556.950 184.050 559.050 ;
        RECT 169.950 547.950 172.050 550.050 ;
        RECT 175.950 544.950 178.050 547.050 ;
        RECT 161.400 542.400 165.450 543.450 ;
        RECT 145.950 535.950 148.050 538.050 ;
        RECT 134.400 526.350 135.600 527.100 ;
        RECT 139.950 526.950 142.050 529.050 ;
        RECT 142.950 527.100 145.050 529.200 ;
        RECT 151.950 527.100 154.050 529.200 ;
        RECT 157.950 528.000 160.050 532.050 ;
        RECT 161.400 529.050 162.450 542.400 ;
        RECT 163.950 538.950 166.050 541.050 ;
        RECT 127.950 523.950 130.050 526.050 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 121.950 520.950 124.050 523.050 ;
        RECT 124.950 520.950 127.050 523.050 ;
        RECT 131.400 521.400 132.600 523.650 ;
        RECT 137.400 521.400 138.600 523.650 ;
        RECT 118.950 517.950 121.050 520.050 ;
        RECT 125.400 517.050 126.450 520.950 ;
        RECT 131.400 517.050 132.450 521.400 ;
        RECT 137.400 517.050 138.450 521.400 ;
        RECT 139.950 520.950 142.050 523.050 ;
        RECT 124.950 514.950 127.050 517.050 ;
        RECT 130.950 514.950 133.050 517.050 ;
        RECT 136.950 514.950 139.050 517.050 ;
        RECT 140.400 508.050 141.450 520.950 ;
        RECT 143.400 508.050 144.450 527.100 ;
        RECT 152.400 526.350 153.600 527.100 ;
        RECT 158.400 526.350 159.600 528.000 ;
        RECT 160.950 526.950 163.050 529.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 149.400 522.900 150.600 523.650 ;
        RECT 148.950 520.800 151.050 522.900 ;
        RECT 155.400 522.000 156.600 523.650 ;
        RECT 164.400 523.050 165.450 538.950 ;
        RECT 176.400 529.050 177.450 544.950 ;
        RECT 178.950 529.950 181.050 532.050 ;
        RECT 166.950 528.600 171.000 529.050 ;
        RECT 166.950 526.950 171.600 528.600 ;
        RECT 175.950 526.950 178.050 529.050 ;
        RECT 170.400 526.350 171.600 526.950 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 154.950 514.950 157.050 522.000 ;
        RECT 163.950 520.950 166.050 523.050 ;
        RECT 166.950 520.950 169.050 523.050 ;
        RECT 173.400 522.900 174.600 523.650 ;
        RECT 160.950 517.950 163.050 520.050 ;
        RECT 124.950 505.950 127.050 508.050 ;
        RECT 139.800 505.950 141.900 508.050 ;
        RECT 142.950 505.950 145.050 508.050 ;
        RECT 125.400 496.050 126.450 505.950 ;
        RECT 128.700 501.300 130.800 503.400 ;
        RECT 131.700 501.300 133.800 503.400 ;
        RECT 134.700 501.300 136.800 503.400 ;
        RECT 129.300 497.700 130.500 501.300 ;
        RECT 104.400 493.350 105.600 494.100 ;
        RECT 110.400 493.350 111.600 495.600 ;
        RECT 115.950 493.950 118.050 496.050 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 128.400 495.600 130.500 497.700 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 107.400 488.400 108.600 490.650 ;
        RECT 97.950 478.950 100.050 481.050 ;
        RECT 107.400 466.050 108.450 488.400 ;
        RECT 115.800 487.950 117.900 490.050 ;
        RECT 121.800 487.950 123.900 490.050 ;
        RECT 124.950 487.950 127.050 490.050 ;
        RECT 112.950 484.950 115.050 487.050 ;
        RECT 116.400 486.000 117.600 487.650 ;
        RECT 100.950 463.950 103.050 466.050 ;
        RECT 106.950 463.950 109.050 466.050 ;
        RECT 101.400 451.200 102.450 463.950 ;
        RECT 100.950 449.100 103.050 451.200 ;
        RECT 106.950 450.000 109.050 454.050 ;
        RECT 113.400 453.450 114.450 484.950 ;
        RECT 115.950 481.950 118.050 486.000 ;
        RECT 116.400 472.050 117.450 481.950 ;
        RECT 115.950 469.950 118.050 472.050 ;
        RECT 125.400 469.050 126.450 487.950 ;
        RECT 128.400 476.700 129.900 495.600 ;
        RECT 132.300 484.800 133.500 501.300 ;
        RECT 131.400 482.700 133.500 484.800 ;
        RECT 132.300 476.700 133.500 482.700 ;
        RECT 134.700 479.700 135.900 501.300 ;
        RECT 142.800 500.400 144.900 502.500 ;
        RECT 148.200 501.300 150.300 503.400 ;
        RECT 151.200 501.300 153.300 503.400 ;
        RECT 154.200 501.300 156.300 503.400 ;
        RECT 139.800 493.950 141.900 496.050 ;
        RECT 140.400 492.900 141.600 493.650 ;
        RECT 139.950 490.800 142.050 492.900 ;
        RECT 143.400 489.900 144.300 500.400 ;
        RECT 146.100 494.400 148.200 496.500 ;
        RECT 143.400 487.800 145.500 489.900 ;
        RECT 149.100 489.000 150.300 501.300 ;
        RECT 143.400 481.200 144.300 487.800 ;
        RECT 148.800 486.900 150.900 489.000 ;
        RECT 134.700 477.600 136.800 479.700 ;
        RECT 143.400 479.100 145.500 481.200 ;
        RECT 149.100 479.700 150.300 486.900 ;
        RECT 151.800 483.600 153.300 501.300 ;
        RECT 151.800 481.500 153.900 483.600 ;
        RECT 128.400 474.600 131.400 476.700 ;
        RECT 132.300 474.600 134.400 476.700 ;
        RECT 139.950 475.950 142.050 478.050 ;
        RECT 148.800 477.600 150.900 479.700 ;
        RECT 151.800 476.700 153.300 481.500 ;
        RECT 155.100 479.700 156.300 501.300 ;
        RECT 133.950 469.950 136.050 472.050 ;
        RECT 124.950 466.950 127.050 469.050 ;
        RECT 130.950 460.950 133.050 463.050 ;
        RECT 127.950 457.950 130.050 460.050 ;
        RECT 113.400 452.400 117.450 453.450 ;
        RECT 101.400 448.350 102.600 449.100 ;
        RECT 107.400 448.350 108.600 450.000 ;
        RECT 112.950 448.950 115.050 451.050 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 98.400 443.400 99.600 445.650 ;
        RECT 104.400 444.900 105.600 445.650 ;
        RECT 98.400 436.050 99.450 443.400 ;
        RECT 103.950 442.800 106.050 444.900 ;
        RECT 97.950 433.950 100.050 436.050 ;
        RECT 113.400 424.050 114.450 448.950 ;
        RECT 91.950 421.950 94.050 424.050 ;
        RECT 97.950 421.950 100.050 424.050 ;
        RECT 112.950 421.950 115.050 424.050 ;
        RECT 89.400 417.450 90.600 417.600 ;
        RECT 86.400 416.400 90.600 417.450 ;
        RECT 79.950 400.950 82.050 403.050 ;
        RECT 67.950 394.950 70.050 397.050 ;
        RECT 62.400 374.400 66.450 375.450 ;
        RECT 46.950 371.100 49.050 373.200 ;
        RECT 52.950 371.100 55.050 373.200 ;
        RECT 58.950 371.100 61.050 373.200 ;
        RECT 65.400 372.600 66.450 374.400 ;
        RECT 68.400 373.050 69.450 394.950 ;
        RECT 76.950 373.950 79.050 376.050 ;
        RECT 47.400 334.050 48.450 371.100 ;
        RECT 53.400 370.350 54.600 371.100 ;
        RECT 59.400 370.350 60.600 371.100 ;
        RECT 65.400 370.350 66.600 372.600 ;
        RECT 67.950 370.950 70.050 373.050 ;
        RECT 71.100 370.950 73.200 373.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 64.950 367.950 67.050 370.050 ;
        RECT 71.400 369.900 72.600 370.650 ;
        RECT 70.950 367.800 73.050 369.900 ;
        RECT 77.400 369.450 78.450 373.950 ;
        RECT 80.100 370.950 82.200 373.050 ;
        RECT 80.400 369.450 81.600 370.650 ;
        RECT 77.400 368.400 81.600 369.450 ;
        RECT 56.400 366.000 57.600 367.650 ;
        RECT 55.950 361.950 58.050 366.000 ;
        RECT 62.400 365.400 63.600 367.650 ;
        RECT 62.400 349.050 63.450 365.400 ;
        RECT 67.950 364.950 70.050 367.050 ;
        RECT 61.950 346.950 64.050 349.050 ;
        RECT 68.400 346.050 69.450 364.950 ;
        RECT 86.400 364.050 87.450 416.400 ;
        RECT 89.400 415.350 90.600 416.400 ;
        RECT 89.400 412.950 91.500 415.050 ;
        RECT 94.500 412.950 96.600 415.050 ;
        RECT 95.400 411.450 96.600 412.650 ;
        RECT 98.400 411.900 99.450 421.950 ;
        RECT 111.000 420.900 114.000 421.050 ;
        RECT 111.000 420.450 115.050 420.900 ;
        RECT 110.400 418.950 115.050 420.450 ;
        RECT 110.400 417.600 111.450 418.950 ;
        RECT 112.950 418.800 115.050 418.950 ;
        RECT 116.400 418.050 117.450 452.400 ;
        RECT 121.950 449.100 124.050 451.200 ;
        RECT 128.400 450.600 129.450 457.950 ;
        RECT 131.400 454.050 132.450 460.950 ;
        RECT 130.950 451.950 133.050 454.050 ;
        RECT 134.400 453.600 135.450 469.950 ;
        RECT 136.950 466.950 139.050 469.050 ;
        RECT 137.400 454.050 138.450 466.950 ;
        RECT 140.400 457.050 141.450 475.950 ;
        RECT 142.950 472.950 145.050 475.050 ;
        RECT 151.200 474.600 153.300 476.700 ;
        RECT 154.200 474.600 156.300 479.700 ;
        RECT 157.200 501.300 159.300 503.400 ;
        RECT 157.200 483.600 158.700 501.300 ;
        RECT 157.200 481.500 159.300 483.600 ;
        RECT 157.200 476.700 158.700 481.500 ;
        RECT 157.200 474.600 159.300 476.700 ;
        RECT 139.950 454.950 142.050 457.050 ;
        RECT 134.400 451.350 135.600 453.600 ;
        RECT 136.950 451.950 139.050 454.050 ;
        RECT 122.400 448.350 123.600 449.100 ;
        RECT 128.400 448.350 129.600 450.600 ;
        RECT 133.800 448.950 135.900 451.050 ;
        RECT 139.800 448.950 141.900 451.050 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 127.950 445.950 130.050 448.050 ;
        RECT 118.950 439.950 121.050 445.050 ;
        RECT 125.400 444.900 126.600 445.650 ;
        RECT 124.950 442.800 127.050 444.900 ;
        RECT 130.800 442.950 132.900 445.050 ;
        RECT 133.950 442.950 136.050 445.050 ;
        RECT 131.400 427.050 132.450 442.950 ;
        RECT 134.400 430.050 135.450 442.950 ;
        RECT 139.950 439.950 142.050 442.050 ;
        RECT 133.950 427.950 136.050 430.050 ;
        RECT 124.950 424.950 127.050 427.050 ;
        RECT 130.950 424.950 133.050 427.050 ;
        RECT 125.400 418.050 126.450 424.950 ;
        RECT 110.400 415.350 111.600 417.600 ;
        RECT 115.950 415.950 118.050 418.050 ;
        RECT 121.800 415.950 123.900 418.050 ;
        RECT 124.950 415.950 127.050 418.050 ;
        RECT 127.950 417.000 130.050 421.050 ;
        RECT 136.950 418.800 139.050 420.900 ;
        RECT 106.950 412.950 109.050 415.050 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 107.400 411.900 108.600 412.650 ;
        RECT 97.950 411.450 100.050 411.900 ;
        RECT 95.400 410.400 100.050 411.450 ;
        RECT 97.950 409.800 100.050 410.400 ;
        RECT 106.950 409.800 109.050 411.900 ;
        RECT 113.400 410.400 114.600 412.650 ;
        RECT 113.400 394.050 114.450 410.400 ;
        RECT 112.950 391.950 115.050 394.050 ;
        RECT 89.700 384.300 91.800 386.400 ;
        RECT 90.300 379.500 91.800 384.300 ;
        RECT 89.700 377.400 91.800 379.500 ;
        RECT 85.950 361.950 88.050 364.050 ;
        RECT 90.300 359.700 91.800 377.400 ;
        RECT 89.700 357.600 91.800 359.700 ;
        RECT 92.700 381.300 94.800 386.400 ;
        RECT 95.700 384.300 97.800 386.400 ;
        RECT 114.600 384.300 116.700 386.400 ;
        RECT 117.600 384.300 120.600 386.400 ;
        RECT 122.400 385.050 123.450 415.950 ;
        RECT 128.400 415.350 129.600 417.000 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 131.400 411.900 132.600 412.650 ;
        RECT 137.400 411.900 138.450 418.800 ;
        RECT 130.950 409.800 133.050 411.900 ;
        RECT 136.950 409.800 139.050 411.900 ;
        RECT 130.950 403.950 133.050 406.050 ;
        RECT 92.700 359.700 93.900 381.300 ;
        RECT 95.700 379.500 97.200 384.300 ;
        RECT 98.100 381.300 100.200 383.400 ;
        RECT 95.100 377.400 97.200 379.500 ;
        RECT 95.700 359.700 97.200 377.400 ;
        RECT 98.700 374.100 99.900 381.300 ;
        RECT 103.500 379.800 105.600 381.900 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 112.200 381.300 114.300 383.400 ;
        RECT 98.100 372.000 100.200 374.100 ;
        RECT 104.700 373.200 105.600 379.800 ;
        RECT 98.700 359.700 99.900 372.000 ;
        RECT 103.500 371.100 105.600 373.200 ;
        RECT 100.800 364.500 102.900 366.600 ;
        RECT 104.700 360.600 105.600 371.100 ;
        RECT 107.400 369.600 108.450 379.950 ;
        RECT 107.400 367.350 108.600 369.600 ;
        RECT 107.100 364.950 109.200 367.050 ;
        RECT 92.700 357.600 94.800 359.700 ;
        RECT 95.700 357.600 97.800 359.700 ;
        RECT 98.700 357.600 100.800 359.700 ;
        RECT 104.100 358.500 106.200 360.600 ;
        RECT 113.100 359.700 114.300 381.300 ;
        RECT 115.500 378.300 116.700 384.300 ;
        RECT 115.500 376.200 117.600 378.300 ;
        RECT 115.500 359.700 116.700 376.200 ;
        RECT 119.100 365.400 120.600 384.300 ;
        RECT 121.950 382.950 124.050 385.050 ;
        RECT 131.400 376.200 132.450 403.950 ;
        RECT 121.950 373.950 124.050 376.050 ;
        RECT 130.950 374.100 133.050 376.200 ;
        RECT 118.500 363.300 120.600 365.400 ;
        RECT 118.500 359.700 119.700 363.300 ;
        RECT 112.200 357.600 114.300 359.700 ;
        RECT 115.200 357.600 117.300 359.700 ;
        RECT 118.200 357.600 120.300 359.700 ;
        RECT 112.950 352.950 115.050 355.050 ;
        RECT 67.950 343.950 70.050 346.050 ;
        RECT 76.950 343.950 79.050 346.050 ;
        RECT 80.700 345.300 82.800 347.400 ;
        RECT 56.400 339.450 57.600 339.600 ;
        RECT 56.400 338.400 63.450 339.450 ;
        RECT 56.400 337.350 57.600 338.400 ;
        RECT 62.400 337.200 63.450 338.400 ;
        RECT 52.950 334.950 55.050 337.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 61.950 335.100 64.050 337.200 ;
        RECT 46.950 331.950 49.050 334.050 ;
        RECT 53.400 333.900 54.600 334.650 ;
        RECT 62.400 334.350 63.600 335.100 ;
        RECT 67.950 334.950 70.050 337.050 ;
        RECT 70.950 336.000 73.050 340.050 ;
        RECT 77.400 336.900 78.450 343.950 ;
        RECT 52.950 331.800 55.050 333.900 ;
        RECT 62.100 331.950 64.200 334.050 ;
        RECT 40.950 322.950 43.050 325.050 ;
        RECT 58.950 322.950 61.050 325.050 ;
        RECT 49.950 307.950 52.050 310.050 ;
        RECT 37.950 301.950 40.050 304.050 ;
        RECT 46.950 301.950 49.050 304.050 ;
        RECT 34.950 298.950 37.050 301.050 ;
        RECT 29.400 296.400 34.050 298.050 ;
        RECT 30.000 295.950 34.050 296.400 ;
        RECT 28.950 293.100 31.050 295.200 ;
        RECT 35.400 294.600 36.450 298.950 ;
        RECT 29.400 292.350 30.600 293.100 ;
        RECT 35.400 292.350 36.600 294.600 ;
        RECT 40.950 293.100 43.050 295.200 ;
        RECT 41.400 292.350 42.600 293.100 ;
        RECT 28.950 289.950 31.050 292.050 ;
        RECT 31.950 289.950 34.050 292.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 32.400 288.900 33.600 289.650 ;
        RECT 38.400 288.900 39.600 289.650 ;
        RECT 22.950 286.800 25.050 288.900 ;
        RECT 31.950 286.800 34.050 288.900 ;
        RECT 37.950 286.800 40.050 288.900 ;
        RECT 47.400 274.050 48.450 301.950 ;
        RECT 50.400 295.050 51.450 307.950 ;
        RECT 55.950 298.950 58.050 301.050 ;
        RECT 49.950 292.950 52.050 295.050 ;
        RECT 56.400 294.600 57.450 298.950 ;
        RECT 59.400 295.050 60.450 322.950 ;
        RECT 68.400 310.050 69.450 334.950 ;
        RECT 71.400 334.350 72.600 336.000 ;
        RECT 76.950 334.800 79.050 336.900 ;
        RECT 71.100 331.950 73.200 334.050 ;
        RECT 81.300 327.600 82.800 345.300 ;
        RECT 80.700 325.500 82.800 327.600 ;
        RECT 81.300 320.700 82.800 325.500 ;
        RECT 80.700 318.600 82.800 320.700 ;
        RECT 83.700 345.300 85.800 347.400 ;
        RECT 86.700 345.300 88.800 347.400 ;
        RECT 89.700 345.300 91.800 347.400 ;
        RECT 83.700 323.700 84.900 345.300 ;
        RECT 86.700 327.600 88.200 345.300 ;
        RECT 89.700 333.000 90.900 345.300 ;
        RECT 95.100 344.400 97.200 346.500 ;
        RECT 103.200 345.300 105.300 347.400 ;
        RECT 106.200 345.300 108.300 347.400 ;
        RECT 109.200 345.300 111.300 347.400 ;
        RECT 91.800 338.400 93.900 340.500 ;
        RECT 95.700 333.900 96.600 344.400 ;
        RECT 98.100 337.950 100.200 340.050 ;
        RECT 98.400 336.900 99.600 337.650 ;
        RECT 97.950 334.800 100.050 336.900 ;
        RECT 89.100 330.900 91.200 333.000 ;
        RECT 94.500 331.800 96.600 333.900 ;
        RECT 86.100 325.500 88.200 327.600 ;
        RECT 83.700 318.600 85.800 323.700 ;
        RECT 86.700 320.700 88.200 325.500 ;
        RECT 89.700 323.700 90.900 330.900 ;
        RECT 95.700 325.200 96.600 331.800 ;
        RECT 89.100 321.600 91.200 323.700 ;
        RECT 94.500 323.100 96.600 325.200 ;
        RECT 104.100 323.700 105.300 345.300 ;
        RECT 103.200 321.600 105.300 323.700 ;
        RECT 106.500 328.800 107.700 345.300 ;
        RECT 109.500 341.700 110.700 345.300 ;
        RECT 113.400 343.050 114.450 352.950 ;
        RECT 109.500 339.600 111.600 341.700 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 122.400 340.050 123.450 373.950 ;
        RECT 131.400 373.350 132.600 374.100 ;
        RECT 125.100 370.950 127.200 373.050 ;
        RECT 131.100 370.950 133.200 373.050 ;
        RECT 137.400 369.450 138.450 409.800 ;
        RECT 140.400 403.050 141.450 439.950 ;
        RECT 143.400 421.050 144.450 472.950 ;
        RECT 161.400 471.450 162.450 517.950 ;
        RECT 163.950 517.800 166.050 519.900 ;
        RECT 164.400 510.450 165.450 517.800 ;
        RECT 167.400 514.050 168.450 520.950 ;
        RECT 172.950 520.800 175.050 522.900 ;
        RECT 175.950 520.950 178.050 523.050 ;
        RECT 166.950 511.950 169.050 514.050 ;
        RECT 164.400 509.400 174.450 510.450 ;
        RECT 169.950 505.950 172.050 508.050 ;
        RECT 166.950 491.100 169.050 493.200 ;
        RECT 167.400 490.350 168.600 491.100 ;
        RECT 166.800 487.950 168.900 490.050 ;
        RECT 170.400 475.050 171.450 505.950 ;
        RECT 173.400 505.050 174.450 509.400 ;
        RECT 172.950 502.950 175.050 505.050 ;
        RECT 176.400 502.050 177.450 520.950 ;
        RECT 179.400 514.050 180.450 529.950 ;
        RECT 182.400 529.050 183.450 556.950 ;
        RECT 191.400 547.050 192.450 586.950 ;
        RECT 205.950 580.950 208.050 583.050 ;
        RECT 193.950 571.950 196.050 574.050 ;
        RECT 199.950 572.100 202.050 574.200 ;
        RECT 206.400 573.600 207.450 580.950 ;
        RECT 214.950 577.950 217.050 580.050 ;
        RECT 190.950 544.950 193.050 547.050 ;
        RECT 187.950 532.950 190.050 535.050 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 188.400 528.600 189.450 532.950 ;
        RECT 194.400 532.050 195.450 571.950 ;
        RECT 200.400 571.350 201.600 572.100 ;
        RECT 206.400 571.350 207.600 573.600 ;
        RECT 211.950 571.950 214.050 577.050 ;
        RECT 199.950 568.950 202.050 571.050 ;
        RECT 202.950 568.950 205.050 571.050 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 203.400 566.400 204.600 568.650 ;
        RECT 209.400 567.900 210.600 568.650 ;
        RECT 199.950 538.950 202.050 541.050 ;
        RECT 190.950 530.400 195.450 532.050 ;
        RECT 190.950 529.950 195.000 530.400 ;
        RECT 188.400 526.350 189.600 528.600 ;
        RECT 193.950 527.100 196.050 529.200 ;
        RECT 194.400 526.350 195.600 527.100 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 193.950 523.950 196.050 526.050 ;
        RECT 181.950 520.950 184.050 523.050 ;
        RECT 185.400 521.400 186.600 523.650 ;
        RECT 191.400 522.900 192.600 523.650 ;
        RECT 178.950 511.950 181.050 514.050 ;
        RECT 175.950 499.950 178.050 502.050 ;
        RECT 172.950 496.950 175.050 499.050 ;
        RECT 173.400 492.450 174.450 496.950 ;
        RECT 175.950 492.450 178.050 493.200 ;
        RECT 173.400 491.400 178.050 492.450 ;
        RECT 175.950 491.100 178.050 491.400 ;
        RECT 176.400 490.350 177.600 491.100 ;
        RECT 175.800 487.950 177.900 490.050 ;
        RECT 172.950 484.950 175.050 487.050 ;
        RECT 173.400 478.050 174.450 484.950 ;
        RECT 172.950 475.950 175.050 478.050 ;
        RECT 169.950 472.950 172.050 475.050 ;
        RECT 158.400 470.400 162.450 471.450 ;
        RECT 146.400 462.300 149.400 464.400 ;
        RECT 150.300 462.300 152.400 464.400 ;
        RECT 146.400 443.400 147.900 462.300 ;
        RECT 150.300 456.300 151.500 462.300 ;
        RECT 149.400 454.200 151.500 456.300 ;
        RECT 146.400 441.300 148.500 443.400 ;
        RECT 147.300 437.700 148.500 441.300 ;
        RECT 150.300 437.700 151.500 454.200 ;
        RECT 152.700 459.300 154.800 461.400 ;
        RECT 152.700 437.700 153.900 459.300 ;
        RECT 158.400 456.450 159.450 470.400 ;
        RECT 169.200 462.300 171.300 464.400 ;
        RECT 155.400 455.400 159.450 456.450 ;
        RECT 161.400 457.800 163.500 459.900 ;
        RECT 166.800 459.300 168.900 461.400 ;
        RECT 155.400 448.050 156.450 455.400 ;
        RECT 157.950 451.950 160.050 454.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 158.400 447.600 159.450 451.950 ;
        RECT 161.400 451.200 162.300 457.800 ;
        RECT 167.100 452.100 168.300 459.300 ;
        RECT 169.800 457.500 171.300 462.300 ;
        RECT 172.200 459.300 174.300 464.400 ;
        RECT 169.800 455.400 171.900 457.500 ;
        RECT 161.400 449.100 163.500 451.200 ;
        RECT 166.800 450.000 168.900 452.100 ;
        RECT 158.400 445.350 159.600 447.600 ;
        RECT 157.800 442.950 159.900 445.050 ;
        RECT 161.400 438.600 162.300 449.100 ;
        RECT 164.100 442.500 166.200 444.600 ;
        RECT 146.700 435.600 148.800 437.700 ;
        RECT 149.700 435.600 151.800 437.700 ;
        RECT 152.700 435.600 154.800 437.700 ;
        RECT 160.800 436.500 162.900 438.600 ;
        RECT 167.100 437.700 168.300 450.000 ;
        RECT 169.800 437.700 171.300 455.400 ;
        RECT 173.100 437.700 174.300 459.300 ;
        RECT 166.200 435.600 168.300 437.700 ;
        RECT 169.200 435.600 171.300 437.700 ;
        RECT 172.200 435.600 174.300 437.700 ;
        RECT 175.200 462.300 177.300 464.400 ;
        RECT 175.200 457.500 176.700 462.300 ;
        RECT 175.200 455.400 177.300 457.500 ;
        RECT 175.200 437.700 176.700 455.400 ;
        RECT 175.200 435.600 177.300 437.700 ;
        RECT 157.950 427.950 160.050 430.050 ;
        RECT 142.950 418.950 145.050 421.050 ;
        RECT 145.950 416.100 148.050 418.200 ;
        RECT 152.400 417.450 153.600 417.600 ;
        RECT 154.950 417.450 157.050 421.050 ;
        RECT 152.400 417.000 157.050 417.450 ;
        RECT 152.400 416.400 156.450 417.000 ;
        RECT 146.400 415.350 147.600 416.100 ;
        RECT 152.400 415.350 153.600 416.400 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 142.950 409.950 145.050 412.050 ;
        RECT 149.400 410.400 150.600 412.650 ;
        RECT 143.400 406.050 144.450 409.950 ;
        RECT 149.400 409.050 150.450 410.400 ;
        RECT 149.400 407.400 154.050 409.050 ;
        RECT 150.000 406.950 154.050 407.400 ;
        RECT 142.950 403.950 145.050 406.050 ;
        RECT 148.950 403.950 151.050 406.050 ;
        RECT 139.950 400.950 142.050 403.050 ;
        RECT 149.400 372.600 150.450 403.950 ;
        RECT 151.950 394.950 154.050 397.050 ;
        RECT 152.400 376.050 153.450 394.950 ;
        RECT 158.400 388.050 159.450 427.950 ;
        RECT 175.950 424.950 178.050 427.050 ;
        RECT 160.950 418.950 163.050 421.050 ;
        RECT 161.400 411.900 162.450 418.950 ;
        RECT 169.950 416.100 172.050 418.200 ;
        RECT 170.400 415.350 171.600 416.100 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 167.400 411.900 168.600 412.650 ;
        RECT 160.950 409.800 163.050 411.900 ;
        RECT 166.950 409.800 169.050 411.900 ;
        RECT 161.400 394.050 162.450 409.800 ;
        RECT 160.950 391.950 163.050 394.050 ;
        RECT 157.950 385.950 160.050 388.050 ;
        RECT 163.950 385.950 166.050 388.050 ;
        RECT 154.950 382.950 157.050 385.050 ;
        RECT 151.950 373.950 154.050 376.050 ;
        RECT 155.400 372.600 156.450 382.950 ;
        RECT 160.950 376.950 163.050 379.050 ;
        RECT 149.400 370.350 150.600 372.600 ;
        RECT 155.400 370.350 156.600 372.600 ;
        RECT 134.400 368.400 138.450 369.450 ;
        RECT 127.950 364.950 130.050 367.050 ;
        RECT 124.950 361.950 127.050 364.050 ;
        RECT 106.500 326.700 108.600 328.800 ;
        RECT 106.500 320.700 107.700 326.700 ;
        RECT 110.100 320.700 111.600 339.600 ;
        RECT 121.950 337.950 124.050 340.050 ;
        RECT 125.400 337.050 126.450 361.950 ;
        RECT 128.400 349.050 129.450 364.950 ;
        RECT 130.950 355.950 133.050 358.050 ;
        RECT 127.950 346.950 130.050 349.050 ;
        RECT 127.950 337.950 130.050 340.050 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 116.100 331.950 118.200 334.050 ;
        RECT 122.100 331.950 124.200 334.050 ;
        RECT 122.400 330.900 123.600 331.650 ;
        RECT 128.400 330.900 129.450 337.950 ;
        RECT 121.950 328.800 124.050 330.900 ;
        RECT 127.950 328.800 130.050 330.900 ;
        RECT 86.700 318.600 88.800 320.700 ;
        RECT 105.600 318.600 107.700 320.700 ;
        RECT 108.600 318.600 111.600 320.700 ;
        RECT 67.950 307.950 70.050 310.050 ;
        RECT 80.700 306.300 82.800 308.400 ;
        RECT 67.950 301.950 70.050 304.050 ;
        RECT 56.400 292.350 57.600 294.600 ;
        RECT 58.950 292.950 61.050 295.050 ;
        RECT 62.100 292.950 64.200 295.050 ;
        RECT 52.950 289.950 55.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 62.400 290.400 63.600 292.650 ;
        RECT 49.950 286.950 52.050 289.050 ;
        RECT 53.400 287.400 54.600 289.650 ;
        RECT 62.400 288.450 63.450 290.400 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 68.400 291.450 69.450 301.950 ;
        RECT 81.300 301.500 82.800 306.300 ;
        RECT 80.700 299.400 82.800 301.500 ;
        RECT 71.100 292.950 73.200 295.050 ;
        RECT 71.400 291.450 72.600 292.650 ;
        RECT 68.400 290.400 72.600 291.450 ;
        RECT 59.400 287.400 63.450 288.450 ;
        RECT 50.400 277.050 51.450 286.950 ;
        RECT 53.400 285.450 54.450 287.400 ;
        RECT 59.400 285.450 60.450 287.400 ;
        RECT 53.400 284.400 60.450 285.450 ;
        RECT 49.950 274.950 52.050 277.050 ;
        RECT 55.950 274.950 58.050 277.050 ;
        RECT 46.950 271.950 49.050 274.050 ;
        RECT 23.700 267.300 25.800 269.400 ;
        RECT 8.400 257.400 12.450 258.450 ;
        RECT 5.100 253.950 7.200 256.050 ;
        RECT 5.100 214.950 7.200 217.050 ;
        RECT 5.400 212.400 6.600 214.650 ;
        RECT 5.400 202.050 6.450 212.400 ;
        RECT 11.400 205.050 12.450 257.400 ;
        RECT 14.400 256.350 15.600 258.600 ;
        RECT 19.950 256.800 22.050 258.900 ;
        RECT 14.100 253.950 16.200 256.050 ;
        RECT 24.300 249.600 25.800 267.300 ;
        RECT 23.700 247.500 25.800 249.600 ;
        RECT 24.300 242.700 25.800 247.500 ;
        RECT 23.700 240.600 25.800 242.700 ;
        RECT 26.700 267.300 28.800 269.400 ;
        RECT 29.700 267.300 31.800 269.400 ;
        RECT 32.700 267.300 34.800 269.400 ;
        RECT 26.700 245.700 27.900 267.300 ;
        RECT 29.700 249.600 31.200 267.300 ;
        RECT 32.700 255.000 33.900 267.300 ;
        RECT 38.100 266.400 40.200 268.500 ;
        RECT 46.200 267.300 48.300 269.400 ;
        RECT 49.200 267.300 51.300 269.400 ;
        RECT 52.200 267.300 54.300 269.400 ;
        RECT 34.800 260.400 36.900 262.500 ;
        RECT 38.700 255.900 39.600 266.400 ;
        RECT 41.100 259.950 43.200 262.050 ;
        RECT 41.400 258.900 42.600 259.650 ;
        RECT 40.800 256.800 42.900 258.900 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 32.100 252.900 34.200 255.000 ;
        RECT 37.500 253.800 39.600 255.900 ;
        RECT 29.100 247.500 31.200 249.600 ;
        RECT 26.700 240.600 28.800 245.700 ;
        RECT 29.700 242.700 31.200 247.500 ;
        RECT 32.700 245.700 33.900 252.900 ;
        RECT 38.700 247.200 39.600 253.800 ;
        RECT 44.400 249.450 45.450 256.950 ;
        RECT 32.100 243.600 34.200 245.700 ;
        RECT 37.500 245.100 39.600 247.200 ;
        RECT 41.400 248.400 45.450 249.450 ;
        RECT 29.700 240.600 31.800 242.700 ;
        RECT 23.700 228.300 25.800 230.400 ;
        RECT 24.300 223.500 25.800 228.300 ;
        RECT 23.700 221.400 25.800 223.500 ;
        RECT 19.950 217.950 22.050 220.050 ;
        RECT 14.100 214.950 16.200 217.050 ;
        RECT 14.400 213.900 15.600 214.650 ;
        RECT 13.950 211.800 16.050 213.900 ;
        RECT 10.950 202.950 13.050 205.050 ;
        RECT 16.950 202.950 19.050 205.050 ;
        RECT 4.950 199.950 7.050 202.050 ;
        RECT 1.950 104.100 4.050 106.200 ;
        RECT 1.950 73.950 4.050 76.050 ;
        RECT 2.400 54.900 3.450 73.950 ;
        RECT 1.950 52.800 4.050 54.900 ;
        RECT 5.400 28.200 6.450 199.950 ;
        RECT 10.950 199.800 13.050 201.900 ;
        RECT 11.400 183.600 12.450 199.800 ;
        RECT 17.400 184.050 18.450 202.950 ;
        RECT 11.400 181.350 12.600 183.600 ;
        RECT 16.950 181.950 19.050 184.050 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 14.400 177.900 15.600 178.650 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 20.400 169.050 21.450 217.950 ;
        RECT 24.300 203.700 25.800 221.400 ;
        RECT 23.700 201.600 25.800 203.700 ;
        RECT 26.700 225.300 28.800 230.400 ;
        RECT 29.700 228.300 31.800 230.400 ;
        RECT 26.700 203.700 27.900 225.300 ;
        RECT 29.700 223.500 31.200 228.300 ;
        RECT 32.100 225.300 34.200 227.400 ;
        RECT 29.100 221.400 31.200 223.500 ;
        RECT 29.700 203.700 31.200 221.400 ;
        RECT 32.700 218.100 33.900 225.300 ;
        RECT 37.500 223.800 39.600 225.900 ;
        RECT 32.100 216.000 34.200 218.100 ;
        RECT 38.700 217.200 39.600 223.800 ;
        RECT 41.400 222.450 42.450 248.400 ;
        RECT 47.100 245.700 48.300 267.300 ;
        RECT 46.200 243.600 48.300 245.700 ;
        RECT 49.500 250.800 50.700 267.300 ;
        RECT 52.500 263.700 53.700 267.300 ;
        RECT 52.500 261.600 54.600 263.700 ;
        RECT 49.500 248.700 51.600 250.800 ;
        RECT 49.500 242.700 50.700 248.700 ;
        RECT 53.100 242.700 54.600 261.600 ;
        RECT 48.600 240.600 50.700 242.700 ;
        RECT 51.600 240.600 54.600 242.700 ;
        RECT 48.600 228.300 50.700 230.400 ;
        RECT 51.600 228.300 54.600 230.400 ;
        RECT 46.200 225.300 48.300 227.400 ;
        RECT 41.400 221.400 45.450 222.450 ;
        RECT 40.950 217.950 43.050 220.050 ;
        RECT 32.700 203.700 33.900 216.000 ;
        RECT 37.500 215.100 39.600 217.200 ;
        RECT 34.800 208.500 36.900 210.600 ;
        RECT 38.700 204.600 39.600 215.100 ;
        RECT 41.400 213.600 42.450 217.950 ;
        RECT 44.400 214.050 45.450 221.400 ;
        RECT 41.400 211.350 42.600 213.600 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 41.100 208.950 43.200 211.050 ;
        RECT 26.700 201.600 28.800 203.700 ;
        RECT 29.700 201.600 31.800 203.700 ;
        RECT 32.700 201.600 34.800 203.700 ;
        RECT 38.100 202.500 40.200 204.600 ;
        RECT 47.100 203.700 48.300 225.300 ;
        RECT 49.500 222.300 50.700 228.300 ;
        RECT 49.500 220.200 51.600 222.300 ;
        RECT 49.500 203.700 50.700 220.200 ;
        RECT 53.100 209.400 54.600 228.300 ;
        RECT 52.500 207.300 54.600 209.400 ;
        RECT 52.500 203.700 53.700 207.300 ;
        RECT 46.200 201.600 48.300 203.700 ;
        RECT 49.200 201.600 51.300 203.700 ;
        RECT 52.200 201.600 54.300 203.700 ;
        RECT 49.950 196.950 52.050 199.050 ;
        RECT 50.400 190.050 51.450 196.950 ;
        RECT 56.400 190.050 57.450 274.950 ;
        RECT 62.400 259.050 63.450 287.400 ;
        RECT 65.400 277.050 66.450 289.950 ;
        RECT 64.950 274.950 67.050 277.050 ;
        RECT 71.400 259.050 72.450 290.400 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 70.950 256.950 73.050 259.050 ;
        RECT 59.100 253.950 61.200 256.050 ;
        RECT 65.100 253.950 67.200 256.050 ;
        RECT 70.950 253.800 73.050 255.900 ;
        RECT 65.400 252.900 66.600 253.650 ;
        RECT 64.950 250.800 67.050 252.900 ;
        RECT 65.400 219.600 66.450 250.800 ;
        RECT 65.400 217.350 66.600 219.600 ;
        RECT 59.100 214.950 61.200 217.050 ;
        RECT 65.100 214.950 67.200 217.050 ;
        RECT 61.950 208.950 64.050 211.050 ;
        RECT 58.950 205.950 61.050 208.050 ;
        RECT 31.950 187.950 34.050 190.050 ;
        RECT 32.400 183.600 33.450 187.950 ;
        RECT 37.950 185.100 40.050 190.050 ;
        RECT 46.950 187.950 49.050 190.050 ;
        RECT 49.950 187.950 52.050 190.050 ;
        RECT 55.950 187.950 58.050 190.050 ;
        RECT 32.400 181.350 33.600 183.600 ;
        RECT 37.950 181.950 40.050 184.050 ;
        RECT 38.400 181.350 39.600 181.950 ;
        RECT 28.950 178.950 31.050 181.050 ;
        RECT 31.950 178.950 34.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 29.400 177.900 30.600 178.650 ;
        RECT 28.950 175.800 31.050 177.900 ;
        RECT 35.400 176.400 36.600 178.650 ;
        RECT 41.400 177.900 42.600 178.650 ;
        RECT 35.400 169.050 36.450 176.400 ;
        RECT 40.950 175.800 43.050 177.900 ;
        RECT 19.950 166.950 22.050 169.050 ;
        RECT 34.950 166.950 37.050 169.050 ;
        RECT 31.950 160.950 34.050 163.050 ;
        RECT 16.950 137.100 19.050 139.200 ;
        RECT 32.400 139.050 33.450 160.950 ;
        RECT 43.950 148.950 46.050 151.050 ;
        RECT 23.400 138.450 24.600 138.600 ;
        RECT 23.400 137.400 30.450 138.450 ;
        RECT 17.400 136.350 18.600 137.100 ;
        RECT 23.400 136.350 24.600 137.400 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 10.950 130.950 13.050 133.050 ;
        RECT 14.400 132.000 15.600 133.650 ;
        RECT 20.400 132.900 21.600 133.650 ;
        RECT 11.400 121.050 12.450 130.950 ;
        RECT 13.950 127.950 16.050 132.000 ;
        RECT 19.950 130.800 22.050 132.900 ;
        RECT 29.400 130.050 30.450 137.400 ;
        RECT 31.800 136.950 33.900 139.050 ;
        RECT 34.950 137.100 37.050 139.200 ;
        RECT 40.950 137.100 43.050 139.200 ;
        RECT 44.400 139.050 45.450 148.950 ;
        RECT 35.400 136.350 36.600 137.100 ;
        RECT 41.400 136.350 42.600 137.100 ;
        RECT 43.950 136.950 46.050 139.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 31.950 130.950 34.050 133.050 ;
        RECT 38.400 132.000 39.600 133.650 ;
        RECT 22.950 127.950 25.050 130.050 ;
        RECT 28.950 127.950 31.050 130.050 ;
        RECT 10.950 118.950 13.050 121.050 ;
        RECT 10.950 104.100 13.050 106.200 ;
        RECT 11.400 103.350 12.600 104.100 ;
        RECT 11.400 100.950 13.500 103.050 ;
        RECT 16.800 100.950 18.900 103.050 ;
        RECT 23.400 99.900 24.450 127.950 ;
        RECT 32.400 112.050 33.450 130.950 ;
        RECT 37.950 127.950 40.050 132.000 ;
        RECT 31.950 109.950 34.050 112.050 ;
        RECT 37.950 109.950 40.050 112.050 ;
        RECT 38.400 109.200 39.600 109.950 ;
        RECT 33.900 105.900 36.000 107.700 ;
        RECT 37.800 106.800 39.900 108.900 ;
        RECT 41.100 108.300 43.200 110.400 ;
        RECT 32.400 104.700 41.100 105.900 ;
        RECT 29.100 100.950 31.200 103.050 ;
        RECT 29.400 99.900 30.600 100.650 ;
        RECT 22.950 97.800 25.050 99.900 ;
        RECT 28.950 97.800 31.050 99.900 ;
        RECT 13.950 60.000 16.050 64.050 ;
        RECT 14.400 58.350 15.600 60.000 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 17.400 54.900 18.600 55.650 ;
        RECT 23.400 55.050 24.450 97.800 ;
        RECT 32.400 95.700 33.300 104.700 ;
        RECT 39.000 103.800 41.100 104.700 ;
        RECT 42.000 102.900 42.900 108.300 ;
        RECT 43.950 104.100 46.050 106.200 ;
        RECT 44.400 103.350 45.600 104.100 ;
        RECT 36.000 101.700 42.900 102.900 ;
        RECT 36.000 99.300 36.900 101.700 ;
        RECT 34.800 97.200 36.900 99.300 ;
        RECT 37.800 97.950 39.900 100.050 ;
        RECT 31.500 93.600 33.600 95.700 ;
        RECT 38.400 95.400 39.600 97.650 ;
        RECT 41.700 94.500 42.900 101.700 ;
        RECT 43.800 100.950 45.900 103.050 ;
        RECT 41.100 92.400 43.200 94.500 ;
        RECT 37.950 73.950 40.050 76.050 ;
        RECT 28.950 64.050 31.050 64.200 ;
        RECT 31.950 64.050 34.050 64.200 ;
        RECT 28.950 62.100 34.050 64.050 ;
        RECT 30.000 61.950 33.000 62.100 ;
        RECT 31.950 58.950 34.050 61.050 ;
        RECT 38.400 60.600 39.450 73.950 ;
        RECT 47.400 64.050 48.450 187.950 ;
        RECT 55.950 182.100 58.050 184.200 ;
        RECT 59.400 184.050 60.450 205.950 ;
        RECT 56.400 181.350 57.600 182.100 ;
        RECT 58.950 181.950 61.050 184.050 ;
        RECT 62.400 181.050 63.450 208.950 ;
        RECT 71.400 196.050 72.450 253.800 ;
        RECT 74.400 211.050 75.450 289.950 ;
        RECT 81.300 281.700 82.800 299.400 ;
        RECT 80.700 279.600 82.800 281.700 ;
        RECT 83.700 303.300 85.800 308.400 ;
        RECT 86.700 306.300 88.800 308.400 ;
        RECT 105.600 306.300 107.700 308.400 ;
        RECT 108.600 306.300 111.600 308.400 ;
        RECT 83.700 281.700 84.900 303.300 ;
        RECT 86.700 301.500 88.200 306.300 ;
        RECT 89.100 303.300 91.200 305.400 ;
        RECT 86.100 299.400 88.200 301.500 ;
        RECT 86.700 281.700 88.200 299.400 ;
        RECT 89.700 296.100 90.900 303.300 ;
        RECT 94.500 301.800 96.600 303.900 ;
        RECT 103.200 303.300 105.300 305.400 ;
        RECT 89.100 294.000 91.200 296.100 ;
        RECT 95.700 295.200 96.600 301.800 ;
        RECT 97.950 295.950 100.050 298.050 ;
        RECT 89.700 281.700 90.900 294.000 ;
        RECT 94.500 293.100 96.600 295.200 ;
        RECT 91.800 286.500 93.900 288.600 ;
        RECT 95.700 282.600 96.600 293.100 ;
        RECT 98.400 291.600 99.450 295.950 ;
        RECT 98.400 289.350 99.600 291.600 ;
        RECT 98.100 286.950 100.200 289.050 ;
        RECT 83.700 279.600 85.800 281.700 ;
        RECT 86.700 279.600 88.800 281.700 ;
        RECT 89.700 279.600 91.800 281.700 ;
        RECT 95.100 280.500 97.200 282.600 ;
        RECT 104.100 281.700 105.300 303.300 ;
        RECT 106.500 300.300 107.700 306.300 ;
        RECT 106.500 298.200 108.600 300.300 ;
        RECT 106.500 281.700 107.700 298.200 ;
        RECT 110.100 287.400 111.600 306.300 ;
        RECT 122.400 297.600 123.450 328.800 ;
        RECT 122.400 295.350 123.600 297.600 ;
        RECT 116.100 292.950 118.200 295.050 ;
        RECT 122.100 292.950 124.200 295.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 109.500 285.300 111.600 287.400 ;
        RECT 115.950 286.950 118.050 289.050 ;
        RECT 109.500 281.700 110.700 285.300 ;
        RECT 103.200 279.600 105.300 281.700 ;
        RECT 106.200 279.600 108.300 281.700 ;
        RECT 109.200 279.600 111.300 281.700 ;
        RECT 112.950 277.950 115.050 280.050 ;
        RECT 82.950 274.950 85.050 277.050 ;
        RECT 88.950 274.950 91.050 277.050 ;
        RECT 100.950 274.950 103.050 277.050 ;
        RECT 83.400 261.600 84.450 274.950 ;
        RECT 89.400 261.600 90.450 274.950 ;
        RECT 97.950 271.950 100.050 274.050 ;
        RECT 94.950 265.950 97.050 268.050 ;
        RECT 83.400 259.350 84.600 261.600 ;
        RECT 89.400 259.350 90.600 261.600 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 76.950 253.950 79.050 256.050 ;
        RECT 80.400 254.400 81.600 256.650 ;
        RECT 86.400 255.900 87.600 256.650 ;
        RECT 77.400 241.050 78.450 253.950 ;
        RECT 80.400 250.050 81.450 254.400 ;
        RECT 85.950 253.800 88.050 255.900 ;
        RECT 95.400 252.900 96.450 265.950 ;
        RECT 94.950 250.800 97.050 252.900 ;
        RECT 79.950 247.950 82.050 250.050 ;
        RECT 76.950 238.950 79.050 241.050 ;
        RECT 88.950 232.950 91.050 235.050 ;
        RECT 82.950 229.950 85.050 232.050 ;
        RECT 83.400 216.600 84.450 229.950 ;
        RECT 89.400 217.050 90.450 232.950 ;
        RECT 95.400 223.050 96.450 250.800 ;
        RECT 98.400 250.050 99.450 271.950 ;
        RECT 101.400 262.050 102.450 274.950 ;
        RECT 113.400 271.050 114.450 277.950 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 112.950 268.950 115.050 271.050 ;
        RECT 100.950 259.950 103.050 262.050 ;
        RECT 107.400 261.600 108.450 268.950 ;
        RECT 116.400 268.050 117.450 286.950 ;
        RECT 125.400 286.050 126.450 289.950 ;
        RECT 128.400 289.050 129.450 328.800 ;
        RECT 127.950 286.950 130.050 289.050 ;
        RECT 124.950 283.950 127.050 286.050 ;
        RECT 115.950 265.950 118.050 268.050 ;
        RECT 125.400 262.200 126.450 283.950 ;
        RECT 127.950 283.800 130.050 285.900 ;
        RECT 128.400 264.450 129.450 283.800 ;
        RECT 131.400 274.050 132.450 355.950 ;
        RECT 134.400 286.050 135.450 368.400 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 148.950 367.950 151.050 370.050 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 146.400 366.900 147.600 367.650 ;
        RECT 145.950 364.800 148.050 366.900 ;
        RECT 152.400 365.400 153.600 367.650 ;
        RECT 152.400 349.050 153.450 365.400 ;
        RECT 154.950 361.950 157.050 364.050 ;
        RECT 145.950 346.950 148.050 349.050 ;
        RECT 151.950 346.950 154.050 349.050 ;
        RECT 136.950 339.600 141.000 340.050 ;
        RECT 146.400 339.600 147.450 346.950 ;
        RECT 151.950 343.800 154.050 345.900 ;
        RECT 152.400 340.050 153.450 343.800 ;
        RECT 136.950 337.950 141.600 339.600 ;
        RECT 140.400 337.350 141.600 337.950 ;
        RECT 146.400 337.350 147.600 339.600 ;
        RECT 151.950 337.950 154.050 340.050 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 136.950 331.950 139.050 334.050 ;
        RECT 143.400 333.900 144.600 334.650 ;
        RECT 149.400 333.900 150.600 334.650 ;
        RECT 137.400 295.050 138.450 331.950 ;
        RECT 142.950 328.950 145.050 333.900 ;
        RECT 148.950 331.800 151.050 333.900 ;
        RECT 151.950 328.950 154.050 331.050 ;
        RECT 148.950 325.950 151.050 328.050 ;
        RECT 149.400 304.050 150.450 325.950 ;
        RECT 148.950 301.950 151.050 304.050 ;
        RECT 152.400 301.050 153.450 328.950 ;
        RECT 155.400 328.050 156.450 361.950 ;
        RECT 161.400 346.050 162.450 376.950 ;
        RECT 164.400 364.050 165.450 385.950 ;
        RECT 176.400 379.050 177.450 424.950 ;
        RECT 179.400 418.200 180.450 511.950 ;
        RECT 182.400 504.450 183.450 520.950 ;
        RECT 185.400 507.450 186.450 521.400 ;
        RECT 190.950 520.800 193.050 522.900 ;
        RECT 196.950 520.950 199.050 523.050 ;
        RECT 185.400 506.400 189.450 507.450 ;
        RECT 182.400 503.400 186.450 504.450 ;
        RECT 181.950 499.950 184.050 502.050 ;
        RECT 182.400 475.050 183.450 499.950 ;
        RECT 181.950 472.950 184.050 475.050 ;
        RECT 181.950 463.950 184.050 466.050 ;
        RECT 182.400 454.050 183.450 463.950 ;
        RECT 185.400 460.050 186.450 503.400 ;
        RECT 188.400 496.050 189.450 506.400 ;
        RECT 197.400 499.050 198.450 520.950 ;
        RECT 200.400 520.050 201.450 538.950 ;
        RECT 203.400 529.050 204.450 566.400 ;
        RECT 208.950 565.800 211.050 567.900 ;
        RECT 211.950 565.950 214.050 568.050 ;
        RECT 205.950 562.950 208.050 565.050 ;
        RECT 206.400 553.050 207.450 562.950 ;
        RECT 208.950 562.650 211.050 564.750 ;
        RECT 205.950 550.950 208.050 553.050 ;
        RECT 209.400 550.050 210.450 562.650 ;
        RECT 208.950 547.950 211.050 550.050 ;
        RECT 202.950 526.950 205.050 529.050 ;
        RECT 208.950 527.100 211.050 529.200 ;
        RECT 212.400 529.050 213.450 565.950 ;
        RECT 215.400 559.050 216.450 577.950 ;
        RECT 218.400 571.050 219.450 598.950 ;
        RECT 221.400 577.200 222.450 610.950 ;
        RECT 224.400 580.050 225.450 625.950 ;
        RECT 227.400 619.050 228.450 644.400 ;
        RECT 226.950 616.950 229.050 619.050 ;
        RECT 230.400 613.050 231.450 652.950 ;
        RECT 233.400 636.450 234.450 661.950 ;
        RECT 236.400 658.050 237.450 661.950 ;
        RECT 235.950 655.950 238.050 658.050 ;
        RECT 245.400 655.050 246.450 664.950 ;
        RECT 250.950 658.950 253.050 661.050 ;
        RECT 238.950 650.100 241.050 652.200 ;
        RECT 244.950 651.000 247.050 655.050 ;
        RECT 251.400 652.050 252.450 658.950 ;
        RECT 239.400 649.350 240.600 650.100 ;
        RECT 245.400 649.350 246.600 651.000 ;
        RECT 250.950 649.950 253.050 652.050 ;
        RECT 254.400 649.050 255.450 664.950 ;
        RECT 263.400 663.450 264.450 679.950 ;
        RECT 266.400 676.050 267.450 680.400 ;
        RECT 265.950 673.950 268.050 676.050 ;
        RECT 269.400 664.050 270.450 694.950 ;
        RECT 274.800 682.950 276.900 685.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 275.400 680.400 276.600 682.650 ;
        RECT 272.400 673.050 273.450 679.950 ;
        RECT 271.950 670.950 274.050 673.050 ;
        RECT 275.400 667.050 276.450 680.400 ;
        RECT 274.950 664.950 277.050 667.050 ;
        RECT 278.400 664.050 279.450 712.950 ;
        RECT 280.950 688.950 283.050 691.050 ;
        RECT 281.400 679.050 282.450 688.950 ;
        RECT 280.950 676.950 283.050 679.050 ;
        RECT 284.400 673.050 285.450 716.400 ;
        RECT 302.400 714.450 303.450 722.400 ;
        RECT 305.400 718.050 306.450 728.100 ;
        RECT 314.400 727.350 315.600 729.600 ;
        RECT 320.400 727.350 321.600 729.600 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 317.400 723.900 318.600 724.650 ;
        RECT 323.400 723.900 324.600 724.650 ;
        RECT 307.950 721.800 310.050 723.900 ;
        RECT 316.950 721.800 319.050 723.900 ;
        RECT 322.950 721.800 325.050 723.900 ;
        RECT 304.950 715.950 307.050 718.050 ;
        RECT 308.400 715.050 309.450 721.800 ;
        RECT 325.950 718.950 328.050 721.050 ;
        RECT 326.400 715.050 327.450 718.950 ;
        RECT 307.950 714.450 310.050 715.050 ;
        RECT 302.400 713.400 310.050 714.450 ;
        RECT 307.950 712.950 310.050 713.400 ;
        RECT 325.950 712.950 328.050 715.050 ;
        RECT 329.400 712.050 330.450 739.950 ;
        RECT 335.400 733.050 336.450 761.100 ;
        RECT 338.400 760.050 339.450 823.950 ;
        RECT 377.400 823.050 378.450 832.800 ;
        RECT 383.400 826.050 384.450 844.950 ;
        RECT 389.400 841.200 390.450 883.950 ;
        RECT 395.400 879.450 396.450 884.100 ;
        RECT 398.100 880.950 400.200 883.050 ;
        RECT 403.500 880.950 405.600 883.050 ;
        RECT 398.400 879.450 399.600 880.650 ;
        RECT 395.400 878.400 399.600 879.450 ;
        RECT 388.950 839.100 391.050 841.200 ;
        RECT 394.950 840.000 397.050 844.050 ;
        RECT 403.950 841.950 406.050 844.050 ;
        RECT 389.400 838.350 390.600 839.100 ;
        RECT 395.400 838.350 396.600 840.000 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 394.950 835.950 397.050 838.050 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 392.400 834.900 393.600 835.650 ;
        RECT 391.950 832.800 394.050 834.900 ;
        RECT 398.400 833.400 399.600 835.650 ;
        RECT 382.950 823.950 385.050 826.050 ;
        RECT 376.950 820.950 379.050 823.050 ;
        RECT 373.950 814.950 376.050 817.050 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 349.950 806.100 352.050 808.200 ;
        RECT 355.950 806.100 358.050 808.200 ;
        RECT 364.950 806.100 367.050 808.200 ;
        RECT 374.400 807.600 375.450 814.950 ;
        RECT 398.400 814.050 399.450 833.400 ;
        RECT 400.950 832.950 403.050 835.050 ;
        RECT 385.950 811.950 388.050 814.050 ;
        RECT 397.950 811.950 400.050 814.050 ;
        RECT 381.000 807.600 385.050 808.050 ;
        RECT 341.400 801.900 342.450 805.950 ;
        RECT 350.400 805.350 351.600 806.100 ;
        RECT 356.400 805.350 357.600 806.100 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 347.400 801.900 348.600 802.650 ;
        RECT 340.950 799.800 343.050 801.900 ;
        RECT 346.950 799.800 349.050 801.900 ;
        RECT 353.400 800.400 354.600 802.650 ;
        RECT 359.400 800.400 360.600 802.650 ;
        RECT 353.400 790.050 354.450 800.400 ;
        RECT 352.950 787.950 355.050 790.050 ;
        RECT 349.950 766.950 352.050 769.050 ;
        RECT 340.950 762.600 345.000 763.050 ;
        RECT 350.400 762.600 351.450 766.950 ;
        RECT 340.950 760.950 345.600 762.600 ;
        RECT 344.400 760.350 345.600 760.950 ;
        RECT 350.400 760.350 351.600 762.600 ;
        RECT 355.950 761.100 358.050 763.200 ;
        RECT 359.400 763.050 360.450 800.400 ;
        RECT 361.950 799.950 364.050 802.050 ;
        RECT 362.400 769.050 363.450 799.950 ;
        RECT 365.400 784.050 366.450 806.100 ;
        RECT 374.400 805.350 375.600 807.600 ;
        RECT 380.400 805.950 385.050 807.600 ;
        RECT 380.400 805.350 381.600 805.950 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 371.400 801.900 372.600 802.650 ;
        RECT 370.950 801.450 373.050 801.900 ;
        RECT 368.400 800.400 373.050 801.450 ;
        RECT 377.400 801.000 378.600 802.650 ;
        RECT 368.400 793.050 369.450 800.400 ;
        RECT 370.950 799.800 373.050 800.400 ;
        RECT 376.950 796.950 379.050 801.000 ;
        RECT 386.400 799.050 387.450 811.950 ;
        RECT 401.400 810.450 402.450 832.950 ;
        RECT 404.400 832.050 405.450 841.950 ;
        RECT 406.950 839.100 409.050 841.200 ;
        RECT 410.400 841.050 411.450 895.950 ;
        RECT 413.400 895.050 414.450 908.400 ;
        RECT 416.400 907.050 417.450 911.400 ;
        RECT 421.950 910.950 424.050 913.050 ;
        RECT 425.400 907.050 426.450 917.100 ;
        RECT 431.400 916.350 432.600 917.100 ;
        RECT 437.400 916.350 438.600 917.100 ;
        RECT 430.950 913.950 433.050 916.050 ;
        RECT 433.950 913.950 436.050 916.050 ;
        RECT 436.950 913.950 439.050 916.050 ;
        RECT 439.950 913.950 442.050 916.050 ;
        RECT 434.400 912.900 435.600 913.650 ;
        RECT 433.950 910.800 436.050 912.900 ;
        RECT 440.400 911.400 441.600 913.650 ;
        RECT 440.400 910.050 441.450 911.400 ;
        RECT 442.950 910.950 445.050 913.050 ;
        RECT 439.950 907.950 442.050 910.050 ;
        RECT 415.950 904.950 418.050 907.050 ;
        RECT 424.950 904.950 427.050 907.050 ;
        RECT 430.950 904.950 433.050 907.050 ;
        RECT 436.950 904.950 439.050 907.050 ;
        RECT 415.950 895.950 418.050 898.050 ;
        RECT 412.950 892.950 415.050 895.050 ;
        RECT 416.400 892.050 417.450 895.950 ;
        RECT 415.950 889.950 418.050 892.050 ;
        RECT 415.950 885.000 418.050 888.900 ;
        RECT 416.400 883.350 417.600 885.000 ;
        RECT 421.950 884.100 424.050 886.200 ;
        RECT 422.400 883.350 423.600 884.100 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 421.950 880.950 424.050 883.050 ;
        RECT 424.950 880.950 427.050 883.050 ;
        RECT 419.400 878.400 420.600 880.650 ;
        RECT 425.400 879.000 426.600 880.650 ;
        RECT 419.400 877.050 420.450 878.400 ;
        RECT 418.950 874.950 421.050 877.050 ;
        RECT 424.950 874.950 427.050 879.000 ;
        RECT 419.400 849.450 420.450 874.950 ;
        RECT 431.400 874.050 432.450 904.950 ;
        RECT 437.400 880.050 438.450 904.950 ;
        RECT 440.400 892.050 441.450 907.950 ;
        RECT 443.400 907.050 444.450 910.950 ;
        RECT 442.950 904.950 445.050 907.050 ;
        RECT 446.400 895.050 447.450 917.100 ;
        RECT 448.950 916.950 453.600 918.600 ;
        RECT 457.950 917.100 460.050 919.200 ;
        RECT 452.400 916.350 453.600 916.950 ;
        RECT 458.400 916.350 459.600 917.100 ;
        RECT 451.950 913.950 454.050 916.050 ;
        RECT 454.950 913.950 457.050 916.050 ;
        RECT 457.950 913.950 460.050 916.050 ;
        RECT 455.400 912.900 456.600 913.650 ;
        RECT 454.950 910.800 457.050 912.900 ;
        RECT 464.400 904.050 465.450 928.950 ;
        RECT 472.950 922.950 475.050 925.050 ;
        RECT 496.950 922.950 499.050 925.050 ;
        RECT 473.400 918.600 474.450 922.950 ;
        RECT 497.400 919.200 498.450 922.950 ;
        RECT 473.400 916.350 474.600 918.600 ;
        RECT 478.950 917.100 481.050 919.200 ;
        RECT 484.950 917.100 487.050 919.200 ;
        RECT 496.950 917.100 499.050 919.200 ;
        RECT 503.400 918.600 504.450 928.950 ;
        RECT 479.400 916.350 480.600 917.100 ;
        RECT 469.950 913.950 472.050 916.050 ;
        RECT 472.950 913.950 475.050 916.050 ;
        RECT 475.950 913.950 478.050 916.050 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 470.400 912.000 471.600 913.650 ;
        RECT 469.950 907.950 472.050 912.000 ;
        RECT 476.400 911.400 477.600 913.650 ;
        RECT 476.400 904.050 477.450 911.400 ;
        RECT 478.950 907.950 481.050 910.050 ;
        RECT 463.950 901.950 466.050 904.050 ;
        RECT 475.950 901.950 478.050 904.050 ;
        RECT 445.950 892.950 448.050 895.050 ;
        RECT 469.950 892.950 472.050 895.050 ;
        RECT 439.950 889.950 442.050 892.050 ;
        RECT 470.400 889.050 471.450 892.950 ;
        RECT 475.950 889.950 478.050 892.050 ;
        RECT 439.950 884.100 442.050 886.200 ;
        RECT 448.950 884.100 451.050 886.200 ;
        RECT 454.950 884.100 457.050 886.200 ;
        RECT 469.950 885.000 472.050 889.050 ;
        RECT 440.400 883.350 441.600 884.100 ;
        RECT 449.400 883.350 450.600 884.100 ;
        RECT 440.100 880.950 442.200 883.050 ;
        RECT 443.100 880.950 445.200 883.050 ;
        RECT 448.800 880.950 450.900 883.050 ;
        RECT 451.800 880.950 453.900 883.050 ;
        RECT 436.950 877.950 439.050 880.050 ;
        RECT 443.400 879.900 444.600 880.650 ;
        RECT 442.950 877.800 445.050 879.900 ;
        RECT 452.400 878.400 453.600 880.650 ;
        RECT 452.400 876.450 453.450 878.400 ;
        RECT 455.400 877.050 456.450 884.100 ;
        RECT 470.400 883.350 471.600 885.000 ;
        RECT 466.950 880.950 469.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 467.400 879.000 468.600 880.650 ;
        RECT 449.400 875.400 453.450 876.450 ;
        RECT 449.400 874.050 450.450 875.400 ;
        RECT 454.950 874.950 457.050 877.050 ;
        RECT 466.950 874.950 469.050 879.000 ;
        RECT 430.950 871.950 433.050 874.050 ;
        RECT 448.950 871.950 451.050 874.050 ;
        RECT 436.950 859.950 439.050 862.050 ;
        RECT 427.950 853.950 430.050 856.050 ;
        RECT 421.950 849.450 424.050 850.050 ;
        RECT 419.400 848.400 424.050 849.450 ;
        RECT 421.950 847.950 424.050 848.400 ;
        RECT 407.400 834.450 408.450 839.100 ;
        RECT 409.950 838.950 412.050 841.050 ;
        RECT 415.950 839.100 418.050 841.200 ;
        RECT 422.400 840.600 423.450 847.950 ;
        RECT 416.400 838.350 417.600 839.100 ;
        RECT 422.400 838.350 423.600 840.600 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 415.950 835.950 418.050 838.050 ;
        RECT 418.950 835.950 421.050 838.050 ;
        RECT 421.950 835.950 424.050 838.050 ;
        RECT 409.950 834.450 412.050 834.900 ;
        RECT 407.400 833.400 412.050 834.450 ;
        RECT 409.950 832.800 412.050 833.400 ;
        RECT 413.400 833.400 414.600 835.650 ;
        RECT 419.400 834.000 420.600 835.650 ;
        RECT 403.950 829.950 406.050 832.050 ;
        RECT 406.950 823.950 409.050 826.050 ;
        RECT 401.400 809.400 405.450 810.450 ;
        RECT 388.950 805.950 391.050 808.050 ;
        RECT 397.950 806.100 400.050 808.200 ;
        RECT 404.400 807.600 405.450 809.400 ;
        RECT 407.400 808.050 408.450 823.950 ;
        RECT 389.400 801.900 390.450 805.950 ;
        RECT 398.400 805.350 399.600 806.100 ;
        RECT 404.400 805.350 405.600 807.600 ;
        RECT 406.950 805.950 409.050 808.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 395.400 801.900 396.600 802.650 ;
        RECT 388.950 799.800 391.050 801.900 ;
        RECT 394.950 799.800 397.050 801.900 ;
        RECT 401.400 800.400 402.600 802.650 ;
        RECT 385.950 796.950 388.050 799.050 ;
        RECT 367.950 790.950 370.050 793.050 ;
        RECT 370.950 787.950 373.050 790.050 ;
        RECT 367.950 784.950 370.050 787.050 ;
        RECT 364.950 781.950 367.050 784.050 ;
        RECT 361.950 766.950 364.050 769.050 ;
        RECT 368.400 763.200 369.450 784.950 ;
        RECT 371.400 781.050 372.450 787.950 ;
        RECT 385.950 784.950 388.050 787.050 ;
        RECT 373.950 781.950 376.050 784.050 ;
        RECT 370.950 778.950 373.050 781.050 ;
        RECT 374.400 775.050 375.450 781.950 ;
        RECT 376.950 778.950 379.050 781.050 ;
        RECT 373.950 772.950 376.050 775.050 ;
        RECT 377.400 771.450 378.450 778.950 ;
        RECT 379.950 775.950 382.050 778.050 ;
        RECT 374.400 770.400 378.450 771.450 ;
        RECT 358.950 762.450 361.050 763.050 ;
        RECT 358.950 761.400 363.450 762.450 ;
        RECT 356.400 760.350 357.600 761.100 ;
        RECT 358.950 760.950 361.050 761.400 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 346.950 757.950 349.050 760.050 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 347.400 756.900 348.600 757.650 ;
        RECT 337.950 754.800 340.050 756.900 ;
        RECT 346.950 754.800 349.050 756.900 ;
        RECT 353.400 755.400 354.600 757.650 ;
        RECT 334.950 730.950 337.050 733.050 ;
        RECT 338.400 729.600 339.450 754.800 ;
        RECT 346.950 751.650 349.050 753.750 ;
        RECT 338.400 727.350 339.600 729.600 ;
        RECT 334.950 724.950 337.050 727.050 ;
        RECT 337.950 724.950 340.050 727.050 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 335.400 723.000 336.600 724.650 ;
        RECT 334.950 718.950 337.050 723.000 ;
        RECT 341.400 722.400 342.600 724.650 ;
        RECT 331.950 715.950 334.050 718.050 ;
        RECT 328.950 709.950 331.050 712.050 ;
        RECT 316.950 706.950 319.050 709.050 ;
        RECT 289.950 703.950 292.050 706.050 ;
        RECT 313.950 703.950 316.050 706.050 ;
        RECT 290.400 684.600 291.450 703.950 ;
        RECT 301.950 697.950 304.050 700.050 ;
        RECT 310.950 697.950 313.050 700.050 ;
        RECT 290.400 682.350 291.600 684.600 ;
        RECT 295.800 683.100 297.900 685.200 ;
        RECT 296.400 682.350 297.600 683.100 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 293.400 678.900 294.600 679.650 ;
        RECT 292.950 676.800 295.050 678.900 ;
        RECT 302.400 678.450 303.450 697.950 ;
        RECT 311.400 694.050 312.450 697.950 ;
        RECT 310.950 691.950 313.050 694.050 ;
        RECT 307.950 688.950 310.050 691.050 ;
        RECT 308.400 684.600 309.450 688.950 ;
        RECT 314.400 684.600 315.450 703.950 ;
        RECT 317.400 703.050 318.450 706.950 ;
        RECT 316.950 700.950 319.050 703.050 ;
        RECT 322.950 700.950 325.050 703.050 ;
        RECT 323.400 694.050 324.450 700.950 ;
        RECT 325.950 694.950 328.050 697.050 ;
        RECT 322.950 691.950 325.050 694.050 ;
        RECT 326.400 688.050 327.450 694.950 ;
        RECT 319.950 687.600 324.000 688.050 ;
        RECT 319.950 685.950 324.600 687.600 ;
        RECT 325.950 685.950 328.050 688.050 ;
        RECT 323.400 685.350 324.600 685.950 ;
        RECT 308.400 682.350 309.600 684.600 ;
        RECT 314.400 682.350 315.600 684.600 ;
        RECT 322.800 682.950 324.900 685.050 ;
        RECT 328.800 682.950 330.900 685.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 311.400 678.900 312.600 679.650 ;
        RECT 302.400 677.400 306.450 678.450 ;
        RECT 295.950 675.450 298.050 676.050 ;
        RECT 305.400 675.450 306.450 677.400 ;
        RECT 310.950 676.800 313.050 678.900 ;
        RECT 317.400 678.450 318.600 679.650 ;
        RECT 317.400 677.400 321.450 678.450 ;
        RECT 295.950 674.400 303.450 675.450 ;
        RECT 305.400 674.400 309.450 675.450 ;
        RECT 295.950 673.950 298.050 674.400 ;
        RECT 283.950 670.950 286.050 673.050 ;
        RECT 298.950 670.950 301.050 673.050 ;
        RECT 260.400 662.400 264.450 663.450 ;
        RECT 260.400 652.050 261.450 662.400 ;
        RECT 268.950 661.950 271.050 664.050 ;
        RECT 277.950 661.950 280.050 664.050 ;
        RECT 295.950 661.950 298.050 664.050 ;
        RECT 263.700 657.300 265.800 659.400 ;
        RECT 266.700 657.300 268.800 659.400 ;
        RECT 269.700 657.300 271.800 659.400 ;
        RECT 264.300 653.700 265.500 657.300 ;
        RECT 259.950 649.950 262.050 652.050 ;
        RECT 263.400 651.600 265.500 653.700 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 241.950 646.950 244.050 649.050 ;
        RECT 244.950 646.950 247.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 242.400 644.400 243.600 646.650 ;
        RECT 235.950 636.450 238.050 637.050 ;
        RECT 233.400 635.400 238.050 636.450 ;
        RECT 235.950 634.950 238.050 635.400 ;
        RECT 229.950 610.950 232.050 613.050 ;
        RECT 226.950 605.100 229.050 607.200 ;
        RECT 227.400 604.350 228.600 605.100 ;
        RECT 227.100 601.950 229.200 604.050 ;
        RECT 232.500 601.950 234.600 604.050 ;
        RECT 233.400 599.400 234.600 601.650 ;
        RECT 233.400 595.050 234.450 599.400 ;
        RECT 236.400 598.050 237.450 634.950 ;
        RECT 242.400 622.050 243.450 644.400 ;
        RECT 250.800 643.950 252.900 646.050 ;
        RECT 256.800 643.950 258.900 646.050 ;
        RECT 251.400 641.400 252.600 643.650 ;
        RECT 251.400 637.050 252.450 641.400 ;
        RECT 253.950 640.950 256.050 643.050 ;
        RECT 250.950 634.950 253.050 637.050 ;
        RECT 254.400 633.450 255.450 640.950 ;
        RECT 251.400 632.400 255.450 633.450 ;
        RECT 263.400 632.700 264.900 651.600 ;
        RECT 267.300 640.800 268.500 657.300 ;
        RECT 266.400 638.700 268.500 640.800 ;
        RECT 267.300 632.700 268.500 638.700 ;
        RECT 269.700 635.700 270.900 657.300 ;
        RECT 277.800 656.400 279.900 658.500 ;
        RECT 283.200 657.300 285.300 659.400 ;
        RECT 286.200 657.300 288.300 659.400 ;
        RECT 289.200 657.300 291.300 659.400 ;
        RECT 274.800 649.950 276.900 652.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 275.400 647.400 276.600 649.650 ;
        RECT 272.400 643.050 273.450 646.950 ;
        RECT 271.950 640.950 274.050 643.050 ;
        RECT 269.700 633.600 271.800 635.700 ;
        RECT 241.950 619.950 244.050 622.050 ;
        RECT 244.950 610.950 247.050 613.050 ;
        RECT 245.400 607.200 246.450 610.950 ;
        RECT 251.400 607.200 252.450 632.400 ;
        RECT 263.400 630.600 266.400 632.700 ;
        RECT 267.300 630.600 269.400 632.700 ;
        RECT 271.950 610.950 274.050 613.050 ;
        RECT 244.950 605.100 247.050 607.200 ;
        RECT 250.950 605.100 253.050 607.200 ;
        RECT 259.950 605.100 262.050 607.200 ;
        RECT 265.950 605.100 268.050 607.200 ;
        RECT 272.400 606.600 273.450 610.950 ;
        RECT 275.400 610.050 276.450 647.400 ;
        RECT 278.400 645.900 279.300 656.400 ;
        RECT 281.100 650.400 283.200 652.500 ;
        RECT 278.400 643.800 280.500 645.900 ;
        RECT 284.100 645.000 285.300 657.300 ;
        RECT 278.400 637.200 279.300 643.800 ;
        RECT 283.800 642.900 285.900 645.000 ;
        RECT 278.400 635.100 280.500 637.200 ;
        RECT 284.100 635.700 285.300 642.900 ;
        RECT 286.800 639.600 288.300 657.300 ;
        RECT 286.800 637.500 288.900 639.600 ;
        RECT 283.800 633.600 285.900 635.700 ;
        RECT 286.800 632.700 288.300 637.500 ;
        RECT 290.100 635.700 291.300 657.300 ;
        RECT 286.200 630.600 288.300 632.700 ;
        RECT 289.200 630.600 291.300 635.700 ;
        RECT 292.200 657.300 294.300 659.400 ;
        RECT 292.200 639.600 293.700 657.300 ;
        RECT 292.200 637.500 294.300 639.600 ;
        RECT 292.200 632.700 293.700 637.500 ;
        RECT 292.200 630.600 294.300 632.700 ;
        RECT 280.950 616.950 283.050 619.050 ;
        RECT 274.950 607.950 277.050 610.050 ;
        RECT 245.400 604.350 246.600 605.100 ;
        RECT 251.400 604.350 252.600 605.100 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 250.950 601.950 253.050 604.050 ;
        RECT 248.400 599.400 249.600 601.650 ;
        RECT 248.400 598.050 249.450 599.400 ;
        RECT 253.950 598.950 256.050 601.050 ;
        RECT 235.950 595.950 238.050 598.050 ;
        RECT 248.400 596.400 253.050 598.050 ;
        RECT 249.000 595.950 253.050 596.400 ;
        RECT 232.950 592.950 235.050 595.050 ;
        RECT 223.950 577.950 226.050 580.050 ;
        RECT 220.950 575.100 223.050 577.200 ;
        RECT 220.950 571.950 223.050 574.050 ;
        RECT 221.400 571.350 222.600 571.950 ;
        RECT 236.400 571.050 237.450 595.950 ;
        RECT 241.950 592.950 244.050 595.050 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 221.400 568.950 223.500 571.050 ;
        RECT 226.800 568.950 228.900 571.050 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 227.400 567.900 228.600 568.650 ;
        RECT 217.950 565.800 220.050 567.900 ;
        RECT 214.950 556.950 217.050 559.050 ;
        RECT 218.400 556.050 219.450 565.800 ;
        RECT 220.950 562.950 223.050 565.050 ;
        RECT 217.950 553.950 220.050 556.050 ;
        RECT 221.400 552.450 222.450 562.950 ;
        RECT 226.950 562.800 229.050 567.900 ;
        RECT 232.800 565.950 234.900 568.050 ;
        RECT 238.800 565.950 240.900 568.050 ;
        RECT 233.400 564.900 234.600 565.650 ;
        RECT 232.950 562.800 235.050 564.900 ;
        RECT 223.950 559.950 226.050 562.050 ;
        RECT 218.400 552.000 222.450 552.450 ;
        RECT 218.400 551.400 223.050 552.000 ;
        RECT 214.950 547.950 217.050 550.050 ;
        RECT 209.400 526.350 210.600 527.100 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 202.950 520.950 205.050 523.050 ;
        RECT 206.400 521.400 207.600 523.650 ;
        RECT 199.950 517.950 202.050 520.050 ;
        RECT 199.950 511.950 202.050 514.050 ;
        RECT 196.950 496.950 199.050 499.050 ;
        RECT 187.950 493.950 190.050 496.050 ;
        RECT 190.950 495.600 195.000 496.050 ;
        RECT 200.400 495.600 201.450 511.950 ;
        RECT 203.400 507.450 204.450 520.950 ;
        RECT 206.400 511.050 207.450 521.400 ;
        RECT 211.950 520.950 214.050 523.050 ;
        RECT 208.950 517.950 211.050 520.050 ;
        RECT 205.950 508.950 208.050 511.050 ;
        RECT 203.400 506.400 207.450 507.450 ;
        RECT 206.400 496.050 207.450 506.400 ;
        RECT 190.950 493.950 195.600 495.600 ;
        RECT 194.400 493.350 195.600 493.950 ;
        RECT 200.400 493.350 201.600 495.600 ;
        RECT 205.950 493.950 208.050 496.050 ;
        RECT 187.950 490.800 190.050 492.900 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 188.400 486.450 189.450 490.800 ;
        RECT 197.400 489.900 198.600 490.650 ;
        RECT 196.950 487.800 199.050 489.900 ;
        RECT 203.400 489.000 204.600 490.650 ;
        RECT 188.400 485.400 192.450 486.450 ;
        RECT 187.950 472.950 190.050 475.050 ;
        RECT 184.950 457.950 187.050 460.050 ;
        RECT 181.950 451.950 184.050 454.050 ;
        RECT 184.800 448.950 186.900 451.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 185.400 446.400 186.600 448.650 ;
        RECT 178.950 416.100 181.050 418.200 ;
        RECT 182.400 418.050 183.450 445.950 ;
        RECT 185.400 433.050 186.450 446.400 ;
        RECT 184.950 430.950 187.050 433.050 ;
        RECT 188.400 427.050 189.450 472.950 ;
        RECT 191.400 454.050 192.450 485.400 ;
        RECT 193.950 484.950 196.050 487.050 ;
        RECT 194.400 466.050 195.450 484.950 ;
        RECT 193.950 463.950 196.050 466.050 ;
        RECT 197.400 463.050 198.450 487.800 ;
        RECT 199.950 484.950 202.050 487.050 ;
        RECT 202.950 484.950 205.050 489.000 ;
        RECT 205.950 484.950 208.050 490.050 ;
        RECT 200.400 478.050 201.450 484.950 ;
        RECT 199.950 475.950 202.050 478.050 ;
        RECT 196.950 460.950 199.050 463.050 ;
        RECT 190.950 451.950 193.050 454.050 ;
        RECT 196.950 451.950 199.050 454.050 ;
        RECT 193.800 448.950 195.900 451.050 ;
        RECT 194.400 446.400 195.600 448.650 ;
        RECT 194.400 442.050 195.450 446.400 ;
        RECT 193.950 439.950 196.050 442.050 ;
        RECT 187.950 424.950 190.050 427.050 ;
        RECT 175.950 376.950 178.050 379.050 ;
        RECT 172.950 371.100 175.050 373.200 ;
        RECT 173.400 370.350 174.600 371.100 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 166.800 364.950 168.900 367.050 ;
        RECT 170.400 366.900 171.600 367.650 ;
        RECT 163.950 361.950 166.050 364.050 ;
        RECT 167.400 355.050 168.450 364.950 ;
        RECT 169.950 364.800 172.050 366.900 ;
        RECT 175.950 364.950 178.050 367.050 ;
        RECT 166.950 352.950 169.050 355.050 ;
        RECT 166.950 346.950 169.050 349.050 ;
        RECT 160.950 343.950 163.050 346.050 ;
        RECT 167.400 340.200 168.450 346.950 ;
        RECT 176.400 345.450 177.450 364.950 ;
        RECT 173.400 344.400 177.450 345.450 ;
        RECT 160.950 338.100 163.050 340.200 ;
        RECT 166.950 338.100 169.050 340.200 ;
        RECT 173.400 340.050 174.450 344.400 ;
        RECT 175.950 340.950 178.050 343.050 ;
        RECT 161.400 337.350 162.600 338.100 ;
        RECT 167.400 337.350 168.600 338.100 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 164.400 333.900 165.600 334.650 ;
        RECT 157.950 328.950 160.050 333.900 ;
        RECT 163.950 331.800 166.050 333.900 ;
        RECT 170.400 332.400 171.600 334.650 ;
        RECT 154.950 325.950 157.050 328.050 ;
        RECT 170.400 325.050 171.450 332.400 ;
        RECT 172.950 331.950 175.050 334.050 ;
        RECT 169.950 322.950 172.050 325.050 ;
        RECT 173.400 307.050 174.450 331.950 ;
        RECT 163.950 304.950 166.050 307.050 ;
        RECT 172.950 304.950 175.050 307.050 ;
        RECT 160.950 301.950 163.050 304.050 ;
        RECT 139.950 298.950 142.050 301.050 ;
        RECT 151.950 298.950 154.050 301.050 ;
        RECT 136.950 292.950 139.050 295.050 ;
        RECT 140.400 294.600 141.450 298.950 ;
        RECT 140.400 292.350 141.600 294.600 ;
        RECT 145.950 294.000 148.050 298.050 ;
        RECT 146.400 292.350 147.600 294.000 ;
        RECT 151.950 293.100 154.050 295.200 ;
        RECT 157.950 293.100 160.050 295.200 ;
        RECT 152.400 292.350 153.600 293.100 ;
        RECT 139.950 289.950 142.050 292.050 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 143.400 288.000 144.600 289.650 ;
        RECT 149.400 288.900 150.600 289.650 ;
        RECT 133.950 283.950 136.050 286.050 ;
        RECT 139.950 283.950 142.050 286.050 ;
        RECT 142.950 283.950 145.050 288.000 ;
        RECT 148.950 286.800 151.050 288.900 ;
        RECT 130.950 271.950 133.050 274.050 ;
        RECT 128.400 263.400 132.450 264.450 ;
        RECT 107.400 259.350 108.600 261.600 ;
        RECT 115.950 259.950 118.050 262.050 ;
        RECT 124.950 260.100 127.050 262.200 ;
        RECT 131.400 261.600 132.450 263.400 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 104.400 255.900 105.600 256.650 ;
        RECT 103.950 253.800 106.050 255.900 ;
        RECT 110.400 255.450 111.600 256.650 ;
        RECT 110.400 254.400 114.450 255.450 ;
        RECT 97.950 247.950 100.050 250.050 ;
        RECT 113.400 247.050 114.450 254.400 ;
        RECT 106.950 244.950 109.050 247.050 ;
        RECT 112.950 244.950 115.050 247.050 ;
        RECT 97.950 238.950 100.050 241.050 ;
        RECT 94.950 220.950 97.050 223.050 ;
        RECT 98.400 220.050 99.450 238.950 ;
        RECT 97.950 217.950 100.050 220.050 ;
        RECT 83.400 214.350 84.600 216.600 ;
        RECT 88.950 214.950 91.050 217.050 ;
        RECT 92.100 214.950 94.200 217.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 92.400 213.000 93.600 214.650 ;
        RECT 73.950 208.950 76.050 211.050 ;
        RECT 86.400 210.900 87.600 211.650 ;
        RECT 85.950 208.800 88.050 210.900 ;
        RECT 91.950 208.950 94.050 213.000 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 98.400 213.450 99.450 217.950 ;
        RECT 101.100 214.950 103.200 217.050 ;
        RECT 101.400 213.450 102.600 214.650 ;
        RECT 98.400 212.400 102.600 213.450 ;
        RECT 70.950 193.950 73.050 196.050 ;
        RECT 82.950 190.950 85.050 193.050 ;
        RECT 64.950 187.950 67.050 190.050 ;
        RECT 52.950 178.950 55.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 49.950 175.950 52.050 178.050 ;
        RECT 53.400 177.000 54.600 178.650 ;
        RECT 50.400 169.050 51.450 175.950 ;
        RECT 52.950 172.950 55.050 177.000 ;
        RECT 58.950 175.950 61.050 178.050 ;
        RECT 65.400 177.450 66.450 187.950 ;
        RECT 70.950 183.000 73.050 187.050 ;
        RECT 71.400 181.350 72.600 183.000 ;
        RECT 76.950 182.100 79.050 184.200 ;
        RECT 83.400 184.050 84.450 190.950 ;
        RECT 77.400 181.350 78.600 182.100 ;
        RECT 82.950 181.950 85.050 184.050 ;
        RECT 70.950 178.950 73.050 181.050 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 74.400 177.900 75.600 178.650 ;
        RECT 62.400 177.000 66.450 177.450 ;
        RECT 61.950 176.400 66.450 177.000 ;
        RECT 49.950 166.950 52.050 169.050 ;
        RECT 50.400 163.050 51.450 166.950 ;
        RECT 49.950 160.950 52.050 163.050 ;
        RECT 59.400 151.050 60.450 175.950 ;
        RECT 61.950 175.050 64.050 176.400 ;
        RECT 73.950 175.800 76.050 177.900 ;
        RECT 80.400 177.000 81.600 178.650 ;
        RECT 61.800 174.000 64.050 175.050 ;
        RECT 61.800 172.950 63.900 174.000 ;
        RECT 64.950 172.950 67.050 175.050 ;
        RECT 79.950 172.950 82.050 177.000 ;
        RECT 82.950 172.950 85.050 177.900 ;
        RECT 58.950 148.950 61.050 151.050 ;
        RECT 58.950 137.100 61.050 139.200 ;
        RECT 65.400 139.050 66.450 172.950 ;
        RECT 59.400 136.350 60.600 137.100 ;
        RECT 64.950 136.950 67.050 139.050 ;
        RECT 67.950 137.100 70.050 139.200 ;
        RECT 76.950 137.100 79.050 139.200 ;
        RECT 82.950 137.100 85.050 139.200 ;
        RECT 86.400 138.450 87.450 208.800 ;
        RECT 95.400 199.050 96.450 211.950 ;
        RECT 94.950 196.950 97.050 199.050 ;
        RECT 103.950 187.950 106.050 193.050 ;
        RECT 89.400 186.000 99.450 186.450 ;
        RECT 88.950 185.400 99.450 186.000 ;
        RECT 88.950 181.950 91.050 185.400 ;
        RECT 91.950 182.100 94.050 184.200 ;
        RECT 98.400 183.600 99.450 185.400 ;
        RECT 92.400 181.350 93.600 182.100 ;
        RECT 98.400 181.350 99.600 183.600 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 88.950 175.950 91.050 178.050 ;
        RECT 95.400 176.400 96.600 178.650 ;
        RECT 101.400 176.400 102.600 178.650 ;
        RECT 89.400 169.050 90.450 175.950 ;
        RECT 95.400 169.050 96.450 176.400 ;
        RECT 97.950 172.950 100.050 175.050 ;
        RECT 88.950 166.950 91.050 169.050 ;
        RECT 94.950 166.950 97.050 169.050 ;
        RECT 86.400 137.400 90.450 138.450 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 49.950 130.950 52.050 133.050 ;
        RECT 56.400 132.000 57.600 133.650 ;
        RECT 50.400 64.050 51.450 130.950 ;
        RECT 55.950 127.950 58.050 132.000 ;
        RECT 62.400 131.400 63.600 133.650 ;
        RECT 62.400 124.050 63.450 131.400 ;
        RECT 64.950 127.950 67.050 133.050 ;
        RECT 68.400 127.050 69.450 137.100 ;
        RECT 77.400 136.350 78.600 137.100 ;
        RECT 83.400 136.350 84.600 137.100 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 74.400 132.900 75.600 133.650 ;
        RECT 73.950 130.800 76.050 132.900 ;
        RECT 80.400 132.000 81.600 133.650 ;
        RECT 67.950 124.950 70.050 127.050 ;
        RECT 61.950 121.950 64.050 124.050 ;
        RECT 52.950 118.950 55.050 121.050 ;
        RECT 53.400 106.200 54.450 118.950 ;
        RECT 74.400 106.200 75.450 130.800 ;
        RECT 79.950 127.950 82.050 132.000 ;
        RECT 85.950 130.950 88.050 133.050 ;
        RECT 86.400 112.050 87.450 130.950 ;
        RECT 79.950 109.950 82.050 112.050 ;
        RECT 85.950 109.950 88.050 112.050 ;
        RECT 52.950 104.100 55.050 106.200 ;
        RECT 61.950 104.100 64.050 106.200 ;
        RECT 67.950 104.100 70.050 106.200 ;
        RECT 73.950 104.100 76.050 106.200 ;
        RECT 80.400 105.600 81.450 109.950 ;
        RECT 62.400 103.350 63.600 104.100 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 59.400 98.400 60.600 100.650 ;
        RECT 59.400 94.050 60.450 98.400 ;
        RECT 68.400 94.050 69.450 104.100 ;
        RECT 74.400 103.350 75.600 104.100 ;
        RECT 80.400 103.350 81.600 105.600 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 76.950 100.950 79.050 103.050 ;
        RECT 79.950 100.950 82.050 103.050 ;
        RECT 77.400 99.900 78.600 100.650 ;
        RECT 76.950 97.800 79.050 99.900 ;
        RECT 89.400 99.450 90.450 137.400 ;
        RECT 91.950 137.100 94.050 139.200 ;
        RECT 98.400 138.600 99.450 172.950 ;
        RECT 101.400 172.050 102.450 176.400 ;
        RECT 107.400 175.050 108.450 244.950 ;
        RECT 116.400 235.050 117.450 259.950 ;
        RECT 125.400 259.350 126.600 260.100 ;
        RECT 131.400 259.350 132.600 261.600 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 133.950 256.950 136.050 259.050 ;
        RECT 122.400 254.400 123.600 256.650 ;
        RECT 128.400 254.400 129.600 256.650 ;
        RECT 134.400 254.400 135.600 256.650 ;
        RECT 115.950 232.950 118.050 235.050 ;
        RECT 122.400 232.050 123.450 254.400 ;
        RECT 110.700 228.300 112.800 230.400 ;
        RECT 111.300 223.500 112.800 228.300 ;
        RECT 110.700 221.400 112.800 223.500 ;
        RECT 111.300 203.700 112.800 221.400 ;
        RECT 110.700 201.600 112.800 203.700 ;
        RECT 113.700 225.300 115.800 230.400 ;
        RECT 116.700 228.300 118.800 230.400 ;
        RECT 121.950 229.950 124.050 232.050 ;
        RECT 113.700 203.700 114.900 225.300 ;
        RECT 116.700 223.500 118.200 228.300 ;
        RECT 119.100 225.300 121.200 227.400 ;
        RECT 116.100 221.400 118.200 223.500 ;
        RECT 116.700 203.700 118.200 221.400 ;
        RECT 119.700 218.100 120.900 225.300 ;
        RECT 124.500 223.800 126.600 225.900 ;
        RECT 119.100 216.000 121.200 218.100 ;
        RECT 125.700 217.200 126.600 223.800 ;
        RECT 119.700 203.700 120.900 216.000 ;
        RECT 124.500 215.100 126.600 217.200 ;
        RECT 121.800 208.500 123.900 210.600 ;
        RECT 125.700 204.600 126.600 215.100 ;
        RECT 128.400 213.600 129.450 254.400 ;
        RECT 134.400 244.050 135.450 254.400 ;
        RECT 136.950 253.950 139.050 256.050 ;
        RECT 140.400 255.450 141.450 283.950 ;
        RECT 158.400 283.050 159.450 293.100 ;
        RECT 142.950 280.800 145.050 282.900 ;
        RECT 157.950 280.950 160.050 283.050 ;
        RECT 143.400 262.050 144.450 280.800 ;
        RECT 145.950 274.950 148.050 277.050 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 146.400 261.600 147.450 274.950 ;
        RECT 146.400 259.350 147.600 261.600 ;
        RECT 151.950 260.100 154.050 262.200 ;
        RECT 152.400 259.350 153.600 260.100 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 140.400 254.400 144.450 255.450 ;
        RECT 137.400 250.050 138.450 253.950 ;
        RECT 136.950 247.950 139.050 250.050 ;
        RECT 133.950 241.950 136.050 244.050 ;
        RECT 135.600 228.300 137.700 230.400 ;
        RECT 138.600 228.300 141.600 230.400 ;
        RECT 133.200 225.300 135.300 227.400 ;
        RECT 128.400 211.350 129.600 213.600 ;
        RECT 128.100 208.950 130.200 211.050 ;
        RECT 113.700 201.600 115.800 203.700 ;
        RECT 116.700 201.600 118.800 203.700 ;
        RECT 119.700 201.600 121.800 203.700 ;
        RECT 125.100 202.500 127.200 204.600 ;
        RECT 134.100 203.700 135.300 225.300 ;
        RECT 136.500 222.300 137.700 228.300 ;
        RECT 136.500 220.200 138.600 222.300 ;
        RECT 136.500 203.700 137.700 220.200 ;
        RECT 140.100 209.400 141.600 228.300 ;
        RECT 139.500 207.300 141.600 209.400 ;
        RECT 143.400 208.050 144.450 254.400 ;
        RECT 149.400 254.400 150.600 256.650 ;
        RECT 155.400 255.900 156.600 256.650 ;
        RECT 149.400 232.050 150.450 254.400 ;
        RECT 154.950 253.800 157.050 255.900 ;
        RECT 157.950 247.950 160.050 250.050 ;
        RECT 148.950 229.950 151.050 232.050 ;
        RECT 151.950 219.000 154.050 223.050 ;
        RECT 152.400 217.350 153.600 219.000 ;
        RECT 146.100 214.950 148.200 217.050 ;
        RECT 152.100 214.950 154.200 217.050 ;
        RECT 139.500 203.700 140.700 207.300 ;
        RECT 142.950 205.950 145.050 208.050 ;
        RECT 133.200 201.600 135.300 203.700 ;
        RECT 136.200 201.600 138.300 203.700 ;
        RECT 139.200 201.600 141.300 203.700 ;
        RECT 133.950 196.950 136.050 199.050 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 112.950 190.950 118.050 193.050 ;
        RECT 109.950 187.950 112.050 190.050 ;
        RECT 110.400 184.200 111.450 187.950 ;
        RECT 109.950 182.100 112.050 184.200 ;
        RECT 118.950 183.000 121.050 187.050 ;
        RECT 119.400 181.350 120.600 183.000 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 112.950 175.950 115.050 178.050 ;
        RECT 116.400 176.400 117.600 178.650 ;
        RECT 128.400 178.050 129.450 193.950 ;
        RECT 134.400 183.600 135.450 196.950 ;
        RECT 158.400 196.050 159.450 247.950 ;
        RECT 161.400 238.050 162.450 301.950 ;
        RECT 164.400 295.050 165.450 304.950 ;
        RECT 163.950 292.950 166.050 295.050 ;
        RECT 169.950 294.000 172.050 298.050 ;
        RECT 176.400 294.600 177.450 340.950 ;
        RECT 179.400 340.200 180.450 416.100 ;
        RECT 181.950 415.950 184.050 418.050 ;
        RECT 184.950 417.000 187.050 421.050 ;
        RECT 185.400 415.350 186.600 417.000 ;
        RECT 190.950 416.100 193.050 418.200 ;
        RECT 197.400 418.050 198.450 451.950 ;
        RECT 200.400 424.050 201.450 475.950 ;
        RECT 203.100 448.950 205.200 451.050 ;
        RECT 203.400 447.900 204.600 448.650 ;
        RECT 202.950 445.800 205.050 447.900 ;
        RECT 209.400 442.050 210.450 517.950 ;
        RECT 212.400 499.050 213.450 520.950 ;
        RECT 211.950 496.950 214.050 499.050 ;
        RECT 215.400 495.450 216.450 547.950 ;
        RECT 218.400 544.050 219.450 551.400 ;
        RECT 220.950 547.950 223.050 551.400 ;
        RECT 220.950 544.800 223.050 546.900 ;
        RECT 217.950 541.950 220.050 544.050 ;
        RECT 217.950 529.950 220.050 535.050 ;
        RECT 221.400 528.450 222.450 544.800 ;
        RECT 224.400 544.050 225.450 559.950 ;
        RECT 235.950 553.950 238.050 556.050 ;
        RECT 232.950 550.950 235.050 553.050 ;
        RECT 223.950 541.950 226.050 544.050 ;
        RECT 218.400 527.400 222.450 528.450 ;
        RECT 218.400 498.450 219.450 527.400 ;
        RECT 226.950 527.100 229.050 529.200 ;
        RECT 233.400 529.050 234.450 550.950 ;
        RECT 227.400 526.350 228.600 527.100 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 223.950 523.950 226.050 526.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 220.950 520.950 223.050 523.050 ;
        RECT 224.400 522.900 225.600 523.650 ;
        RECT 221.400 517.050 222.450 520.950 ;
        RECT 223.950 520.800 226.050 522.900 ;
        RECT 230.400 522.000 231.600 523.650 ;
        RECT 229.950 517.950 232.050 522.000 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 220.950 514.950 223.050 517.050 ;
        RECT 226.950 514.950 229.050 517.050 ;
        RECT 218.400 497.400 222.450 498.450 ;
        RECT 212.400 494.400 216.450 495.450 ;
        RECT 221.400 495.600 222.450 497.400 ;
        RECT 227.400 496.050 228.450 514.950 ;
        RECT 233.400 510.450 234.450 520.950 ;
        RECT 230.400 509.400 234.450 510.450 ;
        RECT 230.400 505.050 231.450 509.400 ;
        RECT 229.950 502.950 232.050 505.050 ;
        RECT 212.400 469.050 213.450 494.400 ;
        RECT 221.400 493.350 222.600 495.600 ;
        RECT 226.950 493.950 229.050 496.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 218.400 489.000 219.600 490.650 ;
        RECT 224.400 489.900 225.600 490.650 ;
        RECT 230.400 489.900 231.450 502.950 ;
        RECT 236.400 495.450 237.450 553.950 ;
        RECT 238.950 547.950 241.050 550.050 ;
        RECT 239.400 538.050 240.450 547.950 ;
        RECT 242.400 547.050 243.450 592.950 ;
        RECT 254.400 592.050 255.450 598.950 ;
        RECT 260.400 598.050 261.450 605.100 ;
        RECT 266.400 604.350 267.600 605.100 ;
        RECT 272.400 604.350 273.600 606.600 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 269.400 600.900 270.600 601.650 ;
        RECT 268.950 598.800 271.050 600.900 ;
        RECT 275.400 599.400 276.600 601.650 ;
        RECT 259.950 595.950 262.050 598.050 ;
        RECT 275.400 595.050 276.450 599.400 ;
        RECT 277.950 598.800 280.050 600.900 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 253.950 589.950 256.050 592.050 ;
        RECT 245.700 579.300 247.800 581.400 ;
        RECT 248.700 579.300 250.800 581.400 ;
        RECT 251.700 579.300 253.800 581.400 ;
        RECT 246.300 575.700 247.500 579.300 ;
        RECT 245.400 573.600 247.500 575.700 ;
        RECT 245.400 554.700 246.900 573.600 ;
        RECT 249.300 562.800 250.500 579.300 ;
        RECT 248.400 560.700 250.500 562.800 ;
        RECT 249.300 554.700 250.500 560.700 ;
        RECT 251.700 557.700 252.900 579.300 ;
        RECT 259.800 578.400 261.900 580.500 ;
        RECT 265.200 579.300 267.300 581.400 ;
        RECT 268.200 579.300 270.300 581.400 ;
        RECT 271.200 579.300 273.300 581.400 ;
        RECT 256.800 571.950 258.900 574.050 ;
        RECT 257.400 570.000 258.600 571.650 ;
        RECT 256.950 565.950 259.050 570.000 ;
        RECT 260.400 567.900 261.300 578.400 ;
        RECT 263.100 572.400 265.200 574.500 ;
        RECT 260.400 565.800 262.500 567.900 ;
        RECT 266.100 567.000 267.300 579.300 ;
        RECT 260.400 559.200 261.300 565.800 ;
        RECT 265.800 564.900 267.900 567.000 ;
        RECT 251.700 555.600 253.800 557.700 ;
        RECT 260.400 557.100 262.500 559.200 ;
        RECT 266.100 557.700 267.300 564.900 ;
        RECT 268.800 561.600 270.300 579.300 ;
        RECT 268.800 559.500 270.900 561.600 ;
        RECT 265.800 555.600 267.900 557.700 ;
        RECT 268.800 554.700 270.300 559.500 ;
        RECT 272.100 557.700 273.300 579.300 ;
        RECT 245.400 552.600 248.400 554.700 ;
        RECT 249.300 552.600 251.400 554.700 ;
        RECT 253.950 550.950 256.050 553.050 ;
        RECT 268.200 552.600 270.300 554.700 ;
        RECT 271.200 552.600 273.300 557.700 ;
        RECT 274.200 579.300 276.300 581.400 ;
        RECT 274.200 561.600 275.700 579.300 ;
        RECT 278.400 568.050 279.450 598.800 ;
        RECT 281.400 595.050 282.450 616.950 ;
        RECT 296.400 616.050 297.450 661.950 ;
        RECT 299.400 661.050 300.450 670.950 ;
        RECT 298.950 658.950 301.050 661.050 ;
        RECT 302.400 658.050 303.450 674.400 ;
        RECT 301.950 655.950 304.050 658.050 ;
        RECT 302.400 648.600 303.450 655.950 ;
        RECT 304.950 652.950 307.050 655.050 ;
        RECT 302.400 646.350 303.600 648.600 ;
        RECT 305.400 646.050 306.450 652.950 ;
        RECT 308.400 652.050 309.450 674.400 ;
        RECT 320.400 667.050 321.450 677.400 ;
        RECT 328.950 673.950 331.050 676.050 ;
        RECT 325.950 667.950 328.050 670.050 ;
        RECT 319.950 664.950 322.050 667.050 ;
        RECT 319.950 655.950 322.050 658.050 ;
        RECT 307.950 649.950 310.050 652.050 ;
        RECT 311.400 648.450 312.600 648.600 ;
        RECT 311.400 647.400 315.450 648.450 ;
        RECT 311.400 646.350 312.600 647.400 ;
        RECT 301.800 643.950 303.900 646.050 ;
        RECT 304.950 643.950 307.050 646.050 ;
        RECT 310.800 643.950 312.900 646.050 ;
        RECT 304.950 640.800 307.050 642.900 ;
        RECT 298.950 631.950 301.050 634.050 ;
        RECT 299.400 619.050 300.450 631.950 ;
        RECT 298.950 616.950 301.050 619.050 ;
        RECT 295.950 613.950 298.050 616.050 ;
        RECT 283.950 607.950 286.050 610.050 ;
        RECT 280.950 592.950 283.050 595.050 ;
        RECT 284.400 592.050 285.450 607.950 ;
        RECT 292.950 605.100 295.050 610.050 ;
        RECT 298.950 605.100 301.050 607.200 ;
        RECT 293.400 604.350 294.600 605.100 ;
        RECT 299.400 604.350 300.600 605.100 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 286.950 598.950 289.050 601.050 ;
        RECT 290.400 599.400 291.600 601.650 ;
        RECT 296.400 599.400 297.600 601.650 ;
        RECT 280.800 589.800 282.900 591.900 ;
        RECT 283.950 589.950 286.050 592.050 ;
        RECT 281.400 571.050 282.450 589.800 ;
        RECT 287.400 586.050 288.450 598.950 ;
        RECT 290.400 595.050 291.450 599.400 ;
        RECT 296.400 595.050 297.450 599.400 ;
        RECT 301.950 598.950 304.050 601.050 ;
        RECT 289.950 592.950 292.050 595.050 ;
        RECT 295.950 592.950 298.050 595.050 ;
        RECT 286.950 583.950 289.050 586.050 ;
        RECT 295.950 583.950 298.050 586.050 ;
        RECT 283.950 574.950 286.050 577.050 ;
        RECT 280.950 568.950 283.050 571.050 ;
        RECT 284.400 570.600 285.450 574.950 ;
        RECT 296.400 574.050 297.450 583.950 ;
        RECT 298.950 574.950 301.050 577.050 ;
        RECT 295.950 571.950 298.050 574.050 ;
        RECT 284.400 568.350 285.600 570.600 ;
        RECT 292.950 570.450 295.050 571.200 ;
        RECT 292.950 569.400 297.450 570.450 ;
        RECT 292.950 569.100 295.050 569.400 ;
        RECT 293.400 568.350 294.600 569.100 ;
        RECT 277.950 565.950 280.050 568.050 ;
        RECT 283.800 565.950 285.900 568.050 ;
        RECT 292.800 565.950 294.900 568.050 ;
        RECT 274.200 559.500 276.300 561.600 ;
        RECT 274.200 554.700 275.700 559.500 ;
        RECT 274.200 552.600 276.300 554.700 ;
        RECT 296.400 553.050 297.450 569.400 ;
        RECT 295.950 550.950 298.050 553.050 ;
        RECT 241.950 544.950 244.050 547.050 ;
        RECT 238.950 535.950 241.050 538.050 ;
        RECT 244.950 528.000 247.050 532.050 ;
        RECT 245.400 526.350 246.600 528.000 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 244.950 523.950 247.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 242.400 522.000 243.600 523.650 ;
        RECT 241.950 517.950 244.050 522.000 ;
        RECT 248.400 521.400 249.600 523.650 ;
        RECT 248.400 514.050 249.450 521.400 ;
        RECT 254.400 517.050 255.450 550.950 ;
        RECT 271.950 541.950 274.050 544.050 ;
        RECT 268.950 532.950 271.050 535.050 ;
        RECT 256.950 526.950 259.050 529.050 ;
        RECT 262.950 528.000 265.050 532.050 ;
        RECT 269.400 528.600 270.450 532.950 ;
        RECT 272.400 529.050 273.450 541.950 ;
        RECT 280.950 535.950 283.050 538.050 ;
        RECT 277.950 532.950 280.050 535.050 ;
        RECT 253.950 514.950 256.050 517.050 ;
        RECT 247.950 511.950 250.050 514.050 ;
        RECT 239.400 495.450 240.600 495.600 ;
        RECT 233.400 494.400 240.600 495.450 ;
        RECT 217.950 484.950 220.050 489.000 ;
        RECT 223.950 487.800 226.050 489.900 ;
        RECT 229.950 487.800 232.050 489.900 ;
        RECT 211.950 466.950 214.050 469.050 ;
        RECT 217.950 466.950 220.050 469.050 ;
        RECT 212.100 448.950 214.200 451.050 ;
        RECT 212.400 447.450 213.600 448.650 ;
        RECT 218.400 447.900 219.450 466.950 ;
        RECT 233.400 466.050 234.450 494.400 ;
        RECT 239.400 493.350 240.600 494.400 ;
        RECT 244.950 494.100 247.050 496.200 ;
        RECT 257.400 495.450 258.450 526.950 ;
        RECT 263.400 526.350 264.600 528.000 ;
        RECT 269.400 526.350 270.600 528.600 ;
        RECT 271.950 526.950 274.050 529.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 266.400 522.900 267.600 523.650 ;
        RECT 265.950 520.800 268.050 522.900 ;
        RECT 271.950 514.950 274.050 517.050 ;
        RECT 254.400 494.400 258.450 495.450 ;
        RECT 245.400 493.350 246.600 494.100 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 235.950 487.950 238.050 490.050 ;
        RECT 242.400 489.000 243.600 490.650 ;
        RECT 248.400 489.900 249.600 490.650 ;
        RECT 221.700 462.300 223.800 464.400 ;
        RECT 222.300 457.500 223.800 462.300 ;
        RECT 221.700 455.400 223.800 457.500 ;
        RECT 212.400 446.400 216.450 447.450 ;
        RECT 208.950 439.950 211.050 442.050 ;
        RECT 215.400 439.050 216.450 446.400 ;
        RECT 217.950 445.800 220.050 447.900 ;
        RECT 214.950 436.950 217.050 439.050 ;
        RECT 215.400 433.050 216.450 436.950 ;
        RECT 214.950 430.950 217.050 433.050 ;
        RECT 199.950 421.950 202.050 424.050 ;
        RECT 215.400 421.050 216.450 430.950 ;
        RECT 214.950 418.950 217.050 421.050 ;
        RECT 191.400 415.350 192.600 416.100 ;
        RECT 196.950 415.950 199.050 418.050 ;
        RECT 202.950 415.950 205.050 418.050 ;
        RECT 211.950 416.100 214.050 418.200 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 193.950 412.950 196.050 415.050 ;
        RECT 181.950 409.950 184.050 412.050 ;
        RECT 188.400 410.400 189.600 412.650 ;
        RECT 182.400 373.050 183.450 409.950 ;
        RECT 188.400 406.050 189.450 410.400 ;
        RECT 196.950 409.950 199.050 412.050 ;
        RECT 187.950 403.950 190.050 406.050 ;
        RECT 184.950 394.950 187.050 397.050 ;
        RECT 185.400 391.050 186.450 394.950 ;
        RECT 184.950 388.950 187.050 391.050 ;
        RECT 190.950 379.950 193.050 382.050 ;
        RECT 181.950 370.950 184.050 373.050 ;
        RECT 184.950 371.100 187.050 373.200 ;
        RECT 191.400 372.600 192.450 379.950 ;
        RECT 197.400 376.200 198.450 409.950 ;
        RECT 196.950 374.100 199.050 376.200 ;
        RECT 185.400 370.350 186.600 371.100 ;
        RECT 191.400 370.350 192.600 372.600 ;
        RECT 196.950 370.950 199.050 373.050 ;
        RECT 197.400 370.350 198.600 370.950 ;
        RECT 184.950 367.950 187.050 370.050 ;
        RECT 187.950 367.950 190.050 370.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 188.400 365.400 189.600 367.650 ;
        RECT 194.400 366.000 195.600 367.650 ;
        RECT 188.400 355.050 189.450 365.400 ;
        RECT 193.950 361.950 196.050 366.000 ;
        RECT 187.950 352.950 190.050 355.050 ;
        RECT 199.950 346.950 202.050 349.050 ;
        RECT 190.950 343.950 193.050 346.050 ;
        RECT 178.950 338.100 181.050 340.200 ;
        RECT 184.950 338.100 187.050 340.200 ;
        RECT 191.400 339.600 192.450 343.950 ;
        RECT 185.400 337.350 186.600 338.100 ;
        RECT 191.400 337.350 192.600 339.600 ;
        RECT 196.950 337.950 199.050 340.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 190.950 334.950 193.050 337.050 ;
        RECT 182.400 333.000 183.600 334.650 ;
        RECT 181.950 328.950 184.050 333.000 ;
        RECT 188.400 332.400 189.600 334.650 ;
        RECT 178.950 313.950 181.050 316.050 ;
        RECT 179.400 295.050 180.450 313.950 ;
        RECT 188.400 313.050 189.450 332.400 ;
        RECT 197.400 325.050 198.450 337.950 ;
        RECT 200.400 331.050 201.450 346.950 ;
        RECT 203.400 340.050 204.450 415.950 ;
        RECT 212.400 415.350 213.600 416.100 ;
        RECT 206.400 412.950 208.500 415.050 ;
        RECT 211.500 412.950 213.600 415.050 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 206.400 410.400 207.600 412.650 ;
        RECT 206.400 379.050 207.450 410.400 ;
        RECT 208.950 400.950 211.050 403.050 ;
        RECT 205.950 376.950 208.050 379.050 ;
        RECT 209.400 376.050 210.450 400.950 ;
        RECT 215.400 388.050 216.450 412.950 ;
        RECT 214.950 385.950 217.050 388.050 ;
        RECT 218.400 385.050 219.450 445.800 ;
        RECT 222.300 437.700 223.800 455.400 ;
        RECT 221.700 435.600 223.800 437.700 ;
        RECT 224.700 459.300 226.800 464.400 ;
        RECT 227.700 462.300 229.800 464.400 ;
        RECT 232.950 463.950 235.050 466.050 ;
        RECT 236.400 463.050 237.450 487.950 ;
        RECT 241.950 484.950 244.050 489.000 ;
        RECT 247.950 487.800 250.050 489.900 ;
        RECT 254.400 466.050 255.450 494.400 ;
        RECT 262.950 494.100 265.050 496.200 ;
        RECT 263.400 493.350 264.600 494.100 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 265.950 490.950 268.050 493.050 ;
        RECT 260.400 489.900 261.600 490.650 ;
        RECT 259.950 484.950 262.050 489.900 ;
        RECT 266.400 488.400 267.600 490.650 ;
        RECT 272.400 489.450 273.450 514.950 ;
        RECT 278.400 502.050 279.450 532.950 ;
        RECT 281.400 517.050 282.450 535.950 ;
        RECT 295.950 530.100 298.050 532.200 ;
        RECT 283.950 527.100 286.050 529.200 ;
        RECT 284.400 526.350 285.600 527.100 ;
        RECT 292.950 526.950 295.050 529.050 ;
        RECT 284.100 523.950 286.200 526.050 ;
        RECT 289.500 523.950 291.600 526.050 ;
        RECT 290.400 522.900 291.600 523.650 ;
        RECT 289.950 520.800 292.050 522.900 ;
        RECT 280.950 514.950 283.050 517.050 ;
        RECT 277.950 499.950 280.050 502.050 ;
        RECT 281.400 498.450 282.450 514.950 ;
        RECT 278.400 497.400 282.450 498.450 ;
        RECT 278.400 495.600 279.450 497.400 ;
        RECT 278.400 493.350 279.600 495.600 ;
        RECT 293.400 493.050 294.450 526.950 ;
        RECT 278.400 490.950 280.500 493.050 ;
        RECT 283.800 490.950 285.900 493.050 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 284.400 489.900 285.600 490.650 ;
        RECT 296.400 490.050 297.450 530.100 ;
        RECT 299.400 508.050 300.450 574.950 ;
        RECT 302.400 568.050 303.450 598.950 ;
        RECT 305.400 595.050 306.450 640.800 ;
        RECT 310.950 637.950 313.050 640.050 ;
        RECT 307.950 631.950 310.050 634.050 ;
        RECT 308.400 607.050 309.450 631.950 ;
        RECT 311.400 607.200 312.450 637.950 ;
        RECT 314.400 634.050 315.450 647.400 ;
        RECT 313.950 631.950 316.050 634.050 ;
        RECT 316.950 610.950 319.050 613.050 ;
        RECT 307.950 604.950 310.050 607.050 ;
        RECT 310.950 605.100 313.050 607.200 ;
        RECT 317.400 606.600 318.450 610.950 ;
        RECT 320.400 607.050 321.450 655.950 ;
        RECT 326.400 654.450 327.450 667.950 ;
        RECT 329.400 664.050 330.450 673.950 ;
        RECT 332.400 670.050 333.450 715.950 ;
        RECT 341.400 712.050 342.450 722.400 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 344.400 715.050 345.450 721.800 ;
        RECT 343.950 712.950 346.050 715.050 ;
        RECT 340.950 709.950 343.050 712.050 ;
        RECT 347.400 703.050 348.450 751.650 ;
        RECT 353.400 751.050 354.450 755.400 ;
        RECT 352.950 748.950 355.050 751.050 ;
        RECT 362.400 741.450 363.450 761.400 ;
        RECT 367.950 761.100 370.050 763.200 ;
        RECT 374.400 762.600 375.450 770.400 ;
        RECT 380.400 762.600 381.450 775.950 ;
        RECT 386.400 775.050 387.450 784.950 ;
        RECT 385.950 772.950 388.050 775.050 ;
        RECT 385.950 763.950 388.050 766.050 ;
        RECT 368.400 760.350 369.600 761.100 ;
        RECT 374.400 760.350 375.600 762.600 ;
        RECT 380.400 760.350 381.600 762.600 ;
        RECT 367.950 757.950 370.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 371.400 755.400 372.600 757.650 ;
        RECT 377.400 756.900 378.600 757.650 ;
        RECT 367.950 748.950 370.050 751.050 ;
        RECT 362.400 740.400 366.450 741.450 ;
        RECT 361.950 736.950 364.050 739.050 ;
        RECT 355.950 733.950 358.050 736.050 ;
        RECT 356.400 729.600 357.450 733.950 ;
        RECT 362.400 729.600 363.450 736.950 ;
        RECT 365.400 730.050 366.450 740.400 ;
        RECT 356.400 727.350 357.600 729.600 ;
        RECT 362.400 727.350 363.600 729.600 ;
        RECT 364.950 727.950 367.050 730.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 353.400 722.400 354.600 724.650 ;
        RECT 359.400 723.000 360.600 724.650 ;
        RECT 353.400 718.050 354.450 722.400 ;
        RECT 358.950 718.950 361.050 723.000 ;
        RECT 352.950 715.950 355.050 718.050 ;
        RECT 346.950 700.950 349.050 703.050 ;
        RECT 335.400 696.300 338.400 698.400 ;
        RECT 339.300 696.300 341.400 698.400 ;
        RECT 358.200 696.300 360.300 698.400 ;
        RECT 335.400 677.400 336.900 696.300 ;
        RECT 339.300 690.300 340.500 696.300 ;
        RECT 338.400 688.200 340.500 690.300 ;
        RECT 335.400 675.300 337.500 677.400 ;
        RECT 336.300 671.700 337.500 675.300 ;
        RECT 339.300 671.700 340.500 688.200 ;
        RECT 341.700 693.300 343.800 695.400 ;
        RECT 341.700 671.700 342.900 693.300 ;
        RECT 350.400 691.800 352.500 693.900 ;
        RECT 355.800 693.300 357.900 695.400 ;
        RECT 350.400 685.200 351.300 691.800 ;
        RECT 356.100 686.100 357.300 693.300 ;
        RECT 358.800 691.500 360.300 696.300 ;
        RECT 361.200 693.300 363.300 698.400 ;
        RECT 358.800 689.400 360.900 691.500 ;
        RECT 350.400 683.100 352.500 685.200 ;
        RECT 355.800 684.000 357.900 686.100 ;
        RECT 346.950 680.100 349.050 682.200 ;
        RECT 347.400 679.350 348.600 680.100 ;
        RECT 346.800 676.950 348.900 679.050 ;
        RECT 350.400 672.600 351.300 683.100 ;
        RECT 353.100 676.500 355.200 678.600 ;
        RECT 331.950 667.950 334.050 670.050 ;
        RECT 335.700 669.600 337.800 671.700 ;
        RECT 338.700 669.600 340.800 671.700 ;
        RECT 341.700 669.600 343.800 671.700 ;
        RECT 349.800 670.500 351.900 672.600 ;
        RECT 356.100 671.700 357.300 684.000 ;
        RECT 358.800 671.700 360.300 689.400 ;
        RECT 362.100 671.700 363.300 693.300 ;
        RECT 355.200 669.600 357.300 671.700 ;
        RECT 358.200 669.600 360.300 671.700 ;
        RECT 361.200 669.600 363.300 671.700 ;
        RECT 364.200 696.300 366.300 698.400 ;
        RECT 364.200 691.500 365.700 696.300 ;
        RECT 364.200 689.400 366.300 691.500 ;
        RECT 368.400 691.050 369.450 748.950 ;
        RECT 371.400 745.050 372.450 755.400 ;
        RECT 376.950 754.800 379.050 756.900 ;
        RECT 382.950 754.950 385.050 757.050 ;
        RECT 386.400 756.900 387.450 763.950 ;
        RECT 389.400 763.050 390.450 799.800 ;
        RECT 401.400 796.050 402.450 800.400 ;
        RECT 406.950 799.950 409.050 802.050 ;
        RECT 400.950 793.950 403.050 796.050 ;
        RECT 397.950 778.950 400.050 781.050 ;
        RECT 388.950 760.950 391.050 763.050 ;
        RECT 391.950 762.000 394.050 766.050 ;
        RECT 398.400 762.600 399.450 778.950 ;
        RECT 392.400 760.350 393.600 762.000 ;
        RECT 398.400 760.350 399.600 762.600 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 370.950 742.950 373.050 745.050 ;
        RECT 376.950 739.950 379.050 742.050 ;
        RECT 377.400 730.200 378.450 739.950 ;
        RECT 379.950 736.950 382.050 739.050 ;
        RECT 380.400 733.050 381.450 736.950 ;
        RECT 379.950 730.950 382.050 733.050 ;
        RECT 376.950 728.100 379.050 730.200 ;
        RECT 383.400 729.600 384.450 754.950 ;
        RECT 385.950 754.800 388.050 756.900 ;
        RECT 388.950 754.950 391.050 757.050 ;
        RECT 395.400 756.900 396.600 757.650 ;
        RECT 401.400 756.900 402.600 757.650 ;
        RECT 389.400 730.050 390.450 754.950 ;
        RECT 394.950 754.800 397.050 756.900 ;
        RECT 400.950 754.800 403.050 756.900 ;
        RECT 407.400 751.050 408.450 799.950 ;
        RECT 406.950 748.950 409.050 751.050 ;
        RECT 410.400 745.050 411.450 832.800 ;
        RECT 413.400 823.050 414.450 833.400 ;
        RECT 418.950 829.950 421.050 834.000 ;
        RECT 412.950 820.950 415.050 823.050 ;
        RECT 424.950 817.950 427.050 820.050 ;
        RECT 425.400 808.200 426.450 817.950 ;
        RECT 428.400 811.050 429.450 853.950 ;
        RECT 437.400 840.600 438.450 859.950 ;
        RECT 445.950 844.950 448.050 847.050 ;
        RECT 437.400 838.350 438.600 840.600 ;
        RECT 433.950 835.950 436.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 434.400 834.900 435.600 835.650 ;
        RECT 440.400 834.900 441.600 835.650 ;
        RECT 446.400 834.900 447.450 844.950 ;
        RECT 433.950 834.450 436.050 834.900 ;
        RECT 431.400 833.400 436.050 834.450 ;
        RECT 427.950 808.950 430.050 811.050 ;
        RECT 415.950 806.100 418.050 808.200 ;
        RECT 424.950 806.100 427.050 808.200 ;
        RECT 416.400 802.050 417.450 806.100 ;
        RECT 425.400 805.350 426.600 806.100 ;
        RECT 419.100 802.950 421.200 805.050 ;
        RECT 424.500 802.950 426.600 805.050 ;
        RECT 427.800 802.950 429.900 805.050 ;
        RECT 415.950 799.950 418.050 802.050 ;
        RECT 419.400 800.400 420.600 802.650 ;
        RECT 428.400 801.900 429.600 802.650 ;
        RECT 419.400 796.050 420.450 800.400 ;
        RECT 427.950 799.800 430.050 801.900 ;
        RECT 418.950 793.950 421.050 796.050 ;
        RECT 415.950 784.950 418.050 787.050 ;
        RECT 416.400 762.600 417.450 784.950 ;
        RECT 419.400 784.050 420.450 793.950 ;
        RECT 431.400 793.050 432.450 833.400 ;
        RECT 433.950 832.800 436.050 833.400 ;
        RECT 439.950 832.800 442.050 834.900 ;
        RECT 445.950 832.800 448.050 834.900 ;
        RECT 449.400 832.050 450.450 871.950 ;
        RECT 469.950 868.950 472.050 871.050 ;
        RECT 454.950 853.950 457.050 856.050 ;
        RECT 455.400 840.600 456.450 853.950 ;
        RECT 455.400 838.350 456.600 840.600 ;
        RECT 466.950 839.100 469.050 841.200 ;
        RECT 454.950 835.950 457.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 458.400 834.900 459.600 835.650 ;
        RECT 467.400 835.050 468.450 839.100 ;
        RECT 470.400 835.050 471.450 868.950 ;
        RECT 476.400 868.050 477.450 889.950 ;
        RECT 479.400 885.450 480.450 907.950 ;
        RECT 485.400 895.050 486.450 917.100 ;
        RECT 497.400 916.350 498.600 917.100 ;
        RECT 503.400 916.350 504.600 918.600 ;
        RECT 508.950 917.100 511.050 919.200 ;
        RECT 515.400 918.600 516.450 928.950 ;
        RECT 565.950 919.950 568.050 922.050 ;
        RECT 493.950 913.950 496.050 916.050 ;
        RECT 496.950 913.950 499.050 916.050 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 494.400 911.400 495.600 913.650 ;
        RECT 500.400 911.400 501.600 913.650 ;
        RECT 494.400 895.050 495.450 911.400 ;
        RECT 484.950 892.950 487.050 895.050 ;
        RECT 493.950 892.950 496.050 895.050 ;
        RECT 484.800 888.300 486.900 890.400 ;
        RECT 487.950 889.950 490.050 892.050 ;
        RECT 488.400 889.200 489.600 889.950 ;
        RECT 482.400 885.450 483.600 885.600 ;
        RECT 479.400 884.400 483.600 885.450 ;
        RECT 482.400 883.350 483.600 884.400 ;
        RECT 482.100 880.950 484.200 883.050 ;
        RECT 485.100 882.900 486.000 888.300 ;
        RECT 488.100 886.800 490.200 888.900 ;
        RECT 492.000 885.900 494.100 887.700 ;
        RECT 486.900 884.700 495.600 885.900 ;
        RECT 486.900 883.800 489.000 884.700 ;
        RECT 485.100 881.700 492.000 882.900 ;
        RECT 485.100 874.500 486.300 881.700 ;
        RECT 488.100 877.950 490.200 880.050 ;
        RECT 491.100 879.300 492.000 881.700 ;
        RECT 488.400 875.400 489.600 877.650 ;
        RECT 491.100 877.200 493.200 879.300 ;
        RECT 494.700 875.700 495.600 884.700 ;
        RECT 496.800 880.950 498.900 883.050 ;
        RECT 497.400 879.450 498.600 880.650 ;
        RECT 500.400 879.450 501.450 911.400 ;
        RECT 509.400 904.050 510.450 917.100 ;
        RECT 515.400 916.350 516.600 918.600 ;
        RECT 520.950 917.100 523.050 919.200 ;
        RECT 541.950 917.100 544.050 919.200 ;
        RECT 556.950 917.100 559.050 919.200 ;
        RECT 521.400 916.350 522.600 917.100 ;
        RECT 542.400 916.350 543.600 917.100 ;
        RECT 557.400 916.350 558.600 917.100 ;
        RECT 514.950 913.950 517.050 916.050 ;
        RECT 517.950 913.950 520.050 916.050 ;
        RECT 520.950 913.950 523.050 916.050 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 538.950 913.950 541.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 556.950 913.950 559.050 916.050 ;
        RECT 559.950 913.950 562.050 916.050 ;
        RECT 518.400 912.900 519.600 913.650 ;
        RECT 524.400 912.900 525.600 913.650 ;
        RECT 517.950 910.800 520.050 912.900 ;
        RECT 523.950 907.950 526.050 912.900 ;
        RECT 539.400 911.400 540.600 913.650 ;
        RECT 545.400 912.450 546.600 913.650 ;
        RECT 545.400 911.400 549.450 912.450 ;
        RECT 560.400 912.000 561.600 913.650 ;
        RECT 539.400 904.050 540.450 911.400 ;
        RECT 508.950 901.950 511.050 904.050 ;
        RECT 538.950 901.950 541.050 904.050 ;
        RECT 523.950 895.950 526.050 898.050 ;
        RECT 541.950 895.950 544.050 898.050 ;
        RECT 508.950 885.000 511.050 889.050 ;
        RECT 509.400 883.350 510.600 885.000 ;
        RECT 514.950 884.100 517.050 886.200 ;
        RECT 515.400 883.350 516.600 884.100 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 511.950 880.950 514.050 883.050 ;
        RECT 514.950 880.950 517.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 497.400 878.400 501.450 879.450 ;
        RECT 512.400 879.000 513.600 880.650 ;
        RECT 518.400 879.900 519.600 880.650 ;
        RECT 524.400 879.900 525.450 895.950 ;
        RECT 526.800 884.100 528.900 886.200 ;
        RECT 527.400 880.050 528.450 884.100 ;
        RECT 529.950 883.950 532.050 889.050 ;
        RECT 535.950 884.100 538.050 886.200 ;
        RECT 542.400 885.600 543.450 895.950 ;
        RECT 548.400 895.050 549.450 911.400 ;
        RECT 559.950 907.950 562.050 912.000 ;
        RECT 566.400 895.050 567.450 919.950 ;
        RECT 571.950 918.000 574.050 922.050 ;
        RECT 578.400 918.600 579.450 934.950 ;
        RECT 697.950 925.950 700.050 928.050 ;
        RECT 829.950 925.950 832.050 928.050 ;
        RECT 844.950 925.950 847.050 928.050 ;
        RECT 862.950 925.950 865.050 928.050 ;
        RECT 622.950 922.950 625.050 925.050 ;
        RECT 646.950 922.950 649.050 925.050 ;
        RECT 682.950 922.950 685.050 925.050 ;
        RECT 572.400 916.350 573.600 918.000 ;
        RECT 578.400 916.350 579.600 918.600 ;
        RECT 583.950 917.100 586.050 919.200 ;
        RECT 584.400 916.350 585.600 917.100 ;
        RECT 589.950 916.950 592.050 919.050 ;
        RECT 601.950 917.100 604.050 919.200 ;
        RECT 623.400 918.600 624.450 922.950 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 574.950 913.950 577.050 916.050 ;
        RECT 577.950 913.950 580.050 916.050 ;
        RECT 580.950 913.950 583.050 916.050 ;
        RECT 583.950 913.950 586.050 916.050 ;
        RECT 575.400 912.900 576.600 913.650 ;
        RECT 574.950 910.800 577.050 912.900 ;
        RECT 581.400 912.000 582.600 913.650 ;
        RECT 574.950 909.300 577.050 909.750 ;
        RECT 580.950 909.300 583.050 912.000 ;
        RECT 586.950 910.950 589.050 913.050 ;
        RECT 574.950 908.250 583.050 909.300 ;
        RECT 574.950 907.650 577.050 908.250 ;
        RECT 580.950 907.950 583.050 908.250 ;
        RECT 583.950 907.950 586.050 910.050 ;
        RECT 577.950 895.950 580.050 898.050 ;
        RECT 547.950 892.950 550.050 895.050 ;
        RECT 565.950 892.950 568.050 895.050 ;
        RECT 536.400 883.350 537.600 884.100 ;
        RECT 542.400 883.350 543.600 885.600 ;
        RECT 532.950 880.950 535.050 883.050 ;
        RECT 535.950 880.950 538.050 883.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 484.800 872.400 486.900 874.500 ;
        RECT 494.400 873.600 496.500 875.700 ;
        RECT 511.950 874.950 514.050 879.000 ;
        RECT 517.950 877.800 520.050 879.900 ;
        RECT 523.800 877.800 525.900 879.900 ;
        RECT 526.950 877.950 529.050 880.050 ;
        RECT 533.400 878.400 534.600 880.650 ;
        RECT 539.400 879.900 540.600 880.650 ;
        RECT 475.950 865.950 478.050 868.050 ;
        RECT 533.400 865.050 534.450 878.400 ;
        RECT 538.950 877.800 541.050 879.900 ;
        RECT 539.400 876.450 540.450 877.800 ;
        RECT 536.400 875.400 540.450 876.450 ;
        RECT 511.950 862.950 514.050 865.050 ;
        RECT 532.950 862.950 535.050 865.050 ;
        RECT 475.950 859.950 478.050 862.050 ;
        RECT 472.950 856.950 475.050 859.050 ;
        RECT 473.400 841.050 474.450 856.950 ;
        RECT 476.400 847.050 477.450 859.950 ;
        RECT 475.950 844.950 478.050 847.050 ;
        RECT 472.950 838.950 475.050 841.050 ;
        RECT 475.950 839.100 478.050 841.200 ;
        RECT 481.950 840.000 484.050 844.050 ;
        RECT 476.400 838.350 477.600 839.100 ;
        RECT 482.400 838.350 483.600 840.000 ;
        RECT 490.950 839.100 493.050 841.200 ;
        RECT 496.950 839.100 499.050 841.200 ;
        RECT 502.950 839.100 505.050 841.200 ;
        RECT 475.950 835.950 478.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 457.950 832.800 460.050 834.900 ;
        RECT 466.800 832.950 468.900 835.050 ;
        RECT 469.950 832.950 472.050 835.050 ;
        RECT 472.950 832.950 475.050 835.050 ;
        RECT 479.400 834.900 480.600 835.650 ;
        RECT 448.950 829.950 451.050 832.050 ;
        RECT 454.950 829.950 457.050 832.050 ;
        RECT 439.950 820.950 442.050 823.050 ;
        RECT 433.950 808.950 436.050 811.050 ;
        RECT 430.950 790.950 433.050 793.050 ;
        RECT 431.400 787.050 432.450 790.950 ;
        RECT 430.950 784.950 433.050 787.050 ;
        RECT 418.950 781.950 421.050 784.050 ;
        RECT 424.950 781.950 427.050 784.050 ;
        RECT 421.950 766.950 424.050 769.050 ;
        RECT 422.400 762.600 423.450 766.950 ;
        RECT 425.400 766.050 426.450 781.950 ;
        RECT 430.950 775.950 433.050 778.050 ;
        RECT 424.950 763.950 427.050 766.050 ;
        RECT 416.400 760.350 417.600 762.600 ;
        RECT 422.400 760.350 423.600 762.600 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 418.950 757.950 421.050 760.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 419.400 756.900 420.600 757.650 ;
        RECT 425.400 756.900 426.600 757.650 ;
        RECT 418.950 754.800 421.050 756.900 ;
        RECT 424.950 754.800 427.050 756.900 ;
        RECT 431.400 754.050 432.450 775.950 ;
        RECT 434.400 763.200 435.450 808.950 ;
        RECT 440.400 807.600 441.450 820.950 ;
        RECT 445.950 814.950 448.050 817.050 ;
        RECT 446.400 807.600 447.450 814.950 ;
        RECT 440.400 805.350 441.600 807.600 ;
        RECT 446.400 805.350 447.600 807.600 ;
        RECT 439.950 802.950 442.050 805.050 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 445.950 802.950 448.050 805.050 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 443.400 801.900 444.600 802.650 ;
        RECT 442.950 799.800 445.050 801.900 ;
        RECT 449.400 800.400 450.600 802.650 ;
        RECT 455.400 801.450 456.450 829.950 ;
        RECT 473.400 829.050 474.450 832.950 ;
        RECT 478.950 832.800 481.050 834.900 ;
        RECT 485.400 833.400 486.600 835.650 ;
        RECT 485.400 831.450 486.450 833.400 ;
        RECT 482.400 830.400 486.450 831.450 ;
        RECT 472.950 826.950 475.050 829.050 ;
        RECT 472.950 820.950 475.050 823.050 ;
        RECT 463.950 806.100 466.050 808.200 ;
        RECT 464.400 805.350 465.600 806.100 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 466.950 802.950 469.050 805.050 ;
        RECT 452.400 800.400 456.450 801.450 ;
        RECT 461.400 800.400 462.600 802.650 ;
        RECT 467.400 801.000 468.600 802.650 ;
        RECT 443.400 796.050 444.450 799.800 ;
        RECT 439.800 793.950 441.900 796.050 ;
        RECT 442.950 793.950 445.050 796.050 ;
        RECT 436.950 790.950 439.050 793.050 ;
        RECT 433.950 761.100 436.050 763.200 ;
        RECT 437.400 763.050 438.450 790.950 ;
        RECT 440.400 787.050 441.450 793.950 ;
        RECT 449.400 793.050 450.450 800.400 ;
        RECT 448.950 790.950 451.050 793.050 ;
        RECT 439.950 784.950 442.050 787.050 ;
        RECT 448.950 769.950 451.050 772.050 ;
        RECT 445.950 766.950 448.050 769.050 ;
        RECT 434.400 756.900 435.450 761.100 ;
        RECT 436.950 760.950 439.050 763.050 ;
        RECT 439.950 761.100 442.050 763.200 ;
        RECT 446.400 762.600 447.450 766.950 ;
        RECT 449.400 763.050 450.450 769.950 ;
        RECT 440.400 760.350 441.600 761.100 ;
        RECT 446.400 760.350 447.600 762.600 ;
        RECT 448.950 760.950 451.050 763.050 ;
        RECT 439.950 757.950 442.050 760.050 ;
        RECT 442.950 757.950 445.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 433.950 754.800 436.050 756.900 ;
        RECT 436.950 754.950 439.050 757.050 ;
        RECT 443.400 756.000 444.600 757.650 ;
        RECT 430.950 751.950 433.050 754.050 ;
        RECT 409.950 742.950 412.050 745.050 ;
        RECT 400.950 733.950 403.050 736.050 ;
        RECT 377.400 727.350 378.600 728.100 ;
        RECT 383.400 727.350 384.600 729.600 ;
        RECT 388.800 727.950 390.900 730.050 ;
        RECT 391.950 727.950 394.050 730.050 ;
        RECT 401.400 729.600 402.450 733.950 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 385.950 724.950 388.050 727.050 ;
        RECT 374.400 723.900 375.600 724.650 ;
        RECT 373.950 721.800 376.050 723.900 ;
        RECT 380.400 722.400 381.600 724.650 ;
        RECT 386.400 723.000 387.600 724.650 ;
        RECT 380.400 721.050 381.450 722.400 ;
        RECT 376.950 719.550 381.450 721.050 ;
        RECT 376.950 718.950 381.000 719.550 ;
        RECT 382.950 718.950 385.050 721.050 ;
        RECT 385.950 718.950 388.050 723.000 ;
        RECT 388.800 721.950 390.900 724.050 ;
        RECT 376.950 715.800 379.050 717.900 ;
        RECT 364.200 671.700 365.700 689.400 ;
        RECT 367.950 688.950 370.050 691.050 ;
        RECT 373.800 682.950 375.900 685.050 ;
        RECT 370.950 679.950 373.050 682.050 ;
        RECT 374.400 680.400 375.600 682.650 ;
        RECT 377.400 682.050 378.450 715.800 ;
        RECT 383.400 703.050 384.450 718.950 ;
        RECT 382.950 700.950 385.050 703.050 ;
        RECT 382.800 682.950 384.900 685.050 ;
        RECT 364.200 669.600 366.300 671.700 ;
        RECT 371.400 664.050 372.450 679.950 ;
        RECT 328.950 661.950 331.050 664.050 ;
        RECT 357.000 663.450 361.050 664.050 ;
        RECT 356.400 661.950 361.050 663.450 ;
        RECT 370.950 661.950 373.050 664.050 ;
        RECT 340.950 654.450 343.050 655.050 ;
        RECT 323.400 653.400 327.450 654.450 ;
        RECT 332.400 653.400 343.050 654.450 ;
        RECT 311.400 604.350 312.600 605.100 ;
        RECT 317.400 604.350 318.600 606.600 ;
        RECT 319.950 604.950 322.050 607.050 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 313.950 601.950 316.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 314.400 600.900 315.600 601.650 ;
        RECT 313.950 598.800 316.050 600.900 ;
        RECT 319.950 598.950 322.050 601.050 ;
        RECT 316.950 595.950 319.050 598.050 ;
        RECT 304.950 592.950 307.050 595.050 ;
        RECT 310.950 572.100 313.050 574.200 ;
        RECT 317.400 573.450 318.450 595.950 ;
        RECT 320.400 577.050 321.450 598.950 ;
        RECT 319.950 574.950 322.050 577.050 ;
        RECT 317.400 572.400 321.450 573.450 ;
        RECT 311.400 571.350 312.600 572.100 ;
        RECT 307.950 568.950 310.050 571.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 301.950 565.950 304.050 568.050 ;
        RECT 304.950 565.950 307.050 568.050 ;
        RECT 308.400 567.900 309.600 568.650 ;
        RECT 301.950 549.450 304.050 550.050 ;
        RECT 305.400 549.450 306.450 565.950 ;
        RECT 307.950 565.800 310.050 567.900 ;
        RECT 314.400 567.000 315.600 568.650 ;
        RECT 308.400 553.050 309.450 565.800 ;
        RECT 313.950 562.950 316.050 567.000 ;
        RECT 320.400 559.050 321.450 572.400 ;
        RECT 319.950 556.950 322.050 559.050 ;
        RECT 307.950 550.950 310.050 553.050 ;
        RECT 301.950 548.400 306.450 549.450 ;
        RECT 301.950 547.950 304.050 548.400 ;
        RECT 302.400 528.600 303.450 547.950 ;
        RECT 313.800 530.100 315.900 532.200 ;
        RECT 314.400 529.350 315.600 530.100 ;
        RECT 302.400 526.350 303.600 528.600 ;
        RECT 313.800 526.950 315.900 529.050 ;
        RECT 319.800 526.950 321.900 529.050 ;
        RECT 302.100 523.950 304.200 526.050 ;
        RECT 307.500 523.950 309.600 526.050 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 308.400 522.900 309.600 523.650 ;
        RECT 307.950 520.800 310.050 522.900 ;
        RECT 298.950 505.950 301.050 508.050 ;
        RECT 304.950 505.950 307.050 508.050 ;
        RECT 299.100 490.950 301.200 493.050 ;
        RECT 269.400 488.400 273.450 489.450 ;
        RECT 266.400 481.050 267.450 488.400 ;
        RECT 265.950 478.950 268.050 481.050 ;
        RECT 266.400 469.050 267.450 478.950 ;
        RECT 265.950 466.950 268.050 469.050 ;
        RECT 238.950 463.950 241.050 466.050 ;
        RECT 224.700 437.700 225.900 459.300 ;
        RECT 227.700 457.500 229.200 462.300 ;
        RECT 230.100 459.300 232.200 461.400 ;
        RECT 235.950 460.950 238.050 463.050 ;
        RECT 227.100 455.400 229.200 457.500 ;
        RECT 227.700 437.700 229.200 455.400 ;
        RECT 230.700 452.100 231.900 459.300 ;
        RECT 235.500 457.800 237.600 459.900 ;
        RECT 230.100 450.000 232.200 452.100 ;
        RECT 236.700 451.200 237.600 457.800 ;
        RECT 230.700 437.700 231.900 450.000 ;
        RECT 235.500 449.100 237.600 451.200 ;
        RECT 239.400 451.050 240.450 463.950 ;
        RECT 246.600 462.300 248.700 464.400 ;
        RECT 249.600 462.300 252.600 464.400 ;
        RECT 253.950 463.950 256.050 466.050 ;
        RECT 259.950 463.950 262.050 466.050 ;
        RECT 244.200 459.300 246.300 461.400 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 232.800 442.500 234.900 444.600 ;
        RECT 236.700 438.600 237.600 449.100 ;
        RECT 238.950 448.950 241.050 451.050 ;
        RECT 239.400 447.450 240.600 447.600 ;
        RECT 242.400 447.450 243.450 454.950 ;
        RECT 239.400 446.400 243.450 447.450 ;
        RECT 239.400 445.350 240.600 446.400 ;
        RECT 239.100 442.950 241.200 445.050 ;
        RECT 224.700 435.600 226.800 437.700 ;
        RECT 227.700 435.600 229.800 437.700 ;
        RECT 230.700 435.600 232.800 437.700 ;
        RECT 236.100 436.500 238.200 438.600 ;
        RECT 245.100 437.700 246.300 459.300 ;
        RECT 247.500 456.300 248.700 462.300 ;
        RECT 247.500 454.200 249.600 456.300 ;
        RECT 247.500 437.700 248.700 454.200 ;
        RECT 251.100 443.400 252.600 462.300 ;
        RECT 260.400 454.050 261.450 463.950 ;
        RECT 259.950 451.950 262.050 454.050 ;
        RECT 262.950 453.000 265.050 457.050 ;
        RECT 269.400 454.050 270.450 488.400 ;
        RECT 283.950 487.800 286.050 489.900 ;
        RECT 295.950 487.950 298.050 490.050 ;
        RECT 299.400 489.000 300.600 490.650 ;
        RECT 284.400 472.050 285.450 487.800 ;
        RECT 298.950 484.950 301.050 489.000 ;
        RECT 305.400 487.050 306.450 505.950 ;
        RECT 308.400 505.050 309.450 520.800 ;
        RECT 307.950 502.950 310.050 505.050 ;
        RECT 304.950 484.950 307.050 487.050 ;
        RECT 271.950 469.950 274.050 472.050 ;
        RECT 283.950 469.950 286.050 472.050 ;
        RECT 272.400 457.050 273.450 469.950 ;
        RECT 311.400 469.050 312.450 523.950 ;
        RECT 323.400 502.050 324.450 653.400 ;
        RECT 332.400 651.600 333.450 653.400 ;
        RECT 340.950 652.950 343.050 653.400 ;
        RECT 346.950 652.950 349.050 655.050 ;
        RECT 332.400 649.350 333.600 651.600 ;
        RECT 337.950 650.100 340.050 652.200 ;
        RECT 338.400 649.350 339.600 650.100 ;
        RECT 328.950 646.950 331.050 649.050 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 329.400 645.900 330.600 646.650 ;
        RECT 328.950 643.800 331.050 645.900 ;
        RECT 328.950 631.950 331.050 634.050 ;
        RECT 325.950 613.950 328.050 616.050 ;
        RECT 326.400 601.050 327.450 613.950 ;
        RECT 329.400 607.050 330.450 631.950 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 347.400 627.450 348.450 652.950 ;
        RECT 356.400 651.600 357.450 661.950 ;
        RECT 374.400 661.050 375.450 680.400 ;
        RECT 376.950 679.950 379.050 682.050 ;
        RECT 383.400 681.450 384.600 682.650 ;
        RECT 380.400 680.400 384.600 681.450 ;
        RECT 376.950 676.800 379.050 678.900 ;
        RECT 373.950 658.950 376.050 661.050 ;
        RECT 377.400 652.050 378.450 676.800 ;
        RECT 356.400 649.350 357.600 651.600 ;
        RECT 376.950 649.950 379.050 652.050 ;
        RECT 352.950 646.950 355.050 649.050 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 373.950 646.950 376.050 649.050 ;
        RECT 353.400 644.400 354.600 646.650 ;
        RECT 374.400 644.400 375.600 646.650 ;
        RECT 353.400 634.050 354.450 644.400 ;
        RECT 361.950 640.950 364.050 643.050 ;
        RECT 352.950 631.950 355.050 634.050 ;
        RECT 347.400 626.400 351.450 627.450 ;
        RECT 328.950 604.950 331.050 607.050 ;
        RECT 334.950 605.100 337.050 607.200 ;
        RECT 335.400 604.350 336.600 605.100 ;
        RECT 331.950 601.950 334.050 604.050 ;
        RECT 334.950 601.950 337.050 604.050 ;
        RECT 325.950 598.950 328.050 601.050 ;
        RECT 332.400 600.900 333.600 601.650 ;
        RECT 331.950 598.800 334.050 600.900 ;
        RECT 337.950 598.950 340.050 601.050 ;
        RECT 325.950 595.800 328.050 597.900 ;
        RECT 326.400 574.050 327.450 595.800 ;
        RECT 331.950 589.950 334.050 592.050 ;
        RECT 325.950 571.950 328.050 574.050 ;
        RECT 332.400 573.600 333.450 589.950 ;
        RECT 338.400 574.200 339.450 598.950 ;
        RECT 341.400 595.050 342.450 625.950 ;
        RECT 350.400 606.600 351.450 626.400 ;
        RECT 350.400 604.350 351.600 606.600 ;
        RECT 355.950 605.100 358.050 607.200 ;
        RECT 356.400 604.350 357.600 605.100 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 347.400 600.000 348.600 601.650 ;
        RECT 346.950 595.950 349.050 600.000 ;
        RECT 353.400 599.400 354.600 601.650 ;
        RECT 353.400 595.050 354.450 599.400 ;
        RECT 358.950 597.450 361.050 601.050 ;
        RECT 362.400 600.450 363.450 640.950 ;
        RECT 374.400 634.050 375.450 644.400 ;
        RECT 380.400 643.050 381.450 680.400 ;
        RECT 389.400 679.050 390.450 721.950 ;
        RECT 392.400 721.050 393.450 727.950 ;
        RECT 401.400 727.350 402.600 729.600 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 404.400 723.900 405.600 724.650 ;
        RECT 403.950 721.800 406.050 723.900 ;
        RECT 391.950 718.950 394.050 721.050 ;
        RECT 394.950 718.950 397.050 721.050 ;
        RECT 395.400 715.050 396.450 718.950 ;
        RECT 394.950 712.950 397.050 715.050 ;
        RECT 391.950 709.950 394.050 712.050 ;
        RECT 392.400 685.200 393.450 709.950 ;
        RECT 391.950 683.100 394.050 685.200 ;
        RECT 397.950 683.100 400.050 685.200 ;
        RECT 388.950 676.950 391.050 679.050 ;
        RECT 392.400 664.050 393.450 683.100 ;
        RECT 398.400 682.350 399.600 683.100 ;
        RECT 397.950 679.950 400.050 682.050 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 401.400 678.900 402.600 679.650 ;
        RECT 400.950 676.800 403.050 678.900 ;
        RECT 403.950 673.950 406.050 676.050 ;
        RECT 400.950 670.950 403.050 673.050 ;
        RECT 401.400 664.050 402.450 670.950 ;
        RECT 404.400 670.050 405.450 673.950 ;
        RECT 410.400 673.050 411.450 742.950 ;
        RECT 433.950 733.950 436.050 736.050 ;
        RECT 412.950 730.950 415.050 733.050 ;
        RECT 413.400 715.050 414.450 730.950 ;
        RECT 421.950 728.100 424.050 730.200 ;
        RECT 422.400 727.350 423.600 728.100 ;
        RECT 418.950 724.950 421.050 727.050 ;
        RECT 421.950 724.950 424.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 419.400 723.900 420.600 724.650 ;
        RECT 418.950 721.800 421.050 723.900 ;
        RECT 425.400 722.400 426.600 724.650 ;
        RECT 412.950 712.950 415.050 715.050 ;
        RECT 419.400 712.050 420.450 721.800 ;
        RECT 425.400 718.050 426.450 722.400 ;
        RECT 424.950 715.950 427.050 718.050 ;
        RECT 418.950 709.950 421.050 712.050 ;
        RECT 434.400 711.450 435.450 733.950 ;
        RECT 437.400 730.050 438.450 754.950 ;
        RECT 442.950 751.950 445.050 756.000 ;
        RECT 452.400 751.050 453.450 800.400 ;
        RECT 461.400 796.050 462.450 800.400 ;
        RECT 466.950 796.950 469.050 801.000 ;
        RECT 469.950 799.950 472.050 802.050 ;
        RECT 460.950 793.950 463.050 796.050 ;
        RECT 466.950 784.950 469.050 787.050 ;
        RECT 457.950 766.950 460.050 769.050 ;
        RECT 454.950 760.950 457.050 763.050 ;
        RECT 458.400 762.600 459.450 766.950 ;
        RECT 467.400 762.600 468.450 784.950 ;
        RECT 470.400 772.050 471.450 799.950 ;
        RECT 473.400 799.050 474.450 820.950 ;
        RECT 482.400 811.050 483.450 830.400 ;
        RECT 484.950 826.950 487.050 829.050 ;
        RECT 485.400 811.050 486.450 826.950 ;
        RECT 491.400 820.050 492.450 839.100 ;
        RECT 497.400 838.350 498.600 839.100 ;
        RECT 503.400 838.350 504.600 839.100 ;
        RECT 496.950 835.950 499.050 838.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 493.950 829.950 496.050 835.050 ;
        RECT 500.400 834.900 501.600 835.650 ;
        RECT 499.950 832.800 502.050 834.900 ;
        RECT 506.400 833.400 507.600 835.650 ;
        RECT 487.800 817.950 489.900 820.050 ;
        RECT 490.950 817.950 493.050 820.050 ;
        RECT 488.400 814.050 489.450 817.950 ;
        RECT 487.950 811.950 490.050 814.050 ;
        RECT 481.950 808.950 484.050 811.050 ;
        RECT 484.950 808.950 487.050 811.050 ;
        RECT 475.950 805.950 478.050 808.050 ;
        RECT 485.400 807.600 486.450 808.950 ;
        RECT 472.950 796.950 475.050 799.050 ;
        RECT 476.400 798.450 477.450 805.950 ;
        RECT 485.400 805.350 486.600 807.600 ;
        RECT 490.950 806.100 493.050 808.200 ;
        RECT 499.950 806.100 502.050 808.200 ;
        RECT 506.400 808.050 507.450 833.400 ;
        RECT 512.400 825.450 513.450 862.950 ;
        RECT 533.400 850.050 534.450 862.950 ;
        RECT 532.950 847.950 535.050 850.050 ;
        RECT 536.400 846.450 537.450 875.400 ;
        RECT 544.950 871.950 547.050 874.050 ;
        RECT 545.400 859.050 546.450 871.950 ;
        RECT 548.400 868.050 549.450 892.950 ;
        RECT 559.950 884.100 562.050 886.200 ;
        RECT 560.400 883.350 561.600 884.100 ;
        RECT 571.950 883.950 574.050 886.050 ;
        RECT 578.400 885.600 579.450 895.950 ;
        RECT 584.400 885.600 585.450 907.950 ;
        RECT 587.400 901.050 588.450 910.950 ;
        RECT 590.400 910.050 591.450 916.950 ;
        RECT 602.400 916.350 603.600 917.100 ;
        RECT 623.400 916.350 624.600 918.600 ;
        RECT 631.950 916.950 634.050 919.050 ;
        RECT 637.950 917.100 640.050 919.200 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 601.950 913.950 604.050 916.050 ;
        RECT 604.950 913.950 607.050 916.050 ;
        RECT 616.950 913.950 619.050 916.050 ;
        RECT 619.950 913.950 622.050 916.050 ;
        RECT 622.950 913.950 625.050 916.050 ;
        RECT 625.950 913.950 628.050 916.050 ;
        RECT 605.400 912.900 606.600 913.650 ;
        RECT 620.400 912.900 621.600 913.650 ;
        RECT 626.400 912.900 627.600 913.650 ;
        RECT 632.400 912.900 633.450 916.950 ;
        RECT 638.400 916.350 639.600 917.100 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 640.950 913.950 643.050 916.050 ;
        RECT 604.950 910.800 607.050 912.900 ;
        RECT 619.950 910.800 622.050 912.900 ;
        RECT 625.950 910.800 628.050 912.900 ;
        RECT 631.950 910.800 634.050 912.900 ;
        RECT 641.400 911.400 642.600 913.650 ;
        RECT 647.400 913.050 648.450 922.950 ;
        RECT 676.950 917.100 679.050 919.200 ;
        RECT 683.400 918.600 684.450 922.950 ;
        RECT 677.400 916.350 678.600 917.100 ;
        RECT 683.400 916.350 684.600 918.600 ;
        RECT 688.950 917.100 691.050 919.200 ;
        RECT 698.400 918.600 699.450 925.950 ;
        RECT 712.950 922.950 715.050 925.050 ;
        RECT 718.950 922.950 721.050 925.050 ;
        RECT 751.950 922.950 754.050 925.050 ;
        RECT 769.950 922.950 772.050 925.050 ;
        RECT 778.950 922.950 781.050 925.050 ;
        RECT 784.950 924.450 787.050 925.050 ;
        RECT 790.950 924.450 793.050 925.050 ;
        RECT 784.950 923.400 793.050 924.450 ;
        RECT 784.950 922.950 787.050 923.400 ;
        RECT 790.950 922.950 793.050 923.400 ;
        RECT 656.400 913.950 658.500 916.050 ;
        RECT 661.500 913.950 663.600 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 676.950 913.950 679.050 916.050 ;
        RECT 679.950 913.950 682.050 916.050 ;
        RECT 682.950 913.950 685.050 916.050 ;
        RECT 589.950 907.950 592.050 910.050 ;
        RECT 595.950 904.950 598.050 907.050 ;
        RECT 586.950 898.950 589.050 901.050 ;
        RECT 556.950 880.950 559.050 883.050 ;
        RECT 559.950 880.950 562.050 883.050 ;
        RECT 562.950 880.950 565.050 883.050 ;
        RECT 557.400 879.450 558.600 880.650 ;
        RECT 554.400 878.400 558.600 879.450 ;
        RECT 554.400 874.050 555.450 878.400 ;
        RECT 565.950 874.950 568.050 877.050 ;
        RECT 553.950 871.950 556.050 874.050 ;
        RECT 547.950 865.950 550.050 868.050 ;
        RECT 566.400 865.050 567.450 874.950 ;
        RECT 565.950 862.950 568.050 865.050 ;
        RECT 572.400 859.050 573.450 883.950 ;
        RECT 578.400 883.350 579.600 885.600 ;
        RECT 584.400 883.350 585.600 885.600 ;
        RECT 577.950 880.950 580.050 883.050 ;
        RECT 580.950 880.950 583.050 883.050 ;
        RECT 583.950 880.950 586.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 581.400 879.000 582.600 880.650 ;
        RECT 587.400 879.900 588.600 880.650 ;
        RECT 580.950 874.950 583.050 879.000 ;
        RECT 586.950 877.800 589.050 879.900 ;
        RECT 596.400 877.050 597.450 904.950 ;
        RECT 610.950 898.950 613.050 901.050 ;
        RECT 604.950 889.950 607.050 892.050 ;
        RECT 605.400 886.200 606.450 889.950 ;
        RECT 604.950 884.100 607.050 886.200 ;
        RECT 611.400 885.600 612.450 898.950 ;
        RECT 628.950 889.950 631.050 892.050 ;
        RECT 605.400 883.350 606.600 884.100 ;
        RECT 611.400 883.350 612.600 885.600 ;
        RECT 616.950 884.100 619.050 886.200 ;
        RECT 622.950 884.100 625.050 886.200 ;
        RECT 629.400 885.600 630.450 889.950 ;
        RECT 632.400 889.050 633.450 910.800 ;
        RECT 641.400 898.050 642.450 911.400 ;
        RECT 646.950 910.950 649.050 913.050 ;
        RECT 656.400 912.900 657.600 913.650 ;
        RECT 647.400 907.050 648.450 910.950 ;
        RECT 655.950 910.800 658.050 912.900 ;
        RECT 674.400 911.400 675.600 913.650 ;
        RECT 680.400 912.900 681.600 913.650 ;
        RECT 689.400 913.050 690.450 917.100 ;
        RECT 698.400 916.350 699.600 918.600 ;
        RECT 703.950 917.100 706.050 919.200 ;
        RECT 704.400 916.350 705.600 917.100 ;
        RECT 697.950 913.950 700.050 916.050 ;
        RECT 700.950 913.950 703.050 916.050 ;
        RECT 703.950 913.950 706.050 916.050 ;
        RECT 706.950 913.950 709.050 916.050 ;
        RECT 646.950 904.950 649.050 907.050 ;
        RECT 674.400 904.050 675.450 911.400 ;
        RECT 679.950 910.800 682.050 912.900 ;
        RECT 688.950 910.950 691.050 913.050 ;
        RECT 701.400 912.900 702.600 913.650 ;
        RECT 673.950 901.950 676.050 904.050 ;
        RECT 680.400 898.050 681.450 910.800 ;
        RECT 640.950 895.950 643.050 898.050 ;
        RECT 679.950 895.950 682.050 898.050 ;
        RECT 640.950 889.950 643.050 892.050 ;
        RECT 649.950 889.950 652.050 892.050 ;
        RECT 631.950 886.950 634.050 889.050 ;
        RECT 637.950 886.950 640.050 889.050 ;
        RECT 601.950 880.950 604.050 883.050 ;
        RECT 604.950 880.950 607.050 883.050 ;
        RECT 607.950 880.950 610.050 883.050 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 602.400 878.400 603.600 880.650 ;
        RECT 608.400 878.400 609.600 880.650 ;
        RECT 595.950 874.950 598.050 877.050 ;
        RECT 586.950 871.950 589.050 874.050 ;
        RECT 583.950 865.950 586.050 868.050 ;
        RECT 544.950 856.950 547.050 859.050 ;
        RECT 565.950 856.950 568.050 859.050 ;
        RECT 571.950 856.950 574.050 859.050 ;
        RECT 533.400 845.400 537.450 846.450 ;
        RECT 523.950 839.100 526.050 841.200 ;
        RECT 524.400 838.350 525.600 839.100 ;
        RECT 520.950 835.950 523.050 838.050 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 527.400 834.900 528.600 835.650 ;
        RECT 526.950 832.800 529.050 834.900 ;
        RECT 533.400 832.050 534.450 845.400 ;
        RECT 538.950 839.100 541.050 841.200 ;
        RECT 545.400 841.050 546.450 856.950 ;
        RECT 566.400 850.050 567.450 856.950 ;
        RECT 547.950 847.950 550.050 850.050 ;
        RECT 539.400 838.350 540.600 839.100 ;
        RECT 544.950 838.950 547.050 841.050 ;
        RECT 538.950 835.950 541.050 838.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 542.400 835.050 543.600 835.650 ;
        RECT 542.400 833.400 547.050 835.050 ;
        RECT 543.000 832.950 547.050 833.400 ;
        RECT 548.400 832.050 549.450 847.950 ;
        RECT 562.800 847.800 564.900 849.900 ;
        RECT 565.950 847.950 568.050 850.050 ;
        RECT 563.400 844.050 564.450 847.800 ;
        RECT 572.400 847.050 573.450 856.950 ;
        RECT 571.950 844.950 574.050 847.050 ;
        RECT 580.950 844.950 583.050 847.050 ;
        RECT 562.950 841.950 565.050 844.050 ;
        RECT 553.950 839.100 556.050 841.200 ;
        RECT 559.950 839.100 562.050 841.200 ;
        RECT 574.950 840.000 577.050 844.050 ;
        RECT 581.400 840.600 582.450 844.950 ;
        RECT 584.400 841.050 585.450 865.950 ;
        RECT 587.400 862.050 588.450 871.950 ;
        RECT 589.950 862.950 592.050 865.050 ;
        RECT 586.950 859.950 589.050 862.050 ;
        RECT 554.400 838.350 555.600 839.100 ;
        RECT 560.400 838.350 561.600 839.100 ;
        RECT 575.400 838.350 576.600 840.000 ;
        RECT 581.400 838.350 582.600 840.600 ;
        RECT 583.950 838.950 586.050 841.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 556.950 835.950 559.050 838.050 ;
        RECT 559.950 835.950 562.050 838.050 ;
        RECT 571.950 835.950 574.050 838.050 ;
        RECT 574.950 835.950 577.050 838.050 ;
        RECT 577.950 835.950 580.050 838.050 ;
        RECT 580.950 835.950 583.050 838.050 ;
        RECT 550.950 832.950 553.050 835.050 ;
        RECT 557.400 834.000 558.600 835.650 ;
        RECT 526.950 829.650 529.050 831.750 ;
        RECT 532.950 829.950 535.050 832.050 ;
        RECT 547.950 829.950 550.050 832.050 ;
        RECT 512.400 824.400 516.450 825.450 ;
        RECT 508.950 814.950 511.050 817.050 ;
        RECT 491.400 805.350 492.600 806.100 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 482.400 801.000 483.600 802.650 ;
        RECT 488.400 801.900 489.600 802.650 ;
        RECT 476.400 797.400 480.450 798.450 ;
        RECT 473.400 790.050 474.450 796.950 ;
        RECT 475.950 793.950 478.050 796.050 ;
        RECT 472.950 787.950 475.050 790.050 ;
        RECT 469.950 769.950 472.050 772.050 ;
        RECT 451.950 748.950 454.050 751.050 ;
        RECT 455.400 742.050 456.450 760.950 ;
        RECT 458.400 760.350 459.600 762.600 ;
        RECT 467.400 760.350 468.600 762.600 ;
        RECT 458.100 757.950 460.200 760.050 ;
        RECT 461.400 757.950 463.500 760.050 ;
        RECT 466.800 757.950 468.900 760.050 ;
        RECT 461.400 755.400 462.600 757.650 ;
        RECT 461.400 745.050 462.450 755.400 ;
        RECT 460.950 742.950 463.050 745.050 ;
        RECT 454.950 739.950 457.050 742.050 ;
        RECT 448.950 733.950 451.050 736.050 ;
        RECT 436.950 727.950 439.050 730.050 ;
        RECT 442.950 728.100 445.050 730.200 ;
        RECT 449.400 729.600 450.450 733.950 ;
        RECT 443.400 727.350 444.600 728.100 ;
        RECT 449.400 727.350 450.600 729.600 ;
        RECT 454.950 727.950 457.050 730.050 ;
        RECT 463.950 728.100 466.050 730.200 ;
        RECT 439.950 724.950 442.050 727.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 440.400 723.900 441.600 724.650 ;
        RECT 446.400 723.900 447.600 724.650 ;
        RECT 439.950 721.800 442.050 723.900 ;
        RECT 445.950 721.800 448.050 723.900 ;
        RECT 441.000 720.450 445.050 721.050 ;
        RECT 440.400 718.950 445.050 720.450 ;
        RECT 436.950 711.450 439.050 712.050 ;
        RECT 434.400 710.400 439.050 711.450 ;
        RECT 436.950 709.950 439.050 710.400 ;
        RECT 424.950 706.950 427.050 709.050 ;
        RECT 421.950 700.950 424.050 703.050 ;
        RECT 422.400 694.050 423.450 700.950 ;
        RECT 425.400 700.050 426.450 706.950 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 421.950 691.950 424.050 694.050 ;
        RECT 424.950 684.000 427.050 688.050 ;
        RECT 433.950 685.950 436.050 688.050 ;
        RECT 425.400 682.350 426.600 684.000 ;
        RECT 418.950 679.950 421.050 682.050 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 427.950 679.950 430.050 682.050 ;
        RECT 412.950 673.950 415.050 679.050 ;
        RECT 422.400 678.900 423.600 679.650 ;
        RECT 428.400 678.900 429.600 679.650 ;
        RECT 421.950 676.800 424.050 678.900 ;
        RECT 427.950 676.800 430.050 678.900 ;
        RECT 434.400 673.050 435.450 685.950 ;
        RECT 409.950 670.950 412.050 673.050 ;
        RECT 418.950 670.950 421.050 673.050 ;
        RECT 433.950 670.950 436.050 673.050 ;
        RECT 403.950 667.950 406.050 670.050 ;
        RECT 412.950 664.950 415.050 667.050 ;
        RECT 391.950 661.950 394.050 664.050 ;
        RECT 397.800 661.950 399.900 664.050 ;
        RECT 400.950 661.950 403.050 664.050 ;
        RECT 409.950 661.950 412.050 664.050 ;
        RECT 388.950 650.100 391.050 652.200 ;
        RECT 389.400 649.350 390.600 650.100 ;
        RECT 385.950 646.950 388.050 649.050 ;
        RECT 388.950 646.950 391.050 649.050 ;
        RECT 391.950 646.950 394.050 649.050 ;
        RECT 386.400 645.000 387.600 646.650 ;
        RECT 379.950 640.950 382.050 643.050 ;
        RECT 385.950 640.950 388.050 645.000 ;
        RECT 392.400 644.400 393.600 646.650 ;
        RECT 398.400 645.450 399.450 661.950 ;
        RECT 400.950 649.950 403.050 652.050 ;
        RECT 410.400 651.600 411.450 661.950 ;
        RECT 413.400 661.050 414.450 664.950 ;
        RECT 415.950 661.950 418.050 664.050 ;
        RECT 412.950 658.950 415.050 661.050 ;
        RECT 416.400 651.600 417.450 661.950 ;
        RECT 419.400 661.050 420.450 670.950 ;
        RECT 421.950 667.950 424.050 670.050 ;
        RECT 422.400 661.050 423.450 667.950 ;
        RECT 418.950 658.950 421.050 661.050 ;
        RECT 421.950 658.950 424.050 661.050 ;
        RECT 424.950 658.950 427.050 661.050 ;
        RECT 401.400 645.900 402.450 649.950 ;
        RECT 410.400 649.350 411.600 651.600 ;
        RECT 416.400 649.350 417.600 651.600 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 421.950 646.950 424.050 649.050 ;
        RECT 407.400 645.900 408.600 646.650 ;
        RECT 395.400 644.400 399.450 645.450 ;
        RECT 392.400 640.050 393.450 644.400 ;
        RECT 391.950 637.950 394.050 640.050 ;
        RECT 373.950 631.950 376.050 634.050 ;
        RECT 391.950 631.950 394.050 634.050 ;
        RECT 364.950 628.950 367.050 631.050 ;
        RECT 365.400 607.050 366.450 628.950 ;
        RECT 367.950 619.950 370.050 622.050 ;
        RECT 364.950 604.950 367.050 607.050 ;
        RECT 368.400 606.600 369.450 619.950 ;
        RECT 392.400 610.200 393.450 631.950 ;
        RECT 395.400 631.050 396.450 644.400 ;
        RECT 400.950 643.800 403.050 645.900 ;
        RECT 406.950 643.800 409.050 645.900 ;
        RECT 413.400 644.400 414.600 646.650 ;
        RECT 397.950 640.950 400.050 643.050 ;
        RECT 398.400 634.050 399.450 640.950 ;
        RECT 413.400 640.050 414.450 644.400 ;
        RECT 412.950 637.950 415.050 640.050 ;
        RECT 397.950 633.450 400.050 634.050 ;
        RECT 397.950 632.400 402.450 633.450 ;
        RECT 397.950 631.950 400.050 632.400 ;
        RECT 394.950 628.950 397.050 631.050 ;
        RECT 397.950 610.950 400.050 613.050 ;
        RECT 391.950 608.100 394.050 610.200 ;
        RECT 368.400 604.350 369.600 606.600 ;
        RECT 373.950 605.100 376.050 607.200 ;
        RECT 374.400 604.350 375.600 605.100 ;
        RECT 382.950 604.950 388.050 607.050 ;
        RECT 391.950 604.950 394.050 607.050 ;
        RECT 398.400 606.600 399.450 610.950 ;
        RECT 401.400 607.050 402.450 632.400 ;
        RECT 409.950 628.950 412.050 631.050 ;
        RECT 403.950 622.950 406.050 625.050 ;
        RECT 392.400 604.350 393.600 604.950 ;
        RECT 398.400 604.350 399.600 606.600 ;
        RECT 400.950 604.950 403.050 607.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 376.950 601.950 379.050 604.050 ;
        RECT 371.400 600.900 372.600 601.650 ;
        RECT 377.400 601.050 378.600 601.650 ;
        RECT 362.400 599.400 366.450 600.450 ;
        RECT 356.400 597.000 361.050 597.450 ;
        RECT 356.400 596.400 360.450 597.000 ;
        RECT 340.950 592.950 343.050 595.050 ;
        RECT 352.950 592.950 355.050 595.050 ;
        RECT 349.950 589.950 352.050 592.050 ;
        RECT 346.950 580.950 349.050 583.050 ;
        RECT 343.950 577.950 346.050 580.050 ;
        RECT 332.400 571.350 333.600 573.600 ;
        RECT 337.950 572.100 340.050 574.200 ;
        RECT 338.400 571.350 339.600 572.100 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 325.950 565.950 328.050 568.050 ;
        RECT 329.400 567.900 330.600 568.650 ;
        RECT 326.400 562.050 327.450 565.950 ;
        RECT 328.950 565.800 331.050 567.900 ;
        RECT 335.400 567.000 336.600 568.650 ;
        RECT 334.950 562.950 337.050 567.000 ;
        RECT 340.950 565.950 343.050 568.050 ;
        RECT 325.950 559.950 328.050 562.050 ;
        RECT 341.400 556.050 342.450 565.950 ;
        RECT 340.950 553.950 343.050 556.050 ;
        RECT 344.400 544.050 345.450 577.950 ;
        RECT 347.400 556.050 348.450 580.950 ;
        RECT 350.400 574.050 351.450 589.950 ;
        RECT 356.400 583.050 357.450 596.400 ;
        RECT 355.950 580.950 358.050 583.050 ;
        RECT 358.950 577.950 361.050 580.050 ;
        RECT 349.950 571.950 352.050 574.050 ;
        RECT 352.950 572.100 355.050 574.200 ;
        RECT 359.400 573.600 360.450 577.950 ;
        RECT 365.400 574.050 366.450 599.400 ;
        RECT 370.950 598.800 373.050 600.900 ;
        RECT 377.400 598.950 382.050 601.050 ;
        RECT 382.950 600.450 385.050 603.900 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 389.400 600.900 390.600 601.650 ;
        RECT 395.400 600.900 396.600 601.650 ;
        RECT 382.950 600.000 387.450 600.450 ;
        RECT 383.400 599.400 387.450 600.000 ;
        RECT 377.400 592.050 378.450 598.950 ;
        RECT 386.400 597.450 387.450 599.400 ;
        RECT 388.950 598.800 391.050 600.900 ;
        RECT 394.950 598.800 397.050 600.900 ;
        RECT 404.400 598.050 405.450 622.950 ;
        RECT 410.400 613.050 411.450 628.950 ;
        RECT 413.400 616.050 414.450 637.950 ;
        RECT 418.950 634.950 421.050 637.050 ;
        RECT 412.950 613.950 415.050 616.050 ;
        RECT 409.950 610.950 412.050 613.050 ;
        RECT 413.400 610.050 414.450 613.950 ;
        RECT 419.400 613.050 420.450 634.950 ;
        RECT 422.400 622.050 423.450 646.950 ;
        RECT 425.400 645.450 426.450 658.950 ;
        RECT 433.950 651.000 436.050 655.050 ;
        RECT 434.400 649.350 435.600 651.000 ;
        RECT 428.100 646.950 430.200 649.050 ;
        RECT 433.500 646.950 435.600 649.050 ;
        RECT 428.400 645.450 429.600 646.650 ;
        RECT 425.400 644.400 429.600 645.450 ;
        RECT 424.950 640.950 427.050 643.050 ;
        RECT 421.950 619.950 424.050 622.050 ;
        RECT 418.950 610.950 421.050 613.050 ;
        RECT 425.400 610.050 426.450 640.950 ;
        RECT 437.400 633.450 438.450 709.950 ;
        RECT 440.400 637.050 441.450 718.950 ;
        RECT 446.400 718.050 447.450 721.800 ;
        RECT 455.400 721.050 456.450 727.950 ;
        RECT 464.400 727.350 465.600 728.100 ;
        RECT 461.100 724.950 463.200 727.050 ;
        RECT 464.400 724.950 466.500 727.050 ;
        RECT 469.800 724.950 471.900 727.050 ;
        RECT 461.400 723.900 462.600 724.650 ;
        RECT 460.950 721.800 463.050 723.900 ;
        RECT 470.400 722.400 471.600 724.650 ;
        RECT 448.950 718.950 451.050 721.050 ;
        RECT 454.950 718.950 457.050 721.050 ;
        RECT 445.950 715.950 448.050 718.050 ;
        RECT 442.950 714.450 445.050 715.050 ;
        RECT 449.400 714.450 450.450 718.950 ;
        RECT 470.400 715.050 471.450 722.400 ;
        RECT 442.950 713.400 450.450 714.450 ;
        RECT 442.950 712.950 445.050 713.400 ;
        RECT 469.950 712.950 472.050 715.050 ;
        RECT 473.400 712.050 474.450 787.950 ;
        RECT 476.400 778.050 477.450 793.950 ;
        RECT 479.400 793.050 480.450 797.400 ;
        RECT 481.950 796.950 484.050 801.000 ;
        RECT 487.950 799.800 490.050 801.900 ;
        RECT 494.400 800.400 495.600 802.650 ;
        RECT 478.950 790.950 481.050 793.050 ;
        RECT 475.950 775.950 478.050 778.050 ;
        RECT 478.950 769.950 481.050 772.050 ;
        RECT 479.400 763.200 480.450 769.950 ;
        RECT 494.400 766.050 495.450 800.400 ;
        RECT 496.950 784.950 499.050 787.050 ;
        RECT 493.950 763.950 496.050 766.050 ;
        RECT 478.950 761.100 481.050 763.200 ;
        RECT 484.950 761.100 487.050 763.200 ;
        RECT 493.950 762.450 496.050 762.900 ;
        RECT 497.400 762.450 498.450 784.950 ;
        RECT 500.400 784.050 501.450 806.100 ;
        RECT 505.950 805.950 508.050 808.050 ;
        RECT 509.400 807.600 510.450 814.950 ;
        RECT 515.400 807.600 516.450 824.400 ;
        RECT 523.950 817.950 526.050 820.050 ;
        RECT 520.950 808.950 523.050 814.050 ;
        RECT 509.400 805.350 510.600 807.600 ;
        RECT 515.400 805.350 516.600 807.600 ;
        RECT 508.950 802.950 511.050 805.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 505.950 799.950 508.050 802.050 ;
        RECT 512.400 801.000 513.600 802.650 ;
        RECT 518.400 802.050 519.600 802.650 ;
        RECT 499.950 781.950 502.050 784.050 ;
        RECT 500.400 769.050 501.450 781.950 ;
        RECT 506.400 771.450 507.450 799.950 ;
        RECT 508.950 796.950 511.050 799.050 ;
        RECT 511.950 796.950 514.050 801.000 ;
        RECT 518.400 800.400 523.050 802.050 ;
        RECT 519.000 799.950 523.050 800.400 ;
        RECT 514.950 796.950 517.050 799.050 ;
        RECT 509.400 790.050 510.450 796.950 ;
        RECT 508.950 787.950 511.050 790.050 ;
        RECT 515.400 787.050 516.450 796.950 ;
        RECT 520.950 796.800 523.050 798.900 ;
        RECT 521.400 793.050 522.450 796.800 ;
        RECT 520.950 790.950 523.050 793.050 ;
        RECT 517.950 789.900 522.000 790.050 ;
        RECT 517.950 787.950 523.050 789.900 ;
        RECT 520.950 787.800 523.050 787.950 ;
        RECT 514.950 784.950 517.050 787.050 ;
        RECT 520.950 784.800 523.050 786.900 ;
        RECT 517.950 772.950 520.050 775.050 ;
        RECT 508.950 771.450 511.050 772.050 ;
        RECT 506.400 770.400 511.050 771.450 ;
        RECT 508.950 769.950 511.050 770.400 ;
        RECT 499.950 766.950 502.050 769.050 ;
        RECT 505.950 766.800 508.050 768.900 ;
        RECT 493.950 761.400 498.450 762.450 ;
        RECT 506.400 762.450 507.450 766.800 ;
        RECT 509.400 766.050 510.450 769.950 ;
        RECT 508.950 763.950 511.050 766.050 ;
        RECT 518.400 762.600 519.450 772.950 ;
        RECT 521.400 769.050 522.450 784.800 ;
        RECT 524.400 781.050 525.450 817.950 ;
        RECT 523.950 778.950 526.050 781.050 ;
        RECT 527.400 778.050 528.450 829.650 ;
        RECT 551.400 820.050 552.450 832.950 ;
        RECT 556.950 829.950 559.050 834.000 ;
        RECT 562.950 832.950 565.050 835.050 ;
        RECT 572.400 833.400 573.600 835.650 ;
        RECT 578.400 834.900 579.600 835.650 ;
        RECT 563.400 826.050 564.450 832.950 ;
        RECT 568.950 826.950 571.050 829.050 ;
        RECT 562.950 823.950 565.050 826.050 ;
        RECT 550.800 817.950 552.900 820.050 ;
        RECT 529.950 811.950 532.050 814.050 ;
        RECT 559.950 811.950 562.050 814.050 ;
        RECT 530.400 808.050 531.450 811.950 ;
        RECT 532.950 811.050 535.050 811.200 ;
        RECT 535.950 811.050 538.050 811.200 ;
        RECT 532.950 809.100 538.050 811.050 ;
        RECT 534.000 808.950 537.000 809.100 ;
        RECT 529.950 805.950 532.050 808.050 ;
        RECT 535.950 805.950 538.050 808.050 ;
        RECT 541.950 807.000 544.050 811.050 ;
        RECT 536.400 805.350 537.600 805.950 ;
        RECT 542.400 805.350 543.600 807.000 ;
        RECT 550.950 806.100 553.050 808.200 ;
        RECT 560.400 807.600 561.450 811.950 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 544.950 802.950 547.050 805.050 ;
        RECT 533.400 801.000 534.600 802.650 ;
        RECT 539.400 801.900 540.600 802.650 ;
        RECT 532.950 796.950 535.050 801.000 ;
        RECT 538.950 799.800 541.050 801.900 ;
        RECT 545.400 801.000 546.600 802.650 ;
        RECT 544.950 798.450 547.050 801.000 ;
        RECT 542.400 797.400 547.050 798.450 ;
        RECT 529.950 784.950 532.050 790.050 ;
        RECT 526.950 775.950 529.050 778.050 ;
        RECT 532.950 775.950 535.050 778.050 ;
        RECT 529.950 772.950 532.050 775.050 ;
        RECT 520.950 766.950 523.050 769.050 ;
        RECT 506.400 761.400 510.450 762.450 ;
        RECT 479.400 760.350 480.600 761.100 ;
        RECT 485.400 760.350 486.600 761.100 ;
        RECT 493.950 760.800 496.050 761.400 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 481.950 757.950 484.050 760.050 ;
        RECT 484.950 757.950 487.050 760.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 482.400 755.400 483.600 757.650 ;
        RECT 488.400 757.050 489.600 757.650 ;
        RECT 494.400 757.050 495.450 760.800 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 502.950 757.950 505.050 760.050 ;
        RECT 488.400 755.400 493.050 757.050 ;
        RECT 478.950 751.950 481.050 754.050 ;
        RECT 475.950 728.100 478.050 730.200 ;
        RECT 457.950 709.950 460.050 712.050 ;
        RECT 472.950 709.950 475.050 712.050 ;
        RECT 454.950 706.950 457.050 709.050 ;
        RECT 442.950 703.950 445.050 706.050 ;
        RECT 448.950 703.950 451.050 706.050 ;
        RECT 443.400 684.600 444.450 703.950 ;
        RECT 449.400 700.050 450.450 703.950 ;
        RECT 448.950 697.950 451.050 700.050 ;
        RECT 451.950 694.950 454.050 697.050 ;
        RECT 452.400 685.200 453.450 694.950 ;
        RECT 455.400 694.050 456.450 706.950 ;
        RECT 454.950 691.950 457.050 694.050 ;
        RECT 443.400 682.350 444.600 684.600 ;
        RECT 451.950 683.100 454.050 685.200 ;
        RECT 452.400 682.350 453.600 683.100 ;
        RECT 443.100 679.950 445.200 682.050 ;
        RECT 446.400 679.950 448.500 682.050 ;
        RECT 451.800 679.950 453.900 682.050 ;
        RECT 446.400 677.400 447.600 679.650 ;
        RECT 455.400 679.050 456.450 691.950 ;
        RECT 442.950 673.950 445.050 676.050 ;
        RECT 439.950 634.950 442.050 637.050 ;
        RECT 443.400 634.050 444.450 673.950 ;
        RECT 446.400 673.050 447.450 677.400 ;
        RECT 454.950 676.950 457.050 679.050 ;
        RECT 445.950 670.950 448.050 673.050 ;
        RECT 447.000 666.450 451.050 667.050 ;
        RECT 446.400 666.000 451.050 666.450 ;
        RECT 445.950 664.950 451.050 666.000 ;
        RECT 445.950 661.950 448.050 664.950 ;
        RECT 448.950 646.950 451.050 649.050 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 452.400 645.000 453.600 646.650 ;
        RECT 451.950 640.950 454.050 645.000 ;
        RECT 454.950 643.950 457.050 646.050 ;
        RECT 448.950 634.950 451.050 637.050 ;
        RECT 437.400 632.400 441.450 633.450 ;
        RECT 433.950 613.950 436.050 616.050 ;
        RECT 427.950 610.950 430.050 613.050 ;
        RECT 406.950 607.950 409.050 610.050 ;
        RECT 412.950 607.950 415.050 610.050 ;
        RECT 386.400 596.400 390.450 597.450 ;
        RECT 376.950 589.950 379.050 592.050 ;
        RECT 385.950 577.950 388.050 580.050 ;
        RECT 353.400 571.350 354.600 572.100 ;
        RECT 359.400 571.350 360.600 573.600 ;
        RECT 364.950 571.950 367.050 574.050 ;
        RECT 367.950 571.950 370.050 574.050 ;
        RECT 376.950 572.100 379.050 574.200 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 355.950 568.950 358.050 571.050 ;
        RECT 358.950 568.950 361.050 571.050 ;
        RECT 361.950 568.950 364.050 571.050 ;
        RECT 356.400 566.400 357.600 568.650 ;
        RECT 362.400 567.900 363.600 568.650 ;
        RECT 356.400 564.300 357.450 566.400 ;
        RECT 361.950 565.800 364.050 567.900 ;
        RECT 364.950 565.950 367.050 568.050 ;
        RECT 368.400 567.900 369.450 571.950 ;
        RECT 377.400 571.350 378.600 572.100 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 376.950 568.950 379.050 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 361.950 564.300 364.050 564.750 ;
        RECT 356.400 563.250 364.050 564.300 ;
        RECT 346.950 553.950 349.050 556.050 ;
        RECT 356.400 550.050 357.450 563.250 ;
        RECT 361.950 562.650 364.050 563.250 ;
        RECT 365.400 550.050 366.450 565.950 ;
        RECT 367.950 565.800 370.050 567.900 ;
        RECT 374.400 567.000 375.600 568.650 ;
        RECT 373.950 562.950 376.050 567.000 ;
        RECT 380.400 566.400 381.600 568.650 ;
        RECT 380.400 565.050 381.450 566.400 ;
        RECT 382.950 565.950 385.050 568.050 ;
        RECT 379.950 564.450 382.050 565.050 ;
        RECT 377.400 563.400 382.050 564.450 ;
        RECT 367.950 550.950 370.050 553.050 ;
        RECT 355.800 547.950 357.900 550.050 ;
        RECT 358.950 547.950 361.050 550.050 ;
        RECT 364.950 547.950 367.050 550.050 ;
        RECT 326.400 540.300 329.400 542.400 ;
        RECT 330.300 540.300 332.400 542.400 ;
        RECT 337.950 541.950 340.050 544.050 ;
        RECT 343.950 541.950 346.050 544.050 ;
        RECT 326.400 521.400 327.900 540.300 ;
        RECT 330.300 534.300 331.500 540.300 ;
        RECT 329.400 532.200 331.500 534.300 ;
        RECT 326.400 519.300 328.500 521.400 ;
        RECT 327.300 515.700 328.500 519.300 ;
        RECT 330.300 515.700 331.500 532.200 ;
        RECT 332.700 537.300 334.800 539.400 ;
        RECT 332.700 515.700 333.900 537.300 ;
        RECT 338.400 525.600 339.450 541.950 ;
        RECT 349.200 540.300 351.300 542.400 ;
        RECT 341.400 535.800 343.500 537.900 ;
        RECT 346.800 537.300 348.900 539.400 ;
        RECT 341.400 529.200 342.300 535.800 ;
        RECT 347.100 530.100 348.300 537.300 ;
        RECT 349.800 535.500 351.300 540.300 ;
        RECT 352.200 537.300 354.300 542.400 ;
        RECT 349.800 533.400 351.900 535.500 ;
        RECT 341.400 527.100 343.500 529.200 ;
        RECT 346.800 528.000 348.900 530.100 ;
        RECT 338.400 523.350 339.600 525.600 ;
        RECT 337.800 520.950 339.900 523.050 ;
        RECT 341.400 516.600 342.300 527.100 ;
        RECT 344.100 520.500 346.200 522.600 ;
        RECT 326.700 513.600 328.800 515.700 ;
        RECT 329.700 513.600 331.800 515.700 ;
        RECT 332.700 513.600 334.800 515.700 ;
        RECT 340.800 514.500 342.900 516.600 ;
        RECT 347.100 515.700 348.300 528.000 ;
        RECT 349.800 515.700 351.300 533.400 ;
        RECT 353.100 515.700 354.300 537.300 ;
        RECT 346.200 513.600 348.300 515.700 ;
        RECT 349.200 513.600 351.300 515.700 ;
        RECT 352.200 513.600 354.300 515.700 ;
        RECT 355.200 540.300 357.300 542.400 ;
        RECT 355.200 535.500 356.700 540.300 ;
        RECT 355.200 533.400 357.300 535.500 ;
        RECT 355.200 515.700 356.700 533.400 ;
        RECT 355.200 513.600 357.300 515.700 ;
        RECT 349.950 508.950 352.050 511.050 ;
        RECT 322.950 499.950 325.050 502.050 ;
        RECT 343.950 499.950 346.050 502.050 ;
        RECT 317.100 490.950 319.200 493.050 ;
        RECT 337.800 490.950 339.900 493.050 ;
        RECT 344.400 487.050 345.450 499.950 ;
        RECT 343.950 484.950 346.050 487.050 ;
        RECT 334.950 475.950 337.050 478.050 ;
        RECT 310.950 466.950 313.050 469.050 ;
        RECT 316.950 466.950 319.050 469.050 ;
        RECT 284.400 462.300 287.400 464.400 ;
        RECT 288.300 462.300 290.400 464.400 ;
        RECT 307.200 462.300 309.300 464.400 ;
        RECT 271.950 454.950 274.050 457.050 ;
        RECT 263.400 451.350 264.600 453.000 ;
        RECT 268.950 451.950 271.050 454.050 ;
        RECT 272.400 453.600 273.450 454.950 ;
        RECT 272.400 451.350 273.600 453.600 ;
        RECT 257.100 448.950 259.200 451.050 ;
        RECT 263.100 448.950 265.200 451.050 ;
        RECT 271.800 448.950 273.900 451.050 ;
        RECT 277.800 448.950 279.900 451.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 250.500 441.300 252.600 443.400 ;
        RECT 250.500 437.700 251.700 441.300 ;
        RECT 244.200 435.600 246.300 437.700 ;
        RECT 247.200 435.600 249.300 437.700 ;
        RECT 250.200 435.600 252.300 437.700 ;
        RECT 250.950 427.950 253.050 430.050 ;
        RECT 232.950 424.950 235.050 427.050 ;
        RECT 229.950 415.950 232.050 418.050 ;
        RECT 226.800 412.950 228.900 415.050 ;
        RECT 230.400 412.050 231.450 415.950 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 229.950 406.800 232.050 408.900 ;
        RECT 223.950 394.950 226.050 397.050 ;
        RECT 220.950 385.950 223.050 388.050 ;
        RECT 217.950 382.950 220.050 385.050 ;
        RECT 217.950 376.950 220.050 379.050 ;
        RECT 208.950 373.950 211.050 376.050 ;
        RECT 205.950 370.950 208.050 373.050 ;
        RECT 211.950 371.100 214.050 373.200 ;
        RECT 218.400 373.050 219.450 376.950 ;
        RECT 206.400 358.050 207.450 370.950 ;
        RECT 212.400 370.350 213.600 371.100 ;
        RECT 217.950 370.950 220.050 373.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 215.400 366.450 216.600 367.650 ;
        RECT 221.400 366.450 222.450 385.950 ;
        RECT 215.400 365.400 222.450 366.450 ;
        RECT 211.950 361.950 214.050 364.050 ;
        RECT 217.950 361.950 220.050 364.050 ;
        RECT 220.950 361.950 223.050 364.050 ;
        RECT 212.400 358.050 213.450 361.950 ;
        RECT 205.950 355.950 208.050 358.050 ;
        RECT 211.950 355.950 214.050 358.050 ;
        RECT 208.950 349.950 211.050 352.050 ;
        RECT 202.950 337.950 205.050 340.050 ;
        RECT 209.400 339.600 210.450 349.950 ;
        RECT 218.400 346.050 219.450 361.950 ;
        RECT 217.950 343.950 220.050 346.050 ;
        RECT 209.400 337.350 210.600 339.600 ;
        RECT 217.950 337.950 220.050 340.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 206.400 332.400 207.600 334.650 ;
        RECT 212.400 333.000 213.600 334.650 ;
        RECT 199.950 328.950 202.050 331.050 ;
        RECT 206.400 328.050 207.450 332.400 ;
        RECT 211.950 328.950 214.050 333.000 ;
        RECT 205.950 325.950 208.050 328.050 ;
        RECT 196.950 322.950 199.050 325.050 ;
        RECT 205.950 322.800 208.050 324.900 ;
        RECT 187.950 310.950 190.050 313.050 ;
        RECT 181.950 295.950 184.050 298.050 ;
        RECT 187.950 297.450 192.000 298.050 ;
        RECT 187.950 295.950 192.450 297.450 ;
        RECT 170.400 292.350 171.600 294.000 ;
        RECT 176.400 292.350 177.600 294.600 ;
        RECT 178.950 292.950 181.050 295.050 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 167.400 287.400 168.600 289.650 ;
        RECT 173.400 288.900 174.600 289.650 ;
        RECT 167.400 262.200 168.450 287.400 ;
        RECT 172.950 286.800 175.050 288.900 ;
        RECT 182.400 273.450 183.450 295.950 ;
        RECT 191.400 294.600 192.450 295.950 ;
        RECT 191.400 292.350 192.600 294.600 ;
        RECT 199.950 292.950 202.050 295.050 ;
        RECT 206.400 294.450 207.450 322.800 ;
        RECT 214.950 319.950 217.050 322.050 ;
        RECT 203.400 293.400 207.450 294.450 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 188.400 287.400 189.600 289.650 ;
        RECT 194.400 288.900 195.600 289.650 ;
        RECT 200.400 288.900 201.450 292.950 ;
        RECT 188.400 277.050 189.450 287.400 ;
        RECT 193.950 286.800 196.050 288.900 ;
        RECT 199.950 286.800 202.050 288.900 ;
        RECT 187.950 274.950 190.050 277.050 ;
        RECT 182.400 272.400 186.450 273.450 ;
        RECT 181.950 268.950 184.050 271.050 ;
        RECT 172.950 265.950 175.050 268.050 ;
        RECT 166.950 261.450 169.050 262.200 ;
        RECT 164.400 260.400 169.050 261.450 ;
        RECT 164.400 255.900 165.450 260.400 ;
        RECT 166.950 260.100 169.050 260.400 ;
        RECT 173.400 261.600 174.450 265.950 ;
        RECT 173.400 259.350 174.600 261.600 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 170.400 255.900 171.600 256.650 ;
        RECT 176.400 255.900 177.600 256.650 ;
        RECT 182.400 255.900 183.450 268.950 ;
        RECT 185.400 262.050 186.450 272.400 ;
        RECT 196.950 268.950 199.050 271.050 ;
        RECT 184.950 259.950 187.050 262.050 ;
        RECT 190.950 260.100 193.050 262.200 ;
        RECT 197.400 261.600 198.450 268.950 ;
        RECT 200.400 262.050 201.450 286.800 ;
        RECT 203.400 271.050 204.450 293.400 ;
        RECT 211.950 293.100 214.050 295.200 ;
        RECT 215.400 295.050 216.450 319.950 ;
        RECT 218.400 310.050 219.450 337.950 ;
        RECT 221.400 316.050 222.450 361.950 ;
        RECT 224.400 361.050 225.450 394.950 ;
        RECT 230.400 373.200 231.450 406.800 ;
        RECT 233.400 379.050 234.450 424.950 ;
        RECT 247.950 418.950 250.050 421.050 ;
        RECT 244.800 412.950 246.900 415.050 ;
        RECT 245.400 411.450 246.600 412.650 ;
        RECT 248.400 411.450 249.450 418.950 ;
        RECT 245.400 410.400 249.450 411.450 ;
        RECT 251.400 409.050 252.450 427.950 ;
        RECT 253.950 418.800 256.050 420.900 ;
        RECT 250.950 406.950 253.050 409.050 ;
        RECT 254.400 406.050 255.450 418.800 ;
        RECT 260.400 418.050 261.450 445.950 ;
        RECT 269.400 427.050 270.450 445.950 ;
        RECT 274.950 442.950 277.050 445.050 ;
        RECT 275.400 430.050 276.450 442.950 ;
        RECT 274.950 427.950 277.050 430.050 ;
        RECT 268.950 424.950 271.050 427.050 ;
        RECT 275.400 421.050 276.450 427.950 ;
        RECT 259.950 415.950 262.050 418.050 ;
        RECT 265.950 417.000 268.050 421.050 ;
        RECT 274.950 418.950 277.050 421.050 ;
        RECT 281.400 420.450 282.450 445.950 ;
        RECT 284.400 443.400 285.900 462.300 ;
        RECT 288.300 456.300 289.500 462.300 ;
        RECT 287.400 454.200 289.500 456.300 ;
        RECT 284.400 441.300 286.500 443.400 ;
        RECT 285.300 437.700 286.500 441.300 ;
        RECT 288.300 437.700 289.500 454.200 ;
        RECT 290.700 459.300 292.800 461.400 ;
        RECT 290.700 437.700 291.900 459.300 ;
        RECT 299.400 457.800 301.500 459.900 ;
        RECT 304.800 459.300 306.900 461.400 ;
        RECT 299.400 451.200 300.300 457.800 ;
        RECT 305.100 452.100 306.300 459.300 ;
        RECT 307.800 457.500 309.300 462.300 ;
        RECT 310.200 459.300 312.300 464.400 ;
        RECT 307.800 455.400 309.900 457.500 ;
        RECT 299.400 449.100 301.500 451.200 ;
        RECT 304.800 450.000 306.900 452.100 ;
        RECT 295.950 446.100 298.050 448.200 ;
        RECT 296.400 445.350 297.600 446.100 ;
        RECT 295.800 442.950 297.900 445.050 ;
        RECT 299.400 438.600 300.300 449.100 ;
        RECT 302.100 442.500 304.200 444.600 ;
        RECT 284.700 435.600 286.800 437.700 ;
        RECT 287.700 435.600 289.800 437.700 ;
        RECT 290.700 435.600 292.800 437.700 ;
        RECT 298.800 436.500 300.900 438.600 ;
        RECT 305.100 437.700 306.300 450.000 ;
        RECT 307.800 437.700 309.300 455.400 ;
        RECT 311.100 437.700 312.300 459.300 ;
        RECT 304.200 435.600 306.300 437.700 ;
        RECT 307.200 435.600 309.300 437.700 ;
        RECT 310.200 435.600 312.300 437.700 ;
        RECT 313.200 462.300 315.300 464.400 ;
        RECT 313.200 457.500 314.700 462.300 ;
        RECT 313.200 455.400 315.300 457.500 ;
        RECT 313.200 437.700 314.700 455.400 ;
        RECT 313.200 435.600 315.300 437.700 ;
        RECT 304.950 430.950 307.050 433.050 ;
        RECT 281.400 419.400 285.450 420.450 ;
        RECT 266.400 415.350 267.600 417.000 ;
        RECT 274.800 415.800 276.900 417.900 ;
        RECT 284.400 417.600 285.450 419.400 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 263.400 410.400 264.600 412.650 ;
        RECT 269.400 411.900 270.600 412.650 ;
        RECT 253.950 403.950 256.050 406.050 ;
        RECT 263.400 400.050 264.450 410.400 ;
        RECT 268.950 409.800 271.050 411.900 ;
        RECT 271.950 403.950 274.050 409.050 ;
        RECT 262.950 397.950 265.050 400.050 ;
        RECT 271.950 385.950 274.050 388.050 ;
        RECT 241.950 382.950 244.050 385.050 ;
        RECT 232.950 376.950 235.050 379.050 ;
        RECT 229.950 371.100 232.050 373.200 ;
        RECT 235.950 371.100 238.050 376.050 ;
        RECT 230.400 370.350 231.600 371.100 ;
        RECT 236.400 370.350 237.600 371.100 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 232.950 367.950 235.050 370.050 ;
        RECT 235.950 367.950 238.050 370.050 ;
        RECT 233.400 366.000 234.600 367.650 ;
        RECT 226.950 361.950 229.050 364.050 ;
        RECT 232.950 361.950 235.050 366.000 ;
        RECT 223.950 358.950 226.050 361.050 ;
        RECT 227.400 349.050 228.450 361.950 ;
        RECT 229.950 349.950 232.050 352.050 ;
        RECT 230.400 349.050 231.450 349.950 ;
        RECT 226.950 346.950 229.050 349.050 ;
        RECT 230.400 346.950 235.050 349.050 ;
        RECT 230.400 339.600 231.450 346.950 ;
        RECT 242.400 340.200 243.450 382.950 ;
        RECT 247.950 371.100 250.050 373.200 ;
        RECT 248.400 370.350 249.600 371.100 ;
        RECT 256.950 370.950 259.050 373.050 ;
        RECT 265.950 371.100 268.050 373.200 ;
        RECT 272.400 372.600 273.450 385.950 ;
        RECT 275.400 373.200 276.450 415.800 ;
        RECT 284.400 415.350 285.600 417.600 ;
        RECT 289.950 417.000 292.050 421.050 ;
        RECT 305.400 420.450 306.450 430.950 ;
        RECT 313.950 427.950 316.050 430.050 ;
        RECT 302.400 419.400 306.450 420.450 ;
        RECT 302.400 417.600 303.450 419.400 ;
        RECT 290.400 415.350 291.600 417.000 ;
        RECT 302.400 415.350 303.600 417.600 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 302.400 412.950 304.500 415.050 ;
        RECT 307.800 412.950 309.900 415.050 ;
        RECT 277.950 409.800 280.050 411.900 ;
        RECT 281.400 411.000 282.600 412.650 ;
        RECT 278.400 403.050 279.450 409.800 ;
        RECT 280.950 406.950 283.050 411.000 ;
        RECT 287.400 410.400 288.600 412.650 ;
        RECT 308.400 410.400 309.600 412.650 ;
        RECT 287.400 406.050 288.450 410.400 ;
        RECT 286.950 403.950 289.050 406.050 ;
        RECT 277.950 400.950 280.050 403.050 ;
        RECT 287.400 400.050 288.450 403.950 ;
        RECT 286.950 397.950 289.050 400.050 ;
        RECT 295.950 385.950 298.050 388.050 ;
        RECT 280.950 379.950 283.050 382.050 ;
        RECT 277.950 376.950 280.050 379.050 ;
        RECT 247.950 367.950 250.050 370.050 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 251.400 366.900 252.600 367.650 ;
        RECT 257.400 366.900 258.450 370.950 ;
        RECT 266.400 370.350 267.600 371.100 ;
        RECT 272.400 370.350 273.600 372.600 ;
        RECT 274.950 371.100 277.050 373.200 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 263.400 366.900 264.600 367.650 ;
        RECT 269.400 366.900 270.600 367.650 ;
        RECT 250.950 364.800 253.050 366.900 ;
        RECT 256.950 364.800 259.050 366.900 ;
        RECT 262.950 364.800 265.050 366.900 ;
        RECT 268.950 364.800 271.050 366.900 ;
        RECT 278.400 355.050 279.450 376.950 ;
        RECT 281.400 367.050 282.450 379.950 ;
        RECT 289.950 371.100 292.050 373.200 ;
        RECT 296.400 372.600 297.450 385.950 ;
        RECT 301.950 382.950 304.050 385.050 ;
        RECT 290.400 370.350 291.600 371.100 ;
        RECT 296.400 370.350 297.600 372.600 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 295.950 367.950 298.050 370.050 ;
        RECT 280.950 364.950 283.050 367.050 ;
        RECT 287.400 365.400 288.600 367.650 ;
        RECT 293.400 365.400 294.600 367.650 ;
        RECT 287.400 361.050 288.450 365.400 ;
        RECT 286.800 358.950 288.900 361.050 ;
        RECT 289.950 358.950 292.050 361.050 ;
        RECT 253.950 352.950 256.050 355.050 ;
        RECT 259.950 352.950 262.050 355.050 ;
        RECT 277.950 352.950 280.050 355.050 ;
        RECT 250.950 340.950 253.050 343.050 ;
        RECT 230.400 337.350 231.600 339.600 ;
        RECT 235.950 337.950 238.050 340.050 ;
        RECT 241.950 338.100 244.050 340.200 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 229.950 334.950 232.050 337.050 ;
        RECT 227.400 332.400 228.600 334.650 ;
        RECT 220.950 313.950 223.050 316.050 ;
        RECT 217.950 307.950 220.050 310.050 ;
        RECT 227.400 297.450 228.450 332.400 ;
        RECT 236.400 328.050 237.450 337.950 ;
        RECT 242.400 337.350 243.600 338.100 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 245.400 332.400 246.600 334.650 ;
        RECT 235.950 325.950 238.050 328.050 ;
        RECT 245.400 322.050 246.450 332.400 ;
        RECT 244.950 319.950 247.050 322.050 ;
        RECT 251.400 319.050 252.450 340.950 ;
        RECT 254.400 331.050 255.450 352.950 ;
        RECT 260.400 339.600 261.450 352.950 ;
        RECT 268.950 349.950 271.050 352.050 ;
        RECT 260.400 337.350 261.600 339.600 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 263.400 332.400 264.600 334.650 ;
        RECT 253.950 328.950 256.050 331.050 ;
        RECT 259.950 319.950 262.050 322.050 ;
        RECT 250.950 316.950 253.050 319.050 ;
        RECT 238.950 307.950 241.050 310.050 ;
        RECT 253.950 307.950 256.050 310.050 ;
        RECT 235.950 301.950 238.050 304.050 ;
        RECT 229.950 298.950 232.050 301.050 ;
        RECT 224.400 296.400 228.450 297.450 ;
        RECT 212.400 292.350 213.600 293.100 ;
        RECT 214.950 292.950 217.050 295.050 ;
        RECT 217.950 292.950 220.050 295.050 ;
        RECT 224.400 294.600 225.450 296.400 ;
        RECT 230.400 294.600 231.450 298.950 ;
        RECT 236.400 295.050 237.450 301.950 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 209.400 287.400 210.600 289.650 ;
        RECT 209.400 283.050 210.450 287.400 ;
        RECT 218.400 283.050 219.450 292.950 ;
        RECT 224.400 292.350 225.600 294.600 ;
        RECT 230.400 292.350 231.600 294.600 ;
        RECT 235.950 292.950 238.050 295.050 ;
        RECT 223.950 289.950 226.050 292.050 ;
        RECT 226.950 289.950 229.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 220.950 286.950 223.050 289.050 ;
        RECT 227.400 287.400 228.600 289.650 ;
        RECT 233.400 287.400 234.600 289.650 ;
        RECT 208.950 280.950 211.050 283.050 ;
        RECT 217.950 280.950 220.050 283.050 ;
        RECT 221.400 277.050 222.450 286.950 ;
        RECT 227.400 283.050 228.450 287.400 ;
        RECT 226.950 280.950 229.050 283.050 ;
        RECT 220.950 274.950 223.050 277.050 ;
        RECT 214.950 271.950 217.050 274.050 ;
        RECT 202.950 270.450 205.050 271.050 ;
        RECT 202.950 269.400 207.450 270.450 ;
        RECT 202.950 268.950 205.050 269.400 ;
        RECT 202.950 265.800 205.050 267.900 ;
        RECT 191.400 259.350 192.600 260.100 ;
        RECT 197.400 259.350 198.600 261.600 ;
        RECT 199.950 259.950 202.050 262.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 196.950 256.950 199.050 259.050 ;
        RECT 188.400 255.900 189.600 256.650 ;
        RECT 163.950 253.800 166.050 255.900 ;
        RECT 169.950 253.800 172.050 255.900 ;
        RECT 175.950 253.800 178.050 255.900 ;
        RECT 181.950 253.800 184.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 194.400 254.400 195.600 256.650 ;
        RECT 164.400 247.050 165.450 253.800 ;
        RECT 194.400 250.050 195.450 254.400 ;
        RECT 199.950 253.950 202.050 256.050 ;
        RECT 193.950 247.950 196.050 250.050 ;
        RECT 163.950 244.950 166.050 247.050 ;
        RECT 160.950 235.950 163.050 238.050 ;
        RECT 200.400 223.050 201.450 253.950 ;
        RECT 203.400 226.050 204.450 265.800 ;
        RECT 206.400 261.450 207.450 269.400 ;
        RECT 215.400 261.600 216.450 271.950 ;
        RECT 221.400 261.600 222.450 274.950 ;
        RECT 223.950 271.950 226.050 274.050 ;
        RECT 209.400 261.450 210.600 261.600 ;
        RECT 206.400 260.400 210.600 261.450 ;
        RECT 209.400 259.350 210.600 260.400 ;
        RECT 215.400 259.350 216.600 261.600 ;
        RECT 221.400 259.350 222.600 261.600 ;
        RECT 224.400 261.450 225.450 271.950 ;
        RECT 227.400 265.050 228.450 280.950 ;
        RECT 226.950 262.950 229.050 265.050 ;
        RECT 233.400 261.450 234.450 287.400 ;
        RECT 239.400 274.050 240.450 307.950 ;
        RECT 247.950 293.100 250.050 295.200 ;
        RECT 254.400 294.600 255.450 307.950 ;
        RECT 248.400 292.350 249.600 293.100 ;
        RECT 254.400 292.350 255.600 294.600 ;
        RECT 244.950 289.950 247.050 292.050 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 245.400 288.900 246.600 289.650 ;
        RECT 244.950 286.800 247.050 288.900 ;
        RECT 251.400 287.400 252.600 289.650 ;
        RECT 260.400 288.900 261.450 319.950 ;
        RECT 263.400 303.450 264.450 332.400 ;
        RECT 269.400 307.050 270.450 349.950 ;
        RECT 280.950 346.950 283.050 349.050 ;
        RECT 274.950 342.450 277.050 346.050 ;
        RECT 272.400 342.000 277.050 342.450 ;
        RECT 272.400 341.400 276.450 342.000 ;
        RECT 272.400 322.050 273.450 341.400 ;
        RECT 281.400 339.600 282.450 346.950 ;
        RECT 290.400 342.450 291.450 358.950 ;
        RECT 293.400 352.050 294.450 365.400 ;
        RECT 298.950 364.950 301.050 367.050 ;
        RECT 299.400 358.050 300.450 364.950 ;
        RECT 298.950 355.950 301.050 358.050 ;
        RECT 292.950 349.950 295.050 352.050 ;
        RECT 302.400 346.050 303.450 382.950 ;
        RECT 304.950 376.950 307.050 379.050 ;
        RECT 305.400 373.050 306.450 376.950 ;
        RECT 308.400 376.050 309.450 410.400 ;
        RECT 314.400 408.900 315.450 427.950 ;
        RECT 313.950 406.800 316.050 408.900 ;
        RECT 317.400 406.050 318.450 466.950 ;
        RECT 325.950 454.950 328.050 457.050 ;
        RECT 322.800 448.950 324.900 451.050 ;
        RECT 323.400 446.400 324.600 448.650 ;
        RECT 323.400 442.050 324.450 446.400 ;
        RECT 322.950 439.950 325.050 442.050 ;
        RECT 323.400 424.050 324.450 439.950 ;
        RECT 326.400 430.050 327.450 454.950 ;
        RECT 331.800 448.950 333.900 451.050 ;
        RECT 332.400 447.000 333.600 448.650 ;
        RECT 331.950 444.450 334.050 447.000 ;
        RECT 335.400 444.450 336.450 475.950 ;
        RECT 350.400 469.050 351.450 508.950 ;
        RECT 355.800 490.950 357.900 493.050 ;
        RECT 356.400 489.900 357.600 490.650 ;
        RECT 355.950 487.800 358.050 489.900 ;
        RECT 359.400 478.050 360.450 547.950 ;
        RECT 361.950 541.950 364.050 544.050 ;
        RECT 362.400 535.050 363.450 541.950 ;
        RECT 368.400 541.050 369.450 550.950 ;
        RECT 367.950 538.950 370.050 541.050 ;
        RECT 361.950 532.950 364.050 535.050 ;
        RECT 364.800 526.950 366.900 529.050 ;
        RECT 365.400 524.400 366.600 526.650 ;
        RECT 361.950 517.950 364.050 520.050 ;
        RECT 362.400 490.050 363.450 517.950 ;
        RECT 365.400 508.050 366.450 524.400 ;
        RECT 368.400 514.050 369.450 538.950 ;
        RECT 373.800 526.950 375.900 529.050 ;
        RECT 374.400 525.450 375.600 526.650 ;
        RECT 377.400 525.450 378.450 563.400 ;
        RECT 379.950 562.950 382.050 563.400 ;
        RECT 379.950 553.950 382.050 556.050 ;
        RECT 374.400 524.400 378.450 525.450 ;
        RECT 374.400 514.050 375.450 524.400 ;
        RECT 367.950 511.950 370.050 514.050 ;
        RECT 373.950 511.950 376.050 514.050 ;
        RECT 364.950 505.950 367.050 508.050 ;
        RECT 367.950 499.950 370.050 502.050 ;
        RECT 364.950 494.100 367.050 496.200 ;
        RECT 361.950 487.950 364.050 490.050 ;
        RECT 358.950 475.950 361.050 478.050 ;
        RECT 349.950 466.950 352.050 469.050 ;
        RECT 353.400 462.300 356.400 464.400 ;
        RECT 357.300 462.300 359.400 464.400 ;
        RECT 340.950 453.000 343.050 457.050 ;
        RECT 341.400 451.350 342.600 453.000 ;
        RECT 340.800 448.950 342.900 451.050 ;
        RECT 346.800 448.950 348.900 451.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 331.950 443.400 336.450 444.450 ;
        RECT 331.950 442.950 334.050 443.400 ;
        RECT 340.950 442.950 343.050 445.050 ;
        RECT 325.950 427.950 328.050 430.050 ;
        RECT 322.950 421.950 325.050 424.050 ;
        RECT 322.950 416.100 325.050 418.200 ;
        RECT 323.400 415.350 324.600 416.100 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 319.950 409.950 322.050 412.050 ;
        RECT 326.400 410.400 327.600 412.650 ;
        RECT 316.950 403.950 319.050 406.050 ;
        RECT 313.950 388.950 316.050 391.050 ;
        RECT 314.400 376.050 315.450 388.950 ;
        RECT 320.400 385.050 321.450 409.950 ;
        RECT 322.950 397.950 325.050 400.050 ;
        RECT 319.950 382.950 322.050 385.050 ;
        RECT 307.950 373.950 310.050 376.050 ;
        RECT 313.950 373.950 316.050 376.050 ;
        RECT 319.950 373.950 322.050 376.050 ;
        RECT 304.950 370.950 307.050 373.050 ;
        RECT 308.400 372.600 309.450 373.950 ;
        RECT 314.400 372.600 315.450 373.950 ;
        RECT 308.400 370.350 309.600 372.600 ;
        RECT 314.400 370.350 315.600 372.600 ;
        RECT 307.950 367.950 310.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 311.400 365.400 312.600 367.650 ;
        RECT 311.400 361.050 312.450 365.400 ;
        RECT 320.400 364.050 321.450 373.950 ;
        RECT 323.400 373.050 324.450 397.950 ;
        RECT 326.400 397.050 327.450 410.400 ;
        RECT 331.800 409.950 333.900 412.050 ;
        RECT 337.800 409.950 339.900 412.050 ;
        RECT 332.400 408.900 333.600 409.650 ;
        RECT 331.950 406.800 334.050 408.900 ;
        RECT 341.400 403.050 342.450 442.950 ;
        RECT 344.400 436.050 345.450 445.950 ;
        RECT 353.400 443.400 354.900 462.300 ;
        RECT 357.300 456.300 358.500 462.300 ;
        RECT 356.400 454.200 358.500 456.300 ;
        RECT 353.400 441.300 355.500 443.400 ;
        RECT 354.300 437.700 355.500 441.300 ;
        RECT 357.300 437.700 358.500 454.200 ;
        RECT 359.700 459.300 361.800 461.400 ;
        RECT 359.700 437.700 360.900 459.300 ;
        RECT 361.950 454.950 364.050 457.050 ;
        RECT 362.400 447.450 363.450 454.950 ;
        RECT 365.400 451.050 366.450 494.100 ;
        RECT 368.400 463.050 369.450 499.950 ;
        RECT 376.950 494.100 379.050 496.200 ;
        RECT 377.400 493.350 378.600 494.100 ;
        RECT 371.100 490.950 373.200 493.050 ;
        RECT 376.500 490.950 378.600 493.050 ;
        RECT 371.400 489.000 372.600 490.650 ;
        RECT 370.950 484.950 373.050 489.000 ;
        RECT 380.400 478.050 381.450 553.950 ;
        RECT 383.400 496.050 384.450 565.950 ;
        RECT 382.950 493.950 385.050 496.050 ;
        RECT 379.950 475.950 382.050 478.050 ;
        RECT 367.950 460.950 370.050 463.050 ;
        RECT 376.200 462.300 378.300 464.400 ;
        RECT 368.400 457.800 370.500 459.900 ;
        RECT 373.800 459.300 375.900 461.400 ;
        RECT 368.400 451.200 369.300 457.800 ;
        RECT 374.100 452.100 375.300 459.300 ;
        RECT 376.800 457.500 378.300 462.300 ;
        RECT 379.200 459.300 381.300 464.400 ;
        RECT 376.800 455.400 378.900 457.500 ;
        RECT 364.950 448.950 367.050 451.050 ;
        RECT 368.400 449.100 370.500 451.200 ;
        RECT 373.800 450.000 375.900 452.100 ;
        RECT 365.400 447.450 366.600 447.600 ;
        RECT 362.400 446.400 366.600 447.450 ;
        RECT 365.400 445.350 366.600 446.400 ;
        RECT 364.800 442.950 366.900 445.050 ;
        RECT 368.400 438.600 369.300 449.100 ;
        RECT 371.100 442.500 373.200 444.600 ;
        RECT 343.950 433.950 346.050 436.050 ;
        RECT 353.700 435.600 355.800 437.700 ;
        RECT 356.700 435.600 358.800 437.700 ;
        RECT 359.700 435.600 361.800 437.700 ;
        RECT 367.800 436.500 369.900 438.600 ;
        RECT 374.100 437.700 375.300 450.000 ;
        RECT 376.800 437.700 378.300 455.400 ;
        RECT 380.100 437.700 381.300 459.300 ;
        RECT 373.200 435.600 375.300 437.700 ;
        RECT 376.200 435.600 378.300 437.700 ;
        RECT 379.200 435.600 381.300 437.700 ;
        RECT 382.200 462.300 384.300 464.400 ;
        RECT 382.200 457.500 383.700 462.300 ;
        RECT 382.200 455.400 384.300 457.500 ;
        RECT 382.200 437.700 383.700 455.400 ;
        RECT 382.200 435.600 384.300 437.700 ;
        RECT 382.950 430.950 385.050 433.050 ;
        RECT 344.700 423.300 346.800 425.400 ;
        RECT 347.700 423.300 349.800 425.400 ;
        RECT 350.700 423.300 352.800 425.400 ;
        RECT 345.300 419.700 346.500 423.300 ;
        RECT 344.400 417.600 346.500 419.700 ;
        RECT 340.950 400.950 343.050 403.050 ;
        RECT 344.400 398.700 345.900 417.600 ;
        RECT 348.300 406.800 349.500 423.300 ;
        RECT 347.400 404.700 349.500 406.800 ;
        RECT 348.300 398.700 349.500 404.700 ;
        RECT 350.700 401.700 351.900 423.300 ;
        RECT 358.800 422.400 360.900 424.500 ;
        RECT 364.200 423.300 366.300 425.400 ;
        RECT 367.200 423.300 369.300 425.400 ;
        RECT 370.200 423.300 372.300 425.400 ;
        RECT 355.800 415.950 357.900 418.050 ;
        RECT 356.400 414.000 357.600 415.650 ;
        RECT 355.950 409.950 358.050 414.000 ;
        RECT 359.400 411.900 360.300 422.400 ;
        RECT 362.100 416.400 364.200 418.500 ;
        RECT 359.400 409.800 361.500 411.900 ;
        RECT 365.100 411.000 366.300 423.300 ;
        RECT 359.400 403.200 360.300 409.800 ;
        RECT 364.800 408.900 366.900 411.000 ;
        RECT 350.700 399.600 352.800 401.700 ;
        RECT 359.400 401.100 361.500 403.200 ;
        RECT 365.100 401.700 366.300 408.900 ;
        RECT 367.800 405.600 369.300 423.300 ;
        RECT 367.800 403.500 369.900 405.600 ;
        RECT 364.800 399.600 366.900 401.700 ;
        RECT 367.800 398.700 369.300 403.500 ;
        RECT 371.100 401.700 372.300 423.300 ;
        RECT 325.950 394.950 328.050 397.050 ;
        RECT 344.400 396.600 347.400 398.700 ;
        RECT 348.300 396.600 350.400 398.700 ;
        RECT 367.200 396.600 369.300 398.700 ;
        RECT 370.200 396.600 372.300 401.700 ;
        RECT 373.200 423.300 375.300 425.400 ;
        RECT 383.400 424.050 384.450 430.950 ;
        RECT 373.200 405.600 374.700 423.300 ;
        RECT 382.950 421.950 385.050 424.050 ;
        RECT 376.950 418.950 379.050 421.050 ;
        RECT 373.200 403.500 375.300 405.600 ;
        RECT 373.200 398.700 374.700 403.500 ;
        RECT 373.200 396.600 375.300 398.700 ;
        RECT 377.400 397.050 378.450 418.950 ;
        RECT 383.400 414.600 384.450 421.950 ;
        RECT 383.400 412.350 384.600 414.600 ;
        RECT 386.400 412.050 387.450 577.950 ;
        RECT 389.400 568.050 390.450 596.400 ;
        RECT 391.950 595.950 394.050 598.050 ;
        RECT 397.950 595.950 400.050 598.050 ;
        RECT 403.950 595.950 406.050 598.050 ;
        RECT 392.400 589.050 393.450 595.950 ;
        RECT 391.950 586.950 394.050 589.050 ;
        RECT 398.400 586.050 399.450 595.950 ;
        RECT 403.950 592.800 406.050 594.900 ;
        RECT 391.950 583.800 394.050 585.900 ;
        RECT 397.950 583.950 400.050 586.050 ;
        RECT 392.400 574.050 393.450 583.800 ;
        RECT 404.400 574.200 405.450 592.800 ;
        RECT 391.950 571.950 394.050 574.050 ;
        RECT 397.950 572.100 400.050 574.200 ;
        RECT 403.950 572.100 406.050 574.200 ;
        RECT 398.400 571.350 399.600 572.100 ;
        RECT 394.950 568.950 397.050 571.050 ;
        RECT 397.950 568.950 400.050 571.050 ;
        RECT 400.950 568.950 403.050 571.050 ;
        RECT 388.950 565.950 391.050 568.050 ;
        RECT 395.400 566.400 396.600 568.650 ;
        RECT 401.400 566.400 402.600 568.650 ;
        RECT 395.400 565.050 396.450 566.400 ;
        RECT 394.950 564.450 397.050 565.050 ;
        RECT 394.950 563.400 399.450 564.450 ;
        RECT 394.950 562.950 397.050 563.400 ;
        RECT 388.950 544.950 391.050 547.050 ;
        RECT 389.400 522.450 390.450 544.950 ;
        RECT 398.400 529.200 399.450 563.400 ;
        RECT 401.400 532.050 402.450 566.400 ;
        RECT 403.950 559.950 406.050 562.050 ;
        RECT 400.950 529.950 403.050 532.050 ;
        RECT 397.950 527.100 400.050 529.200 ;
        RECT 404.400 528.450 405.450 559.950 ;
        RECT 407.400 538.050 408.450 607.950 ;
        RECT 415.950 606.000 418.050 610.050 ;
        RECT 424.950 607.950 427.050 610.050 ;
        RECT 416.400 604.350 417.600 606.000 ;
        RECT 421.950 605.100 424.050 607.200 ;
        RECT 422.400 604.350 423.600 605.100 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 415.950 601.950 418.050 604.050 ;
        RECT 418.950 601.950 421.050 604.050 ;
        RECT 421.950 601.950 424.050 604.050 ;
        RECT 409.950 598.950 412.050 601.050 ;
        RECT 413.400 599.400 414.600 601.650 ;
        RECT 419.400 599.400 420.600 601.650 ;
        RECT 410.400 594.450 411.450 598.950 ;
        RECT 413.400 595.050 414.450 599.400 ;
        RECT 412.800 594.450 414.900 595.050 ;
        RECT 410.400 593.400 414.900 594.450 ;
        RECT 412.800 592.950 414.900 593.400 ;
        RECT 415.950 592.950 418.050 595.050 ;
        RECT 409.950 583.950 412.050 586.050 ;
        RECT 410.400 580.050 411.450 583.950 ;
        RECT 416.400 583.050 417.450 592.950 ;
        RECT 419.400 586.050 420.450 599.400 ;
        RECT 424.950 598.950 427.050 601.050 ;
        RECT 418.950 583.950 421.050 586.050 ;
        RECT 415.950 580.950 418.050 583.050 ;
        RECT 409.950 577.950 412.050 580.050 ;
        RECT 416.400 577.050 417.450 580.950 ;
        RECT 415.950 574.950 418.050 577.050 ;
        RECT 412.950 572.100 415.050 574.200 ;
        RECT 418.950 572.100 421.050 574.200 ;
        RECT 425.400 574.050 426.450 598.950 ;
        RECT 428.400 595.050 429.450 610.950 ;
        RECT 434.400 606.600 435.450 613.950 ;
        RECT 440.400 607.200 441.450 632.400 ;
        RECT 442.950 631.950 445.050 634.050 ;
        RECT 434.400 604.350 435.600 606.600 ;
        RECT 439.950 605.100 442.050 607.200 ;
        RECT 445.950 605.100 448.050 607.200 ;
        RECT 440.400 604.350 441.600 605.100 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 436.950 601.950 439.050 604.050 ;
        RECT 439.950 601.950 442.050 604.050 ;
        RECT 437.400 600.900 438.600 601.650 ;
        RECT 436.950 598.800 439.050 600.900 ;
        RECT 427.950 592.950 430.050 595.050 ;
        RECT 436.950 592.950 439.050 595.050 ;
        RECT 430.950 589.950 433.050 592.050 ;
        RECT 413.400 571.350 414.600 572.100 ;
        RECT 419.400 571.350 420.600 572.100 ;
        RECT 424.950 571.950 427.050 574.050 ;
        RECT 431.400 571.050 432.450 589.950 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 418.950 568.950 421.050 571.050 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 409.950 565.950 412.050 568.050 ;
        RECT 416.400 567.900 417.600 568.650 ;
        RECT 410.400 553.050 411.450 565.950 ;
        RECT 415.950 565.800 418.050 567.900 ;
        RECT 422.400 566.400 423.600 568.650 ;
        RECT 418.950 562.950 421.050 565.050 ;
        RECT 419.400 559.050 420.450 562.950 ;
        RECT 418.950 556.950 421.050 559.050 ;
        RECT 422.400 553.050 423.450 566.400 ;
        RECT 427.800 565.950 429.900 568.050 ;
        RECT 433.800 565.950 435.900 568.050 ;
        RECT 428.400 563.400 429.600 565.650 ;
        RECT 428.400 556.050 429.450 563.400 ;
        RECT 430.950 562.950 433.050 565.050 ;
        RECT 427.950 553.950 430.050 556.050 ;
        RECT 409.950 550.950 412.050 553.050 ;
        RECT 421.950 550.950 424.050 553.050 ;
        RECT 409.950 541.950 412.050 544.050 ;
        RECT 431.400 543.450 432.450 562.950 ;
        RECT 433.950 550.950 436.050 553.050 ;
        RECT 434.400 544.050 435.450 550.950 ;
        RECT 437.400 547.050 438.450 592.950 ;
        RECT 446.400 592.050 447.450 605.100 ;
        RECT 449.400 601.050 450.450 634.950 ;
        RECT 455.400 610.050 456.450 643.950 ;
        RECT 458.400 637.050 459.450 709.950 ;
        RECT 476.400 709.050 477.450 728.100 ;
        RECT 479.400 727.050 480.450 751.950 ;
        RECT 482.400 742.050 483.450 755.400 ;
        RECT 489.000 754.950 493.050 755.400 ;
        RECT 493.950 754.950 496.050 757.050 ;
        RECT 503.400 755.400 504.600 757.650 ;
        RECT 496.950 751.950 499.050 754.050 ;
        RECT 481.950 739.950 484.050 742.050 ;
        RECT 487.950 728.100 490.050 730.200 ;
        RECT 488.400 727.350 489.600 728.100 ;
        RECT 478.950 724.950 481.050 727.050 ;
        RECT 484.950 724.950 487.050 727.050 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 485.400 722.400 486.600 724.650 ;
        RECT 497.400 724.050 498.450 751.950 ;
        RECT 503.400 745.050 504.450 755.400 ;
        RECT 505.950 754.950 508.050 757.050 ;
        RECT 509.400 756.450 510.450 761.400 ;
        RECT 518.400 760.350 519.600 762.600 ;
        RECT 523.950 761.100 526.050 763.200 ;
        RECT 524.400 760.350 525.600 761.100 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 509.400 755.400 513.450 756.450 ;
        RECT 515.400 756.000 516.600 757.650 ;
        RECT 506.400 748.050 507.450 754.950 ;
        RECT 505.950 745.950 508.050 748.050 ;
        RECT 502.950 742.950 505.050 745.050 ;
        RECT 499.950 736.950 502.050 739.050 ;
        RECT 500.400 730.050 501.450 736.950 ;
        RECT 512.400 736.050 513.450 755.400 ;
        RECT 514.950 751.950 517.050 756.000 ;
        RECT 521.400 755.400 522.600 757.650 ;
        RECT 521.400 751.050 522.450 755.400 ;
        RECT 520.950 748.950 523.050 751.050 ;
        RECT 520.950 745.800 523.050 747.900 ;
        RECT 511.950 733.950 514.050 736.050 ;
        RECT 499.950 727.950 502.050 730.050 ;
        RECT 505.950 728.100 508.050 730.200 ;
        RECT 511.950 728.100 514.050 730.200 ;
        RECT 506.400 727.350 507.600 728.100 ;
        RECT 512.400 727.350 513.600 728.100 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 503.400 724.050 504.600 724.650 ;
        RECT 485.400 718.050 486.450 722.400 ;
        RECT 496.950 721.950 499.050 724.050 ;
        RECT 499.950 722.400 504.600 724.050 ;
        RECT 509.400 723.900 510.600 724.650 ;
        RECT 499.950 721.950 504.000 722.400 ;
        RECT 508.950 721.800 511.050 723.900 ;
        RECT 515.400 722.400 516.600 724.650 ;
        RECT 521.400 723.900 522.450 745.800 ;
        RECT 530.400 742.050 531.450 772.950 ;
        RECT 529.950 739.950 532.050 742.050 ;
        RECT 526.950 736.950 529.050 739.050 ;
        RECT 527.400 729.600 528.450 736.950 ;
        RECT 533.400 730.200 534.450 775.950 ;
        RECT 542.400 769.050 543.450 797.400 ;
        RECT 544.950 796.950 547.050 797.400 ;
        RECT 551.400 777.450 552.450 806.100 ;
        RECT 560.400 805.350 561.600 807.600 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 569.400 801.450 570.450 826.950 ;
        RECT 572.400 817.050 573.450 833.400 ;
        RECT 577.950 832.800 580.050 834.900 ;
        RECT 587.400 834.450 588.450 859.950 ;
        RECT 590.400 856.050 591.450 862.950 ;
        RECT 602.400 859.050 603.450 878.400 ;
        RECT 601.950 856.950 604.050 859.050 ;
        RECT 589.950 853.950 592.050 856.050 ;
        RECT 589.950 847.950 592.050 850.050 ;
        RECT 601.950 847.950 604.050 850.050 ;
        RECT 590.400 841.200 591.450 847.950 ;
        RECT 589.950 839.100 592.050 841.200 ;
        RECT 595.950 839.100 598.050 841.200 ;
        RECT 602.400 840.600 603.450 847.950 ;
        RECT 608.400 841.050 609.450 878.400 ;
        RECT 610.950 850.950 613.050 853.050 ;
        RECT 584.400 833.400 588.450 834.450 ;
        RECT 584.400 829.050 585.450 833.400 ;
        RECT 583.950 826.950 586.050 829.050 ;
        RECT 571.950 814.950 574.050 817.050 ;
        RECT 586.950 810.450 589.050 811.050 ;
        RECT 590.400 810.450 591.450 839.100 ;
        RECT 596.400 838.350 597.600 839.100 ;
        RECT 602.400 838.350 603.600 840.600 ;
        RECT 607.950 838.950 610.050 841.050 ;
        RECT 595.950 835.950 598.050 838.050 ;
        RECT 598.950 835.950 601.050 838.050 ;
        RECT 601.950 835.950 604.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 599.400 833.400 600.600 835.650 ;
        RECT 599.400 826.050 600.450 833.400 ;
        RECT 598.950 823.950 601.050 826.050 ;
        RECT 601.950 811.950 604.050 814.050 ;
        RECT 586.950 809.400 591.450 810.450 ;
        RECT 586.950 808.950 589.050 809.400 ;
        RECT 577.950 806.100 580.050 808.200 ;
        RECT 578.400 805.350 579.600 806.100 ;
        RECT 583.950 805.950 586.050 808.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 575.400 801.900 576.600 802.650 ;
        RECT 569.400 800.400 573.450 801.450 ;
        RECT 553.950 796.950 556.050 799.050 ;
        RECT 554.400 790.050 555.450 796.950 ;
        RECT 553.950 787.950 556.050 790.050 ;
        RECT 559.950 781.950 562.050 784.050 ;
        RECT 568.950 781.950 571.050 784.050 ;
        RECT 556.950 778.950 559.050 781.050 ;
        RECT 551.400 776.400 555.450 777.450 ;
        RECT 541.950 766.950 544.050 769.050 ;
        RECT 544.950 762.000 547.050 766.050 ;
        RECT 545.400 760.350 546.600 762.000 ;
        RECT 550.950 760.950 553.050 763.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 542.400 756.900 543.600 757.650 ;
        RECT 541.950 754.800 544.050 756.900 ;
        RECT 547.950 754.950 550.050 757.050 ;
        RECT 548.400 745.050 549.450 754.950 ;
        RECT 551.400 748.050 552.450 760.950 ;
        RECT 550.950 745.950 553.050 748.050 ;
        RECT 547.950 742.950 550.050 745.050 ;
        RECT 554.400 732.450 555.450 776.400 ;
        RECT 557.400 763.050 558.450 778.950 ;
        RECT 560.400 772.050 561.450 781.950 ;
        RECT 559.950 769.950 562.050 772.050 ;
        RECT 565.950 766.950 568.050 769.050 ;
        RECT 556.950 762.600 561.000 763.050 ;
        RECT 566.400 762.600 567.450 766.950 ;
        RECT 569.400 766.050 570.450 781.950 ;
        RECT 568.950 763.950 571.050 766.050 ;
        RECT 572.400 763.050 573.450 800.400 ;
        RECT 574.950 799.800 577.050 801.900 ;
        RECT 574.950 787.950 577.050 790.050 ;
        RECT 556.950 760.950 561.600 762.600 ;
        RECT 560.400 760.350 561.600 760.950 ;
        RECT 566.400 760.350 567.600 762.600 ;
        RECT 571.950 760.950 574.050 763.050 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 562.950 757.950 565.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 563.400 755.400 564.600 757.650 ;
        RECT 569.400 757.050 570.600 757.650 ;
        RECT 563.400 742.050 564.450 755.400 ;
        RECT 569.400 754.950 574.050 757.050 ;
        RECT 562.950 739.950 565.050 742.050 ;
        RECT 554.400 731.400 558.450 732.450 ;
        RECT 527.400 727.350 528.600 729.600 ;
        RECT 532.950 728.100 535.050 730.200 ;
        RECT 541.950 728.100 544.050 730.200 ;
        RECT 547.950 728.100 550.050 730.200 ;
        RECT 533.400 727.350 534.600 728.100 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 530.400 723.900 531.600 724.650 ;
        RECT 515.400 718.050 516.450 722.400 ;
        RECT 520.950 721.800 523.050 723.900 ;
        RECT 529.950 721.800 532.050 723.900 ;
        RECT 536.400 722.400 537.600 724.650 ;
        RECT 484.950 715.950 487.050 718.050 ;
        RECT 514.950 715.950 517.050 718.050 ;
        RECT 521.400 715.050 522.450 721.800 ;
        RECT 520.950 712.950 523.050 715.050 ;
        RECT 496.950 709.950 499.050 712.050 ;
        RECT 475.950 706.950 478.050 709.050 ;
        RECT 475.950 697.950 478.050 700.050 ;
        RECT 469.950 691.950 472.050 694.050 ;
        RECT 463.950 683.100 466.050 685.200 ;
        RECT 470.400 684.600 471.450 691.950 ;
        RECT 476.400 685.200 477.450 697.950 ;
        RECT 497.400 694.050 498.450 709.950 ;
        RECT 536.400 703.050 537.450 722.400 ;
        RECT 538.950 721.950 541.050 724.050 ;
        RECT 539.400 718.050 540.450 721.950 ;
        RECT 538.950 715.950 541.050 718.050 ;
        RECT 542.400 712.050 543.450 728.100 ;
        RECT 548.400 727.350 549.600 728.100 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 550.950 712.950 553.050 715.050 ;
        RECT 541.950 709.950 544.050 712.050 ;
        RECT 535.950 700.950 538.050 703.050 ;
        RECT 520.950 697.950 523.050 700.050 ;
        RECT 526.950 697.950 529.050 700.050 ;
        RECT 514.950 694.950 517.050 697.050 ;
        RECT 496.950 691.950 499.050 694.050 ;
        RECT 464.400 682.350 465.600 683.100 ;
        RECT 470.400 682.350 471.600 684.600 ;
        RECT 475.950 683.100 478.050 685.200 ;
        RECT 484.950 683.100 487.050 685.200 ;
        RECT 502.950 683.100 505.050 685.200 ;
        RECT 463.950 679.950 466.050 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 460.950 676.950 463.050 679.050 ;
        RECT 467.400 677.400 468.600 679.650 ;
        RECT 461.400 646.050 462.450 676.950 ;
        RECT 467.400 673.050 468.450 677.400 ;
        RECT 476.400 676.050 477.450 683.100 ;
        RECT 485.400 682.350 486.600 683.100 ;
        RECT 503.400 682.350 504.600 683.100 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 478.950 676.950 481.050 679.050 ;
        RECT 500.400 677.400 501.600 679.650 ;
        RECT 506.400 679.050 507.600 679.650 ;
        RECT 515.400 679.050 516.450 694.950 ;
        RECT 521.400 694.050 522.450 697.950 ;
        RECT 520.950 691.950 523.050 694.050 ;
        RECT 527.400 684.600 528.450 697.950 ;
        RECT 527.400 682.350 528.600 684.600 ;
        RECT 520.950 679.950 523.050 682.050 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 506.400 677.400 511.050 679.050 ;
        RECT 475.950 673.950 478.050 676.050 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 479.400 667.050 480.450 676.950 ;
        RECT 500.400 673.050 501.450 677.400 ;
        RECT 507.000 676.950 511.050 677.400 ;
        RECT 514.950 676.950 517.050 679.050 ;
        RECT 524.400 677.400 525.600 679.650 ;
        RECT 530.400 678.900 531.600 679.650 ;
        RECT 499.950 670.950 502.050 673.050 ;
        RECT 524.400 670.050 525.450 677.400 ;
        RECT 529.950 676.800 532.050 678.900 ;
        RECT 536.400 670.050 537.450 700.950 ;
        RECT 542.400 684.600 543.450 709.950 ;
        RECT 542.400 682.350 543.600 684.600 ;
        RECT 542.100 679.950 544.200 682.050 ;
        RECT 547.500 679.950 549.600 682.050 ;
        RECT 548.400 677.400 549.600 679.650 ;
        RECT 523.950 667.950 526.050 670.050 ;
        RECT 535.950 667.950 538.050 670.050 ;
        RECT 544.950 667.950 547.050 670.050 ;
        RECT 478.950 664.950 481.050 667.050 ;
        RECT 484.950 664.950 487.050 667.050 ;
        RECT 469.950 650.100 472.050 652.200 ;
        RECT 470.400 649.350 471.600 650.100 ;
        RECT 475.950 649.950 478.050 655.050 ;
        RECT 478.950 652.950 481.050 655.050 ;
        RECT 466.950 646.950 469.050 649.050 ;
        RECT 469.950 646.950 472.050 649.050 ;
        RECT 472.950 646.950 475.050 649.050 ;
        RECT 460.950 643.950 463.050 646.050 ;
        RECT 467.400 644.400 468.600 646.650 ;
        RECT 473.400 644.400 474.600 646.650 ;
        RECT 457.950 634.950 460.050 637.050 ;
        RECT 467.400 634.050 468.450 644.400 ;
        RECT 469.950 640.800 472.050 642.900 ;
        RECT 457.950 631.800 460.050 633.900 ;
        RECT 460.950 631.950 463.050 634.050 ;
        RECT 463.950 631.950 469.050 634.050 ;
        RECT 458.400 613.050 459.450 631.800 ;
        RECT 457.950 610.950 460.050 613.050 ;
        RECT 454.950 607.950 457.050 610.050 ;
        RECT 458.400 606.600 459.450 610.950 ;
        RECT 458.400 604.350 459.600 606.600 ;
        RECT 452.400 601.950 454.500 604.050 ;
        RECT 457.800 601.950 459.900 604.050 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 452.400 599.400 453.600 601.650 ;
        RECT 452.400 595.050 453.450 599.400 ;
        RECT 451.950 592.950 454.050 595.050 ;
        RECT 461.400 592.050 462.450 631.950 ;
        RECT 463.950 622.950 466.050 625.050 ;
        RECT 464.400 619.050 465.450 622.950 ;
        RECT 463.950 616.950 466.050 619.050 ;
        RECT 464.100 604.950 466.200 607.050 ;
        RECT 464.400 602.400 465.600 604.650 ;
        RECT 464.400 595.050 465.450 602.400 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 463.950 592.950 466.050 595.050 ;
        RECT 445.950 589.950 448.050 592.050 ;
        RECT 461.400 591.900 465.000 592.050 ;
        RECT 461.400 590.400 466.050 591.900 ;
        RECT 462.000 589.950 466.050 590.400 ;
        RECT 463.950 589.800 466.050 589.950 ;
        RECT 467.400 586.050 468.450 601.950 ;
        RECT 470.400 589.050 471.450 640.800 ;
        RECT 473.400 631.050 474.450 644.400 ;
        RECT 472.950 628.950 475.050 631.050 ;
        RECT 473.100 604.950 475.200 607.050 ;
        RECT 473.400 603.450 474.600 604.650 ;
        RECT 473.400 602.400 477.450 603.450 ;
        RECT 472.950 598.950 475.050 601.050 ;
        RECT 469.950 586.950 472.050 589.050 ;
        RECT 466.950 583.950 469.050 586.050 ;
        RECT 440.700 579.300 442.800 581.400 ;
        RECT 443.700 579.300 445.800 581.400 ;
        RECT 446.700 579.300 448.800 581.400 ;
        RECT 441.300 575.700 442.500 579.300 ;
        RECT 440.400 573.600 442.500 575.700 ;
        RECT 440.400 554.700 441.900 573.600 ;
        RECT 444.300 562.800 445.500 579.300 ;
        RECT 443.400 560.700 445.500 562.800 ;
        RECT 444.300 554.700 445.500 560.700 ;
        RECT 446.700 557.700 447.900 579.300 ;
        RECT 454.800 578.400 456.900 580.500 ;
        RECT 460.200 579.300 462.300 581.400 ;
        RECT 463.200 579.300 465.300 581.400 ;
        RECT 466.200 579.300 468.300 581.400 ;
        RECT 451.800 571.950 453.900 574.050 ;
        RECT 452.400 569.400 453.600 571.650 ;
        RECT 452.400 567.450 453.450 569.400 ;
        RECT 449.400 566.400 453.450 567.450 ;
        RECT 455.400 567.900 456.300 578.400 ;
        RECT 458.100 572.400 460.200 574.500 ;
        RECT 449.400 562.050 450.450 566.400 ;
        RECT 455.400 565.800 457.500 567.900 ;
        RECT 461.100 567.000 462.300 579.300 ;
        RECT 451.950 562.950 454.050 565.050 ;
        RECT 448.950 559.950 451.050 562.050 ;
        RECT 446.700 555.600 448.800 557.700 ;
        RECT 452.400 555.450 453.450 562.950 ;
        RECT 455.400 559.200 456.300 565.800 ;
        RECT 460.800 564.900 462.900 567.000 ;
        RECT 455.400 557.100 457.500 559.200 ;
        RECT 461.100 557.700 462.300 564.900 ;
        RECT 463.800 561.600 465.300 579.300 ;
        RECT 463.800 559.500 465.900 561.600 ;
        RECT 460.800 555.600 462.900 557.700 ;
        RECT 440.400 552.600 443.400 554.700 ;
        RECT 444.300 552.600 446.400 554.700 ;
        RECT 452.400 554.400 456.450 555.450 ;
        RECT 463.800 554.700 465.300 559.500 ;
        RECT 467.100 557.700 468.300 579.300 ;
        RECT 455.400 552.450 456.450 554.400 ;
        RECT 463.200 552.600 465.300 554.700 ;
        RECT 466.200 552.600 468.300 557.700 ;
        RECT 469.200 579.300 471.300 581.400 ;
        RECT 469.200 561.600 470.700 579.300 ;
        RECT 473.400 562.050 474.450 598.950 ;
        RECT 476.400 598.050 477.450 602.400 ;
        RECT 475.950 595.950 478.050 598.050 ;
        RECT 476.400 570.450 477.450 595.950 ;
        RECT 479.400 577.050 480.450 652.950 ;
        RECT 485.400 651.600 486.450 664.950 ;
        RECT 512.700 657.300 514.800 659.400 ;
        RECT 515.700 657.300 517.800 659.400 ;
        RECT 518.700 657.300 520.800 659.400 ;
        RECT 485.400 649.350 486.600 651.600 ;
        RECT 490.950 651.000 493.050 655.050 ;
        RECT 502.950 652.950 505.050 655.050 ;
        RECT 508.950 652.950 511.050 655.050 ;
        RECT 513.300 653.700 514.500 657.300 ;
        RECT 491.400 649.350 492.600 651.000 ;
        RECT 503.400 649.050 504.450 652.950 ;
        RECT 484.950 646.950 487.050 649.050 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 481.950 640.950 484.050 645.900 ;
        RECT 488.400 644.400 489.600 646.650 ;
        RECT 494.400 645.900 495.600 646.650 ;
        RECT 488.400 634.050 489.450 644.400 ;
        RECT 493.950 643.800 496.050 645.900 ;
        RECT 499.800 643.950 501.900 646.050 ;
        RECT 505.800 643.950 507.900 646.050 ;
        RECT 500.400 642.900 501.600 643.650 ;
        RECT 499.950 640.800 502.050 642.900 ;
        RECT 496.950 634.950 499.050 637.050 ;
        RECT 487.950 631.950 490.050 634.050 ;
        RECT 497.400 631.050 498.450 634.950 ;
        RECT 496.950 628.950 499.050 631.050 ;
        RECT 509.400 625.050 510.450 652.950 ;
        RECT 512.400 651.600 514.500 653.700 ;
        RECT 512.400 632.700 513.900 651.600 ;
        RECT 516.300 640.800 517.500 657.300 ;
        RECT 515.400 638.700 517.500 640.800 ;
        RECT 516.300 632.700 517.500 638.700 ;
        RECT 518.700 635.700 519.900 657.300 ;
        RECT 526.800 656.400 528.900 658.500 ;
        RECT 532.200 657.300 534.300 659.400 ;
        RECT 535.200 657.300 537.300 659.400 ;
        RECT 538.200 657.300 540.300 659.400 ;
        RECT 523.800 649.950 525.900 652.050 ;
        RECT 524.400 648.900 525.600 649.650 ;
        RECT 523.950 646.800 526.050 648.900 ;
        RECT 527.400 645.900 528.300 656.400 ;
        RECT 530.100 650.400 532.200 652.500 ;
        RECT 527.400 643.800 529.500 645.900 ;
        RECT 533.100 645.000 534.300 657.300 ;
        RECT 523.950 640.950 526.050 643.050 ;
        RECT 518.700 633.600 520.800 635.700 ;
        RECT 512.400 630.600 515.400 632.700 ;
        RECT 516.300 630.600 518.400 632.700 ;
        RECT 524.400 625.050 525.450 640.950 ;
        RECT 527.400 637.200 528.300 643.800 ;
        RECT 532.800 642.900 534.900 645.000 ;
        RECT 527.400 635.100 529.500 637.200 ;
        RECT 533.100 635.700 534.300 642.900 ;
        RECT 535.800 639.600 537.300 657.300 ;
        RECT 535.800 637.500 537.900 639.600 ;
        RECT 532.800 633.600 534.900 635.700 ;
        RECT 535.800 632.700 537.300 637.500 ;
        RECT 539.100 635.700 540.300 657.300 ;
        RECT 535.200 630.600 537.300 632.700 ;
        RECT 538.200 630.600 540.300 635.700 ;
        RECT 541.200 657.300 543.300 659.400 ;
        RECT 541.200 639.600 542.700 657.300 ;
        RECT 541.200 637.500 543.300 639.600 ;
        RECT 541.200 632.700 542.700 637.500 ;
        RECT 545.400 634.050 546.450 667.950 ;
        RECT 548.400 667.050 549.450 677.400 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 551.400 657.450 552.450 712.950 ;
        RECT 557.400 694.050 558.450 731.400 ;
        RECT 569.400 730.050 570.450 754.950 ;
        RECT 568.950 727.950 571.050 730.050 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 563.400 722.400 564.600 724.650 ;
        RECT 563.400 715.050 564.450 722.400 ;
        RECT 568.950 721.950 571.050 724.050 ;
        RECT 562.950 712.950 565.050 715.050 ;
        RECT 569.400 703.050 570.450 721.950 ;
        RECT 575.400 718.050 576.450 787.950 ;
        RECT 584.400 787.050 585.450 805.950 ;
        RECT 587.400 802.050 588.450 808.950 ;
        RECT 595.950 807.000 598.050 811.050 ;
        RECT 602.400 807.600 603.450 811.950 ;
        RECT 611.400 811.050 612.450 850.950 ;
        RECT 617.400 850.050 618.450 884.100 ;
        RECT 623.400 883.350 624.600 884.100 ;
        RECT 629.400 883.350 630.600 885.600 ;
        RECT 622.950 880.950 625.050 883.050 ;
        RECT 625.950 880.950 628.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 626.400 879.900 627.600 880.650 ;
        RECT 625.950 877.800 628.050 879.900 ;
        RECT 632.400 878.400 633.600 880.650 ;
        RECT 638.400 879.900 639.450 886.950 ;
        RECT 632.400 874.050 633.450 878.400 ;
        RECT 637.950 877.800 640.050 879.900 ;
        RECT 631.950 871.950 634.050 874.050 ;
        RECT 616.950 847.950 619.050 850.050 ;
        RECT 637.950 847.950 640.050 850.050 ;
        RECT 631.950 841.950 634.050 844.050 ;
        RECT 613.950 840.600 618.000 841.050 ;
        RECT 613.950 838.950 618.600 840.600 ;
        RECT 622.950 839.100 625.050 841.200 ;
        RECT 628.950 839.100 631.050 841.200 ;
        RECT 617.400 838.350 618.600 838.950 ;
        RECT 623.400 838.350 624.600 839.100 ;
        RECT 616.950 835.950 619.050 838.050 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 622.950 835.950 625.050 838.050 ;
        RECT 613.950 832.950 616.050 835.050 ;
        RECT 620.400 834.900 621.600 835.650 ;
        RECT 614.400 814.050 615.450 832.950 ;
        RECT 619.950 832.800 622.050 834.900 ;
        RECT 629.400 829.050 630.450 839.100 ;
        RECT 628.950 826.950 631.050 829.050 ;
        RECT 628.950 817.950 631.050 820.050 ;
        RECT 625.950 814.950 628.050 817.050 ;
        RECT 613.950 811.950 616.050 814.050 ;
        RECT 610.950 808.950 613.050 811.050 ;
        RECT 596.400 805.350 597.600 807.000 ;
        RECT 602.400 805.350 603.600 807.600 ;
        RECT 610.950 805.800 613.050 807.900 ;
        RECT 619.950 806.100 622.050 808.200 ;
        RECT 626.400 808.050 627.450 814.950 ;
        RECT 592.950 802.950 595.050 805.050 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 586.950 799.950 589.050 802.050 ;
        RECT 593.400 801.900 594.600 802.650 ;
        RECT 611.400 801.900 612.450 805.800 ;
        RECT 620.400 805.350 621.600 806.100 ;
        RECT 625.950 805.950 628.050 808.050 ;
        RECT 616.950 802.950 619.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 592.950 799.800 595.050 801.900 ;
        RECT 610.950 799.800 613.050 801.900 ;
        RECT 613.950 799.950 616.050 802.050 ;
        RECT 617.400 800.400 618.600 802.650 ;
        RECT 623.400 801.900 624.600 802.650 ;
        RECT 629.400 802.050 630.450 817.950 ;
        RECT 595.950 790.950 598.050 793.050 ;
        RECT 583.950 784.950 586.050 787.050 ;
        RECT 589.950 778.950 592.050 781.050 ;
        RECT 583.950 766.950 586.050 769.050 ;
        RECT 584.400 762.600 585.450 766.950 ;
        RECT 590.400 763.050 591.450 778.950 ;
        RECT 596.400 766.050 597.450 790.950 ;
        RECT 614.400 769.050 615.450 799.950 ;
        RECT 617.400 793.050 618.450 800.400 ;
        RECT 622.950 799.800 625.050 801.900 ;
        RECT 628.950 799.950 631.050 802.050 ;
        RECT 628.950 796.800 631.050 798.900 ;
        RECT 616.950 790.950 619.050 793.050 ;
        RECT 619.950 787.950 622.050 790.050 ;
        RECT 620.400 784.050 621.450 787.950 ;
        RECT 619.950 781.950 622.050 784.050 ;
        RECT 625.950 775.950 628.050 778.050 ;
        RECT 613.950 766.950 616.050 769.050 ;
        RECT 595.950 763.950 598.050 766.050 ;
        RECT 584.400 760.350 585.600 762.600 ;
        RECT 589.950 760.950 592.050 763.050 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 586.950 757.950 589.050 760.050 ;
        RECT 587.400 757.050 588.600 757.650 ;
        RECT 596.400 757.050 597.450 763.950 ;
        RECT 626.400 763.050 627.450 775.950 ;
        RECT 629.400 772.050 630.450 796.800 ;
        RECT 632.400 778.050 633.450 841.950 ;
        RECT 638.400 841.200 639.450 847.950 ;
        RECT 641.400 844.050 642.450 889.950 ;
        RECT 650.400 885.600 651.450 889.950 ;
        RECT 650.400 883.350 651.600 885.600 ;
        RECT 667.950 885.000 670.050 889.050 ;
        RECT 668.400 883.350 669.600 885.000 ;
        RECT 646.950 880.950 649.050 883.050 ;
        RECT 649.950 880.950 652.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 667.950 880.950 670.050 883.050 ;
        RECT 647.400 878.400 648.600 880.650 ;
        RECT 665.400 878.400 666.600 880.650 ;
        RECT 680.400 879.450 681.450 895.950 ;
        RECT 689.400 889.050 690.450 910.950 ;
        RECT 700.950 910.800 703.050 912.900 ;
        RECT 707.400 911.400 708.600 913.650 ;
        RECT 707.400 907.050 708.450 911.400 ;
        RECT 713.400 907.050 714.450 922.950 ;
        RECT 719.400 918.600 720.450 922.950 ;
        RECT 719.400 916.350 720.600 918.600 ;
        RECT 727.950 917.100 730.050 919.200 ;
        RECT 736.950 918.450 739.050 919.200 ;
        RECT 740.400 918.450 741.600 918.600 ;
        RECT 736.950 917.400 741.600 918.450 ;
        RECT 736.950 917.100 739.050 917.400 ;
        RECT 728.400 916.350 729.600 917.100 ;
        RECT 719.100 913.950 721.200 916.050 ;
        RECT 722.400 913.950 724.500 916.050 ;
        RECT 727.800 913.950 729.900 916.050 ;
        RECT 722.400 912.900 723.600 913.650 ;
        RECT 721.950 910.800 724.050 912.900 ;
        RECT 694.950 904.950 697.050 907.050 ;
        RECT 706.950 904.950 709.050 907.050 ;
        RECT 712.950 904.950 715.050 907.050 ;
        RECT 688.950 886.950 691.050 889.050 ;
        RECT 683.100 880.950 685.200 883.050 ;
        RECT 688.500 880.950 690.600 883.050 ;
        RECT 683.400 879.450 684.600 880.650 ;
        RECT 680.400 878.400 684.600 879.450 ;
        RECT 643.950 868.950 646.050 871.050 ;
        RECT 644.400 859.050 645.450 868.950 ;
        RECT 647.400 868.050 648.450 878.400 ;
        RECT 665.400 874.050 666.450 878.400 ;
        RECT 695.400 877.050 696.450 904.950 ;
        RECT 722.400 898.050 723.450 910.800 ;
        RECT 727.950 898.950 730.050 901.050 ;
        RECT 706.950 895.950 709.050 898.050 ;
        RECT 721.950 895.950 724.050 898.050 ;
        RECT 697.950 889.950 700.050 892.050 ;
        RECT 698.400 877.050 699.450 889.950 ;
        RECT 707.400 885.600 708.450 895.950 ;
        RECT 707.400 883.350 708.600 885.600 ;
        RECT 715.950 883.950 718.050 886.050 ;
        RECT 721.950 884.100 724.050 886.200 ;
        RECT 728.400 885.600 729.450 898.950 ;
        RECT 737.400 889.050 738.450 917.100 ;
        RECT 740.400 916.350 741.600 917.400 ;
        RECT 748.950 917.100 751.050 919.200 ;
        RECT 749.400 916.350 750.600 917.100 ;
        RECT 740.100 913.950 742.200 916.050 ;
        RECT 743.400 913.950 745.500 916.050 ;
        RECT 748.800 913.950 750.900 916.050 ;
        RECT 743.400 912.900 744.600 913.650 ;
        RECT 742.950 910.800 745.050 912.900 ;
        RECT 736.950 886.950 739.050 889.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 704.400 878.400 705.600 880.650 ;
        RECT 710.400 878.400 711.600 880.650 ;
        RECT 704.400 877.050 705.450 878.400 ;
        RECT 694.950 874.950 697.050 877.050 ;
        RECT 697.950 874.950 700.050 877.050 ;
        RECT 703.950 874.950 706.050 877.050 ;
        RECT 664.950 871.950 667.050 874.050 ;
        RECT 646.950 865.950 649.050 868.050 ;
        RECT 643.950 856.950 646.050 859.050 ;
        RECT 704.400 847.050 705.450 874.950 ;
        RECT 710.400 868.050 711.450 878.400 ;
        RECT 709.950 865.950 712.050 868.050 ;
        RECT 709.950 856.950 712.050 859.050 ;
        RECT 703.950 844.950 706.050 847.050 ;
        RECT 640.950 841.950 643.050 844.050 ;
        RECT 637.950 839.100 640.050 841.200 ;
        RECT 661.950 839.100 664.050 841.200 ;
        RECT 676.950 839.100 679.050 841.200 ;
        RECT 682.950 839.100 685.050 841.200 ;
        RECT 694.950 839.100 697.050 841.200 ;
        RECT 704.400 840.450 705.600 840.600 ;
        RECT 704.400 839.400 708.450 840.450 ;
        RECT 638.400 838.350 639.600 839.100 ;
        RECT 662.400 838.350 663.600 839.100 ;
        RECT 677.400 838.350 678.600 839.100 ;
        RECT 683.400 838.350 684.600 839.100 ;
        RECT 637.950 835.950 640.050 838.050 ;
        RECT 640.950 835.950 643.050 838.050 ;
        RECT 653.100 835.950 655.200 838.050 ;
        RECT 656.100 835.950 658.200 838.050 ;
        RECT 661.800 835.950 663.900 838.050 ;
        RECT 664.800 835.950 666.900 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 682.950 835.950 685.050 838.050 ;
        RECT 641.400 833.400 642.600 835.650 ;
        RECT 656.400 834.900 657.600 835.650 ;
        RECT 641.400 820.050 642.450 833.400 ;
        RECT 655.800 832.800 657.900 834.900 ;
        RECT 658.950 832.950 661.050 835.050 ;
        RECT 680.400 834.900 681.600 835.650 ;
        RECT 659.400 829.050 660.450 832.950 ;
        RECT 679.950 832.800 682.050 834.900 ;
        RECT 658.950 826.950 661.050 829.050 ;
        RECT 670.950 826.950 673.050 829.050 ;
        RECT 640.950 817.950 643.050 820.050 ;
        RECT 640.950 806.100 643.050 808.200 ;
        RECT 646.950 806.100 649.050 808.200 ;
        RECT 641.400 805.350 642.600 806.100 ;
        RECT 647.400 805.350 648.600 806.100 ;
        RECT 637.950 802.950 640.050 805.050 ;
        RECT 640.950 802.950 643.050 805.050 ;
        RECT 643.950 802.950 646.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 634.950 796.950 637.050 802.050 ;
        RECT 638.400 801.000 639.600 802.650 ;
        RECT 644.400 801.000 645.600 802.650 ;
        RECT 650.400 801.900 651.600 802.650 ;
        RECT 637.950 796.950 640.050 801.000 ;
        RECT 643.950 796.950 646.050 801.000 ;
        RECT 649.950 799.800 652.050 801.900 ;
        RECT 665.400 800.400 666.600 802.650 ;
        RECT 661.950 796.950 664.050 799.050 ;
        RECT 649.950 787.950 652.050 790.050 ;
        RECT 631.950 775.950 634.050 778.050 ;
        RECT 628.950 769.950 631.050 772.050 ;
        RECT 643.950 769.950 646.050 772.050 ;
        RECT 628.950 766.800 631.050 768.900 ;
        RECT 598.950 762.600 603.000 763.050 ;
        RECT 598.950 760.950 603.600 762.600 ;
        RECT 625.950 760.950 628.050 763.050 ;
        RECT 602.400 760.350 603.600 760.950 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 625.950 757.800 628.050 759.900 ;
        RECT 577.950 754.950 580.050 757.050 ;
        RECT 587.400 755.400 592.050 757.050 ;
        RECT 588.000 754.950 592.050 755.400 ;
        RECT 595.950 754.950 598.050 757.050 ;
        RECT 605.400 756.000 606.600 757.650 ;
        RECT 617.400 756.900 618.600 757.650 ;
        RECT 578.400 748.050 579.450 754.950 ;
        RECT 604.950 754.050 607.050 756.000 ;
        RECT 616.950 754.800 619.050 756.900 ;
        RECT 622.950 754.950 625.050 757.050 ;
        RECT 598.950 751.950 601.050 754.050 ;
        RECT 604.800 753.000 607.050 754.050 ;
        RECT 604.800 751.950 606.900 753.000 ;
        RECT 607.950 751.950 610.050 754.050 ;
        RECT 577.950 745.950 580.050 748.050 ;
        RECT 592.950 745.950 595.050 748.050 ;
        RECT 586.950 736.950 589.050 739.050 ;
        RECT 587.400 729.600 588.450 736.950 ;
        RECT 587.400 727.350 588.600 729.600 ;
        RECT 581.100 724.950 583.200 727.050 ;
        RECT 586.500 724.950 588.600 727.050 ;
        RECT 589.800 724.950 591.900 727.050 ;
        RECT 581.400 722.400 582.600 724.650 ;
        RECT 590.400 722.400 591.600 724.650 ;
        RECT 574.950 715.950 577.050 718.050 ;
        RECT 568.950 700.950 571.050 703.050 ;
        RECT 574.950 700.950 577.050 703.050 ;
        RECT 556.950 691.950 559.050 694.050 ;
        RECT 562.950 683.100 565.050 685.200 ;
        RECT 568.950 684.000 571.050 688.050 ;
        RECT 563.400 682.350 564.600 683.100 ;
        RECT 569.400 682.350 570.600 684.000 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 562.950 679.950 565.050 682.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 568.950 679.950 571.050 682.050 ;
        RECT 560.400 678.900 561.600 679.650 ;
        RECT 559.950 676.800 562.050 678.900 ;
        RECT 566.400 677.400 567.600 679.650 ;
        RECT 562.950 673.950 565.050 676.050 ;
        RECT 563.400 667.050 564.450 673.950 ;
        RECT 566.400 669.450 567.450 677.400 ;
        RECT 575.400 676.050 576.450 700.950 ;
        RECT 581.400 688.200 582.450 722.400 ;
        RECT 583.950 718.950 586.050 721.050 ;
        RECT 584.400 703.050 585.450 718.950 ;
        RECT 590.400 715.050 591.450 722.400 ;
        RECT 589.950 712.950 592.050 715.050 ;
        RECT 583.950 700.950 586.050 703.050 ;
        RECT 580.950 686.100 583.050 688.200 ;
        RECT 580.950 682.950 583.050 685.050 ;
        RECT 586.950 684.000 589.050 688.050 ;
        RECT 593.400 685.050 594.450 745.950 ;
        RECT 595.950 742.950 598.050 745.050 ;
        RECT 596.400 688.050 597.450 742.950 ;
        RECT 599.400 721.050 600.450 751.950 ;
        RECT 608.400 739.050 609.450 751.950 ;
        RECT 616.950 745.950 619.050 748.050 ;
        RECT 607.950 736.950 610.050 739.050 ;
        RECT 613.950 733.950 616.050 736.050 ;
        RECT 610.950 730.800 613.050 732.900 ;
        RECT 601.950 728.100 604.050 730.200 ;
        RECT 602.400 727.350 603.600 728.100 ;
        RECT 602.400 724.950 604.500 727.050 ;
        RECT 607.800 724.950 609.900 727.050 ;
        RECT 608.400 723.000 609.600 724.650 ;
        RECT 598.950 718.950 601.050 721.050 ;
        RECT 607.950 718.950 610.050 723.000 ;
        RECT 611.400 720.450 612.450 730.800 ;
        RECT 614.400 724.050 615.450 733.950 ;
        RECT 617.400 733.050 618.450 745.950 ;
        RECT 619.950 736.950 622.050 739.050 ;
        RECT 616.950 730.950 619.050 733.050 ;
        RECT 620.400 729.600 621.450 736.950 ;
        RECT 623.400 733.050 624.450 754.950 ;
        RECT 626.400 739.050 627.450 757.800 ;
        RECT 629.400 748.050 630.450 766.800 ;
        RECT 631.950 761.100 634.050 763.200 ;
        RECT 640.950 762.000 643.050 766.050 ;
        RECT 632.400 760.350 633.600 761.100 ;
        RECT 641.400 760.350 642.600 762.000 ;
        RECT 632.100 757.950 634.200 760.050 ;
        RECT 635.400 757.950 637.500 760.050 ;
        RECT 640.800 757.950 642.900 760.050 ;
        RECT 635.400 755.400 636.600 757.650 ;
        RECT 628.950 745.950 631.050 748.050 ;
        RECT 625.950 736.950 628.050 739.050 ;
        RECT 625.950 733.800 628.050 735.900 ;
        RECT 622.950 730.950 625.050 733.050 ;
        RECT 626.400 729.600 627.450 733.800 ;
        RECT 635.400 730.050 636.450 755.400 ;
        RECT 620.400 727.350 621.600 729.600 ;
        RECT 626.400 727.350 627.600 729.600 ;
        RECT 634.950 727.950 637.050 730.050 ;
        RECT 644.400 729.600 645.450 769.950 ;
        RECT 646.950 763.950 649.050 769.050 ;
        RECT 646.950 760.800 649.050 762.900 ;
        RECT 647.400 745.050 648.450 760.800 ;
        RECT 646.950 742.950 649.050 745.050 ;
        RECT 650.400 742.050 651.450 787.950 ;
        RECT 662.400 787.050 663.450 796.950 ;
        RECT 661.950 784.950 664.050 787.050 ;
        RECT 658.950 772.950 661.050 775.050 ;
        RECT 652.950 766.950 658.050 769.050 ;
        RECT 659.400 765.450 660.450 772.950 ;
        RECT 656.400 764.400 660.450 765.450 ;
        RECT 656.400 763.200 657.450 764.400 ;
        RECT 655.950 761.100 658.050 763.200 ;
        RECT 662.400 762.600 663.450 784.950 ;
        RECT 665.400 781.050 666.450 800.400 ;
        RECT 667.950 799.950 670.050 802.050 ;
        RECT 664.950 778.950 667.050 781.050 ;
        RECT 656.400 760.350 657.600 761.100 ;
        RECT 662.400 760.350 663.600 762.600 ;
        RECT 668.400 760.050 669.450 799.950 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 667.950 757.950 670.050 760.050 ;
        RECT 659.400 755.400 660.600 757.650 ;
        RECT 659.400 754.050 660.450 755.400 ;
        RECT 658.950 751.950 661.050 754.050 ;
        RECT 659.400 748.050 660.450 751.950 ;
        RECT 658.950 745.950 661.050 748.050 ;
        RECT 649.950 739.950 652.050 742.050 ;
        RECT 644.400 727.350 645.600 729.600 ;
        RECT 646.950 727.950 649.050 733.050 ;
        RECT 658.950 728.100 661.050 730.200 ;
        RECT 671.400 729.450 672.450 826.950 ;
        RECT 688.950 823.950 691.050 826.050 ;
        RECT 673.950 811.950 676.050 814.050 ;
        RECT 674.400 808.050 675.450 811.950 ;
        RECT 673.950 805.950 676.050 808.050 ;
        RECT 679.950 806.100 682.050 808.200 ;
        RECT 680.400 805.350 681.600 806.100 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 677.400 801.000 678.600 802.650 ;
        RECT 676.950 796.950 679.050 801.000 ;
        RECT 685.950 799.950 688.050 802.050 ;
        RECT 686.400 796.050 687.450 799.950 ;
        RECT 685.950 793.950 688.050 796.050 ;
        RECT 689.400 789.450 690.450 823.950 ;
        RECT 695.400 823.050 696.450 839.100 ;
        RECT 704.400 838.350 705.600 839.400 ;
        RECT 698.400 835.950 700.500 838.050 ;
        RECT 703.800 835.950 705.900 838.050 ;
        RECT 698.400 834.900 699.600 835.650 ;
        RECT 697.950 832.800 700.050 834.900 ;
        RECT 698.400 829.050 699.450 832.800 ;
        RECT 697.950 826.950 700.050 829.050 ;
        RECT 703.950 826.950 706.050 829.050 ;
        RECT 694.950 820.950 697.050 823.050 ;
        RECT 700.950 820.950 703.050 823.050 ;
        RECT 691.950 817.950 694.050 820.050 ;
        RECT 692.400 808.050 693.450 817.950 ;
        RECT 691.950 805.950 694.050 808.050 ;
        RECT 701.400 807.600 702.450 820.950 ;
        RECT 704.400 814.050 705.450 826.950 ;
        RECT 703.950 811.950 706.050 814.050 ;
        RECT 707.400 808.050 708.450 839.400 ;
        RECT 692.400 801.900 693.450 805.950 ;
        RECT 701.400 805.350 702.600 807.600 ;
        RECT 706.950 805.950 709.050 808.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 698.400 801.900 699.600 802.650 ;
        RECT 691.950 799.800 694.050 801.900 ;
        RECT 697.950 799.800 700.050 801.900 ;
        RECT 704.400 800.400 705.600 802.650 ;
        RECT 710.400 801.450 711.450 856.950 ;
        RECT 716.400 850.050 717.450 883.950 ;
        RECT 722.400 883.350 723.600 884.100 ;
        RECT 728.400 883.350 729.600 885.600 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 725.400 879.000 726.600 880.650 ;
        RECT 731.400 879.900 732.600 880.650 ;
        RECT 737.400 879.900 738.450 886.950 ;
        RECT 743.400 885.600 744.450 910.800 ;
        RECT 743.400 883.350 744.600 885.600 ;
        RECT 748.950 885.000 751.050 889.050 ;
        RECT 752.400 886.050 753.450 922.950 ;
        RECT 763.950 917.100 766.050 919.200 ;
        RECT 770.400 918.600 771.450 922.950 ;
        RECT 764.400 916.350 765.600 917.100 ;
        RECT 770.400 916.350 771.600 918.600 ;
        RECT 763.950 913.950 766.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 769.950 913.950 772.050 916.050 ;
        RECT 772.950 913.950 775.050 916.050 ;
        RECT 767.400 912.900 768.600 913.650 ;
        RECT 766.950 910.800 769.050 912.900 ;
        RECT 773.400 911.400 774.600 913.650 ;
        RECT 779.400 913.050 780.450 922.950 ;
        RECT 787.950 917.100 790.050 919.200 ;
        RECT 795.000 918.600 799.050 919.050 ;
        RECT 788.400 916.350 789.600 917.100 ;
        RECT 794.400 916.950 799.050 918.600 ;
        RECT 799.950 916.950 802.050 919.050 ;
        RECT 802.950 916.950 805.050 919.050 ;
        RECT 808.950 917.100 811.050 919.200 ;
        RECT 817.950 917.100 820.050 919.200 ;
        RECT 823.950 917.100 826.050 919.200 ;
        RECT 830.400 918.600 831.450 925.950 ;
        RECT 845.400 918.600 846.450 925.950 ;
        RECT 850.950 922.950 853.050 925.050 ;
        RECT 851.400 919.200 852.450 922.950 ;
        RECT 794.400 916.350 795.600 916.950 ;
        RECT 784.950 913.950 787.050 916.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 793.950 913.950 796.050 916.050 ;
        RECT 773.400 898.050 774.450 911.400 ;
        RECT 778.950 910.950 781.050 913.050 ;
        RECT 785.400 911.400 786.600 913.650 ;
        RECT 791.400 912.900 792.600 913.650 ;
        RECT 800.400 912.900 801.450 916.950 ;
        RECT 772.950 897.450 775.050 898.050 ;
        RECT 772.950 896.400 777.450 897.450 ;
        RECT 772.950 895.950 775.050 896.400 ;
        RECT 754.950 886.950 757.050 889.050 ;
        RECT 749.400 883.350 750.600 885.000 ;
        RECT 751.950 883.950 754.050 886.050 ;
        RECT 742.950 880.950 745.050 883.050 ;
        RECT 745.950 880.950 748.050 883.050 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 746.400 879.900 747.600 880.650 ;
        RECT 755.400 880.050 756.450 886.950 ;
        RECT 760.950 885.000 763.050 889.050 ;
        RECT 761.400 883.350 762.600 885.000 ;
        RECT 766.950 884.100 769.050 886.200 ;
        RECT 767.400 883.350 768.600 884.100 ;
        RECT 772.950 883.950 775.050 889.050 ;
        RECT 760.950 880.950 763.050 883.050 ;
        RECT 763.950 880.950 766.050 883.050 ;
        RECT 766.950 880.950 769.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 724.950 874.950 727.050 879.000 ;
        RECT 730.950 877.800 733.050 879.900 ;
        RECT 736.950 877.800 739.050 879.900 ;
        RECT 745.950 877.800 748.050 879.900 ;
        RECT 754.950 877.950 757.050 880.050 ;
        RECT 764.400 879.000 765.600 880.650 ;
        RECT 770.400 879.900 771.600 880.650 ;
        RECT 776.400 880.050 777.450 896.400 ;
        RECT 785.400 889.050 786.450 911.400 ;
        RECT 790.950 910.800 793.050 912.900 ;
        RECT 799.950 910.800 802.050 912.900 ;
        RECT 787.950 895.950 790.050 898.050 ;
        RECT 788.400 889.050 789.450 895.950 ;
        RECT 778.950 886.950 781.050 889.050 ;
        RECT 784.800 886.950 786.900 889.050 ;
        RECT 724.950 859.950 727.050 862.050 ;
        RECT 715.950 847.950 718.050 850.050 ;
        RECT 721.950 844.950 724.050 847.050 ;
        RECT 722.400 841.200 723.450 844.950 ;
        RECT 721.950 839.100 724.050 841.200 ;
        RECT 722.400 838.350 723.600 839.100 ;
        RECT 716.400 835.950 718.500 838.050 ;
        RECT 721.800 835.950 723.900 838.050 ;
        RECT 716.400 834.900 717.600 835.650 ;
        RECT 715.950 832.800 718.050 834.900 ;
        RECT 718.950 814.950 721.050 817.050 ;
        RECT 719.400 807.600 720.450 814.950 ;
        RECT 725.400 807.600 726.450 859.950 ;
        RECT 731.400 843.450 732.450 877.800 ;
        RECT 763.950 874.950 766.050 879.000 ;
        RECT 769.950 877.800 772.050 879.900 ;
        RECT 775.950 877.950 778.050 880.050 ;
        RECT 775.950 874.800 778.050 876.900 ;
        RECT 739.950 847.950 742.050 850.050 ;
        RECT 728.400 842.400 732.450 843.450 ;
        RECT 728.400 829.050 729.450 842.400 ;
        RECT 730.950 838.950 733.050 841.050 ;
        RECT 740.400 840.600 741.450 847.950 ;
        RECT 731.400 834.900 732.450 838.950 ;
        RECT 740.400 838.350 741.600 840.600 ;
        RECT 745.950 839.100 748.050 841.200 ;
        RECT 754.950 839.100 757.050 841.200 ;
        RECT 760.950 840.000 763.050 844.050 ;
        RECT 776.400 841.200 777.450 874.800 ;
        RECT 779.400 844.050 780.450 886.950 ;
        RECT 787.950 885.000 790.050 889.050 ;
        RECT 788.400 883.350 789.600 885.000 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 785.400 878.400 786.600 880.650 ;
        RECT 791.400 878.400 792.600 880.650 ;
        RECT 800.400 879.900 801.450 910.800 ;
        RECT 803.400 901.050 804.450 916.950 ;
        RECT 809.400 916.350 810.600 917.100 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 812.400 911.400 813.600 913.650 ;
        RECT 802.950 898.950 805.050 901.050 ;
        RECT 808.950 898.950 811.050 901.050 ;
        RECT 809.400 885.600 810.450 898.950 ;
        RECT 812.400 889.050 813.450 911.400 ;
        RECT 818.400 907.050 819.450 917.100 ;
        RECT 824.400 916.350 825.600 917.100 ;
        RECT 830.400 916.350 831.600 918.600 ;
        RECT 845.400 916.350 846.600 918.600 ;
        RECT 850.950 917.100 853.050 919.200 ;
        RECT 851.400 916.350 852.600 917.100 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 826.950 913.950 829.050 916.050 ;
        RECT 829.950 913.950 832.050 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 844.950 913.950 847.050 916.050 ;
        RECT 847.950 913.950 850.050 916.050 ;
        RECT 850.950 913.950 853.050 916.050 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 827.400 912.900 828.600 913.650 ;
        RECT 833.400 912.900 834.600 913.650 ;
        RECT 848.400 912.900 849.600 913.650 ;
        RECT 826.950 910.800 829.050 912.900 ;
        RECT 832.950 910.800 835.050 912.900 ;
        RECT 841.950 910.800 844.050 912.900 ;
        RECT 817.950 904.950 820.050 907.050 ;
        RECT 835.950 904.950 838.050 910.050 ;
        RECT 832.950 889.950 835.050 892.050 ;
        RECT 811.950 886.950 814.050 889.050 ;
        RECT 809.400 883.350 810.600 885.600 ;
        RECT 814.950 884.100 817.050 886.200 ;
        RECT 815.400 883.350 816.600 884.100 ;
        RECT 820.950 883.950 823.050 886.050 ;
        RECT 826.950 884.100 829.050 886.200 ;
        RECT 833.400 885.600 834.450 889.950 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 806.400 879.900 807.600 880.650 ;
        RECT 812.400 879.900 813.600 880.650 ;
        RECT 821.400 879.900 822.450 883.950 ;
        RECT 827.400 883.350 828.600 884.100 ;
        RECT 833.400 883.350 834.600 885.600 ;
        RECT 826.950 880.950 829.050 883.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 830.400 879.900 831.600 880.650 ;
        RECT 785.400 862.050 786.450 878.400 ;
        RECT 787.950 865.950 790.050 868.050 ;
        RECT 784.950 859.950 787.050 862.050 ;
        RECT 788.400 855.450 789.450 865.950 ;
        RECT 791.400 859.050 792.450 878.400 ;
        RECT 799.950 877.800 802.050 879.900 ;
        RECT 805.950 877.800 808.050 879.900 ;
        RECT 811.950 877.800 814.050 879.900 ;
        RECT 820.950 877.800 823.050 879.900 ;
        RECT 829.950 877.800 832.050 879.900 ;
        RECT 836.400 878.400 837.600 880.650 ;
        RECT 836.400 868.050 837.450 878.400 ;
        RECT 835.950 865.950 838.050 868.050 ;
        RECT 808.950 862.950 811.050 865.050 ;
        RECT 790.950 856.950 793.050 859.050 ;
        RECT 802.950 856.950 805.050 859.050 ;
        RECT 788.400 854.400 792.450 855.450 ;
        RECT 778.950 843.450 781.050 844.050 ;
        RECT 778.950 842.400 783.450 843.450 ;
        RECT 778.950 841.950 781.050 842.400 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 737.400 834.900 738.600 835.650 ;
        RECT 730.950 832.800 733.050 834.900 ;
        RECT 736.950 832.800 739.050 834.900 ;
        RECT 727.950 826.950 730.050 829.050 ;
        RECT 728.400 811.050 729.450 826.950 ;
        RECT 746.400 826.050 747.450 839.100 ;
        RECT 755.400 838.350 756.600 839.100 ;
        RECT 761.400 838.350 762.600 840.000 ;
        RECT 766.950 838.950 769.050 841.050 ;
        RECT 775.950 839.100 778.050 841.200 ;
        RECT 782.400 840.600 783.450 842.400 ;
        RECT 751.950 835.950 754.050 838.050 ;
        RECT 754.950 835.950 757.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 752.400 833.400 753.600 835.650 ;
        RECT 758.400 834.900 759.600 835.650 ;
        RECT 767.400 834.900 768.450 838.950 ;
        RECT 776.400 838.350 777.600 839.100 ;
        RECT 782.400 838.350 783.600 840.600 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 775.950 835.950 778.050 838.050 ;
        RECT 778.950 835.950 781.050 838.050 ;
        RECT 781.950 835.950 784.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 745.950 823.950 748.050 826.050 ;
        RECT 752.400 817.050 753.450 833.400 ;
        RECT 757.950 832.800 760.050 834.900 ;
        RECT 766.950 832.800 769.050 834.900 ;
        RECT 766.950 817.950 769.050 820.050 ;
        RECT 733.950 814.950 736.050 817.050 ;
        RECT 751.950 814.950 754.050 817.050 ;
        RECT 727.950 808.950 730.050 811.050 ;
        RECT 719.400 805.350 720.600 807.600 ;
        RECT 725.400 805.350 726.600 807.600 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 707.400 800.400 711.450 801.450 ;
        RECT 692.400 793.050 693.450 799.800 ;
        RECT 704.400 796.050 705.450 800.400 ;
        RECT 694.950 793.950 700.050 796.050 ;
        RECT 703.950 793.950 706.050 796.050 ;
        RECT 691.950 790.950 694.050 793.050 ;
        RECT 689.400 788.400 693.450 789.450 ;
        RECT 676.950 781.950 679.050 784.050 ;
        RECT 677.400 775.050 678.450 781.950 ;
        RECT 676.950 772.950 679.050 775.050 ;
        RECT 679.950 766.950 682.050 769.050 ;
        RECT 680.400 762.600 681.450 766.950 ;
        RECT 680.400 760.350 681.600 762.600 ;
        RECT 685.950 762.000 688.050 766.050 ;
        RECT 686.400 760.350 687.600 762.000 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 677.400 755.400 678.600 757.650 ;
        RECT 683.400 756.900 684.600 757.650 ;
        RECT 692.400 757.050 693.450 788.400 ;
        RECT 707.400 784.050 708.450 800.400 ;
        RECT 712.950 799.800 715.050 801.900 ;
        RECT 716.400 800.400 717.600 802.650 ;
        RECT 722.400 800.400 723.600 802.650 ;
        RECT 728.400 801.900 729.600 802.650 ;
        RECT 709.950 784.950 712.050 787.050 ;
        RECT 706.950 781.950 709.050 784.050 ;
        RECT 694.950 775.950 697.050 778.050 ;
        RECT 677.400 748.050 678.450 755.400 ;
        RECT 682.950 754.800 685.050 756.900 ;
        RECT 691.950 754.950 694.050 757.050 ;
        RECT 695.400 754.050 696.450 775.950 ;
        RECT 710.400 769.050 711.450 784.950 ;
        RECT 713.400 778.050 714.450 799.800 ;
        RECT 716.400 793.050 717.450 800.400 ;
        RECT 715.950 790.950 718.050 793.050 ;
        RECT 712.950 775.950 715.050 778.050 ;
        RECT 718.950 775.950 721.050 778.050 ;
        RECT 703.950 766.950 706.050 769.050 ;
        RECT 709.950 766.950 712.050 769.050 ;
        RECT 704.400 762.600 705.450 766.950 ;
        RECT 715.950 763.950 718.050 766.050 ;
        RECT 704.400 760.350 705.600 762.600 ;
        RECT 709.950 761.100 712.050 763.200 ;
        RECT 710.400 760.350 711.600 761.100 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 701.400 755.400 702.600 757.650 ;
        RECT 707.400 755.400 708.600 757.650 ;
        RECT 694.950 751.950 697.050 754.050 ;
        RECT 676.950 745.950 679.050 748.050 ;
        RECT 682.950 745.950 685.050 748.050 ;
        RECT 683.400 742.050 684.450 745.950 ;
        RECT 682.950 739.950 685.050 742.050 ;
        RECT 688.950 739.950 691.050 742.050 ;
        RECT 676.950 733.950 679.050 736.050 ;
        RECT 668.400 728.400 672.450 729.450 ;
        RECT 677.400 729.600 678.450 733.950 ;
        RECT 659.400 727.350 660.600 728.100 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 622.950 724.950 625.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 628.950 724.950 631.050 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 613.950 721.950 616.050 724.050 ;
        RECT 623.400 723.000 624.600 724.650 ;
        RECT 629.400 723.000 630.600 724.650 ;
        RECT 611.400 719.400 615.450 720.450 ;
        RECT 598.950 712.950 601.050 715.050 ;
        RECT 595.950 685.950 598.050 688.050 ;
        RECT 581.400 682.350 582.600 682.950 ;
        RECT 587.400 682.350 588.600 684.000 ;
        RECT 592.950 682.950 595.050 685.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 589.950 679.950 592.050 682.050 ;
        RECT 584.400 677.400 585.600 679.650 ;
        RECT 590.400 677.400 591.600 679.650 ;
        RECT 574.950 673.950 577.050 676.050 ;
        RECT 580.950 673.950 583.050 676.050 ;
        RECT 566.400 668.400 570.450 669.450 ;
        RECT 562.950 664.950 565.050 667.050 ;
        RECT 551.400 656.400 555.450 657.450 ;
        RECT 547.950 648.450 550.050 652.050 ;
        RECT 551.400 648.450 552.600 648.600 ;
        RECT 547.950 648.000 552.600 648.450 ;
        RECT 548.400 647.400 552.600 648.000 ;
        RECT 551.400 646.350 552.600 647.400 ;
        RECT 550.800 643.950 552.900 646.050 ;
        RECT 541.200 630.600 543.300 632.700 ;
        RECT 544.950 631.950 547.050 634.050 ;
        RECT 554.400 628.050 555.450 656.400 ;
        RECT 559.950 655.950 562.050 658.050 ;
        RECT 560.400 648.600 561.450 655.950 ;
        RECT 560.400 646.350 561.600 648.600 ;
        RECT 559.800 643.950 561.900 646.050 ;
        RECT 563.400 631.050 564.450 664.950 ;
        RECT 569.400 661.050 570.450 668.400 ;
        RECT 571.950 667.950 574.050 670.050 ;
        RECT 568.950 658.950 571.050 661.050 ;
        RECT 572.400 658.050 573.450 667.950 ;
        RECT 581.400 660.450 582.450 673.950 ;
        RECT 584.400 664.050 585.450 677.400 ;
        RECT 590.400 676.050 591.450 677.400 ;
        RECT 596.400 676.050 597.450 685.950 ;
        RECT 586.950 673.950 589.050 676.050 ;
        RECT 590.400 674.400 595.050 676.050 ;
        RECT 591.000 673.950 595.050 674.400 ;
        RECT 595.950 673.950 598.050 676.050 ;
        RECT 583.950 661.950 586.050 664.050 ;
        RECT 581.400 659.400 585.450 660.450 ;
        RECT 565.950 655.950 568.050 658.050 ;
        RECT 571.950 655.950 574.050 658.050 ;
        RECT 566.400 652.050 567.450 655.950 ;
        RECT 568.950 652.950 571.050 655.050 ;
        RECT 565.950 649.950 568.050 652.050 ;
        RECT 562.950 628.950 565.050 631.050 ;
        RECT 538.950 625.950 541.050 628.050 ;
        RECT 553.950 625.950 556.050 628.050 ;
        RECT 508.950 622.950 511.050 625.050 ;
        RECT 514.950 622.950 517.050 625.050 ;
        RECT 523.950 622.950 526.050 625.050 ;
        RECT 482.700 618.300 484.800 620.400 ;
        RECT 483.300 613.500 484.800 618.300 ;
        RECT 482.700 611.400 484.800 613.500 ;
        RECT 483.300 593.700 484.800 611.400 ;
        RECT 482.700 591.600 484.800 593.700 ;
        RECT 485.700 615.300 487.800 620.400 ;
        RECT 488.700 618.300 490.800 620.400 ;
        RECT 507.600 618.300 509.700 620.400 ;
        RECT 510.600 618.300 513.600 620.400 ;
        RECT 485.700 593.700 486.900 615.300 ;
        RECT 488.700 613.500 490.200 618.300 ;
        RECT 491.100 615.300 493.200 617.400 ;
        RECT 488.100 611.400 490.200 613.500 ;
        RECT 488.700 593.700 490.200 611.400 ;
        RECT 491.700 608.100 492.900 615.300 ;
        RECT 496.500 613.800 498.600 615.900 ;
        RECT 505.200 615.300 507.300 617.400 ;
        RECT 491.100 606.000 493.200 608.100 ;
        RECT 497.700 607.200 498.600 613.800 ;
        RECT 491.700 593.700 492.900 606.000 ;
        RECT 496.500 605.100 498.600 607.200 ;
        RECT 493.800 598.500 495.900 600.600 ;
        RECT 497.700 594.600 498.600 605.100 ;
        RECT 499.950 603.000 502.050 607.050 ;
        RECT 500.400 601.350 501.600 603.000 ;
        RECT 500.100 598.950 502.200 601.050 ;
        RECT 485.700 591.600 487.800 593.700 ;
        RECT 488.700 591.600 490.800 593.700 ;
        RECT 491.700 591.600 493.800 593.700 ;
        RECT 497.100 592.500 499.200 594.600 ;
        RECT 506.100 593.700 507.300 615.300 ;
        RECT 508.500 612.300 509.700 618.300 ;
        RECT 508.500 610.200 510.600 612.300 ;
        RECT 508.500 593.700 509.700 610.200 ;
        RECT 512.100 599.400 513.600 618.300 ;
        RECT 511.500 597.300 513.600 599.400 ;
        RECT 515.400 598.050 516.450 622.950 ;
        RECT 524.400 609.600 525.450 622.950 ;
        RECT 535.950 613.950 538.050 616.050 ;
        RECT 524.400 607.350 525.600 609.600 ;
        RECT 518.100 604.950 520.200 607.050 ;
        RECT 524.100 604.950 526.200 607.050 ;
        RECT 532.950 604.950 535.050 607.050 ;
        RECT 529.950 598.800 532.050 600.900 ;
        RECT 511.500 593.700 512.700 597.300 ;
        RECT 514.950 595.950 517.050 598.050 ;
        RECT 505.200 591.600 507.300 593.700 ;
        RECT 508.200 591.600 510.300 593.700 ;
        RECT 511.200 591.600 513.300 593.700 ;
        RECT 514.950 592.800 517.050 594.900 ;
        RECT 481.950 586.950 484.050 589.050 ;
        RECT 493.950 586.950 496.050 589.050 ;
        RECT 478.950 574.950 481.050 577.050 ;
        RECT 478.950 570.450 481.050 571.200 ;
        RECT 476.400 569.400 481.050 570.450 ;
        RECT 478.950 569.100 481.050 569.400 ;
        RECT 479.400 568.350 480.600 569.100 ;
        RECT 478.800 565.950 480.900 568.050 ;
        RECT 475.950 562.950 478.050 565.050 ;
        RECT 469.200 559.500 471.300 561.600 ;
        RECT 472.950 559.950 475.050 562.050 ;
        RECT 469.200 554.700 470.700 559.500 ;
        RECT 469.200 552.600 471.300 554.700 ;
        RECT 455.400 551.400 459.450 552.450 ;
        RECT 448.950 547.950 451.050 550.050 ;
        RECT 436.950 544.950 439.050 547.050 ;
        RECT 428.400 542.400 432.450 543.450 ;
        RECT 406.950 535.950 409.050 538.050 ;
        RECT 410.400 535.050 411.450 541.950 ;
        RECT 418.950 535.950 421.050 538.050 ;
        RECT 409.950 532.950 412.050 535.050 ;
        RECT 401.400 527.400 405.450 528.450 ;
        RECT 419.400 528.600 420.450 535.950 ;
        RECT 421.950 529.950 424.050 532.050 ;
        RECT 398.400 526.350 399.600 527.100 ;
        RECT 392.400 523.950 394.500 526.050 ;
        RECT 397.800 523.950 399.900 526.050 ;
        RECT 392.400 522.450 393.600 523.650 ;
        RECT 389.400 521.400 393.600 522.450 ;
        RECT 388.950 511.950 391.050 514.050 ;
        RECT 389.400 472.050 390.450 511.950 ;
        RECT 392.400 495.600 393.450 521.400 ;
        RECT 392.400 493.350 393.600 495.600 ;
        RECT 392.400 490.950 394.500 493.050 ;
        RECT 397.800 490.950 399.900 493.050 ;
        RECT 398.400 488.400 399.600 490.650 ;
        RECT 398.400 481.050 399.450 488.400 ;
        RECT 397.950 478.950 400.050 481.050 ;
        RECT 401.400 475.050 402.450 527.400 ;
        RECT 419.400 526.350 420.600 528.600 ;
        RECT 403.950 523.950 406.050 526.050 ;
        RECT 413.400 523.950 415.500 526.050 ;
        RECT 418.800 523.950 420.900 526.050 ;
        RECT 404.400 502.050 405.450 523.950 ;
        RECT 413.400 521.400 414.600 523.650 ;
        RECT 413.400 514.050 414.450 521.400 ;
        RECT 418.950 517.950 421.050 520.050 ;
        RECT 415.950 514.950 418.050 517.050 ;
        RECT 412.950 511.950 415.050 514.050 ;
        RECT 413.400 505.050 414.450 511.950 ;
        RECT 412.950 502.950 415.050 505.050 ;
        RECT 416.400 502.050 417.450 514.950 ;
        RECT 419.400 511.050 420.450 517.950 ;
        RECT 418.950 508.950 421.050 511.050 ;
        RECT 403.950 499.950 406.050 502.050 ;
        RECT 415.950 499.950 418.050 502.050 ;
        RECT 403.950 493.950 406.050 496.050 ;
        RECT 412.950 494.100 415.050 496.200 ;
        RECT 394.950 472.950 397.050 475.050 ;
        RECT 400.950 472.950 403.050 475.050 ;
        RECT 388.950 469.950 391.050 472.050 ;
        RECT 391.800 448.950 393.900 451.050 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 392.400 446.400 393.600 448.650 ;
        RECT 389.400 427.050 390.450 445.950 ;
        RECT 392.400 433.050 393.450 446.400 ;
        RECT 391.950 430.950 394.050 433.050 ;
        RECT 391.950 427.800 394.050 429.900 ;
        RECT 388.950 424.950 391.050 427.050 ;
        RECT 392.400 414.600 393.450 427.800 ;
        RECT 392.400 412.350 393.600 414.600 ;
        RECT 382.800 409.950 384.900 412.050 ;
        RECT 385.950 409.950 388.050 412.050 ;
        RECT 391.800 409.950 393.900 412.050 ;
        RECT 376.950 394.950 379.050 397.050 ;
        RECT 346.950 388.950 349.050 391.050 ;
        RECT 325.950 379.950 328.050 382.050 ;
        RECT 331.950 379.950 334.050 382.050 ;
        RECT 322.950 370.950 325.050 373.050 ;
        RECT 326.400 372.600 327.450 379.950 ;
        RECT 332.400 372.600 333.450 379.950 ;
        RECT 340.950 373.950 343.050 376.050 ;
        RECT 326.400 370.350 327.600 372.600 ;
        RECT 332.400 370.350 333.600 372.600 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 328.950 367.950 331.050 370.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 329.400 366.900 330.600 367.650 ;
        RECT 328.950 364.800 331.050 366.900 ;
        RECT 335.400 365.400 336.600 367.650 ;
        RECT 341.400 366.900 342.450 373.950 ;
        RECT 347.400 372.600 348.450 388.950 ;
        RECT 377.400 379.050 378.450 394.950 ;
        RECT 395.400 391.050 396.450 472.950 ;
        RECT 400.800 448.950 402.900 451.050 ;
        RECT 401.400 447.900 402.600 448.650 ;
        RECT 400.950 447.450 403.050 447.900 ;
        RECT 398.400 446.400 403.050 447.450 ;
        RECT 394.950 388.950 397.050 391.050 ;
        RECT 388.950 385.950 391.050 388.050 ;
        RECT 379.950 379.950 382.050 382.050 ;
        RECT 361.950 378.450 364.050 379.050 ;
        RECT 359.400 377.400 364.050 378.450 ;
        RECT 347.400 370.350 348.600 372.600 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 349.950 367.950 352.050 370.050 ;
        RECT 355.950 367.950 358.050 370.050 ;
        RECT 313.950 361.950 316.050 364.050 ;
        RECT 319.950 361.950 322.050 364.050 ;
        RECT 310.950 358.950 313.050 361.050 ;
        RECT 301.950 343.950 304.050 346.050 ;
        RECT 287.400 341.400 291.450 342.450 ;
        RECT 281.400 337.350 282.600 339.600 ;
        RECT 275.100 334.950 277.200 337.050 ;
        RECT 280.500 334.950 282.600 337.050 ;
        RECT 283.800 334.950 285.900 337.050 ;
        RECT 275.400 333.900 276.600 334.650 ;
        RECT 274.950 331.800 277.050 333.900 ;
        RECT 284.400 333.450 285.600 334.650 ;
        RECT 287.400 333.450 288.450 341.400 ;
        RECT 310.950 340.950 313.050 343.050 ;
        RECT 298.950 338.100 301.050 340.200 ;
        RECT 299.400 337.350 300.600 338.100 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 284.400 332.400 288.450 333.450 ;
        RECT 292.950 331.950 295.050 334.050 ;
        RECT 296.400 332.400 297.600 334.650 ;
        RECT 302.400 332.400 303.600 334.650 ;
        RECT 280.950 322.950 283.050 325.050 ;
        RECT 271.950 319.950 274.050 322.050 ;
        RECT 281.400 310.050 282.450 322.950 ;
        RECT 274.950 307.950 277.050 310.050 ;
        RECT 280.950 307.950 283.050 310.050 ;
        RECT 268.950 304.950 271.050 307.050 ;
        RECT 263.400 302.400 270.450 303.450 ;
        RECT 265.950 300.450 268.050 301.050 ;
        RECT 263.400 299.400 268.050 300.450 ;
        RECT 238.950 271.950 241.050 274.050 ;
        RECT 224.400 260.400 228.450 261.450 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 211.950 256.950 214.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 212.400 255.900 213.600 256.650 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 218.400 254.400 219.600 256.650 ;
        RECT 218.400 250.050 219.450 254.400 ;
        RECT 227.400 250.050 228.450 260.400 ;
        RECT 230.400 260.400 234.450 261.450 ;
        RECT 217.950 247.950 220.050 250.050 ;
        RECT 226.950 247.950 229.050 250.050 ;
        RECT 208.950 229.950 211.050 232.050 ;
        RECT 202.950 223.950 205.050 226.050 ;
        RECT 184.950 220.950 187.050 223.050 ;
        RECT 170.400 211.950 172.500 214.050 ;
        RECT 175.800 211.950 177.900 214.050 ;
        RECT 170.400 210.000 171.600 211.650 ;
        RECT 185.400 210.450 186.450 220.950 ;
        RECT 193.800 220.500 195.900 222.600 ;
        RECT 199.950 220.950 202.050 223.050 ;
        RECT 191.100 211.950 193.200 214.050 ;
        RECT 194.100 213.300 195.300 220.500 ;
        RECT 197.400 217.350 198.600 219.600 ;
        RECT 203.400 219.300 205.500 221.400 ;
        RECT 197.100 214.950 199.200 217.050 ;
        RECT 200.100 215.700 202.200 217.800 ;
        RECT 200.100 213.300 201.000 215.700 ;
        RECT 194.100 212.100 201.000 213.300 ;
        RECT 191.400 210.450 192.600 211.650 ;
        RECT 169.950 205.950 172.050 210.000 ;
        RECT 185.400 209.400 192.600 210.450 ;
        RECT 194.100 206.700 195.000 212.100 ;
        RECT 195.900 210.300 198.000 211.200 ;
        RECT 203.700 210.300 204.600 219.300 ;
        RECT 206.400 216.450 207.600 216.600 ;
        RECT 209.400 216.450 210.450 229.950 ;
        RECT 230.400 226.050 231.450 260.400 ;
        RECT 238.950 260.100 241.050 262.200 ;
        RECT 245.400 262.050 246.450 286.800 ;
        RECT 251.400 283.050 252.450 287.400 ;
        RECT 259.950 286.800 262.050 288.900 ;
        RECT 250.950 280.950 253.050 283.050 ;
        RECT 259.950 274.950 262.050 277.050 ;
        RECT 247.950 268.950 250.050 271.050 ;
        RECT 239.400 259.350 240.600 260.100 ;
        RECT 244.950 259.950 247.050 262.050 ;
        RECT 235.950 256.950 238.050 259.050 ;
        RECT 238.950 256.950 241.050 259.050 ;
        RECT 241.950 256.950 244.050 259.050 ;
        RECT 236.400 256.050 237.600 256.650 ;
        RECT 232.950 254.400 237.600 256.050 ;
        RECT 242.400 255.000 243.600 256.650 ;
        RECT 232.950 253.950 237.000 254.400 ;
        RECT 241.950 250.950 244.050 255.000 ;
        RECT 244.950 253.950 247.050 256.050 ;
        RECT 235.950 247.950 238.050 250.050 ;
        RECT 214.950 223.950 217.050 226.050 ;
        RECT 229.950 223.950 232.050 226.050 ;
        RECT 206.400 215.400 210.450 216.450 ;
        RECT 206.400 214.350 207.600 215.400 ;
        RECT 205.800 211.950 207.900 214.050 ;
        RECT 195.900 209.100 204.600 210.300 ;
        RECT 193.800 204.600 195.900 206.700 ;
        RECT 197.100 206.100 199.200 208.200 ;
        RECT 201.000 207.300 203.100 209.100 ;
        RECT 197.400 203.550 198.600 205.800 ;
        RECT 181.950 196.950 184.050 199.050 ;
        RECT 187.950 196.950 190.050 199.050 ;
        RECT 157.950 193.950 160.050 196.050 ;
        RECT 154.950 190.950 157.050 193.050 ;
        RECT 169.950 190.950 172.050 193.050 ;
        RECT 148.950 184.950 151.050 187.050 ;
        RECT 134.400 181.350 135.600 183.600 ;
        RECT 139.950 182.100 142.050 184.200 ;
        RECT 140.400 181.350 141.600 182.100 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 106.950 172.950 109.050 175.050 ;
        RECT 100.950 169.950 103.050 172.050 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 92.400 130.050 93.450 137.100 ;
        RECT 98.400 136.350 99.600 138.600 ;
        RECT 103.950 137.100 106.050 139.200 ;
        RECT 110.400 139.050 111.450 166.950 ;
        RECT 104.400 136.350 105.600 137.100 ;
        RECT 109.950 136.950 112.050 139.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 101.400 131.400 102.600 133.650 ;
        RECT 107.400 132.900 108.600 133.650 ;
        RECT 113.400 133.050 114.450 175.950 ;
        RECT 116.400 172.050 117.450 176.400 ;
        RECT 127.950 175.950 130.050 178.050 ;
        RECT 137.400 177.000 138.600 178.650 ;
        RECT 143.400 177.900 144.600 178.650 ;
        RECT 136.950 172.950 139.050 177.000 ;
        RECT 142.950 175.800 145.050 177.900 ;
        RECT 149.400 175.050 150.450 184.950 ;
        RECT 155.400 183.600 156.450 190.950 ;
        RECT 170.400 187.050 171.450 190.950 ;
        RECT 169.800 184.950 171.900 187.050 ;
        RECT 155.400 181.350 156.600 183.600 ;
        RECT 160.950 182.100 163.050 184.200 ;
        RECT 161.400 181.350 162.600 182.100 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 160.950 178.950 163.050 181.050 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 158.400 177.900 159.600 178.650 ;
        RECT 157.950 175.800 160.050 177.900 ;
        RECT 164.400 177.000 165.600 178.650 ;
        RECT 148.950 172.950 151.050 175.050 ;
        RECT 115.950 169.950 118.050 172.050 ;
        RECT 136.950 154.950 139.050 157.050 ;
        RECT 115.950 137.100 118.050 139.200 ;
        RECT 124.950 137.100 127.050 139.200 ;
        RECT 130.950 138.000 133.050 142.050 ;
        RECT 91.950 127.950 94.050 130.050 ;
        RECT 101.400 129.450 102.450 131.400 ;
        RECT 106.950 130.800 109.050 132.900 ;
        RECT 112.950 130.950 115.050 133.050 ;
        RECT 98.400 128.400 102.450 129.450 ;
        RECT 98.400 105.600 99.450 128.400 ;
        RECT 109.950 121.950 112.050 124.050 ;
        RECT 98.400 103.350 99.600 105.600 ;
        RECT 103.950 104.100 106.050 106.200 ;
        RECT 104.400 103.350 105.600 104.100 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 103.950 100.950 106.050 103.050 ;
        RECT 95.400 99.900 96.600 100.650 ;
        RECT 86.400 98.400 90.450 99.450 ;
        RECT 58.950 91.950 61.050 94.050 ;
        RECT 67.950 91.950 70.050 94.050 ;
        RECT 86.400 70.050 87.450 98.400 ;
        RECT 94.950 97.800 97.050 99.900 ;
        RECT 101.400 98.400 102.600 100.650 ;
        RECT 88.950 94.950 91.050 97.050 ;
        RECT 85.950 67.950 88.050 70.050 ;
        RECT 85.950 64.800 88.050 66.900 ;
        RECT 43.950 61.950 46.050 64.050 ;
        RECT 46.950 61.950 49.050 64.050 ;
        RECT 49.950 61.950 52.050 64.050 ;
        RECT 32.400 58.350 33.600 58.950 ;
        RECT 38.400 58.350 39.600 60.600 ;
        RECT 28.950 55.950 31.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 16.950 52.800 19.050 54.900 ;
        RECT 22.950 52.950 25.050 55.050 ;
        RECT 29.400 54.900 30.600 55.650 ;
        RECT 28.950 52.800 31.050 54.900 ;
        RECT 35.400 53.400 36.600 55.650 ;
        RECT 35.400 34.050 36.450 53.400 ;
        RECT 34.950 31.950 37.050 34.050 ;
        RECT 44.400 28.200 45.450 61.950 ;
        RECT 48.000 60.900 51.000 61.050 ;
        RECT 46.950 60.600 51.000 60.900 ;
        RECT 46.950 58.950 51.600 60.600 ;
        RECT 55.950 60.000 58.050 64.050 ;
        RECT 64.950 61.950 67.050 64.050 ;
        RECT 46.950 58.800 49.050 58.950 ;
        RECT 50.400 58.350 51.600 58.950 ;
        RECT 56.400 58.350 57.600 60.000 ;
        RECT 49.950 55.950 52.050 58.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 53.400 53.400 54.600 55.650 ;
        RECT 59.400 54.900 60.600 55.650 ;
        RECT 53.400 49.050 54.450 53.400 ;
        RECT 58.950 52.800 61.050 54.900 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 52.950 46.950 55.050 49.050 ;
        RECT 4.950 26.100 7.050 28.200 ;
        RECT 13.950 26.100 16.050 28.200 ;
        RECT 37.950 26.100 40.050 28.200 ;
        RECT 43.950 26.100 46.050 28.200 ;
        RECT 55.950 26.100 58.050 28.200 ;
        RECT 14.400 25.350 15.600 26.100 ;
        RECT 38.400 25.350 39.600 26.100 ;
        RECT 56.400 25.350 57.600 26.100 ;
        RECT 14.400 22.950 16.500 25.050 ;
        RECT 19.800 22.950 21.900 25.050 ;
        RECT 32.100 22.950 34.200 25.050 ;
        RECT 37.500 22.950 39.600 25.050 ;
        RECT 50.100 22.950 52.200 25.050 ;
        RECT 55.500 22.950 57.600 25.050 ;
        RECT 62.400 22.050 63.450 52.950 ;
        RECT 65.400 28.200 66.450 61.950 ;
        RECT 67.950 58.950 70.050 61.050 ;
        RECT 76.950 59.100 79.050 61.200 ;
        RECT 68.400 54.900 69.450 58.950 ;
        RECT 77.400 58.350 78.600 59.100 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 74.400 54.900 75.600 55.650 ;
        RECT 67.950 52.800 70.050 54.900 ;
        RECT 73.950 52.800 76.050 54.900 ;
        RECT 80.400 53.400 81.600 55.650 ;
        RECT 86.400 54.900 87.450 64.800 ;
        RECT 89.400 61.050 90.450 94.950 ;
        RECT 101.400 88.050 102.450 98.400 ;
        RECT 110.400 94.050 111.450 121.950 ;
        RECT 116.400 106.050 117.450 137.100 ;
        RECT 125.400 136.350 126.600 137.100 ;
        RECT 131.400 136.350 132.600 138.000 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 118.950 130.950 121.050 133.050 ;
        RECT 122.400 131.400 123.600 133.650 ;
        RECT 128.400 132.000 129.600 133.650 ;
        RECT 119.400 118.050 120.450 130.950 ;
        RECT 122.400 127.050 123.450 131.400 ;
        RECT 127.950 127.950 130.050 132.000 ;
        RECT 121.950 124.950 124.050 127.050 ;
        RECT 118.950 115.950 121.050 118.050 ;
        RECT 115.950 103.950 118.050 106.050 ;
        RECT 121.950 104.100 124.050 106.200 ;
        RECT 137.400 106.050 138.450 154.950 ;
        RECT 145.950 137.100 148.050 139.200 ;
        RECT 151.950 137.100 154.050 139.200 ;
        RECT 146.400 136.350 147.600 137.100 ;
        RECT 152.400 136.350 153.600 137.100 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 139.950 130.950 142.050 133.050 ;
        RECT 143.400 131.400 144.600 133.650 ;
        RECT 149.400 132.000 150.600 133.650 ;
        RECT 140.400 124.050 141.450 130.950 ;
        RECT 139.950 121.950 142.050 124.050 ;
        RECT 143.400 118.050 144.450 131.400 ;
        RECT 148.950 127.950 151.050 132.000 ;
        RECT 158.400 127.050 159.450 175.800 ;
        RECT 163.950 172.950 166.050 177.000 ;
        RECT 170.400 175.050 171.450 184.950 ;
        RECT 182.400 183.600 183.450 196.950 ;
        RECT 182.400 181.350 183.600 183.600 ;
        RECT 178.950 178.950 181.050 181.050 ;
        RECT 181.950 178.950 184.050 181.050 ;
        RECT 179.400 177.000 180.600 178.650 ;
        RECT 169.950 172.950 172.050 175.050 ;
        RECT 178.950 172.950 181.050 177.000 ;
        RECT 163.950 166.950 166.050 169.050 ;
        RECT 160.950 148.950 163.050 151.050 ;
        RECT 161.400 130.050 162.450 148.950 ;
        RECT 164.400 132.450 165.450 166.950 ;
        RECT 169.800 142.500 171.900 144.600 ;
        RECT 167.100 133.950 169.200 136.050 ;
        RECT 170.100 135.300 171.300 142.500 ;
        RECT 173.400 139.350 174.600 141.600 ;
        RECT 179.400 141.300 181.500 143.400 ;
        RECT 173.100 136.950 175.200 139.050 ;
        RECT 176.100 137.700 178.200 139.800 ;
        RECT 176.100 135.300 177.000 137.700 ;
        RECT 170.100 134.100 177.000 135.300 ;
        RECT 167.400 132.450 168.600 133.650 ;
        RECT 164.400 131.400 168.600 132.450 ;
        RECT 160.950 127.950 163.050 130.050 ;
        RECT 170.100 128.700 171.000 134.100 ;
        RECT 171.900 132.300 174.000 133.200 ;
        RECT 179.700 132.300 180.600 141.300 ;
        RECT 188.400 139.200 189.450 196.950 ;
        RECT 197.400 193.050 198.450 203.550 ;
        RECT 209.400 202.050 210.450 215.400 ;
        RECT 215.400 210.450 216.450 223.950 ;
        RECT 221.100 220.500 223.200 222.600 ;
        RECT 218.100 211.950 220.200 214.050 ;
        RECT 221.100 213.900 222.000 220.500 ;
        RECT 230.100 220.200 232.200 222.300 ;
        RECT 224.400 217.350 225.600 219.600 ;
        RECT 223.800 214.950 225.900 217.050 ;
        RECT 228.000 213.900 230.100 214.200 ;
        RECT 221.100 213.000 230.100 213.900 ;
        RECT 218.400 210.450 219.600 211.650 ;
        RECT 215.400 209.400 219.600 210.450 ;
        RECT 208.950 199.950 211.050 202.050 ;
        RECT 196.950 190.950 199.050 193.050 ;
        RECT 215.400 190.050 216.450 209.400 ;
        RECT 221.100 207.900 222.000 213.000 ;
        RECT 228.000 212.100 230.100 213.000 ;
        RECT 222.900 211.200 225.000 212.100 ;
        RECT 222.900 210.000 230.100 211.200 ;
        RECT 228.000 209.100 230.100 210.000 ;
        RECT 220.500 205.800 222.600 207.900 ;
        RECT 223.800 206.100 225.900 208.200 ;
        RECT 231.000 207.600 231.900 220.200 ;
        RECT 232.950 215.100 235.050 217.200 ;
        RECT 233.400 214.350 234.600 215.100 ;
        RECT 232.800 211.950 234.900 214.050 ;
        RECT 236.400 208.050 237.450 247.950 ;
        RECT 241.950 223.950 244.050 226.050 ;
        RECT 238.950 217.950 241.050 220.050 ;
        RECT 224.400 203.550 225.600 205.800 ;
        RECT 230.400 205.500 232.500 207.600 ;
        RECT 235.950 205.950 238.050 208.050 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 205.950 187.950 208.050 190.050 ;
        RECT 214.950 187.950 217.050 190.050 ;
        RECT 196.950 182.100 199.050 184.200 ;
        RECT 197.400 181.350 198.600 182.100 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 194.400 177.000 195.600 178.650 ;
        RECT 193.950 172.950 196.050 177.000 ;
        RECT 200.400 176.400 201.600 178.650 ;
        RECT 200.400 169.050 201.450 176.400 ;
        RECT 206.400 175.050 207.450 187.950 ;
        RECT 208.950 181.950 211.050 184.050 ;
        RECT 218.400 183.600 219.450 199.950 ;
        RECT 224.400 199.050 225.450 203.550 ;
        RECT 223.950 196.950 226.050 199.050 ;
        RECT 223.950 187.950 226.050 190.050 ;
        RECT 224.400 183.600 225.450 187.950 ;
        RECT 209.400 177.900 210.450 181.950 ;
        RECT 218.400 181.350 219.600 183.600 ;
        RECT 224.400 181.350 225.600 183.600 ;
        RECT 229.950 181.950 232.050 184.050 ;
        RECT 236.400 183.600 237.450 205.950 ;
        RECT 239.400 186.450 240.450 217.950 ;
        RECT 242.400 217.200 243.450 223.950 ;
        RECT 245.400 220.050 246.450 253.950 ;
        RECT 248.400 253.050 249.450 268.950 ;
        RECT 260.400 264.450 261.450 274.950 ;
        RECT 263.400 271.050 264.450 299.400 ;
        RECT 265.950 298.950 268.050 299.400 ;
        RECT 266.400 294.600 267.450 298.950 ;
        RECT 269.400 298.050 270.450 302.400 ;
        RECT 268.950 295.950 271.050 298.050 ;
        RECT 275.400 294.600 276.450 307.950 ;
        RECT 266.400 292.350 267.600 294.600 ;
        RECT 275.400 294.450 276.600 294.600 ;
        RECT 275.400 293.400 279.450 294.450 ;
        RECT 275.400 292.350 276.600 293.400 ;
        RECT 266.100 289.950 268.200 292.050 ;
        RECT 271.500 289.950 273.600 292.050 ;
        RECT 274.800 289.950 276.900 292.050 ;
        RECT 272.400 288.900 273.600 289.650 ;
        RECT 271.950 286.800 274.050 288.900 ;
        RECT 268.950 283.950 271.050 286.050 ;
        RECT 262.950 268.950 265.050 271.050 ;
        RECT 260.400 263.400 264.450 264.450 ;
        RECT 256.950 260.100 259.050 262.200 ;
        RECT 263.400 261.600 264.450 263.400 ;
        RECT 257.400 259.350 258.600 260.100 ;
        RECT 263.400 259.350 264.600 261.600 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 259.950 256.950 262.050 259.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 250.950 253.950 253.050 256.050 ;
        RECT 254.400 255.000 255.600 256.650 ;
        RECT 260.400 255.900 261.600 256.650 ;
        RECT 269.400 255.900 270.450 283.950 ;
        RECT 278.400 283.050 279.450 293.400 ;
        RECT 277.950 280.950 280.050 283.050 ;
        RECT 281.400 268.050 282.450 307.950 ;
        RECT 293.400 307.050 294.450 331.950 ;
        RECT 296.400 328.050 297.450 332.400 ;
        RECT 298.950 328.950 301.050 331.050 ;
        RECT 295.950 325.950 298.050 328.050 ;
        RECT 296.400 316.050 297.450 325.950 ;
        RECT 299.400 322.050 300.450 328.950 ;
        RECT 302.400 325.050 303.450 332.400 ;
        RECT 301.950 322.950 304.050 325.050 ;
        RECT 298.950 319.950 301.050 322.050 ;
        RECT 303.000 321.450 307.050 322.050 ;
        RECT 302.400 319.950 307.050 321.450 ;
        RECT 295.950 313.950 298.050 316.050 ;
        RECT 302.400 313.050 303.450 319.950 ;
        RECT 304.950 316.800 307.050 318.900 ;
        RECT 301.950 310.950 304.050 313.050 ;
        RECT 286.950 304.950 289.050 307.050 ;
        RECT 292.950 304.950 295.050 307.050 ;
        RECT 301.950 304.950 304.050 307.050 ;
        RECT 283.950 301.950 286.050 304.050 ;
        RECT 284.400 288.900 285.450 301.950 ;
        RECT 287.400 295.050 288.450 304.950 ;
        RECT 293.400 298.050 294.450 304.950 ;
        RECT 302.400 298.050 303.450 304.950 ;
        RECT 305.400 301.050 306.450 316.800 ;
        RECT 308.400 307.050 309.450 337.950 ;
        RECT 311.400 310.050 312.450 340.950 ;
        RECT 314.400 340.050 315.450 361.950 ;
        RECT 316.950 358.950 319.050 361.050 ;
        RECT 317.400 343.050 318.450 358.950 ;
        RECT 325.950 352.950 328.050 355.050 ;
        RECT 316.950 340.950 319.050 343.050 ;
        RECT 313.950 337.950 316.050 340.050 ;
        RECT 319.950 338.100 322.050 340.200 ;
        RECT 326.400 340.050 327.450 352.950 ;
        RECT 335.400 352.050 336.450 365.400 ;
        RECT 340.950 364.800 343.050 366.900 ;
        RECT 350.400 365.400 351.600 367.650 ;
        RECT 350.400 361.050 351.450 365.400 ;
        RECT 349.950 358.950 352.050 361.050 ;
        RECT 340.950 352.950 343.050 355.050 ;
        RECT 334.950 349.950 337.050 352.050 ;
        RECT 320.400 337.350 321.600 338.100 ;
        RECT 325.950 337.950 328.050 340.050 ;
        RECT 331.950 337.950 334.050 340.050 ;
        RECT 341.400 339.600 342.450 352.950 ;
        RECT 352.950 349.950 355.050 352.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 322.950 334.950 325.050 337.050 ;
        RECT 313.950 331.950 316.050 334.050 ;
        RECT 317.400 333.000 318.600 334.650 ;
        RECT 323.400 333.900 324.600 334.650 ;
        RECT 310.950 307.950 313.050 310.050 ;
        RECT 307.950 304.950 310.050 307.050 ;
        RECT 304.950 298.950 307.050 301.050 ;
        RECT 292.950 295.950 295.050 298.050 ;
        RECT 301.950 295.950 304.050 298.050 ;
        RECT 286.950 292.950 289.050 295.050 ;
        RECT 293.400 294.600 294.450 295.950 ;
        RECT 293.400 292.350 294.600 294.600 ;
        RECT 298.950 293.100 301.050 295.200 ;
        RECT 299.400 292.350 300.600 293.100 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 298.950 289.950 301.050 292.050 ;
        RECT 283.950 286.800 286.050 288.900 ;
        RECT 286.950 286.950 289.050 289.050 ;
        RECT 290.400 287.400 291.600 289.650 ;
        RECT 296.400 287.400 297.600 289.650 ;
        RECT 274.950 265.950 277.050 268.050 ;
        RECT 280.950 265.950 283.050 268.050 ;
        RECT 271.950 259.950 274.050 265.050 ;
        RECT 275.400 261.600 276.450 265.950 ;
        RECT 275.400 259.350 276.600 261.600 ;
        RECT 280.950 260.100 283.050 262.200 ;
        RECT 287.400 262.050 288.450 286.950 ;
        RECT 290.400 277.050 291.450 287.400 ;
        RECT 296.400 283.050 297.450 287.400 ;
        RECT 301.950 286.950 304.050 289.050 ;
        RECT 295.950 280.950 298.050 283.050 ;
        RECT 289.950 274.950 292.050 277.050 ;
        RECT 302.400 265.050 303.450 286.950 ;
        RECT 289.950 262.950 292.050 265.050 ;
        RECT 281.400 259.350 282.600 260.100 ;
        RECT 286.950 259.950 289.050 262.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 247.950 250.950 250.050 253.050 ;
        RECT 248.400 223.050 249.450 250.950 ;
        RECT 247.950 220.950 250.050 223.050 ;
        RECT 244.950 217.950 247.050 220.050 ;
        RECT 241.950 216.450 244.050 217.200 ;
        RECT 251.400 216.600 252.450 253.950 ;
        RECT 253.950 250.950 256.050 255.000 ;
        RECT 259.950 253.800 262.050 255.900 ;
        RECT 268.950 253.800 271.050 255.900 ;
        RECT 271.950 253.950 274.050 256.050 ;
        RECT 278.400 255.900 279.600 256.650 ;
        RECT 256.950 229.950 259.050 232.050 ;
        RECT 245.400 216.450 246.600 216.600 ;
        RECT 241.950 215.400 246.600 216.450 ;
        RECT 241.950 215.100 244.050 215.400 ;
        RECT 245.400 214.350 246.600 215.400 ;
        RECT 251.400 214.350 252.600 216.600 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 241.950 208.950 244.050 211.050 ;
        RECT 248.400 209.400 249.600 211.650 ;
        RECT 242.400 190.050 243.450 208.950 ;
        RECT 248.400 204.450 249.450 209.400 ;
        RECT 245.400 203.400 249.450 204.450 ;
        RECT 241.950 187.950 244.050 190.050 ;
        RECT 239.400 185.400 243.450 186.450 ;
        RECT 242.400 183.600 243.450 185.400 ;
        RECT 245.400 184.050 246.450 203.400 ;
        RECT 247.950 199.950 250.050 202.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 215.400 177.900 216.600 178.650 ;
        RECT 208.950 175.800 211.050 177.900 ;
        RECT 214.950 175.800 217.050 177.900 ;
        RECT 221.400 177.000 222.600 178.650 ;
        RECT 205.950 172.950 208.050 175.050 ;
        RECT 220.950 172.950 223.050 177.000 ;
        RECT 199.950 166.950 202.050 169.050 ;
        RECT 230.400 157.050 231.450 181.950 ;
        RECT 236.400 181.350 237.600 183.600 ;
        RECT 242.400 181.350 243.600 183.600 ;
        RECT 244.950 181.950 247.050 184.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 239.400 177.900 240.600 178.650 ;
        RECT 238.950 175.800 241.050 177.900 ;
        RECT 229.950 154.950 232.050 157.050 ;
        RECT 199.950 145.950 202.050 148.050 ;
        RECT 208.950 145.950 211.050 148.050 ;
        RECT 193.950 142.950 196.050 145.050 ;
        RECT 181.950 137.100 184.050 139.200 ;
        RECT 187.950 137.100 190.050 139.200 ;
        RECT 194.400 138.600 195.450 142.950 ;
        RECT 200.400 138.600 201.450 145.950 ;
        RECT 182.400 136.350 183.600 137.100 ;
        RECT 194.400 136.350 195.600 138.600 ;
        RECT 200.400 136.350 201.600 138.600 ;
        RECT 181.800 133.950 183.900 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 171.900 131.100 180.600 132.300 ;
        RECT 197.400 131.400 198.600 133.650 ;
        RECT 203.400 131.400 204.600 133.650 ;
        RECT 209.400 132.900 210.450 145.950 ;
        RECT 217.950 137.100 220.050 139.200 ;
        RECT 235.950 137.100 238.050 139.200 ;
        RECT 241.950 137.100 244.050 139.200 ;
        RECT 218.400 136.350 219.600 137.100 ;
        RECT 236.400 136.350 237.600 137.100 ;
        RECT 242.400 136.350 243.600 137.100 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 232.950 133.950 235.050 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 215.400 132.900 216.600 133.650 ;
        RECT 157.950 124.950 160.050 127.050 ;
        RECT 169.800 126.600 171.900 128.700 ;
        RECT 173.100 128.100 175.200 130.200 ;
        RECT 177.000 129.300 179.100 131.100 ;
        RECT 173.400 125.550 174.600 127.800 ;
        RECT 148.950 121.950 151.050 124.050 ;
        RECT 142.950 115.950 145.050 118.050 ;
        RECT 149.400 112.050 150.450 121.950 ;
        RECT 173.400 121.050 174.450 125.550 ;
        RECT 175.950 124.950 178.050 127.050 ;
        RECT 172.950 118.950 175.050 121.050 ;
        RECT 142.950 109.950 145.050 112.050 ;
        RECT 148.950 109.950 151.050 112.050 ;
        RECT 122.400 103.350 123.600 104.100 ;
        RECT 130.950 103.950 133.050 106.050 ;
        RECT 136.950 103.950 139.050 106.050 ;
        RECT 143.400 105.600 144.450 109.950 ;
        RECT 149.400 105.600 150.450 109.950 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 121.950 100.950 124.050 103.050 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 119.400 99.000 120.600 100.650 ;
        RECT 125.400 99.000 126.600 100.650 ;
        RECT 118.950 94.950 121.050 99.000 ;
        RECT 124.950 94.950 127.050 99.000 ;
        RECT 109.950 91.950 112.050 94.050 ;
        RECT 100.950 85.950 103.050 88.050 ;
        RECT 100.950 67.950 103.050 70.050 ;
        RECT 127.950 67.950 130.050 70.050 ;
        RECT 88.950 58.950 91.050 61.050 ;
        RECT 94.950 59.100 97.050 61.200 ;
        RECT 101.400 60.600 102.450 67.950 ;
        RECT 106.950 61.950 109.050 64.050 ;
        RECT 115.950 63.450 118.050 64.200 ;
        RECT 115.950 62.400 123.450 63.450 ;
        RECT 115.950 62.100 118.050 62.400 ;
        RECT 95.400 58.350 96.600 59.100 ;
        RECT 101.400 58.350 102.600 60.600 ;
        RECT 91.950 55.950 94.050 58.050 ;
        RECT 94.950 55.950 97.050 58.050 ;
        RECT 97.950 55.950 100.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 73.950 31.950 76.050 34.050 ;
        RECT 74.400 28.200 75.450 31.950 ;
        RECT 64.950 26.100 67.050 28.200 ;
        RECT 73.950 26.100 76.050 28.200 ;
        RECT 74.400 25.350 75.600 26.100 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 61.950 19.950 64.050 22.050 ;
        RECT 71.400 21.900 72.600 22.650 ;
        RECT 80.400 22.050 81.450 53.400 ;
        RECT 85.950 52.800 88.050 54.900 ;
        RECT 88.950 52.950 91.050 55.050 ;
        RECT 92.400 54.900 93.600 55.650 ;
        RECT 70.950 19.800 73.050 21.900 ;
        RECT 79.950 19.950 82.050 22.050 ;
        RECT 86.400 16.050 87.450 52.800 ;
        RECT 89.400 27.600 90.450 52.950 ;
        RECT 91.950 52.800 94.050 54.900 ;
        RECT 98.400 53.400 99.600 55.650 ;
        RECT 98.400 34.050 99.450 53.400 ;
        RECT 107.400 34.050 108.450 61.950 ;
        RECT 109.950 58.950 112.050 61.050 ;
        RECT 115.950 58.950 118.050 61.050 ;
        RECT 122.400 60.600 123.450 62.400 ;
        RECT 110.400 49.050 111.450 58.950 ;
        RECT 116.400 58.350 117.600 58.950 ;
        RECT 122.400 58.350 123.600 60.600 ;
        RECT 115.950 55.950 118.050 58.050 ;
        RECT 118.950 55.950 121.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 119.400 54.900 120.600 55.650 ;
        RECT 118.950 52.800 121.050 54.900 ;
        RECT 109.950 46.950 112.050 49.050 ;
        RECT 128.400 40.050 129.450 67.950 ;
        RECT 131.400 67.050 132.450 103.950 ;
        RECT 143.400 103.350 144.600 105.600 ;
        RECT 149.400 103.350 150.600 105.600 ;
        RECT 154.950 104.100 157.050 106.200 ;
        RECT 163.950 104.100 166.050 106.200 ;
        RECT 169.950 104.100 172.050 106.200 ;
        RECT 176.400 106.050 177.450 124.950 ;
        RECT 178.950 115.950 181.050 118.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 140.400 99.000 141.600 100.650 ;
        RECT 139.950 94.950 142.050 99.000 ;
        RECT 146.400 98.400 147.600 100.650 ;
        RECT 146.400 97.050 147.450 98.400 ;
        RECT 155.400 97.050 156.450 104.100 ;
        RECT 164.400 103.350 165.600 104.100 ;
        RECT 170.400 103.350 171.600 104.100 ;
        RECT 175.950 103.950 178.050 106.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 161.400 98.400 162.600 100.650 ;
        RECT 167.400 98.400 168.600 100.650 ;
        RECT 173.400 99.900 174.600 100.650 ;
        RECT 179.400 99.900 180.450 115.950 ;
        RECT 184.950 109.950 187.050 112.050 ;
        RECT 193.950 109.950 196.050 112.050 ;
        RECT 185.400 105.600 186.450 109.950 ;
        RECT 185.400 103.350 186.600 105.600 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 188.400 99.900 189.600 100.650 ;
        RECT 194.400 100.050 195.450 109.950 ;
        RECT 145.950 94.950 148.050 97.050 ;
        RECT 154.950 94.950 157.050 97.050 ;
        RECT 146.400 91.050 147.450 94.950 ;
        RECT 161.400 91.050 162.450 98.400 ;
        RECT 167.400 94.050 168.450 98.400 ;
        RECT 172.950 97.800 175.050 99.900 ;
        RECT 178.950 97.800 181.050 99.900 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 193.950 97.950 196.050 100.050 ;
        RECT 166.950 91.950 169.050 94.050 ;
        RECT 145.950 88.950 148.050 91.050 ;
        RECT 151.950 88.950 154.050 91.050 ;
        RECT 160.950 88.950 163.050 91.050 ;
        RECT 148.950 73.950 151.050 76.050 ;
        RECT 130.950 64.950 133.050 67.050 ;
        RECT 136.950 59.100 139.050 61.200 ;
        RECT 142.950 59.100 145.050 61.200 ;
        RECT 137.400 58.350 138.600 59.100 ;
        RECT 143.400 58.350 144.600 59.100 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 134.400 54.000 135.600 55.650 ;
        RECT 133.950 49.950 136.050 54.000 ;
        RECT 140.400 53.400 141.600 55.650 ;
        RECT 140.400 43.050 141.450 53.400 ;
        RECT 139.950 40.950 142.050 43.050 ;
        RECT 127.950 37.950 130.050 40.050 ;
        RECT 97.950 31.950 100.050 34.050 ;
        RECT 106.950 31.950 109.050 34.050 ;
        RECT 118.950 31.950 121.050 34.050 ;
        RECT 89.400 25.350 90.600 27.600 ;
        RECT 109.950 26.100 112.050 28.200 ;
        RECT 110.400 25.350 111.600 26.100 ;
        RECT 89.400 22.950 91.500 25.050 ;
        RECT 94.800 22.950 96.900 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 107.400 21.900 108.600 22.650 ;
        RECT 106.950 19.800 109.050 21.900 ;
        RECT 113.400 20.400 114.600 22.650 ;
        RECT 119.400 21.900 120.450 31.950 ;
        RECT 124.950 27.000 127.050 31.050 ;
        RECT 149.400 30.450 150.450 73.950 ;
        RECT 152.400 52.050 153.450 88.950 ;
        RECT 197.400 76.050 198.450 131.400 ;
        RECT 199.950 124.950 202.050 127.050 ;
        RECT 200.400 106.050 201.450 124.950 ;
        RECT 203.400 124.050 204.450 131.400 ;
        RECT 208.950 130.800 211.050 132.900 ;
        RECT 214.950 130.800 217.050 132.900 ;
        RECT 229.950 130.950 232.050 133.050 ;
        RECT 233.400 131.400 234.600 133.650 ;
        RECT 239.400 132.900 240.600 133.650 ;
        RECT 202.950 121.950 205.050 124.050 ;
        RECT 217.950 115.950 220.050 118.050 ;
        RECT 208.950 109.950 211.050 112.050 ;
        RECT 199.950 103.950 202.050 106.050 ;
        RECT 202.950 104.100 205.050 106.200 ;
        RECT 209.400 105.600 210.450 109.950 ;
        RECT 203.400 103.350 204.600 104.100 ;
        RECT 209.400 103.350 210.600 105.600 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 199.950 97.950 202.050 100.050 ;
        RECT 206.400 99.000 207.600 100.650 ;
        RECT 212.400 99.900 213.600 100.650 ;
        RECT 218.400 99.900 219.450 115.950 ;
        RECT 230.400 112.050 231.450 130.950 ;
        RECT 233.400 127.050 234.450 131.400 ;
        RECT 238.950 130.800 241.050 132.900 ;
        RECT 232.950 124.950 235.050 127.050 ;
        RECT 235.950 112.950 238.050 115.050 ;
        RECT 229.950 109.950 232.050 112.050 ;
        RECT 226.950 104.100 229.050 106.200 ;
        RECT 227.400 103.350 228.600 104.100 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 224.400 99.900 225.600 100.650 ;
        RECT 196.950 73.950 199.050 76.050 ;
        RECT 200.400 66.450 201.450 97.950 ;
        RECT 205.950 94.950 208.050 99.000 ;
        RECT 211.950 97.800 214.050 99.900 ;
        RECT 212.400 79.050 213.450 97.800 ;
        RECT 217.950 94.950 220.050 99.900 ;
        RECT 223.950 97.800 226.050 99.900 ;
        RECT 230.400 98.400 231.600 100.650 ;
        RECT 230.400 79.050 231.450 98.400 ;
        RECT 211.950 76.950 214.050 79.050 ;
        RECT 229.950 76.950 232.050 79.050 ;
        RECT 202.950 67.950 205.050 70.050 ;
        RECT 197.400 65.400 201.450 66.450 ;
        RECT 197.400 64.050 198.450 65.400 ;
        RECT 196.950 61.950 199.050 64.050 ;
        RECT 157.950 59.100 160.050 61.200 ;
        RECT 163.950 59.100 166.050 61.200 ;
        RECT 175.950 59.100 178.050 61.200 ;
        RECT 158.400 58.350 159.600 59.100 ;
        RECT 164.400 58.350 165.600 59.100 ;
        RECT 176.400 58.350 177.600 59.100 ;
        RECT 184.950 58.950 187.050 61.050 ;
        RECT 197.400 60.600 198.450 61.950 ;
        RECT 203.400 60.600 204.450 67.950 ;
        RECT 223.950 64.950 226.050 67.050 ;
        RECT 211.950 61.950 214.050 64.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 154.950 52.950 157.050 55.050 ;
        RECT 161.400 53.400 162.600 55.650 ;
        RECT 151.950 49.950 154.050 52.050 ;
        RECT 155.400 49.050 156.450 52.950 ;
        RECT 154.950 46.950 157.050 49.050 ;
        RECT 161.400 40.050 162.450 53.400 ;
        RECT 166.950 52.950 169.050 55.050 ;
        RECT 179.400 54.900 180.600 55.650 ;
        RECT 167.400 43.050 168.450 52.950 ;
        RECT 178.950 52.800 181.050 54.900 ;
        RECT 181.950 46.950 184.050 49.050 ;
        RECT 166.950 40.950 169.050 43.050 ;
        RECT 160.950 37.950 163.050 40.050 ;
        RECT 154.950 31.950 157.050 34.050 ;
        RECT 163.950 31.950 166.050 34.050 ;
        RECT 146.400 29.400 150.450 30.450 ;
        RECT 125.400 25.350 126.600 27.000 ;
        RECT 130.950 26.100 133.050 28.200 ;
        RECT 131.400 25.350 132.600 26.100 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 113.400 16.050 114.450 20.400 ;
        RECT 118.950 19.800 121.050 21.900 ;
        RECT 128.400 20.400 129.600 22.650 ;
        RECT 134.400 21.000 135.600 22.650 ;
        RECT 128.400 16.050 129.450 20.400 ;
        RECT 133.950 16.950 136.050 21.000 ;
        RECT 146.400 19.050 147.450 29.400 ;
        RECT 155.400 27.600 156.450 31.950 ;
        RECT 155.400 25.350 156.600 27.600 ;
        RECT 149.100 22.950 151.200 25.050 ;
        RECT 154.500 22.950 156.600 25.050 ;
        RECT 157.800 22.950 159.900 25.050 ;
        RECT 149.400 20.400 150.600 22.650 ;
        RECT 158.400 20.400 159.600 22.650 ;
        RECT 164.400 21.900 165.450 31.950 ;
        RECT 175.950 26.100 178.050 28.200 ;
        RECT 182.400 27.600 183.450 46.950 ;
        RECT 185.400 46.050 186.450 58.950 ;
        RECT 197.400 58.350 198.600 60.600 ;
        RECT 203.400 58.350 204.600 60.600 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 194.400 54.900 195.600 55.650 ;
        RECT 200.400 54.900 201.600 55.650 ;
        RECT 212.400 54.900 213.450 61.950 ;
        RECT 217.950 60.000 220.050 64.050 ;
        RECT 224.400 60.600 225.450 64.950 ;
        RECT 236.400 64.050 237.450 112.950 ;
        RECT 244.950 109.950 247.050 112.050 ;
        RECT 238.950 103.950 241.050 106.050 ;
        RECT 245.400 105.600 246.450 109.950 ;
        RECT 248.400 109.050 249.450 199.950 ;
        RECT 257.400 190.050 258.450 229.950 ;
        RECT 272.400 223.050 273.450 253.950 ;
        RECT 277.950 253.800 280.050 255.900 ;
        RECT 284.400 254.400 285.600 256.650 ;
        RECT 284.400 238.050 285.450 254.400 ;
        RECT 277.950 235.950 280.050 238.050 ;
        RECT 283.950 235.950 286.050 238.050 ;
        RECT 265.950 220.950 268.050 223.050 ;
        RECT 271.950 220.950 274.050 223.050 ;
        RECT 266.400 216.600 267.450 220.950 ;
        RECT 266.400 214.350 267.600 216.600 ;
        RECT 271.950 216.000 274.050 219.900 ;
        RECT 278.400 217.050 279.450 235.950 ;
        RECT 290.400 232.050 291.450 262.950 ;
        RECT 298.950 261.000 301.050 265.050 ;
        RECT 301.950 262.950 304.050 265.050 ;
        RECT 305.400 262.050 306.450 298.950 ;
        RECT 314.400 298.050 315.450 331.950 ;
        RECT 316.950 325.950 319.050 333.000 ;
        RECT 322.950 331.800 325.050 333.900 ;
        RECT 321.000 327.450 325.050 328.050 ;
        RECT 320.400 325.950 325.050 327.450 ;
        RECT 328.950 325.950 331.050 328.050 ;
        RECT 320.400 324.450 321.450 325.950 ;
        RECT 317.400 323.400 321.450 324.450 ;
        RECT 317.400 316.050 318.450 323.400 ;
        RECT 325.950 319.950 328.050 325.050 ;
        RECT 325.950 316.800 328.050 318.900 ;
        RECT 316.950 313.950 319.050 316.050 ;
        RECT 326.400 310.050 327.450 316.800 ;
        RECT 329.400 316.050 330.450 325.950 ;
        RECT 332.400 325.050 333.450 337.950 ;
        RECT 341.400 337.350 342.600 339.600 ;
        RECT 346.950 338.100 349.050 340.200 ;
        RECT 353.400 340.050 354.450 349.950 ;
        RECT 347.400 337.350 348.600 338.100 ;
        RECT 352.950 337.950 355.050 340.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 338.400 333.000 339.600 334.650 ;
        RECT 337.950 328.950 340.050 333.000 ;
        RECT 344.400 332.400 345.600 334.650 ;
        RECT 350.400 333.450 351.600 334.650 ;
        RECT 350.400 332.400 354.450 333.450 ;
        RECT 331.950 322.950 334.050 325.050 ;
        RECT 334.950 319.950 340.050 322.050 ;
        RECT 328.950 313.950 331.050 316.050 ;
        RECT 322.800 307.950 324.900 310.050 ;
        RECT 325.950 307.950 328.050 310.050 ;
        RECT 340.950 307.950 343.050 310.050 ;
        RECT 310.950 294.000 313.050 298.050 ;
        RECT 313.950 295.950 316.050 298.050 ;
        RECT 311.400 292.350 312.600 294.000 ;
        RECT 316.950 293.100 319.050 295.200 ;
        RECT 323.400 295.050 324.450 307.950 ;
        RECT 325.800 301.950 327.900 304.050 ;
        RECT 328.950 301.950 331.050 304.050 ;
        RECT 317.400 292.350 318.600 293.100 ;
        RECT 322.950 292.950 325.050 295.050 ;
        RECT 326.400 292.050 327.450 301.950 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 319.950 289.950 322.050 292.050 ;
        RECT 325.950 289.950 328.050 292.050 ;
        RECT 314.400 288.900 315.600 289.650 ;
        RECT 320.400 289.050 321.600 289.650 ;
        RECT 313.950 286.800 316.050 288.900 ;
        RECT 320.400 287.400 325.050 289.050 ;
        RECT 321.000 286.950 325.050 287.400 ;
        RECT 325.950 286.800 328.050 288.900 ;
        RECT 310.950 283.950 313.050 286.050 ;
        RECT 307.950 274.950 310.050 277.050 ;
        RECT 299.400 259.350 300.600 261.000 ;
        RECT 304.950 259.950 307.050 262.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 292.950 253.950 295.050 256.050 ;
        RECT 296.400 255.900 297.600 256.650 ;
        RECT 302.400 256.050 303.600 256.650 ;
        RECT 289.950 229.950 292.050 232.050 ;
        RECT 280.950 220.950 283.050 223.050 ;
        RECT 272.400 214.350 273.600 216.000 ;
        RECT 277.950 214.950 280.050 217.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 269.400 209.400 270.600 211.650 ;
        RECT 275.400 210.000 276.600 211.650 ;
        RECT 281.400 210.900 282.450 220.950 ;
        RECT 293.400 220.050 294.450 253.950 ;
        RECT 295.950 253.800 298.050 255.900 ;
        RECT 302.400 254.400 307.050 256.050 ;
        RECT 303.000 253.950 307.050 254.400 ;
        RECT 308.400 247.050 309.450 274.950 ;
        RECT 307.950 244.950 310.050 247.050 ;
        RECT 301.950 241.950 304.050 244.050 ;
        RECT 298.950 220.950 301.050 223.050 ;
        RECT 283.950 217.950 289.050 220.050 ;
        RECT 292.950 219.450 295.050 220.050 ;
        RECT 292.950 218.400 297.450 219.450 ;
        RECT 292.950 217.950 295.050 218.400 ;
        RECT 296.400 216.600 297.450 218.400 ;
        RECT 287.400 216.450 288.600 216.600 ;
        RECT 284.400 215.400 288.600 216.450 ;
        RECT 250.950 187.950 253.050 190.050 ;
        RECT 256.950 187.950 259.050 190.050 ;
        RECT 262.950 187.950 265.050 190.050 ;
        RECT 251.400 130.050 252.450 187.950 ;
        RECT 256.950 182.100 259.050 184.200 ;
        RECT 263.400 183.600 264.450 187.950 ;
        RECT 269.400 184.050 270.450 209.400 ;
        RECT 274.950 205.950 277.050 210.000 ;
        RECT 280.950 208.800 283.050 210.900 ;
        RECT 284.400 202.050 285.450 215.400 ;
        RECT 287.400 214.350 288.600 215.400 ;
        RECT 296.400 214.350 297.600 216.600 ;
        RECT 287.100 211.950 289.200 214.050 ;
        RECT 290.400 211.950 292.500 214.050 ;
        RECT 295.800 211.950 297.900 214.050 ;
        RECT 290.400 210.900 291.600 211.650 ;
        RECT 289.950 208.800 292.050 210.900 ;
        RECT 283.950 199.950 286.050 202.050 ;
        RECT 299.400 190.050 300.450 220.950 ;
        RECT 302.400 211.050 303.450 241.950 ;
        RECT 304.950 217.950 307.050 220.050 ;
        RECT 301.950 208.950 304.050 211.050 ;
        RECT 305.400 205.050 306.450 217.950 ;
        RECT 311.400 216.600 312.450 283.950 ;
        RECT 326.400 277.050 327.450 286.800 ;
        RECT 325.950 274.950 328.050 277.050 ;
        RECT 329.400 274.050 330.450 301.950 ;
        RECT 334.950 293.100 337.050 295.200 ;
        RECT 341.400 294.600 342.450 307.950 ;
        RECT 335.400 292.350 336.600 293.100 ;
        RECT 341.400 292.350 342.600 294.600 ;
        RECT 344.400 294.450 345.450 332.400 ;
        RECT 353.400 316.050 354.450 332.400 ;
        RECT 356.400 325.050 357.450 367.950 ;
        RECT 359.400 333.900 360.450 377.400 ;
        RECT 361.950 376.950 364.050 377.400 ;
        RECT 376.950 376.950 379.050 379.050 ;
        RECT 362.400 372.600 363.450 376.950 ;
        RECT 362.400 370.350 363.600 372.600 ;
        RECT 370.950 371.100 373.050 373.200 ;
        RECT 371.400 370.350 372.600 371.100 ;
        RECT 362.100 367.950 364.200 370.050 ;
        RECT 367.500 367.950 369.600 370.050 ;
        RECT 370.800 367.950 372.900 370.050 ;
        RECT 368.400 366.900 369.600 367.650 ;
        RECT 367.950 364.800 370.050 366.900 ;
        RECT 368.400 340.200 369.450 364.800 ;
        RECT 373.950 355.950 376.050 358.050 ;
        RECT 367.950 338.100 370.050 340.200 ;
        RECT 374.400 339.600 375.450 355.950 ;
        RECT 380.400 340.050 381.450 379.950 ;
        RECT 389.400 372.600 390.450 385.950 ;
        RECT 394.950 376.950 397.050 379.050 ;
        RECT 395.400 373.200 396.450 376.950 ;
        RECT 389.400 370.350 390.600 372.600 ;
        RECT 394.800 371.100 396.900 373.200 ;
        RECT 398.400 373.050 399.450 446.400 ;
        RECT 400.950 445.800 403.050 446.400 ;
        RECT 404.400 444.450 405.450 493.950 ;
        RECT 413.400 493.350 414.600 494.100 ;
        RECT 409.950 490.950 412.050 493.050 ;
        RECT 412.950 490.950 415.050 493.050 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 410.400 489.000 411.600 490.650 ;
        RECT 409.950 484.950 412.050 489.000 ;
        RECT 416.400 488.400 417.600 490.650 ;
        RECT 416.400 481.050 417.450 488.400 ;
        RECT 415.950 478.950 418.050 481.050 ;
        RECT 422.400 469.050 423.450 529.950 ;
        RECT 428.400 520.050 429.450 542.400 ;
        RECT 433.950 541.950 436.050 544.050 ;
        RECT 436.800 535.950 438.900 538.050 ;
        RECT 439.950 535.950 442.050 538.050 ;
        RECT 437.400 528.600 438.450 535.950 ;
        RECT 440.400 532.050 441.450 535.950 ;
        RECT 439.950 529.950 442.050 532.050 ;
        RECT 437.400 526.350 438.600 528.600 ;
        RECT 442.950 527.100 445.050 529.200 ;
        RECT 443.400 526.350 444.600 527.100 ;
        RECT 433.950 523.950 436.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 434.400 521.400 435.600 523.650 ;
        RECT 440.400 522.900 441.600 523.650 ;
        RECT 434.400 520.050 435.450 521.400 ;
        RECT 439.950 520.800 442.050 522.900 ;
        RECT 427.950 517.950 430.050 520.050 ;
        RECT 433.950 517.950 436.050 520.050 ;
        RECT 427.950 505.950 430.050 508.050 ;
        RECT 428.400 502.050 429.450 505.950 ;
        RECT 434.400 505.050 435.450 517.950 ;
        RECT 433.950 502.950 436.050 505.050 ;
        RECT 439.950 502.950 442.050 505.050 ;
        RECT 427.950 499.950 430.050 502.050 ;
        RECT 433.950 499.800 436.050 501.900 ;
        RECT 424.950 493.950 427.050 496.050 ;
        RECT 434.400 495.600 435.450 499.800 ;
        RECT 440.400 495.600 441.450 502.950 ;
        RECT 425.400 489.450 426.450 493.950 ;
        RECT 434.400 493.350 435.600 495.600 ;
        RECT 440.400 493.350 441.600 495.600 ;
        RECT 430.950 490.950 433.050 493.050 ;
        RECT 433.950 490.950 436.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 446.400 492.450 447.600 492.600 ;
        RECT 449.400 492.450 450.450 547.950 ;
        RECT 454.950 544.950 457.050 547.050 ;
        RECT 451.950 538.950 454.050 541.050 ;
        RECT 452.400 508.050 453.450 538.950 ;
        RECT 455.400 511.050 456.450 544.950 ;
        RECT 458.400 528.600 459.450 551.400 ;
        RECT 476.400 547.050 477.450 562.950 ;
        RECT 482.400 547.050 483.450 586.950 ;
        RECT 487.950 583.950 490.050 586.050 ;
        RECT 484.950 574.950 487.050 577.050 ;
        RECT 485.400 571.050 486.450 574.950 ;
        RECT 484.950 568.950 487.050 571.050 ;
        RECT 488.400 570.600 489.450 583.950 ;
        RECT 488.400 570.450 489.600 570.600 ;
        RECT 488.400 569.400 492.450 570.450 ;
        RECT 488.400 568.350 489.600 569.400 ;
        RECT 487.800 565.950 489.900 568.050 ;
        RECT 484.950 562.950 487.050 565.050 ;
        RECT 485.400 550.050 486.450 562.950 ;
        RECT 487.950 559.950 490.050 562.050 ;
        RECT 484.950 547.950 487.050 550.050 ;
        RECT 475.950 544.950 478.050 547.050 ;
        RECT 481.950 544.950 484.050 547.050 ;
        RECT 476.400 541.050 477.450 544.950 ;
        RECT 475.950 538.950 478.050 541.050 ;
        RECT 483.000 537.450 487.050 538.050 ;
        RECT 482.400 535.950 487.050 537.450 ;
        RECT 458.400 526.350 459.600 528.600 ;
        RECT 466.950 527.100 469.050 529.200 ;
        RECT 482.400 528.600 483.450 535.950 ;
        RECT 458.100 523.950 460.200 526.050 ;
        RECT 463.500 523.950 465.600 526.050 ;
        RECT 464.400 521.400 465.600 523.650 ;
        RECT 454.950 508.950 457.050 511.050 ;
        RECT 451.950 505.950 454.050 508.050 ;
        RECT 455.400 492.600 456.450 508.950 ;
        RECT 464.400 508.050 465.450 521.400 ;
        RECT 467.400 520.050 468.450 527.100 ;
        RECT 482.400 526.350 483.600 528.600 ;
        RECT 484.950 527.100 487.050 529.200 ;
        RECT 476.400 523.950 478.500 526.050 ;
        RECT 481.800 523.950 483.900 526.050 ;
        RECT 476.400 521.400 477.600 523.650 ;
        RECT 466.950 517.950 469.050 520.050 ;
        RECT 476.400 514.050 477.450 521.400 ;
        RECT 475.950 511.950 478.050 514.050 ;
        RECT 485.400 511.050 486.450 527.100 ;
        RECT 488.400 517.050 489.450 559.950 ;
        RECT 491.400 556.050 492.450 569.400 ;
        RECT 490.950 553.950 493.050 556.050 ;
        RECT 491.400 538.050 492.450 553.950 ;
        RECT 494.400 553.050 495.450 586.950 ;
        RECT 502.950 580.950 505.050 583.050 ;
        RECT 496.950 572.100 499.050 574.200 ;
        RECT 493.950 550.950 496.050 553.050 ;
        RECT 497.400 544.050 498.450 572.100 ;
        RECT 499.950 565.800 502.050 567.900 ;
        RECT 496.950 541.950 499.050 544.050 ;
        RECT 500.400 538.050 501.450 565.800 ;
        RECT 503.400 559.050 504.450 580.950 ;
        RECT 505.950 572.100 508.050 574.200 ;
        RECT 506.400 571.350 507.600 572.100 ;
        RECT 506.400 568.950 508.500 571.050 ;
        RECT 511.800 568.950 513.900 571.050 ;
        RECT 512.400 566.400 513.600 568.650 ;
        RECT 502.950 556.950 505.050 559.050 ;
        RECT 508.950 547.950 511.050 550.050 ;
        RECT 505.950 541.950 508.050 544.050 ;
        RECT 490.800 535.950 492.900 538.050 ;
        RECT 493.950 535.950 499.050 538.050 ;
        RECT 499.950 535.950 502.050 538.050 ;
        RECT 493.950 527.100 496.050 529.200 ;
        RECT 500.400 528.600 501.450 535.950 ;
        RECT 506.400 532.200 507.450 541.950 ;
        RECT 509.400 541.050 510.450 547.950 ;
        RECT 512.400 544.050 513.450 566.400 ;
        RECT 511.950 541.950 514.050 544.050 ;
        RECT 508.950 538.950 511.050 541.050 ;
        RECT 505.950 530.100 508.050 532.200 ;
        RECT 506.400 529.350 507.600 530.100 ;
        RECT 494.400 526.350 495.600 527.100 ;
        RECT 500.400 526.350 501.600 528.600 ;
        RECT 505.800 526.950 507.900 529.050 ;
        RECT 511.800 526.950 513.900 529.050 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 497.400 522.900 498.600 523.650 ;
        RECT 496.950 520.800 499.050 522.900 ;
        RECT 508.950 520.950 511.050 523.050 ;
        RECT 487.950 514.950 490.050 517.050 ;
        RECT 496.950 514.950 499.050 517.050 ;
        RECT 484.950 508.950 487.050 511.050 ;
        RECT 457.950 505.950 460.050 508.050 ;
        RECT 463.950 505.950 466.050 508.050 ;
        RECT 458.400 493.050 459.450 505.950 ;
        RECT 460.950 499.950 463.050 502.050 ;
        RECT 464.700 501.300 466.800 503.400 ;
        RECT 446.400 491.400 453.450 492.450 ;
        RECT 431.400 489.450 432.600 490.650 ;
        RECT 425.400 488.400 432.600 489.450 ;
        RECT 437.400 488.400 438.600 490.650 ;
        RECT 446.400 490.350 447.600 491.400 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 421.950 466.950 424.050 469.050 ;
        RECT 425.400 466.050 426.450 484.950 ;
        RECT 437.400 481.050 438.450 488.400 ;
        RECT 446.100 487.950 448.200 490.050 ;
        RECT 436.950 478.950 439.050 481.050 ;
        RECT 433.800 475.950 435.900 478.050 ;
        RECT 412.950 463.950 415.050 466.050 ;
        RECT 424.950 463.950 427.050 466.050 ;
        RECT 409.950 457.950 412.050 460.050 ;
        RECT 401.400 443.400 405.450 444.450 ;
        RECT 395.400 370.350 396.600 371.100 ;
        RECT 397.950 370.950 400.050 373.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 394.950 367.950 397.050 370.050 ;
        RECT 382.950 364.950 385.050 367.050 ;
        RECT 386.400 365.400 387.600 367.650 ;
        RECT 392.400 365.400 393.600 367.650 ;
        RECT 401.400 367.050 402.450 443.400 ;
        RECT 410.400 418.200 411.450 457.950 ;
        RECT 413.400 457.050 414.450 463.950 ;
        RECT 412.950 454.950 415.050 457.050 ;
        RECT 416.400 450.450 417.600 450.600 ;
        RECT 413.400 449.400 417.600 450.450 ;
        RECT 413.400 424.050 414.450 449.400 ;
        RECT 416.400 448.350 417.600 449.400 ;
        RECT 416.100 445.950 418.200 448.050 ;
        RECT 421.500 445.950 423.600 448.050 ;
        RECT 422.400 444.450 423.600 445.650 ;
        RECT 425.400 444.450 426.450 463.950 ;
        RECT 428.100 448.950 430.200 451.050 ;
        RECT 422.400 443.400 426.450 444.450 ;
        RECT 428.400 446.400 429.600 448.650 ;
        RECT 434.400 447.900 435.450 475.950 ;
        RECT 452.400 475.050 453.450 491.400 ;
        RECT 455.400 490.350 456.600 492.600 ;
        RECT 457.950 490.950 460.050 493.050 ;
        RECT 455.100 487.950 457.200 490.050 ;
        RECT 451.950 472.950 454.050 475.050 ;
        RECT 461.400 471.450 462.450 499.950 ;
        RECT 465.300 483.600 466.800 501.300 ;
        RECT 464.700 481.500 466.800 483.600 ;
        RECT 465.300 476.700 466.800 481.500 ;
        RECT 464.700 474.600 466.800 476.700 ;
        RECT 467.700 501.300 469.800 503.400 ;
        RECT 470.700 501.300 472.800 503.400 ;
        RECT 473.700 501.300 475.800 503.400 ;
        RECT 467.700 479.700 468.900 501.300 ;
        RECT 470.700 483.600 472.200 501.300 ;
        RECT 473.700 489.000 474.900 501.300 ;
        RECT 479.100 500.400 481.200 502.500 ;
        RECT 487.200 501.300 489.300 503.400 ;
        RECT 490.200 501.300 492.300 503.400 ;
        RECT 493.200 501.300 495.300 503.400 ;
        RECT 475.800 494.400 477.900 496.500 ;
        RECT 479.700 489.900 480.600 500.400 ;
        RECT 482.100 493.950 484.200 496.050 ;
        RECT 482.400 492.900 483.600 493.650 ;
        RECT 481.950 490.800 484.050 492.900 ;
        RECT 473.100 486.900 475.200 489.000 ;
        RECT 478.500 487.800 480.600 489.900 ;
        RECT 470.100 481.500 472.200 483.600 ;
        RECT 467.700 474.600 469.800 479.700 ;
        RECT 470.700 476.700 472.200 481.500 ;
        RECT 473.700 479.700 474.900 486.900 ;
        RECT 479.700 481.200 480.600 487.800 ;
        RECT 473.100 477.600 475.200 479.700 ;
        RECT 478.500 479.100 480.600 481.200 ;
        RECT 488.100 479.700 489.300 501.300 ;
        RECT 487.200 477.600 489.300 479.700 ;
        RECT 490.500 484.800 491.700 501.300 ;
        RECT 493.500 497.700 494.700 501.300 ;
        RECT 493.500 495.600 495.600 497.700 ;
        RECT 490.500 482.700 492.600 484.800 ;
        RECT 490.500 476.700 491.700 482.700 ;
        RECT 494.100 476.700 495.600 495.600 ;
        RECT 497.400 484.050 498.450 514.950 ;
        RECT 509.400 495.450 510.450 520.950 ;
        RECT 509.400 494.400 513.450 495.450 ;
        RECT 500.100 487.950 502.200 490.050 ;
        RECT 506.100 487.950 508.200 490.050 ;
        RECT 506.400 486.900 507.600 487.650 ;
        RECT 512.400 486.900 513.450 494.400 ;
        RECT 515.400 489.450 516.450 592.800 ;
        RECT 517.950 589.950 520.050 592.050 ;
        RECT 518.400 586.050 519.450 589.950 ;
        RECT 517.950 583.950 520.050 586.050 ;
        RECT 526.950 579.450 529.050 580.050 ;
        RECT 530.400 579.450 531.450 598.800 ;
        RECT 533.400 592.050 534.450 604.950 ;
        RECT 536.400 595.050 537.450 613.950 ;
        RECT 539.400 607.050 540.450 625.950 ;
        RECT 565.950 613.950 568.050 616.050 ;
        RECT 538.950 604.950 541.050 607.050 ;
        RECT 544.950 605.100 547.050 610.050 ;
        RECT 550.950 605.100 553.050 607.200 ;
        RECT 556.950 605.100 559.050 607.200 ;
        RECT 562.950 606.000 565.050 610.050 ;
        RECT 566.400 609.450 567.450 613.950 ;
        RECT 569.400 613.050 570.450 652.950 ;
        RECT 574.950 650.100 577.050 655.050 ;
        RECT 575.400 649.350 576.600 650.100 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 578.400 644.400 579.600 646.650 ;
        RECT 578.400 640.050 579.450 644.400 ;
        RECT 577.950 637.950 580.050 640.050 ;
        RECT 577.950 628.950 580.050 631.050 ;
        RECT 574.950 622.950 577.050 625.050 ;
        RECT 571.950 616.950 574.050 619.050 ;
        RECT 568.950 610.950 571.050 613.050 ;
        RECT 572.400 609.450 573.450 616.950 ;
        RECT 566.400 608.400 573.450 609.450 ;
        RECT 575.400 609.600 576.450 622.950 ;
        RECT 578.400 616.050 579.450 628.950 ;
        RECT 577.950 613.950 580.050 616.050 ;
        RECT 569.400 606.600 570.450 608.400 ;
        RECT 575.400 607.350 576.600 609.600 ;
        RECT 545.400 604.350 546.600 605.100 ;
        RECT 551.400 604.350 552.600 605.100 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 601.950 547.050 604.050 ;
        RECT 547.950 601.950 550.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 538.950 598.950 541.050 601.050 ;
        RECT 542.400 600.000 543.600 601.650 ;
        RECT 535.950 592.950 538.050 595.050 ;
        RECT 532.950 589.950 535.050 592.050 ;
        RECT 526.950 578.400 531.450 579.450 ;
        RECT 539.400 579.450 540.450 598.950 ;
        RECT 541.950 595.950 544.050 600.000 ;
        RECT 548.400 599.400 549.600 601.650 ;
        RECT 557.400 601.050 558.450 605.100 ;
        RECT 563.400 604.350 564.600 606.000 ;
        RECT 569.400 604.350 570.600 606.600 ;
        RECT 574.800 604.950 576.900 607.050 ;
        RECT 580.800 604.950 582.900 607.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 541.950 592.800 544.050 594.900 ;
        RECT 542.400 586.050 543.450 592.800 ;
        RECT 548.400 592.050 549.450 599.400 ;
        RECT 556.950 598.950 559.050 601.050 ;
        RECT 566.400 600.900 567.600 601.650 ;
        RECT 565.950 598.800 568.050 600.900 ;
        RECT 571.950 598.950 574.050 601.050 ;
        RECT 577.950 600.450 580.050 604.050 ;
        RECT 575.400 600.000 580.050 600.450 ;
        RECT 575.400 599.400 579.450 600.000 ;
        RECT 547.950 589.950 550.050 592.050 ;
        RECT 541.950 583.950 544.050 586.050 ;
        RECT 553.950 583.950 556.050 586.050 ;
        RECT 565.950 583.950 568.050 586.050 ;
        RECT 554.400 580.050 555.450 583.950 ;
        RECT 539.400 578.400 543.450 579.450 ;
        RECT 526.950 577.950 529.050 578.400 ;
        RECT 520.950 571.950 523.050 574.050 ;
        RECT 527.400 573.600 528.450 577.950 ;
        RECT 521.400 547.050 522.450 571.950 ;
        RECT 527.400 571.350 528.600 573.600 ;
        RECT 532.950 572.100 535.050 574.200 ;
        RECT 533.400 571.350 534.600 572.100 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 530.400 567.900 531.600 568.650 ;
        RECT 536.400 568.050 537.600 568.650 ;
        RECT 529.950 565.800 532.050 567.900 ;
        RECT 536.400 566.400 541.050 568.050 ;
        RECT 537.000 565.950 541.050 566.400 ;
        RECT 530.400 562.050 531.450 565.800 ;
        RECT 542.400 562.050 543.450 578.400 ;
        RECT 553.950 577.950 556.050 580.050 ;
        RECT 544.950 571.950 547.050 577.050 ;
        RECT 550.950 572.100 553.050 574.200 ;
        RECT 566.400 573.600 567.450 583.950 ;
        RECT 572.400 573.600 573.450 598.950 ;
        RECT 575.400 589.050 576.450 599.400 ;
        RECT 584.400 598.050 585.450 659.400 ;
        RECT 587.400 652.050 588.450 673.950 ;
        RECT 595.950 661.950 598.050 664.050 ;
        RECT 586.950 649.950 589.050 652.050 ;
        RECT 596.400 651.600 597.450 661.950 ;
        RECT 599.400 661.050 600.450 712.950 ;
        RECT 607.950 697.950 610.050 700.050 ;
        RECT 608.400 691.050 609.450 697.950 ;
        RECT 607.950 688.950 610.050 691.050 ;
        RECT 608.400 684.600 609.450 688.950 ;
        RECT 608.400 682.350 609.600 684.600 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 607.950 679.950 610.050 682.050 ;
        RECT 605.400 678.900 606.600 679.650 ;
        RECT 604.950 673.950 607.050 678.900 ;
        RECT 614.400 678.450 615.450 719.400 ;
        RECT 616.950 718.950 619.050 721.050 ;
        RECT 619.950 718.950 622.050 721.050 ;
        RECT 622.950 718.950 625.050 723.000 ;
        RECT 628.950 718.950 631.050 723.000 ;
        RECT 634.950 718.950 637.050 724.050 ;
        RECT 641.400 722.400 642.600 724.650 ;
        RECT 641.400 721.050 642.450 722.400 ;
        RECT 646.950 721.950 649.050 724.050 ;
        RECT 656.400 723.900 657.600 724.650 ;
        RECT 637.950 719.400 642.450 721.050 ;
        RECT 637.950 718.950 642.000 719.400 ;
        RECT 617.400 697.050 618.450 718.950 ;
        RECT 620.400 715.050 621.450 718.950 ;
        RECT 619.950 712.950 622.050 715.050 ;
        RECT 647.400 712.050 648.450 721.950 ;
        RECT 655.950 721.800 658.050 723.900 ;
        RECT 662.400 722.400 663.600 724.650 ;
        RECT 662.400 715.050 663.450 722.400 ;
        RECT 664.950 721.950 667.050 724.050 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 637.950 709.950 640.050 712.050 ;
        RECT 646.950 709.950 649.050 712.050 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 616.950 694.950 619.050 697.050 ;
        RECT 611.400 677.400 615.450 678.450 ;
        RECT 617.400 678.450 618.450 694.950 ;
        RECT 622.950 683.100 625.050 685.200 ;
        RECT 629.400 684.600 630.450 697.950 ;
        RECT 623.400 682.350 624.600 683.100 ;
        RECT 629.400 682.350 630.600 684.600 ;
        RECT 634.950 683.100 637.050 685.200 ;
        RECT 638.400 685.050 639.450 709.950 ;
        RECT 652.950 706.950 655.050 709.050 ;
        RECT 646.950 703.950 649.050 706.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 625.950 679.950 628.050 682.050 ;
        RECT 628.950 679.950 631.050 682.050 ;
        RECT 626.400 678.900 627.600 679.650 ;
        RECT 635.400 679.050 636.450 683.100 ;
        RECT 637.950 682.950 640.050 685.050 ;
        RECT 640.950 683.100 643.050 685.200 ;
        RECT 647.400 684.600 648.450 703.950 ;
        RECT 641.400 682.350 642.600 683.100 ;
        RECT 647.400 682.350 648.600 684.600 ;
        RECT 640.950 679.950 643.050 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 617.400 677.400 621.450 678.450 ;
        RECT 598.950 658.950 601.050 661.050 ;
        RECT 607.950 658.950 610.050 661.050 ;
        RECT 596.400 649.350 597.600 651.600 ;
        RECT 601.950 650.100 604.050 652.200 ;
        RECT 602.400 649.350 603.600 650.100 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 598.950 646.950 601.050 649.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 593.400 645.900 594.600 646.650 ;
        RECT 592.950 643.800 595.050 645.900 ;
        RECT 599.400 644.400 600.600 646.650 ;
        RECT 608.400 645.900 609.450 658.950 ;
        RECT 599.400 640.050 600.450 644.400 ;
        RECT 607.950 643.800 610.050 645.900 ;
        RECT 598.950 637.950 601.050 640.050 ;
        RECT 611.400 631.050 612.450 677.400 ;
        RECT 620.400 651.600 621.450 677.400 ;
        RECT 625.950 676.800 628.050 678.900 ;
        RECT 631.950 676.950 634.050 679.050 ;
        RECT 634.950 676.950 637.050 679.050 ;
        RECT 644.400 677.400 645.600 679.650 ;
        RECT 620.400 649.350 621.600 651.600 ;
        RECT 628.950 650.100 631.050 652.200 ;
        RECT 616.950 646.950 619.050 649.050 ;
        RECT 619.950 646.950 622.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 617.400 644.400 618.600 646.650 ;
        RECT 623.400 644.400 624.600 646.650 ;
        RECT 617.400 642.450 618.450 644.400 ;
        RECT 617.400 641.400 621.450 642.450 ;
        RECT 620.400 634.050 621.450 641.400 ;
        RECT 623.400 637.050 624.450 644.400 ;
        RECT 629.400 643.050 630.450 650.100 ;
        RECT 628.950 640.950 631.050 643.050 ;
        RECT 632.400 640.050 633.450 676.950 ;
        RECT 644.400 670.050 645.450 677.400 ;
        RECT 643.950 667.950 646.050 670.050 ;
        RECT 649.950 661.950 652.050 664.050 ;
        RECT 637.950 650.100 640.050 652.200 ;
        RECT 643.950 651.000 646.050 655.050 ;
        RECT 638.400 649.350 639.600 650.100 ;
        RECT 644.400 649.350 645.600 651.000 ;
        RECT 637.950 646.950 640.050 649.050 ;
        RECT 640.950 646.950 643.050 649.050 ;
        RECT 643.950 646.950 646.050 649.050 ;
        RECT 641.400 645.900 642.600 646.650 ;
        RECT 650.400 645.900 651.450 661.950 ;
        RECT 653.400 658.050 654.450 706.950 ;
        RECT 655.950 700.950 658.050 703.050 ;
        RECT 656.400 679.050 657.450 700.950 ;
        RECT 665.400 700.050 666.450 721.950 ;
        RECT 668.400 709.050 669.450 728.400 ;
        RECT 677.400 727.350 678.600 729.600 ;
        RECT 682.950 728.100 685.050 730.200 ;
        RECT 683.400 727.350 684.600 728.100 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 674.400 722.400 675.600 724.650 ;
        RECT 680.400 722.400 681.600 724.650 ;
        RECT 667.950 706.950 670.050 709.050 ;
        RECT 664.950 697.950 667.050 700.050 ;
        RECT 661.950 694.950 664.050 697.050 ;
        RECT 662.400 684.600 663.450 694.950 ;
        RECT 674.400 691.050 675.450 722.400 ;
        RECT 680.400 715.050 681.450 722.400 ;
        RECT 685.950 721.950 688.050 724.050 ;
        RECT 679.950 712.950 682.050 715.050 ;
        RECT 686.400 697.050 687.450 721.950 ;
        RECT 685.950 694.950 688.050 697.050 ;
        RECT 676.950 691.950 679.050 694.050 ;
        RECT 673.950 688.950 676.050 691.050 ;
        RECT 662.400 682.350 663.600 684.600 ;
        RECT 667.950 683.100 670.050 685.200 ;
        RECT 668.400 682.350 669.600 683.100 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 664.950 679.950 667.050 682.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 655.950 676.950 658.050 679.050 ;
        RECT 665.400 678.900 666.600 679.650 ;
        RECT 664.950 676.800 667.050 678.900 ;
        RECT 667.950 670.950 670.050 673.050 ;
        RECT 652.950 655.950 655.050 658.050 ;
        RECT 652.950 652.800 655.050 654.900 ;
        RECT 640.950 643.800 643.050 645.900 ;
        RECT 649.950 643.800 652.050 645.900 ;
        RECT 653.400 643.050 654.450 652.800 ;
        RECT 661.950 651.000 664.050 655.050 ;
        RECT 668.400 652.050 669.450 670.950 ;
        RECT 677.400 664.050 678.450 691.950 ;
        RECT 682.950 683.100 685.050 685.200 ;
        RECT 689.400 685.050 690.450 739.950 ;
        RECT 701.400 736.050 702.450 755.400 ;
        RECT 707.400 751.050 708.450 755.400 ;
        RECT 712.950 754.950 715.050 757.050 ;
        RECT 706.950 748.950 709.050 751.050 ;
        RECT 703.950 742.950 706.050 745.050 ;
        RECT 700.950 733.950 703.050 736.050 ;
        RECT 691.950 727.950 694.050 733.050 ;
        RECT 697.950 728.100 700.050 730.200 ;
        RECT 704.400 729.600 705.450 742.950 ;
        RECT 709.950 730.950 712.050 733.050 ;
        RECT 698.400 727.350 699.600 728.100 ;
        RECT 704.400 727.350 705.600 729.600 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 695.400 723.900 696.600 724.650 ;
        RECT 694.950 721.800 697.050 723.900 ;
        RECT 701.400 722.400 702.600 724.650 ;
        RECT 695.400 706.050 696.450 721.800 ;
        RECT 701.400 718.050 702.450 722.400 ;
        RECT 706.950 721.950 709.050 724.050 ;
        RECT 700.950 715.950 703.050 718.050 ;
        RECT 694.950 703.950 697.050 706.050 ;
        RECT 695.400 688.050 696.450 703.950 ;
        RECT 707.400 694.050 708.450 721.950 ;
        RECT 710.400 715.050 711.450 730.950 ;
        RECT 713.400 730.050 714.450 754.950 ;
        RECT 716.400 751.050 717.450 763.950 ;
        RECT 715.950 748.950 718.050 751.050 ;
        RECT 719.400 733.050 720.450 775.950 ;
        RECT 722.400 769.050 723.450 800.400 ;
        RECT 727.950 799.800 730.050 801.900 ;
        RECT 734.400 793.050 735.450 814.950 ;
        RECT 752.400 811.050 753.450 814.950 ;
        RECT 742.950 807.000 745.050 811.050 ;
        RECT 751.950 808.950 754.050 811.050 ;
        RECT 743.400 805.350 744.600 807.000 ;
        RECT 748.950 805.950 751.050 808.050 ;
        RECT 757.950 807.000 760.050 811.050 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 736.950 799.950 739.050 802.050 ;
        RECT 740.400 800.400 741.600 802.650 ;
        RECT 737.400 796.050 738.450 799.950 ;
        RECT 736.950 793.950 739.050 796.050 ;
        RECT 733.950 790.950 736.050 793.050 ;
        RECT 740.400 787.050 741.450 800.400 ;
        RECT 745.950 796.950 748.050 799.050 ;
        RECT 739.950 784.950 742.050 787.050 ;
        RECT 742.950 772.950 745.050 775.050 ;
        RECT 724.950 769.950 727.050 772.050 ;
        RECT 721.950 766.950 724.050 769.050 ;
        RECT 725.400 766.050 726.450 769.950 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 727.950 761.100 730.050 766.050 ;
        RECT 733.950 761.100 736.050 763.200 ;
        RECT 739.950 761.100 742.050 763.200 ;
        RECT 728.400 760.350 729.600 761.100 ;
        RECT 734.400 760.350 735.600 761.100 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 733.950 757.950 736.050 760.050 ;
        RECT 725.400 755.400 726.600 757.650 ;
        RECT 731.400 755.400 732.600 757.650 ;
        RECT 740.400 757.050 741.450 761.100 ;
        RECT 721.950 742.950 724.050 745.050 ;
        RECT 718.950 730.950 721.050 733.050 ;
        RECT 722.400 730.050 723.450 742.950 ;
        RECT 725.400 730.050 726.450 755.400 ;
        RECT 727.950 751.950 730.050 754.050 ;
        RECT 728.400 730.050 729.450 751.950 ;
        RECT 731.400 751.050 732.450 755.400 ;
        RECT 739.950 754.950 742.050 757.050 ;
        RECT 730.950 748.950 733.050 751.050 ;
        RECT 733.950 733.950 736.050 736.050 ;
        RECT 712.950 729.450 715.050 730.050 ;
        RECT 716.400 729.450 717.600 729.600 ;
        RECT 712.950 728.400 717.600 729.450 ;
        RECT 712.950 727.950 715.050 728.400 ;
        RECT 716.400 727.350 717.600 728.400 ;
        RECT 721.950 727.950 724.050 730.050 ;
        RECT 724.800 727.950 726.900 730.050 ;
        RECT 727.950 727.950 730.050 730.050 ;
        RECT 734.400 729.600 735.450 733.950 ;
        RECT 734.400 727.350 735.600 729.600 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 724.950 724.800 727.050 726.900 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 712.950 721.950 715.050 724.050 ;
        RECT 719.400 723.900 720.600 724.650 ;
        RECT 709.950 712.950 712.050 715.050 ;
        RECT 706.950 691.950 709.050 694.050 ;
        RECT 694.950 685.950 697.050 688.050 ;
        RECT 683.400 682.350 684.600 683.100 ;
        RECT 688.950 682.950 691.050 685.050 ;
        RECT 691.950 682.950 694.050 685.050 ;
        RECT 697.950 682.950 700.050 685.050 ;
        RECT 700.950 683.100 703.050 685.200 ;
        RECT 709.950 684.000 712.050 688.050 ;
        RECT 713.400 685.050 714.450 721.950 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 721.950 715.950 724.050 718.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 686.400 678.900 687.600 679.650 ;
        RECT 692.400 678.900 693.450 682.950 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 685.950 676.800 688.050 678.900 ;
        RECT 691.950 676.800 694.050 678.900 ;
        RECT 679.950 664.950 682.050 667.050 ;
        RECT 676.950 661.950 679.050 664.050 ;
        RECT 670.950 658.950 673.050 661.050 ;
        RECT 662.400 649.350 663.600 651.000 ;
        RECT 667.950 649.950 670.050 652.050 ;
        RECT 658.950 646.950 661.050 649.050 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 659.400 644.400 660.600 646.650 ;
        RECT 665.400 645.900 666.600 646.650 ;
        RECT 637.950 640.950 640.050 643.050 ;
        RECT 643.950 640.950 646.050 643.050 ;
        RECT 652.950 640.950 655.050 643.050 ;
        RECT 631.950 637.950 634.050 640.050 ;
        RECT 622.950 634.950 625.050 637.050 ;
        RECT 619.950 631.950 622.050 634.050 ;
        RECT 610.950 628.950 613.050 631.050 ;
        RECT 587.400 618.300 590.400 620.400 ;
        RECT 591.300 618.300 593.400 620.400 ;
        RECT 610.200 618.300 612.300 620.400 ;
        RECT 587.400 599.400 588.900 618.300 ;
        RECT 591.300 612.300 592.500 618.300 ;
        RECT 590.400 610.200 592.500 612.300 ;
        RECT 583.950 595.950 586.050 598.050 ;
        RECT 587.400 597.300 589.500 599.400 ;
        RECT 574.950 586.950 577.050 589.050 ;
        RECT 551.400 571.350 552.600 572.100 ;
        RECT 566.400 571.350 567.600 573.600 ;
        RECT 572.400 571.350 573.600 573.600 ;
        RECT 580.950 571.950 583.050 577.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 559.950 568.950 562.050 571.050 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 548.400 567.900 549.600 568.650 ;
        RECT 547.950 565.800 550.050 567.900 ;
        RECT 554.400 566.400 555.600 568.650 ;
        RECT 554.400 562.050 555.450 566.400 ;
        RECT 529.950 559.950 532.050 562.050 ;
        RECT 541.950 559.950 544.050 562.050 ;
        RECT 553.950 559.950 556.050 562.050 ;
        RECT 532.950 553.950 535.050 556.050 ;
        RECT 520.950 544.950 523.050 547.050 ;
        RECT 518.400 540.300 521.400 542.400 ;
        RECT 522.300 540.300 524.400 542.400 ;
        RECT 533.400 541.050 534.450 553.950 ;
        RECT 560.400 550.050 561.450 568.950 ;
        RECT 580.950 568.800 583.050 570.900 ;
        RECT 569.400 567.900 570.600 568.650 ;
        RECT 575.400 568.050 576.600 568.650 ;
        RECT 568.950 565.800 571.050 567.900 ;
        RECT 575.400 566.400 580.050 568.050 ;
        RECT 576.000 565.950 580.050 566.400 ;
        RECT 569.400 559.050 570.450 565.800 ;
        RECT 581.400 559.050 582.450 568.800 ;
        RECT 568.950 556.950 571.050 559.050 ;
        RECT 580.950 556.950 583.050 559.050 ;
        RECT 568.950 553.800 571.050 555.900 ;
        RECT 559.950 547.950 562.050 550.050 ;
        RECT 565.950 547.950 568.050 550.050 ;
        RECT 550.950 544.950 553.050 547.050 ;
        RECT 518.400 521.400 519.900 540.300 ;
        RECT 522.300 534.300 523.500 540.300 ;
        RECT 521.400 532.200 523.500 534.300 ;
        RECT 518.400 519.300 520.500 521.400 ;
        RECT 519.300 515.700 520.500 519.300 ;
        RECT 522.300 515.700 523.500 532.200 ;
        RECT 524.700 537.300 526.800 539.400 ;
        RECT 532.950 538.950 535.050 541.050 ;
        RECT 541.200 540.300 543.300 542.400 ;
        RECT 524.700 515.700 525.900 537.300 ;
        RECT 533.400 535.800 535.500 537.900 ;
        RECT 538.800 537.300 540.900 539.400 ;
        RECT 533.400 529.200 534.300 535.800 ;
        RECT 539.100 530.100 540.300 537.300 ;
        RECT 541.800 535.500 543.300 540.300 ;
        RECT 544.200 537.300 546.300 542.400 ;
        RECT 541.800 533.400 543.900 535.500 ;
        RECT 529.950 525.000 532.050 529.050 ;
        RECT 533.400 527.100 535.500 529.200 ;
        RECT 538.800 528.000 540.900 530.100 ;
        RECT 530.400 523.350 531.600 525.000 ;
        RECT 529.800 520.950 531.900 523.050 ;
        RECT 533.400 516.600 534.300 527.100 ;
        RECT 536.100 520.500 538.200 522.600 ;
        RECT 518.700 513.600 520.800 515.700 ;
        RECT 521.700 513.600 523.800 515.700 ;
        RECT 524.700 513.600 526.800 515.700 ;
        RECT 532.800 514.500 534.900 516.600 ;
        RECT 539.100 515.700 540.300 528.000 ;
        RECT 541.800 515.700 543.300 533.400 ;
        RECT 545.100 515.700 546.300 537.300 ;
        RECT 538.200 513.600 540.300 515.700 ;
        RECT 541.200 513.600 543.300 515.700 ;
        RECT 544.200 513.600 546.300 515.700 ;
        RECT 547.200 540.300 549.300 542.400 ;
        RECT 547.200 535.500 548.700 540.300 ;
        RECT 547.200 533.400 549.300 535.500 ;
        RECT 547.200 515.700 548.700 533.400 ;
        RECT 551.400 529.050 552.450 544.950 ;
        RECT 550.950 526.950 553.050 529.050 ;
        RECT 556.800 526.950 558.900 529.050 ;
        RECT 553.950 522.450 556.050 526.050 ;
        RECT 557.400 525.450 558.600 526.650 ;
        RECT 560.400 525.450 561.450 547.950 ;
        RECT 566.400 541.050 567.450 547.950 ;
        RECT 565.950 538.950 568.050 541.050 ;
        RECT 565.800 526.950 567.900 529.050 ;
        RECT 557.400 524.400 561.450 525.450 ;
        RECT 566.400 524.400 567.600 526.650 ;
        RECT 553.950 522.000 558.450 522.450 ;
        RECT 554.400 521.400 558.450 522.000 ;
        RECT 547.200 513.600 549.300 515.700 ;
        RECT 535.950 508.950 538.050 511.050 ;
        RECT 529.950 505.950 532.050 508.050 ;
        RECT 523.950 495.000 526.050 499.050 ;
        RECT 530.400 495.600 531.450 505.950 ;
        RECT 524.400 493.350 525.600 495.000 ;
        RECT 530.400 493.350 531.600 495.600 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 526.950 490.950 529.050 493.050 ;
        RECT 529.950 490.950 532.050 493.050 ;
        RECT 521.400 489.900 522.600 490.650 ;
        RECT 527.400 489.900 528.600 490.650 ;
        RECT 515.400 488.400 519.450 489.450 ;
        RECT 505.950 484.800 508.050 486.900 ;
        RECT 511.950 484.800 514.050 486.900 ;
        RECT 496.950 481.950 499.050 484.050 ;
        RECT 470.700 474.600 472.800 476.700 ;
        RECT 489.600 474.600 491.700 476.700 ;
        RECT 492.600 474.600 495.600 476.700 ;
        RECT 461.400 470.400 465.450 471.450 ;
        RECT 442.950 466.950 445.050 469.050 ;
        RECT 437.100 448.950 439.200 451.050 ;
        RECT 422.400 430.050 423.450 443.400 ;
        RECT 421.950 427.950 424.050 430.050 ;
        RECT 428.400 424.050 429.450 446.400 ;
        RECT 433.950 445.800 436.050 447.900 ;
        RECT 437.400 446.400 438.600 448.650 ;
        RECT 430.950 439.950 433.050 442.050 ;
        RECT 412.950 421.950 415.050 424.050 ;
        RECT 427.950 421.950 430.050 424.050 ;
        RECT 409.950 416.100 412.050 418.200 ;
        RECT 410.400 415.350 411.600 416.100 ;
        RECT 415.950 415.950 418.050 418.050 ;
        RECT 431.400 417.600 432.450 439.950 ;
        RECT 434.400 439.050 435.450 445.800 ;
        RECT 433.950 436.950 436.050 439.050 ;
        RECT 437.400 433.050 438.450 446.400 ;
        RECT 436.950 430.950 439.050 433.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 407.400 411.900 408.600 412.650 ;
        RECT 406.950 409.800 409.050 411.900 ;
        RECT 409.950 388.950 412.050 391.050 ;
        RECT 410.400 372.600 411.450 388.950 ;
        RECT 416.400 388.050 417.450 415.950 ;
        RECT 431.400 415.350 432.600 417.600 ;
        RECT 425.100 412.950 427.200 415.050 ;
        RECT 430.500 412.950 432.600 415.050 ;
        RECT 425.400 411.900 426.600 412.650 ;
        RECT 424.950 409.800 427.050 411.900 ;
        RECT 421.950 403.950 424.050 406.050 ;
        RECT 422.400 400.050 423.450 403.950 ;
        RECT 421.950 397.950 424.050 400.050 ;
        RECT 415.950 385.950 418.050 388.050 ;
        RECT 410.400 370.350 411.600 372.600 ;
        RECT 418.950 371.100 421.050 373.200 ;
        RECT 419.400 370.350 420.600 371.100 ;
        RECT 410.100 367.950 412.200 370.050 ;
        RECT 415.500 367.950 417.600 370.050 ;
        RECT 418.800 367.950 420.900 370.050 ;
        RECT 368.400 337.350 369.600 338.100 ;
        RECT 374.400 337.350 375.600 339.600 ;
        RECT 379.950 337.950 382.050 340.050 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 358.950 331.800 361.050 333.900 ;
        RECT 361.950 331.950 364.050 334.050 ;
        RECT 365.400 333.900 366.600 334.650 ;
        RECT 371.400 333.900 372.600 334.650 ;
        RECT 362.400 328.050 363.450 331.950 ;
        RECT 364.950 331.800 367.050 333.900 ;
        RECT 370.950 331.800 373.050 333.900 ;
        RECT 377.400 333.000 378.600 334.650 ;
        RECT 361.950 325.950 364.050 328.050 ;
        RECT 355.950 322.950 358.050 325.050 ;
        RECT 352.950 313.950 355.050 316.050 ;
        RECT 356.400 304.050 357.450 322.950 ;
        RECT 365.400 304.050 366.450 331.800 ;
        RECT 367.950 328.950 370.050 331.050 ;
        RECT 368.400 316.050 369.450 328.950 ;
        RECT 367.950 313.950 370.050 316.050 ;
        RECT 371.400 313.050 372.450 331.800 ;
        RECT 373.950 328.950 376.050 331.050 ;
        RECT 376.950 328.950 379.050 333.000 ;
        RECT 383.400 331.050 384.450 364.950 ;
        RECT 386.400 361.050 387.450 365.400 ;
        RECT 392.400 361.050 393.450 365.400 ;
        RECT 400.950 364.950 403.050 367.050 ;
        RECT 416.400 366.900 417.600 367.650 ;
        RECT 415.950 364.800 418.050 366.900 ;
        RECT 385.950 358.950 388.050 361.050 ;
        RECT 391.950 358.950 394.050 361.050 ;
        RECT 406.950 358.950 409.050 361.050 ;
        RECT 397.950 343.950 400.050 346.050 ;
        RECT 388.950 338.100 391.050 340.200 ;
        RECT 389.400 337.350 390.600 338.100 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 392.400 332.400 393.600 334.650 ;
        RECT 382.950 328.950 385.050 331.050 ;
        RECT 388.950 328.950 391.050 331.050 ;
        RECT 370.950 310.950 373.050 313.050 ;
        RECT 370.950 304.950 373.050 307.050 ;
        RECT 355.950 301.950 358.050 304.050 ;
        RECT 364.950 301.950 367.050 304.050 ;
        RECT 355.800 298.200 357.900 300.300 ;
        RECT 364.800 298.500 366.900 300.600 ;
        RECT 353.400 294.450 354.600 294.600 ;
        RECT 344.400 293.400 348.450 294.450 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 338.400 288.900 339.600 289.650 ;
        RECT 337.950 286.800 340.050 288.900 ;
        RECT 313.950 271.950 316.050 274.050 ;
        RECT 328.950 271.950 331.050 274.050 ;
        RECT 314.400 262.050 315.450 271.950 ;
        RECT 328.950 268.800 331.050 270.900 ;
        RECT 313.950 259.950 316.050 262.050 ;
        RECT 316.950 260.100 319.050 265.050 ;
        RECT 322.950 261.000 325.050 265.050 ;
        RECT 329.400 261.600 330.450 268.800 ;
        RECT 347.400 265.050 348.450 293.400 ;
        RECT 350.400 293.400 354.600 294.450 ;
        RECT 334.950 262.950 337.050 265.050 ;
        RECT 346.950 262.950 349.050 265.050 ;
        RECT 317.400 259.350 318.600 260.100 ;
        RECT 323.400 259.350 324.600 261.000 ;
        RECT 329.400 259.350 330.600 261.600 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 320.400 254.400 321.600 256.650 ;
        RECT 326.400 255.900 327.600 256.650 ;
        RECT 335.400 255.900 336.450 262.950 ;
        RECT 343.950 260.100 346.050 262.200 ;
        RECT 350.400 261.600 351.450 293.400 ;
        RECT 353.400 292.350 354.600 293.400 ;
        RECT 353.100 289.950 355.200 292.050 ;
        RECT 356.100 285.600 357.000 298.200 ;
        RECT 362.400 295.350 363.600 297.600 ;
        RECT 362.100 292.950 364.200 295.050 ;
        RECT 357.900 291.900 360.000 292.200 ;
        RECT 366.000 291.900 366.900 298.500 ;
        RECT 357.900 291.000 366.900 291.900 ;
        RECT 357.900 290.100 360.000 291.000 ;
        RECT 363.000 289.200 365.100 290.100 ;
        RECT 357.900 288.000 365.100 289.200 ;
        RECT 357.900 287.100 360.000 288.000 ;
        RECT 355.500 283.500 357.600 285.600 ;
        RECT 362.100 284.100 364.200 286.200 ;
        RECT 366.000 285.900 366.900 291.000 ;
        RECT 367.800 289.950 369.900 292.050 ;
        RECT 368.400 288.900 369.600 289.650 ;
        RECT 367.950 286.800 370.050 288.900 ;
        RECT 365.400 283.800 367.500 285.900 ;
        RECT 362.400 281.550 363.600 283.800 ;
        RECT 358.950 274.950 361.050 277.050 ;
        RECT 344.400 259.350 345.600 260.100 ;
        RECT 350.400 259.350 351.600 261.600 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 347.400 255.900 348.600 256.650 ;
        RECT 314.400 223.050 315.450 253.950 ;
        RECT 320.400 244.050 321.450 254.400 ;
        RECT 325.950 253.800 328.050 255.900 ;
        RECT 334.950 253.800 337.050 255.900 ;
        RECT 346.950 253.800 349.050 255.900 ;
        RECT 353.400 255.000 354.600 256.650 ;
        RECT 359.400 255.900 360.450 274.950 ;
        RECT 362.400 262.050 363.450 281.550 ;
        RECT 371.400 277.050 372.450 304.950 ;
        RECT 374.400 283.050 375.450 328.950 ;
        RECT 376.950 325.800 379.050 327.900 ;
        RECT 377.400 295.050 378.450 325.800 ;
        RECT 379.950 301.950 382.050 304.050 ;
        RECT 380.400 295.200 381.450 301.950 ;
        RECT 376.950 292.950 379.050 295.050 ;
        RECT 379.950 293.100 382.050 295.200 ;
        RECT 385.950 293.100 388.050 295.200 ;
        RECT 389.400 294.450 390.450 328.950 ;
        RECT 392.400 298.050 393.450 332.400 ;
        RECT 398.400 331.050 399.450 343.950 ;
        RECT 407.400 340.200 408.450 358.950 ;
        RECT 416.400 358.050 417.450 364.800 ;
        RECT 415.950 355.950 418.050 358.050 ;
        RECT 406.950 338.100 409.050 340.200 ;
        RECT 412.950 338.100 415.050 340.200 ;
        RECT 422.400 340.050 423.450 397.950 ;
        RECT 425.400 366.900 426.450 409.800 ;
        RECT 443.400 406.050 444.450 466.950 ;
        RECT 446.700 462.300 448.800 464.400 ;
        RECT 447.300 457.500 448.800 462.300 ;
        RECT 446.700 455.400 448.800 457.500 ;
        RECT 447.300 437.700 448.800 455.400 ;
        RECT 446.700 435.600 448.800 437.700 ;
        RECT 449.700 459.300 451.800 464.400 ;
        RECT 452.700 462.300 454.800 464.400 ;
        RECT 449.700 437.700 450.900 459.300 ;
        RECT 452.700 457.500 454.200 462.300 ;
        RECT 455.100 459.300 457.200 461.400 ;
        RECT 452.100 455.400 454.200 457.500 ;
        RECT 452.700 437.700 454.200 455.400 ;
        RECT 455.700 452.100 456.900 459.300 ;
        RECT 460.500 457.800 462.600 459.900 ;
        RECT 455.100 450.000 457.200 452.100 ;
        RECT 461.700 451.200 462.600 457.800 ;
        RECT 455.700 437.700 456.900 450.000 ;
        RECT 460.500 449.100 462.600 451.200 ;
        RECT 457.800 442.500 459.900 444.600 ;
        RECT 461.700 438.600 462.600 449.100 ;
        RECT 464.400 447.600 465.450 470.400 ;
        RECT 478.950 466.950 481.050 469.050 ;
        RECT 471.600 462.300 473.700 464.400 ;
        RECT 474.600 462.300 477.600 464.400 ;
        RECT 469.200 459.300 471.300 461.400 ;
        RECT 464.400 445.350 465.600 447.600 ;
        RECT 464.100 442.950 466.200 445.050 ;
        RECT 449.700 435.600 451.800 437.700 ;
        RECT 452.700 435.600 454.800 437.700 ;
        RECT 455.700 435.600 457.800 437.700 ;
        RECT 461.100 436.500 463.200 438.600 ;
        RECT 470.100 437.700 471.300 459.300 ;
        RECT 472.500 456.300 473.700 462.300 ;
        RECT 472.500 454.200 474.600 456.300 ;
        RECT 472.500 437.700 473.700 454.200 ;
        RECT 476.100 443.400 477.600 462.300 ;
        RECT 479.400 460.050 480.450 466.950 ;
        RECT 478.950 457.950 481.050 460.050 ;
        RECT 502.950 457.950 505.050 460.050 ;
        RECT 475.500 441.300 477.600 443.400 ;
        RECT 475.500 437.700 476.700 441.300 ;
        RECT 469.200 435.600 471.300 437.700 ;
        RECT 472.200 435.600 474.300 437.700 ;
        RECT 475.200 435.600 477.300 437.700 ;
        RECT 457.950 430.950 460.050 433.050 ;
        RECT 445.950 421.950 448.050 424.050 ;
        RECT 446.400 417.600 447.450 421.950 ;
        RECT 446.400 415.350 447.600 417.600 ;
        RECT 454.950 416.100 457.050 418.200 ;
        RECT 446.400 412.950 448.500 415.050 ;
        RECT 451.800 412.950 453.900 415.050 ;
        RECT 452.400 411.900 453.600 412.650 ;
        RECT 451.950 409.800 454.050 411.900 ;
        RECT 442.950 403.950 445.050 406.050 ;
        RECT 442.950 400.800 445.050 402.900 ;
        RECT 430.950 376.950 433.050 379.050 ;
        RECT 431.400 372.600 432.450 376.950 ;
        RECT 431.400 370.350 432.600 372.600 ;
        RECT 436.950 371.100 439.050 373.200 ;
        RECT 437.400 370.350 438.600 371.100 ;
        RECT 443.400 370.050 444.450 400.800 ;
        RECT 455.400 379.050 456.450 416.100 ;
        RECT 458.400 391.050 459.450 430.950 ;
        RECT 479.400 420.450 480.450 457.950 ;
        RECT 487.950 452.100 490.050 454.200 ;
        RECT 488.400 451.350 489.600 452.100 ;
        RECT 482.100 448.950 484.200 451.050 ;
        RECT 488.100 448.950 490.200 451.050 ;
        RECT 503.400 439.050 504.450 457.950 ;
        RECT 506.400 454.200 507.450 484.800 ;
        RECT 514.950 472.950 517.050 475.050 ;
        RECT 505.950 452.100 508.050 454.200 ;
        RECT 511.950 449.100 514.050 451.200 ;
        RECT 512.400 448.350 513.600 449.100 ;
        RECT 506.400 445.950 508.500 448.050 ;
        RECT 511.800 445.950 513.900 448.050 ;
        RECT 506.400 443.400 507.600 445.650 ;
        RECT 484.950 436.950 487.050 439.050 ;
        RECT 502.950 436.950 505.050 439.050 ;
        RECT 476.400 419.400 480.450 420.450 ;
        RECT 466.950 416.100 469.050 418.200 ;
        RECT 467.400 415.350 468.600 416.100 ;
        RECT 463.950 412.950 466.050 415.050 ;
        RECT 466.950 412.950 469.050 415.050 ;
        RECT 464.400 411.900 465.600 412.650 ;
        RECT 463.950 409.800 466.050 411.900 ;
        RECT 457.950 388.950 460.050 391.050 ;
        RECT 454.950 376.950 457.050 379.050 ;
        RECT 448.950 371.100 451.050 373.200 ;
        RECT 455.400 372.600 456.450 376.950 ;
        RECT 449.400 370.350 450.600 371.100 ;
        RECT 455.400 370.350 456.600 372.600 ;
        RECT 430.950 367.950 433.050 370.050 ;
        RECT 433.950 367.950 436.050 370.050 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 442.950 367.950 445.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 424.950 364.800 427.050 366.900 ;
        RECT 434.400 365.400 435.600 367.650 ;
        RECT 427.950 346.950 430.050 349.050 ;
        RECT 428.400 346.050 429.450 346.950 ;
        RECT 424.950 343.950 429.450 346.050 ;
        RECT 434.400 345.450 435.450 365.400 ;
        RECT 443.400 345.450 444.450 367.950 ;
        RECT 452.400 365.400 453.600 367.650 ;
        RECT 458.400 366.900 459.600 367.650 ;
        RECT 452.400 349.050 453.450 365.400 ;
        RECT 457.950 364.800 460.050 366.900 ;
        RECT 464.400 358.050 465.450 409.800 ;
        RECT 466.950 382.950 469.050 385.050 ;
        RECT 467.400 366.900 468.450 382.950 ;
        RECT 476.400 372.600 477.450 419.400 ;
        RECT 485.400 418.200 486.450 436.950 ;
        RECT 499.950 433.950 502.050 436.050 ;
        RECT 500.400 418.200 501.450 433.950 ;
        RECT 506.400 424.050 507.450 443.400 ;
        RECT 515.400 442.050 516.450 472.950 ;
        RECT 518.400 463.050 519.450 488.400 ;
        RECT 520.950 487.800 523.050 489.900 ;
        RECT 526.950 487.800 529.050 489.900 ;
        RECT 527.400 478.050 528.450 487.800 ;
        RECT 532.950 478.950 535.050 481.050 ;
        RECT 526.950 475.950 529.050 478.050 ;
        RECT 533.400 469.050 534.450 478.950 ;
        RECT 532.950 466.950 535.050 469.050 ;
        RECT 517.950 460.950 520.050 463.050 ;
        RECT 532.950 457.950 535.050 460.050 ;
        RECT 523.950 454.950 526.050 457.050 ;
        RECT 514.950 439.950 517.050 442.050 ;
        RECT 505.950 421.950 508.050 424.050 ;
        RECT 484.950 416.100 487.050 418.200 ;
        RECT 499.950 416.100 502.050 418.200 ;
        RECT 515.400 417.600 516.450 439.950 ;
        RECT 485.400 415.350 486.600 416.100 ;
        RECT 500.400 415.350 501.600 416.100 ;
        RECT 515.400 415.350 516.600 417.600 ;
        RECT 479.100 412.950 481.200 415.050 ;
        RECT 484.500 412.950 486.600 415.050 ;
        RECT 487.800 412.950 489.900 415.050 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 515.400 412.950 517.500 415.050 ;
        RECT 520.800 412.950 522.900 415.050 ;
        RECT 479.400 411.900 480.600 412.650 ;
        RECT 478.950 409.800 481.050 411.900 ;
        RECT 488.400 410.400 489.600 412.650 ;
        RECT 503.400 410.400 504.600 412.650 ;
        RECT 521.400 411.000 522.600 412.650 ;
        RECT 488.400 373.200 489.450 410.400 ;
        RECT 503.400 403.050 504.450 410.400 ;
        RECT 520.950 406.950 523.050 411.000 ;
        RECT 524.400 403.050 525.450 454.950 ;
        RECT 533.400 450.600 534.450 457.950 ;
        RECT 533.400 448.350 534.600 450.600 ;
        RECT 527.400 445.950 529.500 448.050 ;
        RECT 532.800 445.950 534.900 448.050 ;
        RECT 527.400 444.900 528.600 445.650 ;
        RECT 526.950 442.800 529.050 444.900 ;
        RECT 536.400 436.050 537.450 508.950 ;
        RECT 547.950 494.100 550.050 496.200 ;
        RECT 548.400 493.350 549.600 494.100 ;
        RECT 544.950 490.950 547.050 493.050 ;
        RECT 547.950 490.950 550.050 493.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 545.400 489.900 546.600 490.650 ;
        RECT 544.950 487.800 547.050 489.900 ;
        RECT 551.400 488.400 552.600 490.650 ;
        RECT 551.400 484.050 552.450 488.400 ;
        RECT 541.950 481.950 544.050 484.050 ;
        RECT 550.950 481.950 553.050 484.050 ;
        RECT 538.950 463.950 541.050 466.050 ;
        RECT 535.950 435.450 538.050 436.050 ;
        RECT 533.400 434.400 538.050 435.450 ;
        RECT 529.950 418.950 532.050 421.050 ;
        RECT 502.950 400.950 505.050 403.050 ;
        RECT 508.950 400.950 511.050 403.050 ;
        RECT 523.950 400.950 526.050 403.050 ;
        RECT 505.950 385.950 508.050 388.050 ;
        RECT 476.400 370.350 477.600 372.600 ;
        RECT 481.950 371.100 484.050 373.200 ;
        RECT 487.950 371.100 490.050 373.200 ;
        RECT 493.950 371.100 496.050 373.200 ;
        RECT 499.950 371.100 502.050 373.200 ;
        RECT 482.400 370.350 483.600 371.100 ;
        RECT 494.400 370.350 495.600 371.100 ;
        RECT 500.400 370.350 501.600 371.100 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 473.400 366.900 474.600 367.650 ;
        RECT 479.400 366.900 480.600 367.650 ;
        RECT 466.950 364.800 469.050 366.900 ;
        RECT 472.950 364.800 475.050 366.900 ;
        RECT 478.950 364.800 481.050 366.900 ;
        RECT 497.400 365.400 498.600 367.650 ;
        RECT 463.950 355.950 466.050 358.050 ;
        RECT 451.950 346.950 454.050 349.050 ;
        RECT 497.400 346.050 498.450 365.400 ;
        RECT 434.400 344.400 438.450 345.450 ;
        RECT 407.400 337.350 408.600 338.100 ;
        RECT 413.400 337.350 414.600 338.100 ;
        RECT 418.950 337.950 421.050 340.050 ;
        RECT 421.950 337.950 424.050 340.050 ;
        RECT 428.400 339.600 429.450 343.950 ;
        RECT 403.950 334.950 406.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 409.950 334.950 412.050 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 404.400 332.400 405.600 334.650 ;
        RECT 410.400 333.000 411.600 334.650 ;
        RECT 397.950 328.950 400.050 331.050 ;
        RECT 404.400 328.050 405.450 332.400 ;
        RECT 409.950 328.950 412.050 333.000 ;
        RECT 415.950 331.950 418.050 334.050 ;
        RECT 403.950 325.950 406.050 328.050 ;
        RECT 416.400 325.050 417.450 331.950 ;
        RECT 397.950 322.950 400.050 325.050 ;
        RECT 415.950 322.950 418.050 325.050 ;
        RECT 391.950 295.950 394.050 298.050 ;
        RECT 398.400 294.600 399.450 322.950 ;
        RECT 416.400 298.050 417.450 322.950 ;
        RECT 419.400 319.050 420.450 337.950 ;
        RECT 428.400 337.350 429.600 339.600 ;
        RECT 433.950 339.000 436.050 343.050 ;
        RECT 437.400 340.050 438.450 344.400 ;
        RECT 440.400 344.400 444.450 345.450 ;
        RECT 434.400 337.350 435.600 339.000 ;
        RECT 436.950 337.950 439.050 340.050 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 425.400 333.900 426.600 334.650 ;
        RECT 424.950 331.800 427.050 333.900 ;
        RECT 431.400 332.400 432.600 334.650 ;
        RECT 431.400 328.050 432.450 332.400 ;
        RECT 430.950 325.950 433.050 328.050 ;
        RECT 418.950 316.950 421.050 319.050 ;
        RECT 418.950 310.950 421.050 313.050 ;
        RECT 389.400 293.400 393.450 294.450 ;
        RECT 380.400 292.350 381.600 293.100 ;
        RECT 386.400 292.350 387.600 293.100 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 376.950 286.950 379.050 289.050 ;
        RECT 383.400 288.900 384.600 289.650 ;
        RECT 373.950 280.950 376.050 283.050 ;
        RECT 377.400 280.050 378.450 286.950 ;
        RECT 382.950 286.800 385.050 288.900 ;
        RECT 376.950 277.950 379.050 280.050 ;
        RECT 370.950 274.950 373.050 277.050 ;
        RECT 370.950 271.800 373.050 273.900 ;
        RECT 371.400 268.050 372.450 271.800 ;
        RECT 383.400 271.050 384.450 286.800 ;
        RECT 382.950 268.950 385.050 271.050 ;
        RECT 370.950 265.950 373.050 268.050 ;
        RECT 392.400 267.450 393.450 293.400 ;
        RECT 398.400 292.350 399.600 294.600 ;
        RECT 403.950 293.100 406.050 298.050 ;
        RECT 415.950 295.950 418.050 298.050 ;
        RECT 419.400 294.600 420.450 310.950 ;
        RECT 404.400 292.350 405.600 293.100 ;
        RECT 419.400 292.350 420.600 294.600 ;
        RECT 424.950 293.100 427.050 295.200 ;
        RECT 425.400 292.350 426.600 293.100 ;
        RECT 397.950 289.950 400.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 401.400 288.900 402.600 289.650 ;
        RECT 416.400 288.900 417.600 289.650 ;
        RECT 400.950 286.800 403.050 288.900 ;
        RECT 415.950 286.800 418.050 288.900 ;
        RECT 422.400 287.400 423.600 289.650 ;
        RECT 431.400 289.050 432.450 325.950 ;
        RECT 440.400 307.050 441.450 344.400 ;
        RECT 454.950 343.950 457.050 346.050 ;
        RECT 472.950 343.950 475.050 346.050 ;
        RECT 487.950 343.950 490.050 346.050 ;
        RECT 496.800 343.950 498.900 346.050 ;
        RECT 499.950 345.450 502.050 346.050 ;
        RECT 499.950 344.400 504.450 345.450 ;
        RECT 499.950 343.950 502.050 344.400 ;
        RECT 442.950 340.950 445.050 343.050 ;
        RECT 443.400 313.050 444.450 340.950 ;
        RECT 448.950 339.000 451.050 343.050 ;
        RECT 455.400 339.600 456.450 343.950 ;
        RECT 449.400 337.350 450.600 339.000 ;
        RECT 455.400 337.350 456.600 339.600 ;
        RECT 463.950 338.100 466.050 340.200 ;
        RECT 473.400 339.600 474.450 343.950 ;
        RECT 448.950 334.950 451.050 337.050 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 452.400 332.400 453.600 334.650 ;
        RECT 458.400 333.000 459.600 334.650 ;
        RECT 452.400 319.050 453.450 332.400 ;
        RECT 457.950 328.950 460.050 333.000 ;
        RECT 451.950 316.950 454.050 319.050 ;
        RECT 442.950 310.950 445.050 313.050 ;
        RECT 439.950 304.950 442.050 307.050 ;
        RECT 451.950 304.950 454.050 307.050 ;
        RECT 457.950 304.950 460.050 307.050 ;
        RECT 442.950 298.950 445.050 301.050 ;
        RECT 443.400 294.600 444.450 298.950 ;
        RECT 443.400 292.350 444.600 294.600 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 415.950 277.950 418.050 280.050 ;
        RECT 392.400 265.200 393.600 267.450 ;
        RECT 361.950 259.950 364.050 262.050 ;
        RECT 367.950 261.000 370.050 265.050 ;
        RECT 368.400 259.350 369.600 261.000 ;
        RECT 373.950 259.950 376.050 262.050 ;
        RECT 387.900 261.900 390.000 263.700 ;
        RECT 391.800 262.800 393.900 264.900 ;
        RECT 395.100 264.300 397.200 266.400 ;
        RECT 386.400 260.700 395.100 261.900 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 347.400 244.050 348.450 253.800 ;
        RECT 352.950 250.950 355.050 255.000 ;
        RECT 358.950 253.800 361.050 255.900 ;
        RECT 365.400 254.400 366.600 256.650 ;
        RECT 365.400 253.050 366.450 254.400 ;
        RECT 361.950 251.400 366.450 253.050 ;
        RECT 361.950 250.950 366.000 251.400 ;
        RECT 319.950 241.950 322.050 244.050 ;
        RECT 346.950 241.950 349.050 244.050 ;
        RECT 320.400 238.050 321.450 241.950 ;
        RECT 319.950 235.950 322.050 238.050 ;
        RECT 340.950 229.950 343.050 232.050 ;
        RECT 313.950 220.950 316.050 223.050 ;
        RECT 334.950 220.950 337.050 223.050 ;
        RECT 311.400 214.350 312.600 216.600 ;
        RECT 316.950 216.000 319.050 220.050 ;
        RECT 335.400 216.600 336.450 220.950 ;
        RECT 341.400 216.600 342.450 229.950 ;
        RECT 317.400 214.350 318.600 216.000 ;
        RECT 335.400 214.350 336.600 216.600 ;
        RECT 341.400 214.350 342.600 216.600 ;
        RECT 346.950 214.950 349.050 217.050 ;
        RECT 361.950 215.100 364.050 217.200 ;
        RECT 374.400 216.450 375.450 259.950 ;
        RECT 383.100 256.950 385.200 259.050 ;
        RECT 383.400 255.450 384.600 256.650 ;
        RECT 380.400 254.400 384.600 255.450 ;
        RECT 380.400 232.050 381.450 254.400 ;
        RECT 386.400 251.700 387.300 260.700 ;
        RECT 393.000 259.800 395.100 260.700 ;
        RECT 396.000 258.900 396.900 264.300 ;
        RECT 416.400 261.600 417.450 277.950 ;
        RECT 422.400 274.050 423.450 287.400 ;
        RECT 430.950 286.950 433.050 289.050 ;
        RECT 440.400 288.900 441.600 289.650 ;
        RECT 439.950 286.800 442.050 288.900 ;
        RECT 430.950 280.950 433.050 283.050 ;
        RECT 421.950 271.950 424.050 274.050 ;
        RECT 398.400 261.450 399.600 261.600 ;
        RECT 398.400 260.400 402.450 261.450 ;
        RECT 398.400 259.350 399.600 260.400 ;
        RECT 390.000 257.700 396.900 258.900 ;
        RECT 390.000 255.300 390.900 257.700 ;
        RECT 388.800 253.200 390.900 255.300 ;
        RECT 391.800 253.950 393.900 256.050 ;
        RECT 385.500 249.600 387.600 251.700 ;
        RECT 392.400 251.400 393.600 253.650 ;
        RECT 395.700 250.500 396.900 257.700 ;
        RECT 397.800 256.950 399.900 259.050 ;
        RECT 395.100 248.400 397.200 250.500 ;
        RECT 401.400 250.050 402.450 260.400 ;
        RECT 416.400 259.350 417.600 261.600 ;
        RECT 421.950 260.100 424.050 262.200 ;
        RECT 422.400 259.350 423.600 260.100 ;
        RECT 412.950 256.950 415.050 259.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 419.400 254.400 420.600 256.650 ;
        RECT 431.400 255.450 432.450 280.950 ;
        RECT 452.400 273.450 453.450 304.950 ;
        RECT 458.400 294.600 459.450 304.950 ;
        RECT 464.400 298.050 465.450 338.100 ;
        RECT 473.400 337.350 474.600 339.600 ;
        RECT 478.950 338.100 481.050 340.200 ;
        RECT 479.400 337.350 480.600 338.100 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 466.950 328.950 469.050 334.050 ;
        RECT 476.400 333.000 477.600 334.650 ;
        RECT 475.950 330.450 478.050 333.000 ;
        RECT 482.400 332.400 483.600 334.650 ;
        RECT 475.950 329.400 480.450 330.450 ;
        RECT 475.950 328.950 478.050 329.400 ;
        RECT 466.950 316.950 469.050 319.050 ;
        RECT 463.950 295.950 466.050 298.050 ;
        RECT 458.400 292.350 459.600 294.600 ;
        RECT 464.400 294.450 465.600 294.600 ;
        RECT 467.400 294.450 468.450 316.950 ;
        RECT 469.950 307.950 472.050 310.050 ;
        RECT 464.400 293.400 468.450 294.450 ;
        RECT 464.400 292.350 465.600 293.400 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 449.400 272.400 453.450 273.450 ;
        RECT 461.400 287.400 462.600 289.650 ;
        RECT 436.950 260.100 439.050 262.200 ;
        RECT 445.950 260.100 448.050 262.200 ;
        RECT 437.400 259.350 438.600 260.100 ;
        RECT 434.100 256.950 436.200 259.050 ;
        RECT 437.400 256.950 439.500 259.050 ;
        RECT 442.800 256.950 444.900 259.050 ;
        RECT 434.400 255.450 435.600 256.650 ;
        RECT 431.400 254.400 435.600 255.450 ;
        RECT 443.400 254.400 444.600 256.650 ;
        RECT 400.950 247.950 403.050 250.050 ;
        RECT 419.400 244.050 420.450 254.400 ;
        RECT 424.950 247.950 427.050 250.050 ;
        RECT 418.950 241.950 421.050 244.050 ;
        RECT 421.950 232.950 424.050 235.050 ;
        RECT 379.950 229.950 382.050 232.050 ;
        RECT 418.950 229.950 421.050 232.050 ;
        RECT 371.400 215.400 375.450 216.450 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 314.400 210.900 315.600 211.650 ;
        RECT 313.950 208.800 316.050 210.900 ;
        RECT 320.400 209.400 321.600 211.650 ;
        RECT 304.950 202.950 307.050 205.050 ;
        RECT 313.950 202.950 316.050 205.050 ;
        RECT 301.950 190.950 304.050 193.050 ;
        RECT 286.950 187.950 289.050 190.050 ;
        RECT 298.950 187.950 301.050 190.050 ;
        RECT 257.400 181.350 258.600 182.100 ;
        RECT 263.400 181.350 264.600 183.600 ;
        RECT 268.950 181.950 271.050 184.050 ;
        RECT 277.950 182.100 280.050 184.200 ;
        RECT 278.400 181.350 279.600 182.100 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 260.400 176.400 261.600 178.650 ;
        RECT 260.400 148.050 261.450 176.400 ;
        RECT 265.950 175.950 268.050 178.050 ;
        RECT 268.950 177.450 271.050 180.900 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 277.950 178.950 280.050 181.050 ;
        RECT 280.950 178.950 283.050 181.050 ;
        RECT 275.400 177.450 276.600 178.650 ;
        RECT 281.400 177.900 282.600 178.650 ;
        RECT 287.400 177.900 288.450 187.950 ;
        RECT 292.950 182.100 295.050 184.200 ;
        RECT 293.400 181.350 294.600 182.100 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 296.400 178.050 297.600 178.650 ;
        RECT 268.950 177.000 276.600 177.450 ;
        RECT 269.400 176.400 276.600 177.000 ;
        RECT 266.400 169.050 267.450 175.950 ;
        RECT 280.950 175.800 283.050 177.900 ;
        RECT 286.950 175.800 289.050 177.900 ;
        RECT 296.400 176.400 301.050 178.050 ;
        RECT 302.400 177.900 303.450 190.950 ;
        RECT 304.950 183.600 309.000 184.050 ;
        RECT 314.400 183.600 315.450 202.950 ;
        RECT 320.400 184.050 321.450 209.400 ;
        RECT 325.950 208.800 328.050 210.900 ;
        RECT 332.400 209.400 333.600 211.650 ;
        RECT 338.400 210.900 339.600 211.650 ;
        RECT 347.400 211.050 348.450 214.950 ;
        RECT 362.400 214.350 363.600 215.100 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 364.950 211.950 367.050 214.050 ;
        RECT 304.950 181.950 309.600 183.600 ;
        RECT 308.400 181.350 309.600 181.950 ;
        RECT 314.400 181.350 315.600 183.600 ;
        RECT 319.950 181.950 322.050 184.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 311.400 177.900 312.600 178.650 ;
        RECT 297.000 175.950 301.050 176.400 ;
        RECT 301.950 175.800 304.050 177.900 ;
        RECT 310.950 175.800 313.050 177.900 ;
        RECT 268.950 172.950 271.050 175.050 ;
        RECT 265.950 166.950 268.050 169.050 ;
        RECT 259.950 145.950 262.050 148.050 ;
        RECT 269.400 145.050 270.450 172.950 ;
        RECT 323.400 172.050 324.450 178.950 ;
        RECT 322.950 169.950 325.050 172.050 ;
        RECT 283.950 145.950 286.050 148.050 ;
        RECT 322.950 147.450 325.050 148.050 ;
        RECT 326.400 147.450 327.450 208.800 ;
        RECT 332.400 186.450 333.450 209.400 ;
        RECT 337.950 208.800 340.050 210.900 ;
        RECT 346.950 208.950 349.050 211.050 ;
        RECT 359.400 210.900 360.600 211.650 ;
        RECT 358.950 208.800 361.050 210.900 ;
        RECT 365.400 210.000 366.600 211.650 ;
        RECT 364.950 205.950 367.050 210.000 ;
        RECT 365.400 202.050 366.450 205.950 ;
        RECT 337.950 199.950 340.050 202.050 ;
        RECT 364.950 199.950 367.050 202.050 ;
        RECT 329.400 185.400 333.450 186.450 ;
        RECT 329.400 151.050 330.450 185.400 ;
        RECT 338.400 183.600 339.450 199.950 ;
        RECT 355.950 193.950 358.050 196.050 ;
        RECT 338.400 181.350 339.600 183.600 ;
        RECT 346.950 182.100 349.050 184.200 ;
        RECT 352.950 182.100 355.050 184.200 ;
        RECT 347.400 181.350 348.600 182.100 ;
        RECT 332.400 178.950 334.500 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 340.950 178.950 343.050 181.050 ;
        RECT 347.100 178.950 349.200 181.050 ;
        RECT 332.400 177.900 333.600 178.650 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 341.400 176.400 342.600 178.650 ;
        RECT 334.950 172.950 337.050 175.050 ;
        RECT 331.950 169.950 334.050 172.050 ;
        RECT 328.950 148.950 331.050 151.050 ;
        RECT 322.950 146.400 327.450 147.450 ;
        RECT 322.950 145.950 325.050 146.400 ;
        RECT 268.950 142.950 271.050 145.050 ;
        RECT 256.950 137.100 259.050 139.200 ;
        RECT 269.400 138.450 270.450 142.950 ;
        RECT 266.400 137.400 270.450 138.450 ;
        RECT 257.400 136.350 258.600 137.100 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 260.400 132.000 261.600 133.650 ;
        RECT 266.400 132.900 267.450 137.400 ;
        RECT 271.950 137.100 274.050 139.200 ;
        RECT 277.950 137.100 280.050 139.200 ;
        RECT 284.400 138.600 285.450 145.950 ;
        RECT 313.950 139.950 316.050 142.050 ;
        RECT 272.400 136.350 273.600 137.100 ;
        RECT 278.400 136.350 279.600 137.100 ;
        RECT 284.400 136.350 285.600 138.600 ;
        RECT 289.950 137.100 292.050 139.200 ;
        RECT 295.950 137.100 298.050 139.200 ;
        RECT 301.950 137.100 304.050 139.200 ;
        RECT 310.950 137.100 313.050 139.200 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 274.950 133.950 277.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 275.400 132.900 276.600 133.650 ;
        RECT 250.950 127.950 253.050 130.050 ;
        RECT 259.950 129.450 262.050 132.000 ;
        RECT 265.950 130.800 268.050 132.900 ;
        RECT 274.950 130.800 277.050 132.900 ;
        RECT 281.400 131.400 282.600 133.650 ;
        RECT 290.400 132.450 291.450 137.100 ;
        RECT 296.400 136.350 297.600 137.100 ;
        RECT 302.400 136.350 303.600 137.100 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 299.400 132.900 300.600 133.650 ;
        RECT 305.400 132.900 306.600 133.650 ;
        RECT 290.400 131.400 294.450 132.450 ;
        RECT 257.400 128.400 262.050 129.450 ;
        RECT 251.400 124.050 252.450 127.950 ;
        RECT 250.950 121.950 253.050 124.050 ;
        RECT 250.950 112.950 253.050 115.050 ;
        RECT 247.950 106.950 250.050 109.050 ;
        RECT 251.400 105.600 252.450 112.950 ;
        RECT 257.400 106.050 258.450 128.400 ;
        RECT 259.950 127.950 262.050 128.400 ;
        RECT 266.400 111.450 267.450 130.800 ;
        RECT 281.400 124.050 282.450 131.400 ;
        RECT 280.950 121.950 283.050 124.050 ;
        RECT 293.400 120.450 294.450 131.400 ;
        RECT 298.950 130.800 301.050 132.900 ;
        RECT 304.950 130.800 307.050 132.900 ;
        RECT 293.400 119.400 297.450 120.450 ;
        RECT 266.400 110.400 270.450 111.450 ;
        RECT 259.950 106.950 262.050 109.050 ;
        RECT 239.400 88.050 240.450 103.950 ;
        RECT 245.400 103.350 246.600 105.600 ;
        RECT 251.400 103.350 252.600 105.600 ;
        RECT 256.950 103.950 259.050 106.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 248.400 99.000 249.600 100.650 ;
        RECT 254.400 99.900 255.600 100.650 ;
        RECT 247.950 94.950 250.050 99.000 ;
        RECT 253.950 97.800 256.050 99.900 ;
        RECT 238.950 85.950 241.050 88.050 ;
        RECT 260.400 67.050 261.450 106.950 ;
        RECT 269.400 105.600 270.450 110.400 ;
        RECT 269.400 103.350 270.600 105.600 ;
        RECT 274.950 103.950 277.050 106.050 ;
        RECT 283.950 105.000 286.050 109.050 ;
        RECT 292.950 106.950 295.050 109.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 266.400 99.000 267.600 100.650 ;
        RECT 265.950 94.950 268.050 99.000 ;
        RECT 271.950 88.950 274.050 91.050 ;
        RECT 259.950 64.950 262.050 67.050 ;
        RECT 235.950 61.950 238.050 64.050 ;
        RECT 272.400 61.200 273.450 88.950 ;
        RECT 275.400 79.050 276.450 103.950 ;
        RECT 284.400 103.350 285.600 105.000 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 281.400 98.400 282.600 100.650 ;
        RECT 287.400 98.400 288.600 100.650 ;
        RECT 281.400 97.050 282.450 98.400 ;
        RECT 280.950 94.950 283.050 97.050 ;
        RECT 274.950 76.950 277.050 79.050 ;
        RECT 218.400 58.350 219.600 60.000 ;
        RECT 224.400 58.350 225.600 60.600 ;
        RECT 241.950 59.100 244.050 61.200 ;
        RECT 248.400 60.450 249.600 60.600 ;
        RECT 248.400 59.400 255.450 60.450 ;
        RECT 242.400 58.350 243.600 59.100 ;
        RECT 248.400 58.350 249.600 59.400 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 220.950 55.950 223.050 58.050 ;
        RECT 223.950 55.950 226.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 221.400 54.900 222.600 55.650 ;
        RECT 227.400 54.900 228.600 55.650 ;
        RECT 193.950 52.800 196.050 54.900 ;
        RECT 199.950 52.800 202.050 54.900 ;
        RECT 211.950 52.800 214.050 54.900 ;
        RECT 220.950 52.800 223.050 54.900 ;
        RECT 226.950 52.800 229.050 54.900 ;
        RECT 232.950 54.450 235.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 239.400 54.900 240.600 55.650 ;
        RECT 230.400 54.000 235.050 54.450 ;
        RECT 230.400 53.400 234.450 54.000 ;
        RECT 184.950 43.950 187.050 46.050 ;
        RECT 194.400 34.050 195.450 52.800 ;
        RECT 208.950 49.950 211.050 52.050 ;
        RECT 223.950 49.950 226.050 52.050 ;
        RECT 209.400 46.050 210.450 49.950 ;
        RECT 208.950 43.950 211.050 46.050 ;
        RECT 214.950 43.950 217.050 46.050 ;
        RECT 196.950 37.950 199.050 40.050 ;
        RECT 193.950 31.950 196.050 34.050 ;
        RECT 176.400 25.350 177.600 26.100 ;
        RECT 182.400 25.350 183.600 27.600 ;
        RECT 187.950 26.100 190.050 28.200 ;
        RECT 197.400 27.600 198.450 37.950 ;
        RECT 211.950 31.950 214.050 34.050 ;
        RECT 212.400 27.600 213.450 31.950 ;
        RECT 215.400 31.050 216.450 43.950 ;
        RECT 224.400 37.050 225.450 49.950 ;
        RECT 227.400 40.050 228.450 52.800 ;
        RECT 230.400 49.050 231.450 53.400 ;
        RECT 238.950 52.800 241.050 54.900 ;
        RECT 245.400 54.000 246.600 55.650 ;
        RECT 254.400 55.050 255.450 59.400 ;
        RECT 256.950 59.100 259.050 61.200 ;
        RECT 265.950 59.100 268.050 61.200 ;
        RECT 271.950 59.100 274.050 61.200 ;
        RECT 244.950 49.950 247.050 54.000 ;
        RECT 253.950 52.950 256.050 55.050 ;
        RECT 229.950 46.950 232.050 49.050 ;
        RECT 235.950 46.950 238.050 49.050 ;
        RECT 226.950 37.950 229.050 40.050 ;
        RECT 223.950 34.950 226.050 37.050 ;
        RECT 227.400 34.050 228.450 37.950 ;
        RECT 229.950 34.950 232.050 37.050 ;
        RECT 226.950 31.950 229.050 34.050 ;
        RECT 214.950 28.950 217.050 31.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 181.950 22.950 184.050 25.050 ;
        RECT 173.400 21.900 174.600 22.650 ;
        RECT 145.950 16.950 148.050 19.050 ;
        RECT 149.400 16.050 150.450 20.400 ;
        RECT 85.950 13.950 88.050 16.050 ;
        RECT 112.950 13.950 115.050 16.050 ;
        RECT 127.950 13.950 130.050 16.050 ;
        RECT 148.950 13.950 151.050 16.050 ;
        RECT 113.400 7.050 114.450 13.950 ;
        RECT 158.400 7.050 159.450 20.400 ;
        RECT 163.950 19.800 166.050 21.900 ;
        RECT 172.950 19.800 175.050 21.900 ;
        RECT 179.400 20.400 180.600 22.650 ;
        RECT 188.400 22.050 189.450 26.100 ;
        RECT 197.400 25.350 198.600 27.600 ;
        RECT 212.400 25.350 213.600 27.600 ;
        RECT 217.950 26.100 220.050 28.200 ;
        RECT 218.400 25.350 219.600 26.100 ;
        RECT 223.950 25.950 226.050 28.050 ;
        RECT 230.400 27.450 231.450 34.950 ;
        RECT 232.950 31.950 235.050 34.050 ;
        RECT 227.400 26.400 231.450 27.450 ;
        RECT 233.400 27.600 234.450 31.950 ;
        RECT 236.400 31.050 237.450 46.950 ;
        RECT 254.400 46.050 255.450 52.950 ;
        RECT 257.400 52.050 258.450 59.100 ;
        RECT 266.400 58.350 267.600 59.100 ;
        RECT 272.400 58.350 273.600 59.100 ;
        RECT 277.950 58.950 280.050 61.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 263.400 53.400 264.600 55.650 ;
        RECT 269.400 53.400 270.600 55.650 ;
        RECT 256.950 49.950 259.050 52.050 ;
        RECT 253.950 43.950 256.050 46.050 ;
        RECT 263.400 40.050 264.450 53.400 ;
        RECT 269.400 49.050 270.450 53.400 ;
        RECT 268.950 46.950 271.050 49.050 ;
        RECT 262.950 37.950 265.050 40.050 ;
        RECT 235.950 28.950 238.050 31.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 179.400 16.050 180.450 20.400 ;
        RECT 187.950 19.950 190.050 22.050 ;
        RECT 194.400 21.900 195.600 22.650 ;
        RECT 209.400 21.900 210.600 22.650 ;
        RECT 215.400 21.900 216.600 22.650 ;
        RECT 193.950 19.800 196.050 21.900 ;
        RECT 208.950 19.800 211.050 21.900 ;
        RECT 214.950 19.800 217.050 21.900 ;
        RECT 178.950 13.950 181.050 16.050 ;
        RECT 224.400 13.050 225.450 25.950 ;
        RECT 227.400 21.900 228.450 26.400 ;
        RECT 233.400 25.350 234.600 27.600 ;
        RECT 238.950 26.100 241.050 28.200 ;
        RECT 256.950 26.100 259.050 28.200 ;
        RECT 262.950 26.100 265.050 28.200 ;
        RECT 278.400 27.600 279.450 58.950 ;
        RECT 281.400 31.050 282.450 94.950 ;
        RECT 287.400 94.050 288.450 98.400 ;
        RECT 293.400 97.050 294.450 106.950 ;
        RECT 296.400 97.050 297.450 119.400 ;
        RECT 299.400 106.050 300.450 130.800 ;
        RECT 311.400 124.050 312.450 137.100 ;
        RECT 314.400 133.050 315.450 139.950 ;
        RECT 323.400 138.600 324.450 145.950 ;
        RECT 323.400 136.350 324.600 138.600 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 325.950 133.950 328.050 136.050 ;
        RECT 313.950 130.950 316.050 133.050 ;
        RECT 320.400 131.400 321.600 133.650 ;
        RECT 326.400 131.400 327.600 133.650 ;
        RECT 316.950 124.950 319.050 127.050 ;
        RECT 310.950 121.950 313.050 124.050 ;
        RECT 317.400 106.200 318.450 124.950 ;
        RECT 320.400 121.050 321.450 131.400 ;
        RECT 326.400 127.050 327.450 131.400 ;
        RECT 325.950 124.950 328.050 127.050 ;
        RECT 319.950 118.950 322.050 121.050 ;
        RECT 328.950 120.450 331.050 121.050 ;
        RECT 332.400 120.450 333.450 169.950 ;
        RECT 335.400 127.050 336.450 172.950 ;
        RECT 341.400 172.050 342.450 176.400 ;
        RECT 353.400 175.050 354.450 182.100 ;
        RECT 352.950 172.950 355.050 175.050 ;
        RECT 340.950 169.950 343.050 172.050 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 340.950 138.000 343.050 142.050 ;
        RECT 347.400 138.600 348.450 163.950 ;
        RECT 341.400 136.350 342.600 138.000 ;
        RECT 347.400 136.350 348.600 138.600 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 343.950 133.950 346.050 136.050 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 344.400 131.400 345.600 133.650 ;
        RECT 350.400 132.450 351.600 133.650 ;
        RECT 356.400 132.450 357.450 193.950 ;
        RECT 371.400 193.050 372.450 215.400 ;
        RECT 379.950 215.100 382.050 217.200 ;
        RECT 397.950 215.100 400.050 217.200 ;
        RECT 403.950 215.100 406.050 217.200 ;
        RECT 409.950 215.100 412.050 217.200 ;
        RECT 419.400 216.600 420.450 229.950 ;
        RECT 422.400 223.050 423.450 232.950 ;
        RECT 425.400 229.050 426.450 247.950 ;
        RECT 443.400 244.050 444.450 254.400 ;
        RECT 446.400 247.050 447.450 260.100 ;
        RECT 445.950 244.950 448.050 247.050 ;
        RECT 442.950 241.950 445.050 244.050 ;
        RECT 449.400 241.050 450.450 272.400 ;
        RECT 461.400 271.050 462.450 287.400 ;
        RECT 466.950 271.950 469.050 274.050 ;
        RECT 451.950 268.950 454.050 271.050 ;
        RECT 460.950 268.950 463.050 271.050 ;
        RECT 448.950 238.950 451.050 241.050 ;
        RECT 424.950 226.950 427.050 229.050 ;
        RECT 421.950 220.950 424.050 223.050 ;
        RECT 425.400 216.600 426.450 226.950 ;
        RECT 439.950 223.950 442.050 226.050 ;
        RECT 430.950 220.950 433.050 223.050 ;
        RECT 380.400 214.350 381.600 215.100 ;
        RECT 398.400 214.350 399.600 215.100 ;
        RECT 404.400 214.350 405.600 215.100 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 382.950 211.950 385.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 400.950 211.950 403.050 214.050 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 377.400 209.400 378.600 211.650 ;
        RECT 383.400 209.400 384.600 211.650 ;
        RECT 377.400 202.050 378.450 209.400 ;
        RECT 376.950 201.450 379.050 202.050 ;
        RECT 376.950 200.400 381.450 201.450 ;
        RECT 376.950 199.950 379.050 200.400 ;
        RECT 364.950 190.950 367.050 193.050 ;
        RECT 370.950 190.950 373.050 193.050 ;
        RECT 365.400 183.600 366.450 190.950 ;
        RECT 365.400 181.350 366.600 183.600 ;
        RECT 370.950 182.100 373.050 184.200 ;
        RECT 371.400 181.350 372.600 182.100 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 367.950 178.950 370.050 181.050 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 373.950 178.950 376.050 181.050 ;
        RECT 368.400 176.400 369.600 178.650 ;
        RECT 374.400 177.900 375.600 178.650 ;
        RECT 380.400 177.900 381.450 200.400 ;
        RECT 383.400 184.200 384.450 209.400 ;
        RECT 391.950 208.950 394.050 211.050 ;
        RECT 395.400 210.000 396.600 211.650 ;
        RECT 392.400 184.200 393.450 208.950 ;
        RECT 394.950 205.950 397.050 210.000 ;
        RECT 401.400 209.400 402.600 211.650 ;
        RECT 410.400 211.050 411.450 215.100 ;
        RECT 419.400 214.350 420.600 216.600 ;
        RECT 425.400 214.350 426.600 216.600 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 397.950 190.950 400.050 193.050 ;
        RECT 382.950 182.100 385.050 184.200 ;
        RECT 391.950 182.100 394.050 184.200 ;
        RECT 368.400 175.050 369.450 176.400 ;
        RECT 373.950 175.800 376.050 177.900 ;
        RECT 379.950 175.800 382.050 177.900 ;
        RECT 383.400 175.050 384.450 182.100 ;
        RECT 392.400 181.350 393.600 182.100 ;
        RECT 388.950 178.950 391.050 181.050 ;
        RECT 391.950 178.950 394.050 181.050 ;
        RECT 389.400 177.000 390.600 178.650 ;
        RECT 367.950 172.950 370.050 175.050 ;
        RECT 382.950 172.950 385.050 175.050 ;
        RECT 388.950 172.950 391.050 177.000 ;
        RECT 364.950 169.950 367.050 172.050 ;
        RECT 365.400 138.600 366.450 169.950 ;
        RECT 368.400 139.050 369.450 172.950 ;
        RECT 398.400 157.050 399.450 190.950 ;
        RECT 401.400 184.050 402.450 209.400 ;
        RECT 409.950 208.950 412.050 211.050 ;
        RECT 416.400 210.900 417.600 211.650 ;
        RECT 415.950 208.800 418.050 210.900 ;
        RECT 422.400 210.000 423.600 211.650 ;
        RECT 431.400 210.900 432.450 220.950 ;
        RECT 440.400 216.600 441.450 223.950 ;
        RECT 452.400 217.200 453.450 268.950 ;
        RECT 457.950 260.100 460.050 262.200 ;
        RECT 458.400 259.350 459.600 260.100 ;
        RECT 455.100 256.950 457.200 259.050 ;
        RECT 458.400 256.950 460.500 259.050 ;
        RECT 463.800 256.950 465.900 259.050 ;
        RECT 455.400 254.400 456.600 256.650 ;
        RECT 464.400 255.450 465.600 256.650 ;
        RECT 467.400 255.450 468.450 271.950 ;
        RECT 470.400 262.200 471.450 307.950 ;
        RECT 472.950 295.950 475.050 298.050 ;
        RECT 473.400 288.900 474.450 295.950 ;
        RECT 479.400 295.200 480.450 329.400 ;
        RECT 482.400 301.050 483.450 332.400 ;
        RECT 481.950 298.950 484.050 301.050 ;
        RECT 484.950 298.950 487.050 301.050 ;
        RECT 478.950 293.100 481.050 295.200 ;
        RECT 485.400 294.600 486.450 298.950 ;
        RECT 488.400 298.050 489.450 343.950 ;
        RECT 493.950 338.100 496.050 340.200 ;
        RECT 500.400 339.600 501.450 343.950 ;
        RECT 503.400 340.050 504.450 344.400 ;
        RECT 506.400 340.200 507.450 385.950 ;
        RECT 509.400 363.450 510.450 400.950 ;
        RECT 520.950 382.950 523.050 385.050 ;
        RECT 511.950 371.100 514.050 373.200 ;
        RECT 521.400 372.600 522.450 382.950 ;
        RECT 521.400 372.450 522.600 372.600 ;
        RECT 521.400 371.400 525.450 372.450 ;
        RECT 512.400 370.350 513.600 371.100 ;
        RECT 521.400 370.350 522.600 371.400 ;
        RECT 512.100 367.950 514.200 370.050 ;
        RECT 515.400 367.950 517.500 370.050 ;
        RECT 520.800 367.950 522.900 370.050 ;
        RECT 515.400 365.400 516.600 367.650 ;
        RECT 509.400 362.400 513.450 363.450 ;
        RECT 494.400 337.350 495.600 338.100 ;
        RECT 500.400 337.350 501.600 339.600 ;
        RECT 502.950 337.950 505.050 340.050 ;
        RECT 505.950 338.100 508.050 340.200 ;
        RECT 512.400 339.450 513.450 362.400 ;
        RECT 515.400 361.050 516.450 365.400 ;
        RECT 514.950 358.950 517.050 361.050 ;
        RECT 524.400 352.050 525.450 371.400 ;
        RECT 526.950 364.950 529.050 367.050 ;
        RECT 523.950 349.950 526.050 352.050 ;
        RECT 527.400 346.050 528.450 364.950 ;
        RECT 517.950 343.950 520.050 346.050 ;
        RECT 526.950 343.950 529.050 346.050 ;
        RECT 509.400 339.000 513.450 339.450 ;
        RECT 508.950 338.400 513.450 339.000 ;
        RECT 518.400 339.600 519.450 343.950 ;
        RECT 526.950 340.800 529.050 342.900 ;
        RECT 493.950 334.950 496.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 497.400 333.900 498.600 334.650 ;
        RECT 496.950 331.800 499.050 333.900 ;
        RECT 502.950 331.950 505.050 334.050 ;
        RECT 503.400 310.050 504.450 331.950 ;
        RECT 502.950 307.950 505.050 310.050 ;
        RECT 506.400 301.050 507.450 338.100 ;
        RECT 508.950 334.950 511.050 338.400 ;
        RECT 518.400 337.350 519.600 339.600 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 508.950 331.800 511.050 333.900 ;
        RECT 515.400 332.400 516.600 334.650 ;
        RECT 521.400 334.050 522.600 334.650 ;
        RECT 521.400 332.400 526.050 334.050 ;
        RECT 496.950 298.950 499.050 301.050 ;
        RECT 505.950 298.950 508.050 301.050 ;
        RECT 487.950 295.950 490.050 298.050 ;
        RECT 493.950 295.950 496.050 298.050 ;
        RECT 479.400 292.350 480.600 293.100 ;
        RECT 485.400 292.350 486.600 294.600 ;
        RECT 478.950 289.950 481.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 482.400 288.900 483.600 289.650 ;
        RECT 488.400 289.050 489.600 289.650 ;
        RECT 472.950 286.800 475.050 288.900 ;
        RECT 481.950 286.800 484.050 288.900 ;
        RECT 488.400 287.400 493.050 289.050 ;
        RECT 489.000 286.950 493.050 287.400 ;
        RECT 478.950 265.950 481.050 268.050 ;
        RECT 469.950 260.100 472.050 262.200 ;
        RECT 479.400 261.600 480.450 265.950 ;
        RECT 479.400 259.350 480.600 261.600 ;
        RECT 484.950 260.100 487.050 262.200 ;
        RECT 494.400 261.450 495.450 295.950 ;
        RECT 497.400 288.900 498.450 298.950 ;
        RECT 499.950 292.950 502.050 298.050 ;
        RECT 509.400 297.450 510.450 331.800 ;
        RECT 515.400 330.450 516.450 332.400 ;
        RECT 522.000 331.950 526.050 332.400 ;
        RECT 515.400 329.400 519.450 330.450 ;
        RECT 511.950 310.950 514.050 313.050 ;
        RECT 506.400 296.400 510.450 297.450 ;
        RECT 506.400 294.600 507.450 296.400 ;
        RECT 512.400 294.600 513.450 310.950 ;
        RECT 518.400 304.050 519.450 329.400 ;
        RECT 517.950 301.950 520.050 304.050 ;
        RECT 523.950 295.950 526.050 298.050 ;
        RECT 506.400 292.350 507.600 294.600 ;
        RECT 512.400 292.350 513.600 294.600 ;
        RECT 520.950 292.950 523.050 295.050 ;
        RECT 502.950 289.950 505.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 508.950 289.950 511.050 292.050 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 514.950 289.950 517.050 292.050 ;
        RECT 503.400 288.900 504.600 289.650 ;
        RECT 496.950 286.800 499.050 288.900 ;
        RECT 502.950 286.800 505.050 288.900 ;
        RECT 509.400 287.400 510.600 289.650 ;
        RECT 515.400 288.900 516.600 289.650 ;
        RECT 509.400 277.050 510.450 287.400 ;
        RECT 514.950 286.800 517.050 288.900 ;
        RECT 517.950 286.950 520.050 289.050 ;
        RECT 521.400 288.900 522.450 292.950 ;
        RECT 508.950 274.950 511.050 277.050 ;
        RECT 491.400 260.400 495.450 261.450 ;
        RECT 485.400 259.350 486.600 260.100 ;
        RECT 478.950 256.950 481.050 259.050 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 482.400 255.900 483.600 256.650 ;
        RECT 464.400 254.400 468.450 255.450 ;
        RECT 455.400 226.050 456.450 254.400 ;
        RECT 463.950 244.950 466.050 247.050 ;
        RECT 454.950 223.950 457.050 226.050 ;
        RECT 440.400 214.350 441.600 216.600 ;
        RECT 445.950 215.100 448.050 217.200 ;
        RECT 451.950 215.100 454.050 217.200 ;
        RECT 464.400 217.050 465.450 244.950 ;
        RECT 454.950 216.600 459.000 217.050 ;
        RECT 446.400 214.350 447.600 215.100 ;
        RECT 436.950 211.950 439.050 214.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 437.400 210.900 438.600 211.650 ;
        RECT 421.950 205.950 424.050 210.000 ;
        RECT 430.950 208.800 433.050 210.900 ;
        RECT 436.950 208.800 439.050 210.900 ;
        RECT 443.400 209.400 444.600 211.650 ;
        RECT 452.400 210.900 453.450 215.100 ;
        RECT 454.950 214.950 459.600 216.600 ;
        RECT 463.950 214.950 466.050 217.050 ;
        RECT 458.400 214.350 459.600 214.950 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 439.950 205.950 442.050 208.050 ;
        RECT 406.950 199.950 409.050 202.050 ;
        RECT 400.950 181.950 403.050 184.050 ;
        RECT 407.400 183.600 408.450 199.950 ;
        RECT 412.950 193.950 415.050 196.050 ;
        RECT 413.400 183.600 414.450 193.950 ;
        RECT 421.950 190.950 424.050 193.050 ;
        RECT 418.950 187.950 421.050 190.050 ;
        RECT 407.400 181.350 408.600 183.600 ;
        RECT 413.400 181.350 414.600 183.600 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 404.400 177.900 405.600 178.650 ;
        RECT 410.400 177.900 411.600 178.650 ;
        RECT 403.950 175.800 406.050 177.900 ;
        RECT 409.950 175.800 412.050 177.900 ;
        RECT 404.400 172.050 405.450 175.800 ;
        RECT 403.950 169.950 406.050 172.050 ;
        RECT 410.400 166.050 411.450 175.800 ;
        RECT 409.950 163.950 412.050 166.050 ;
        RECT 397.950 154.950 400.050 157.050 ;
        RECT 412.950 154.950 415.050 157.050 ;
        RECT 398.400 148.050 399.450 154.950 ;
        RECT 400.950 148.950 403.050 151.050 ;
        RECT 370.950 145.950 373.050 148.050 ;
        RECT 376.950 145.950 379.050 148.050 ;
        RECT 397.950 145.950 400.050 148.050 ;
        RECT 365.400 136.350 366.600 138.600 ;
        RECT 367.950 136.950 370.050 139.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 350.400 131.400 357.450 132.450 ;
        RECT 358.800 132.000 360.900 133.050 ;
        RECT 362.400 132.900 363.600 133.650 ;
        RECT 334.950 124.950 337.050 127.050 ;
        RECT 328.950 119.400 333.450 120.450 ;
        RECT 328.950 118.950 331.050 119.400 ;
        RECT 298.950 103.950 301.050 106.050 ;
        RECT 304.950 104.100 307.050 106.200 ;
        RECT 310.950 104.100 313.050 106.200 ;
        RECT 316.950 104.100 319.050 106.200 ;
        RECT 305.400 103.350 306.600 104.100 ;
        RECT 311.400 103.350 312.600 104.100 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 302.400 99.000 303.600 100.650 ;
        RECT 308.400 99.900 309.600 100.650 ;
        RECT 292.950 94.950 295.050 97.050 ;
        RECT 295.950 94.950 298.050 97.050 ;
        RECT 299.400 94.050 300.450 97.950 ;
        RECT 301.950 94.950 304.050 99.000 ;
        RECT 307.950 97.800 310.050 99.900 ;
        RECT 286.950 91.950 289.050 94.050 ;
        RECT 298.950 91.950 301.050 94.050 ;
        RECT 286.950 67.950 289.050 70.050 ;
        RECT 287.400 60.600 288.450 67.950 ;
        RECT 287.400 58.350 288.600 60.600 ;
        RECT 292.950 59.100 295.050 61.200 ;
        RECT 293.400 58.350 294.600 59.100 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 283.950 52.950 286.050 55.050 ;
        RECT 290.400 54.900 291.600 55.650 ;
        RECT 299.400 55.050 300.450 91.950 ;
        RECT 307.950 67.950 310.050 70.050 ;
        RECT 301.950 59.100 304.050 61.200 ;
        RECT 308.400 60.600 309.450 67.950 ;
        RECT 302.400 55.050 303.450 59.100 ;
        RECT 308.400 58.350 309.600 60.600 ;
        RECT 313.950 59.100 316.050 61.200 ;
        RECT 317.400 61.050 318.450 104.100 ;
        RECT 320.400 99.900 321.450 118.950 ;
        RECT 329.400 105.600 330.450 118.950 ;
        RECT 344.400 118.050 345.450 131.400 ;
        RECT 358.800 130.950 361.050 132.000 ;
        RECT 358.950 129.450 361.050 130.950 ;
        RECT 361.950 130.800 364.050 132.900 ;
        RECT 356.400 129.000 361.050 129.450 ;
        RECT 356.400 128.400 360.450 129.000 ;
        RECT 343.950 115.950 346.050 118.050 ;
        RECT 352.950 112.950 355.050 115.050 ;
        RECT 329.400 103.350 330.600 105.600 ;
        RECT 337.950 104.100 340.050 106.200 ;
        RECT 343.950 104.100 346.050 106.200 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 328.950 100.950 331.050 103.050 ;
        RECT 331.950 100.950 334.050 103.050 ;
        RECT 319.950 97.800 322.050 99.900 ;
        RECT 326.400 99.000 327.600 100.650 ;
        RECT 325.950 94.950 328.050 99.000 ;
        RECT 332.400 98.400 333.600 100.650 ;
        RECT 332.400 94.050 333.450 98.400 ;
        RECT 319.950 91.950 322.050 94.050 ;
        RECT 331.950 91.950 334.050 94.050 ;
        RECT 314.400 58.350 315.600 59.100 ;
        RECT 316.950 58.950 319.050 61.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 284.400 34.050 285.450 52.950 ;
        RECT 289.950 52.800 292.050 54.900 ;
        RECT 298.800 52.950 300.900 55.050 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 311.400 54.000 312.600 55.650 ;
        RECT 316.950 54.450 319.050 55.050 ;
        RECT 320.400 54.450 321.450 91.950 ;
        RECT 331.950 82.950 334.050 85.050 ;
        RECT 322.950 59.100 325.050 61.200 ;
        RECT 332.400 60.600 333.450 82.950 ;
        RECT 338.400 70.050 339.450 104.100 ;
        RECT 344.400 103.350 345.600 104.100 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 347.400 99.900 348.600 100.650 ;
        RECT 346.950 97.800 349.050 99.900 ;
        RECT 353.400 91.050 354.450 112.950 ;
        RECT 356.400 100.050 357.450 128.400 ;
        RECT 362.400 124.050 363.450 130.800 ;
        RECT 361.950 121.950 364.050 124.050 ;
        RECT 371.400 109.050 372.450 145.950 ;
        RECT 377.400 138.600 378.450 145.950 ;
        RECT 377.400 136.350 378.600 138.600 ;
        RECT 382.950 138.000 385.050 142.050 ;
        RECT 388.950 139.950 391.050 142.050 ;
        RECT 401.400 141.450 402.450 148.950 ;
        RECT 398.400 140.400 402.450 141.450 ;
        RECT 383.400 136.350 384.600 138.000 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 380.400 132.900 381.600 133.650 ;
        RECT 379.950 130.800 382.050 132.900 ;
        RECT 389.400 121.050 390.450 139.950 ;
        RECT 398.400 139.200 399.450 140.400 ;
        RECT 391.950 136.950 394.050 139.050 ;
        RECT 397.950 137.100 400.050 139.200 ;
        RECT 403.950 138.000 406.050 142.050 ;
        RECT 409.950 139.950 412.050 142.050 ;
        RECT 388.950 120.450 391.050 121.050 ;
        RECT 386.400 119.400 391.050 120.450 ;
        RECT 364.950 105.000 367.050 109.050 ;
        RECT 370.950 106.950 373.050 109.050 ;
        RECT 365.400 103.350 366.600 105.000 ;
        RECT 370.950 103.800 373.050 105.900 ;
        RECT 379.950 104.100 382.050 106.200 ;
        RECT 386.400 106.050 387.450 119.400 ;
        RECT 388.950 118.950 391.050 119.400 ;
        RECT 388.950 106.950 391.050 109.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 355.950 97.950 358.050 100.050 ;
        RECT 362.400 99.900 363.600 100.650 ;
        RECT 361.950 97.800 364.050 99.900 ;
        RECT 371.400 94.050 372.450 103.800 ;
        RECT 380.400 103.350 381.600 104.100 ;
        RECT 385.950 103.950 388.050 106.050 ;
        RECT 376.950 100.950 379.050 103.050 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 377.400 99.900 378.600 100.650 ;
        RECT 383.400 99.900 384.600 100.650 ;
        RECT 376.950 97.800 379.050 99.900 ;
        RECT 382.950 97.800 385.050 99.900 ;
        RECT 370.950 91.950 373.050 94.050 ;
        RECT 352.950 88.950 355.050 91.050 ;
        RECT 346.950 85.950 349.050 88.050 ;
        RECT 340.950 70.950 343.050 73.050 ;
        RECT 337.950 67.950 340.050 70.050 ;
        RECT 310.950 49.950 313.050 54.000 ;
        RECT 316.950 53.400 321.450 54.450 ;
        RECT 316.950 52.950 319.050 53.400 ;
        RECT 286.950 37.950 289.050 40.050 ;
        RECT 310.950 37.950 313.050 40.050 ;
        RECT 283.950 31.950 286.050 34.050 ;
        RECT 280.950 28.950 283.050 31.050 ;
        RECT 287.400 28.050 288.450 37.950 ;
        RECT 239.400 25.350 240.600 26.100 ;
        RECT 257.400 25.350 258.600 26.100 ;
        RECT 263.400 25.350 264.600 26.100 ;
        RECT 278.400 25.350 279.600 27.600 ;
        RECT 286.950 25.950 289.050 28.050 ;
        RECT 292.950 26.100 295.050 28.200 ;
        RECT 311.400 27.600 312.450 37.950 ;
        RECT 317.400 27.600 318.450 52.950 ;
        RECT 319.950 46.950 322.050 51.900 ;
        RECT 293.400 25.350 294.600 26.100 ;
        RECT 311.400 25.350 312.600 27.600 ;
        RECT 317.400 25.350 318.600 27.600 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 307.950 22.950 310.050 25.050 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 236.400 21.900 237.600 22.650 ;
        RECT 226.950 19.800 229.050 21.900 ;
        RECT 235.950 19.800 238.050 21.900 ;
        RECT 242.400 20.400 243.600 22.650 ;
        RECT 254.400 21.900 255.600 22.650 ;
        RECT 242.400 16.050 243.450 20.400 ;
        RECT 253.950 19.800 256.050 21.900 ;
        RECT 260.400 21.000 261.600 22.650 ;
        RECT 275.400 21.900 276.600 22.650 ;
        RECT 244.950 16.950 247.050 19.050 ;
        RECT 259.950 16.950 262.050 21.000 ;
        RECT 274.950 19.800 277.050 21.900 ;
        RECT 241.950 13.950 244.050 16.050 ;
        RECT 223.950 10.950 226.050 13.050 ;
        RECT 238.950 12.450 241.050 13.050 ;
        RECT 245.400 12.450 246.450 16.950 ;
        RECT 284.400 16.050 285.450 22.950 ;
        RECT 290.400 21.900 291.600 22.650 ;
        RECT 296.400 21.900 297.600 22.650 ;
        RECT 308.400 21.900 309.600 22.650 ;
        RECT 314.400 21.900 315.600 22.650 ;
        RECT 289.950 19.800 292.050 21.900 ;
        RECT 295.950 19.800 298.050 21.900 ;
        RECT 307.950 19.800 310.050 21.900 ;
        RECT 313.950 19.800 316.050 21.900 ;
        RECT 296.400 18.450 297.450 19.800 ;
        RECT 293.400 17.400 297.450 18.450 ;
        RECT 293.400 16.050 294.450 17.400 ;
        RECT 319.950 16.950 322.050 21.900 ;
        RECT 283.950 13.950 286.050 16.050 ;
        RECT 289.950 14.400 294.450 16.050 ;
        RECT 289.950 13.950 294.000 14.400 ;
        RECT 323.400 13.050 324.450 59.100 ;
        RECT 332.400 58.350 333.600 60.600 ;
        RECT 338.400 60.450 339.600 60.600 ;
        RECT 341.400 60.450 342.450 70.950 ;
        RECT 347.400 64.050 348.450 85.950 ;
        RECT 355.950 70.950 358.050 73.050 ;
        RECT 346.950 61.950 349.050 64.050 ;
        RECT 338.400 59.400 342.450 60.450 ;
        RECT 338.400 58.350 339.600 59.400 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 329.400 53.400 330.600 55.650 ;
        RECT 335.400 54.900 336.600 55.650 ;
        RECT 347.400 54.900 348.450 61.950 ;
        RECT 356.400 60.600 357.450 70.950 ;
        RECT 371.400 64.050 372.450 91.950 ;
        RECT 389.400 88.050 390.450 106.950 ;
        RECT 392.400 106.200 393.450 136.950 ;
        RECT 398.400 136.350 399.600 137.100 ;
        RECT 404.400 136.350 405.600 138.000 ;
        RECT 397.950 133.950 400.050 136.050 ;
        RECT 400.950 133.950 403.050 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 401.400 131.400 402.600 133.650 ;
        RECT 401.400 127.050 402.450 131.400 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 400.950 124.950 403.050 127.050 ;
        RECT 391.950 104.100 394.050 106.200 ;
        RECT 388.950 85.950 391.050 88.050 ;
        RECT 376.950 76.950 379.050 79.050 ;
        RECT 356.400 58.350 357.600 60.600 ;
        RECT 361.950 60.000 364.050 64.050 ;
        RECT 370.950 63.450 373.050 64.050 ;
        RECT 368.400 62.400 373.050 63.450 ;
        RECT 362.400 58.350 363.600 60.000 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 329.400 39.450 330.450 53.400 ;
        RECT 334.950 52.800 337.050 54.900 ;
        RECT 346.950 52.800 349.050 54.900 ;
        RECT 353.400 53.400 354.600 55.650 ;
        RECT 359.400 54.900 360.600 55.650 ;
        RECT 353.400 49.050 354.450 53.400 ;
        RECT 358.950 52.800 361.050 54.900 ;
        RECT 352.950 46.950 355.050 49.050 ;
        RECT 337.950 40.950 340.050 43.050 ;
        RECT 326.400 38.400 330.450 39.450 ;
        RECT 326.400 34.050 327.450 38.400 ;
        RECT 325.950 31.950 328.050 34.050 ;
        RECT 330.000 33.450 334.050 34.050 ;
        RECT 329.400 31.950 334.050 33.450 ;
        RECT 329.400 28.050 330.450 31.950 ;
        RECT 325.950 25.950 328.050 28.050 ;
        RECT 328.950 25.950 331.050 28.050 ;
        RECT 331.950 27.000 334.050 30.900 ;
        RECT 338.400 27.600 339.450 40.950 ;
        RECT 352.950 34.950 355.050 37.050 ;
        RECT 326.400 21.900 327.450 25.950 ;
        RECT 332.400 25.350 333.600 27.000 ;
        RECT 338.400 25.350 339.600 27.600 ;
        RECT 353.400 27.450 354.450 34.950 ;
        RECT 364.950 31.950 367.050 34.050 ;
        RECT 350.400 26.400 354.450 27.450 ;
        RECT 358.950 27.000 361.050 31.050 ;
        RECT 365.400 27.600 366.450 31.950 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 335.400 21.900 336.600 22.650 ;
        RECT 341.400 22.050 342.600 22.650 ;
        RECT 350.400 22.050 351.450 26.400 ;
        RECT 359.400 25.350 360.600 27.000 ;
        RECT 365.400 25.350 366.600 27.600 ;
        RECT 368.400 27.450 369.450 62.400 ;
        RECT 370.950 61.950 373.050 62.400 ;
        RECT 377.400 60.600 378.450 76.950 ;
        RECT 388.950 67.950 391.050 70.050 ;
        RECT 377.400 58.350 378.600 60.600 ;
        RECT 382.950 59.100 385.050 61.200 ;
        RECT 383.400 58.350 384.600 59.100 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 374.400 53.400 375.600 55.650 ;
        RECT 380.400 53.400 381.600 55.650 ;
        RECT 374.400 31.050 375.450 53.400 ;
        RECT 380.400 49.050 381.450 53.400 ;
        RECT 379.950 46.950 382.050 49.050 ;
        RECT 389.400 46.050 390.450 67.950 ;
        RECT 395.400 67.050 396.450 124.950 ;
        RECT 397.950 121.950 400.050 124.050 ;
        RECT 398.400 115.050 399.450 121.950 ;
        RECT 397.950 112.950 400.050 115.050 ;
        RECT 400.950 109.950 403.050 112.050 ;
        RECT 401.400 106.200 402.450 109.950 ;
        RECT 400.950 104.100 403.050 106.200 ;
        RECT 401.400 103.350 402.600 104.100 ;
        RECT 410.400 103.050 411.450 139.950 ;
        RECT 413.400 130.050 414.450 154.950 ;
        RECT 419.400 142.050 420.450 187.950 ;
        RECT 422.400 151.050 423.450 190.950 ;
        RECT 430.950 182.100 433.050 184.200 ;
        RECT 431.400 181.350 432.600 182.100 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 428.400 176.400 429.600 178.650 ;
        RECT 434.400 177.000 435.600 178.650 ;
        RECT 428.400 172.050 429.450 176.400 ;
        RECT 433.950 172.950 436.050 177.000 ;
        RECT 427.950 169.950 430.050 172.050 ;
        RECT 436.950 171.450 439.050 172.050 ;
        RECT 440.400 171.450 441.450 205.950 ;
        RECT 443.400 193.050 444.450 209.400 ;
        RECT 451.950 208.800 454.050 210.900 ;
        RECT 454.950 208.950 457.050 211.050 ;
        RECT 461.400 210.900 462.600 211.650 ;
        RECT 455.400 199.050 456.450 208.950 ;
        RECT 460.950 208.800 463.050 210.900 ;
        RECT 467.400 205.050 468.450 254.400 ;
        RECT 481.950 253.800 484.050 255.900 ;
        RECT 469.950 226.950 472.050 229.050 ;
        RECT 466.950 202.950 469.050 205.050 ;
        RECT 454.950 196.950 457.050 199.050 ;
        RECT 463.950 196.950 466.050 199.050 ;
        RECT 442.950 190.950 445.050 193.050 ;
        RECT 448.950 187.950 451.050 190.050 ;
        RECT 442.950 181.950 445.050 184.050 ;
        RECT 449.400 183.600 450.450 187.950 ;
        RECT 457.950 186.450 460.050 190.050 ;
        RECT 455.400 186.000 460.050 186.450 ;
        RECT 455.400 185.400 459.450 186.000 ;
        RECT 455.400 183.600 456.450 185.400 ;
        RECT 443.400 175.050 444.450 181.950 ;
        RECT 449.400 181.350 450.600 183.600 ;
        RECT 455.400 181.350 456.600 183.600 ;
        RECT 448.950 178.950 451.050 181.050 ;
        RECT 451.950 178.950 454.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 452.400 177.000 453.600 178.650 ;
        RECT 458.400 177.900 459.600 178.650 ;
        RECT 442.950 172.950 445.050 175.050 ;
        RECT 451.950 172.950 454.050 177.000 ;
        RECT 457.950 175.800 460.050 177.900 ;
        RECT 460.950 175.950 463.050 178.050 ;
        RECT 464.400 177.900 465.450 196.950 ;
        RECT 466.950 190.950 469.050 193.050 ;
        RECT 467.400 178.050 468.450 190.950 ;
        RECT 470.400 187.050 471.450 226.950 ;
        RECT 482.400 226.050 483.450 253.800 ;
        RECT 491.400 253.050 492.450 260.400 ;
        RECT 496.950 260.100 499.050 262.200 ;
        RECT 502.950 260.100 505.050 262.200 ;
        RECT 511.950 260.100 514.050 262.200 ;
        RECT 518.400 261.450 519.450 286.950 ;
        RECT 520.950 286.800 523.050 288.900 ;
        RECT 524.400 271.050 525.450 295.950 ;
        RECT 527.400 295.050 528.450 340.800 ;
        RECT 530.400 340.050 531.450 418.950 ;
        RECT 533.400 373.050 534.450 434.400 ;
        RECT 535.950 433.950 538.050 434.400 ;
        RECT 539.400 423.450 540.450 463.950 ;
        RECT 536.400 422.400 540.450 423.450 ;
        RECT 536.400 417.600 537.450 422.400 ;
        RECT 542.400 421.050 543.450 481.950 ;
        RECT 544.950 478.950 550.050 481.050 ;
        RECT 544.800 460.950 546.900 463.050 ;
        RECT 547.950 460.950 550.050 463.050 ;
        RECT 545.400 444.900 546.450 460.950 ;
        RECT 548.400 451.200 549.450 460.950 ;
        RECT 551.400 460.050 552.450 481.950 ;
        RECT 557.400 474.450 558.450 521.400 ;
        RECT 559.950 517.950 562.050 520.050 ;
        RECT 560.400 511.050 561.450 517.950 ;
        RECT 559.950 508.950 562.050 511.050 ;
        RECT 566.400 510.450 567.450 524.400 ;
        RECT 569.400 514.050 570.450 553.800 ;
        RECT 571.950 550.950 574.050 553.050 ;
        RECT 572.400 529.050 573.450 550.950 ;
        RECT 584.400 532.050 585.450 595.950 ;
        RECT 588.300 593.700 589.500 597.300 ;
        RECT 591.300 593.700 592.500 610.200 ;
        RECT 593.700 615.300 595.800 617.400 ;
        RECT 593.700 593.700 594.900 615.300 ;
        RECT 602.400 613.800 604.500 615.900 ;
        RECT 607.800 615.300 609.900 617.400 ;
        RECT 595.950 610.950 598.050 613.050 ;
        RECT 596.400 604.050 597.450 610.950 ;
        RECT 602.400 607.200 603.300 613.800 ;
        RECT 608.100 608.100 609.300 615.300 ;
        RECT 610.800 613.500 612.300 618.300 ;
        RECT 613.200 615.300 615.300 620.400 ;
        RECT 610.800 611.400 612.900 613.500 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 598.950 603.000 601.050 607.050 ;
        RECT 602.400 605.100 604.500 607.200 ;
        RECT 607.800 606.000 609.900 608.100 ;
        RECT 599.400 601.350 600.600 603.000 ;
        RECT 598.800 598.950 600.900 601.050 ;
        RECT 602.400 594.600 603.300 605.100 ;
        RECT 605.100 598.500 607.200 600.600 ;
        RECT 587.700 591.600 589.800 593.700 ;
        RECT 590.700 591.600 592.800 593.700 ;
        RECT 593.700 591.600 595.800 593.700 ;
        RECT 601.800 592.500 603.900 594.600 ;
        RECT 608.100 593.700 609.300 606.000 ;
        RECT 610.800 593.700 612.300 611.400 ;
        RECT 614.100 593.700 615.300 615.300 ;
        RECT 607.200 591.600 609.300 593.700 ;
        RECT 610.200 591.600 612.300 593.700 ;
        RECT 613.200 591.600 615.300 593.700 ;
        RECT 616.200 618.300 618.300 620.400 ;
        RECT 616.200 613.500 617.700 618.300 ;
        RECT 616.200 611.400 618.300 613.500 ;
        RECT 616.200 593.700 617.700 611.400 ;
        RECT 616.200 591.600 618.300 593.700 ;
        RECT 604.950 586.950 607.050 589.050 ;
        RECT 620.400 588.450 621.450 631.950 ;
        RECT 625.950 628.950 628.050 631.050 ;
        RECT 626.400 612.450 627.450 628.950 ;
        RECT 628.950 625.950 631.050 628.050 ;
        RECT 629.400 616.050 630.450 625.950 ;
        RECT 628.950 613.950 631.050 616.050 ;
        RECT 626.400 611.400 630.450 612.450 ;
        RECT 625.800 604.950 627.900 607.050 ;
        RECT 626.400 602.400 627.600 604.650 ;
        RECT 622.950 598.950 625.050 601.050 ;
        RECT 617.400 587.400 621.450 588.450 ;
        RECT 605.400 583.050 606.450 586.950 ;
        RECT 604.950 580.950 607.050 583.050 ;
        RECT 592.950 573.000 595.050 577.050 ;
        RECT 601.950 574.950 604.050 577.050 ;
        RECT 593.400 571.350 594.600 573.000 ;
        RECT 602.400 571.050 603.450 574.950 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 595.950 568.950 598.050 571.050 ;
        RECT 601.950 568.950 604.050 571.050 ;
        RECT 590.400 567.900 591.600 568.650 ;
        RECT 589.950 565.800 592.050 567.900 ;
        RECT 596.400 567.000 597.600 568.650 ;
        RECT 605.400 568.050 606.450 580.950 ;
        RECT 613.950 577.950 616.050 580.050 ;
        RECT 614.400 573.600 615.450 577.950 ;
        RECT 617.400 577.050 618.450 587.400 ;
        RECT 619.950 583.950 622.050 586.050 ;
        RECT 616.950 574.950 619.050 577.050 ;
        RECT 620.400 574.050 621.450 583.950 ;
        RECT 614.400 571.350 615.600 573.600 ;
        RECT 619.950 571.950 622.050 574.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 595.950 562.950 598.050 567.000 ;
        RECT 598.950 565.800 601.050 567.900 ;
        RECT 604.950 565.950 607.050 568.050 ;
        RECT 611.400 567.900 612.600 568.650 ;
        RECT 610.950 565.800 613.050 567.900 ;
        RECT 617.400 566.400 618.600 568.650 ;
        RECT 592.950 556.950 595.050 559.050 ;
        RECT 574.950 529.950 577.050 532.050 ;
        RECT 583.950 529.950 586.050 532.050 ;
        RECT 571.950 526.950 574.050 529.050 ;
        RECT 571.950 520.800 574.050 522.900 ;
        RECT 568.950 511.950 571.050 514.050 ;
        RECT 563.400 509.400 567.450 510.450 ;
        RECT 563.400 496.200 564.450 509.400 ;
        RECT 568.950 502.950 571.050 505.050 ;
        RECT 562.950 494.100 565.050 496.200 ;
        RECT 569.400 496.050 570.450 502.950 ;
        RECT 563.400 493.350 564.600 494.100 ;
        RECT 568.950 493.950 571.050 496.050 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 566.400 488.400 567.600 490.650 ;
        RECT 566.400 478.050 567.450 488.400 ;
        RECT 568.950 487.950 571.050 490.050 ;
        RECT 565.950 475.950 568.050 478.050 ;
        RECT 554.400 473.400 558.450 474.450 ;
        RECT 550.950 457.950 553.050 460.050 ;
        RECT 554.400 457.050 555.450 473.400 ;
        RECT 553.950 454.950 556.050 457.050 ;
        RECT 569.400 454.050 570.450 487.950 ;
        RECT 572.400 469.050 573.450 520.800 ;
        RECT 575.400 508.050 576.450 529.950 ;
        RECT 577.950 526.950 580.050 529.050 ;
        RECT 587.400 528.450 588.600 528.600 ;
        RECT 587.400 527.400 591.450 528.450 ;
        RECT 578.400 520.050 579.450 526.950 ;
        RECT 587.400 526.350 588.600 527.400 ;
        RECT 581.400 523.950 583.500 526.050 ;
        RECT 586.800 523.950 588.900 526.050 ;
        RECT 581.400 522.900 582.600 523.650 ;
        RECT 580.950 520.800 583.050 522.900 ;
        RECT 577.950 517.950 580.050 520.050 ;
        RECT 586.950 517.950 589.050 520.050 ;
        RECT 580.950 511.950 583.050 514.050 ;
        RECT 577.950 508.950 580.050 511.050 ;
        RECT 574.950 505.950 577.050 508.050 ;
        RECT 578.400 505.050 579.450 508.950 ;
        RECT 581.400 505.050 582.450 511.950 ;
        RECT 587.400 505.050 588.450 517.950 ;
        RECT 574.950 502.800 577.050 504.900 ;
        RECT 577.950 502.950 580.050 505.050 ;
        RECT 580.950 502.950 583.050 505.050 ;
        RECT 586.950 502.950 589.050 505.050 ;
        RECT 575.400 490.050 576.450 502.800 ;
        RECT 590.400 502.050 591.450 527.400 ;
        RECT 593.400 511.050 594.450 556.950 ;
        RECT 599.400 555.450 600.450 565.800 ;
        RECT 601.950 562.950 604.050 565.050 ;
        RECT 596.400 554.400 600.450 555.450 ;
        RECT 596.400 520.050 597.450 554.400 ;
        RECT 602.400 538.050 603.450 562.950 ;
        RECT 610.950 559.950 613.050 562.050 ;
        RECT 601.950 535.950 604.050 538.050 ;
        RECT 598.950 532.950 601.050 535.050 ;
        RECT 595.950 517.950 598.050 520.050 ;
        RECT 595.950 514.800 598.050 516.900 ;
        RECT 592.950 508.950 595.050 511.050 ;
        RECT 592.950 502.950 595.050 505.050 ;
        RECT 589.950 499.950 592.050 502.050 ;
        RECT 577.950 493.950 580.050 496.050 ;
        RECT 586.950 494.100 589.050 496.200 ;
        RECT 574.950 487.950 577.050 490.050 ;
        RECT 578.400 475.050 579.450 493.950 ;
        RECT 587.400 493.350 588.600 494.100 ;
        RECT 581.100 490.950 583.200 493.050 ;
        RECT 586.500 490.950 588.600 493.050 ;
        RECT 589.800 490.950 591.900 493.050 ;
        RECT 581.400 489.900 582.600 490.650 ;
        RECT 580.950 487.800 583.050 489.900 ;
        RECT 590.400 488.400 591.600 490.650 ;
        RECT 580.950 484.650 583.050 486.750 ;
        RECT 586.950 484.950 589.050 487.050 ;
        RECT 577.950 472.950 580.050 475.050 ;
        RECT 578.400 469.050 579.450 472.950 ;
        RECT 571.950 466.950 574.050 469.050 ;
        RECT 577.950 466.950 580.050 469.050 ;
        RECT 574.950 457.950 577.050 460.050 ;
        RECT 562.950 451.950 565.050 454.050 ;
        RECT 568.950 451.950 571.050 454.050 ;
        RECT 547.950 449.100 550.050 451.200 ;
        RECT 556.950 449.100 559.050 451.200 ;
        RECT 548.400 448.350 549.600 449.100 ;
        RECT 557.400 448.350 558.600 449.100 ;
        RECT 548.100 445.950 550.200 448.050 ;
        RECT 553.500 445.950 555.600 448.050 ;
        RECT 556.800 445.950 558.900 448.050 ;
        RECT 554.400 444.900 555.600 445.650 ;
        RECT 544.950 442.800 547.050 444.900 ;
        RECT 553.950 442.800 556.050 444.900 ;
        RECT 541.950 418.950 544.050 421.050 ;
        RECT 536.400 415.350 537.600 417.600 ;
        RECT 536.400 412.950 538.500 415.050 ;
        RECT 541.800 412.950 543.900 415.050 ;
        RECT 542.400 410.400 543.600 412.650 ;
        RECT 538.950 403.950 541.050 406.050 ;
        RECT 539.400 375.450 540.450 403.950 ;
        RECT 542.400 385.050 543.450 410.400 ;
        RECT 545.400 400.050 546.450 442.800 ;
        RECT 556.950 439.950 559.050 442.050 ;
        RECT 557.400 424.050 558.450 439.950 ;
        RECT 559.950 430.950 562.050 433.050 ;
        RECT 556.950 421.950 559.050 424.050 ;
        RECT 560.400 418.200 561.450 430.950 ;
        RECT 563.400 420.450 564.450 451.950 ;
        RECT 569.400 450.600 570.450 451.950 ;
        RECT 575.400 450.600 576.450 457.950 ;
        RECT 578.400 451.050 579.450 466.950 ;
        RECT 569.400 448.350 570.600 450.600 ;
        RECT 575.400 448.350 576.600 450.600 ;
        RECT 577.950 448.950 580.050 451.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 572.400 444.900 573.600 445.650 ;
        RECT 571.950 442.800 574.050 444.900 ;
        RECT 577.950 442.950 580.050 445.050 ;
        RECT 568.950 433.950 571.050 436.050 ;
        RECT 563.400 419.400 567.450 420.450 ;
        RECT 559.950 416.100 562.050 418.200 ;
        RECT 560.400 415.350 561.600 416.100 ;
        RECT 554.100 412.950 556.200 415.050 ;
        RECT 559.500 412.950 561.600 415.050 ;
        RECT 562.800 412.950 564.900 415.050 ;
        RECT 554.400 411.450 555.600 412.650 ;
        RECT 548.400 410.400 555.600 411.450 ;
        RECT 563.400 410.400 564.600 412.650 ;
        RECT 544.950 397.950 547.050 400.050 ;
        RECT 548.400 391.050 549.450 410.400 ;
        RECT 563.400 409.050 564.450 410.400 ;
        RECT 553.950 406.950 556.050 409.050 ;
        RECT 562.950 406.950 565.050 409.050 ;
        RECT 550.950 394.950 553.050 397.050 ;
        RECT 547.950 388.950 550.050 391.050 ;
        RECT 541.950 382.950 544.050 385.050 ;
        RECT 544.950 379.950 547.050 382.050 ;
        RECT 545.400 376.050 546.450 379.950 ;
        RECT 551.400 379.050 552.450 394.950 ;
        RECT 550.950 376.950 553.050 379.050 ;
        RECT 539.400 374.400 543.450 375.450 ;
        RECT 532.950 370.950 535.050 373.050 ;
        RECT 535.950 371.100 538.050 373.200 ;
        RECT 542.400 372.600 543.450 374.400 ;
        RECT 544.950 373.950 547.050 376.050 ;
        RECT 536.400 370.350 537.600 371.100 ;
        RECT 542.400 370.350 543.600 372.600 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 532.950 364.950 535.050 367.050 ;
        RECT 539.400 365.400 540.600 367.650 ;
        RECT 545.400 366.900 546.600 367.650 ;
        RECT 551.400 366.900 552.450 376.950 ;
        RECT 554.400 370.050 555.450 406.950 ;
        RECT 563.400 388.050 564.450 406.950 ;
        RECT 566.400 394.050 567.450 419.400 ;
        RECT 565.950 391.950 568.050 394.050 ;
        RECT 562.950 385.950 565.050 388.050 ;
        RECT 569.400 378.450 570.450 433.950 ;
        RECT 578.400 430.050 579.450 442.950 ;
        RECT 581.400 441.450 582.450 484.650 ;
        RECT 583.950 460.950 586.050 463.050 ;
        RECT 584.400 444.450 585.450 460.950 ;
        RECT 587.400 460.050 588.450 484.950 ;
        RECT 590.400 484.050 591.450 488.400 ;
        RECT 593.400 487.050 594.450 502.950 ;
        RECT 596.400 490.050 597.450 514.800 ;
        RECT 599.400 508.050 600.450 532.950 ;
        RECT 602.400 528.600 603.450 535.950 ;
        RECT 602.400 526.350 603.600 528.600 ;
        RECT 602.100 523.950 604.200 526.050 ;
        RECT 607.500 523.950 609.600 526.050 ;
        RECT 608.400 521.400 609.600 523.650 ;
        RECT 601.950 517.950 604.050 520.050 ;
        RECT 598.950 505.950 601.050 508.050 ;
        RECT 602.400 501.450 603.450 517.950 ;
        RECT 608.400 514.050 609.450 521.400 ;
        RECT 607.950 511.950 610.050 514.050 ;
        RECT 599.400 500.400 603.450 501.450 ;
        RECT 595.950 487.950 598.050 490.050 ;
        RECT 599.400 489.450 600.450 500.400 ;
        RECT 604.950 494.100 607.050 496.200 ;
        RECT 611.400 495.600 612.450 559.950 ;
        RECT 617.400 558.450 618.450 566.400 ;
        RECT 619.950 565.950 622.050 568.050 ;
        RECT 614.400 557.400 618.450 558.450 ;
        RECT 614.400 547.050 615.450 557.400 ;
        RECT 620.400 553.050 621.450 565.950 ;
        RECT 623.400 556.050 624.450 598.950 ;
        RECT 626.400 586.050 627.450 602.400 ;
        RECT 625.950 583.950 628.050 586.050 ;
        RECT 629.400 582.450 630.450 611.400 ;
        RECT 638.400 607.200 639.450 640.950 ;
        RECT 640.950 625.950 643.050 628.050 ;
        RECT 634.800 604.950 636.900 607.050 ;
        RECT 637.950 605.100 640.050 607.200 ;
        RECT 635.400 603.000 636.600 604.650 ;
        RECT 634.950 598.950 637.050 603.000 ;
        RECT 626.400 581.400 630.450 582.450 ;
        RECT 626.400 574.050 627.450 581.400 ;
        RECT 631.950 577.950 634.050 580.050 ;
        RECT 632.400 574.200 633.450 577.950 ;
        RECT 625.950 571.950 628.050 574.050 ;
        RECT 631.950 572.100 634.050 574.200 ;
        RECT 632.400 571.350 633.600 572.100 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 629.400 566.400 630.600 568.650 ;
        RECT 638.400 567.450 639.450 605.100 ;
        RECT 641.400 601.050 642.450 625.950 ;
        RECT 640.950 598.950 643.050 601.050 ;
        RECT 644.400 595.050 645.450 640.950 ;
        RECT 649.950 625.950 652.050 628.050 ;
        RECT 650.400 619.050 651.450 625.950 ;
        RECT 649.950 616.950 652.050 619.050 ;
        RECT 659.400 610.050 660.450 644.400 ;
        RECT 664.950 643.800 667.050 645.900 ;
        RECT 661.950 640.950 664.050 643.050 ;
        RECT 658.950 607.950 661.050 610.050 ;
        RECT 652.950 605.100 655.050 607.200 ;
        RECT 653.400 604.350 654.600 605.100 ;
        RECT 658.950 604.800 661.050 606.900 ;
        RECT 649.950 601.950 652.050 604.050 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 650.400 599.400 651.600 601.650 ;
        RECT 643.950 592.950 646.050 595.050 ;
        RECT 650.400 583.050 651.450 599.400 ;
        RECT 652.950 586.950 655.050 589.050 ;
        RECT 649.950 580.950 652.050 583.050 ;
        RECT 646.950 573.000 649.050 577.050 ;
        RECT 653.400 573.600 654.450 586.950 ;
        RECT 647.400 571.350 648.600 573.000 ;
        RECT 653.400 571.350 654.600 573.600 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 644.400 567.900 645.600 568.650 ;
        RECT 635.400 566.400 639.450 567.450 ;
        RECT 622.950 553.950 625.050 556.050 ;
        RECT 619.950 550.950 622.050 553.050 ;
        RECT 625.950 550.950 628.050 553.050 ;
        RECT 613.950 544.950 616.050 547.050 ;
        RECT 614.400 523.050 615.450 544.950 ;
        RECT 619.950 538.950 622.050 541.050 ;
        RECT 620.400 528.600 621.450 538.950 ;
        RECT 626.400 532.050 627.450 550.950 ;
        RECT 629.400 544.050 630.450 566.400 ;
        RECT 628.950 541.950 631.050 544.050 ;
        RECT 628.950 532.950 631.050 535.050 ;
        RECT 625.950 529.950 628.050 532.050 ;
        RECT 629.400 528.600 630.450 532.950 ;
        RECT 620.400 528.450 621.600 528.600 ;
        RECT 617.400 527.400 621.600 528.450 ;
        RECT 613.950 520.950 616.050 523.050 ;
        RECT 617.400 517.050 618.450 527.400 ;
        RECT 620.400 526.350 621.600 527.400 ;
        RECT 629.400 526.350 630.600 528.600 ;
        RECT 631.950 527.100 634.050 529.200 ;
        RECT 620.100 523.950 622.200 526.050 ;
        RECT 625.500 523.950 627.600 526.050 ;
        RECT 628.800 523.950 630.900 526.050 ;
        RECT 626.400 521.400 627.600 523.650 ;
        RECT 616.950 514.950 619.050 517.050 ;
        RECT 626.400 514.050 627.450 521.400 ;
        RECT 625.950 511.950 628.050 514.050 ;
        RECT 622.950 508.950 625.050 511.050 ;
        RECT 605.400 493.350 606.600 494.100 ;
        RECT 611.400 493.350 612.600 495.600 ;
        RECT 619.950 493.950 622.050 496.050 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 599.400 488.400 603.450 489.450 ;
        RECT 592.950 484.950 595.050 487.050 ;
        RECT 589.950 481.950 592.050 484.050 ;
        RECT 602.400 468.450 603.450 488.400 ;
        RECT 608.400 488.400 609.600 490.650 ;
        RECT 614.400 488.400 615.600 490.650 ;
        RECT 608.400 478.050 609.450 488.400 ;
        RECT 614.400 484.050 615.450 488.400 ;
        RECT 616.950 487.800 619.050 489.900 ;
        RECT 613.950 483.450 616.050 484.050 ;
        RECT 611.400 482.400 616.050 483.450 ;
        RECT 607.950 477.450 610.050 478.050 ;
        RECT 599.400 467.400 603.450 468.450 ;
        RECT 605.400 476.400 610.050 477.450 ;
        RECT 586.950 457.950 589.050 460.050 ;
        RECT 586.950 450.600 591.000 451.050 ;
        RECT 586.950 448.950 591.600 450.600 ;
        RECT 590.400 448.350 591.600 448.950 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 593.400 444.900 594.600 445.650 ;
        RECT 584.400 443.400 588.450 444.450 ;
        RECT 581.400 440.400 585.450 441.450 ;
        RECT 577.950 427.950 580.050 430.050 ;
        RECT 571.950 421.950 574.050 424.050 ;
        RECT 566.400 377.400 570.450 378.450 ;
        RECT 559.950 376.050 562.050 376.200 ;
        RECT 559.950 374.100 565.050 376.050 ;
        RECT 561.000 373.950 565.050 374.100 ;
        RECT 559.950 370.950 562.050 373.050 ;
        RECT 566.400 372.600 567.450 377.400 ;
        RECT 560.400 370.350 561.600 370.950 ;
        RECT 566.400 370.350 567.600 372.600 ;
        RECT 568.950 370.950 571.050 376.050 ;
        RECT 553.950 367.950 556.050 370.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 533.400 355.050 534.450 364.950 ;
        RECT 532.950 352.950 535.050 355.050 ;
        RECT 539.400 348.450 540.450 365.400 ;
        RECT 544.950 364.800 547.050 366.900 ;
        RECT 550.950 364.800 553.050 366.900 ;
        RECT 547.950 358.950 550.050 361.050 ;
        RECT 541.950 352.950 544.050 355.050 ;
        RECT 536.400 347.400 540.450 348.450 ;
        RECT 536.400 343.050 537.450 347.400 ;
        RECT 538.950 343.950 541.050 346.050 ;
        RECT 535.950 340.950 538.050 343.050 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 532.950 338.100 535.050 340.200 ;
        RECT 539.400 339.600 540.450 343.950 ;
        RECT 542.400 343.050 543.450 352.950 ;
        RECT 544.950 349.950 547.050 352.050 ;
        RECT 541.950 340.950 544.050 343.050 ;
        RECT 533.400 337.350 534.600 338.100 ;
        RECT 539.400 337.350 540.600 339.600 ;
        RECT 545.400 339.450 546.450 349.950 ;
        RECT 548.400 349.050 549.450 358.950 ;
        RECT 550.950 355.950 553.050 358.050 ;
        RECT 547.950 346.950 550.050 349.050 ;
        RECT 551.400 340.050 552.450 355.950 ;
        RECT 554.400 349.050 555.450 367.950 ;
        RECT 563.400 365.400 564.600 367.650 ;
        RECT 563.400 355.050 564.450 365.400 ;
        RECT 572.400 358.050 573.450 421.950 ;
        RECT 574.950 415.950 577.050 418.050 ;
        RECT 584.400 417.600 585.450 440.400 ;
        RECT 575.400 406.050 576.450 415.950 ;
        RECT 584.400 415.350 585.600 417.600 ;
        RECT 578.100 412.950 580.200 415.050 ;
        RECT 583.500 412.950 585.600 415.050 ;
        RECT 578.400 410.400 579.600 412.650 ;
        RECT 574.950 403.950 577.050 406.050 ;
        RECT 574.950 391.950 577.050 394.050 ;
        RECT 575.400 376.050 576.450 391.950 ;
        RECT 578.400 391.050 579.450 410.400 ;
        RECT 587.400 409.050 588.450 443.400 ;
        RECT 592.950 442.800 595.050 444.900 ;
        RECT 593.400 439.050 594.450 442.800 ;
        RECT 595.950 439.950 598.050 442.050 ;
        RECT 592.950 436.950 595.050 439.050 ;
        RECT 596.400 427.050 597.450 439.950 ;
        RECT 599.400 436.050 600.450 467.400 ;
        RECT 601.950 451.950 604.050 454.050 ;
        RECT 602.400 442.050 603.450 451.950 ;
        RECT 605.400 451.050 606.450 476.400 ;
        RECT 607.950 475.950 610.050 476.400 ;
        RECT 611.400 453.450 612.450 482.400 ;
        RECT 613.950 481.950 616.050 482.400 ;
        RECT 613.950 472.950 616.050 475.050 ;
        RECT 614.400 457.050 615.450 472.950 ;
        RECT 617.400 463.050 618.450 487.800 ;
        RECT 620.400 469.050 621.450 493.950 ;
        RECT 623.400 484.050 624.450 508.950 ;
        RECT 626.400 496.050 627.450 511.950 ;
        RECT 632.400 511.050 633.450 527.100 ;
        RECT 631.950 508.950 634.050 511.050 ;
        RECT 635.400 499.050 636.450 566.400 ;
        RECT 643.950 565.800 646.050 567.900 ;
        RECT 650.400 567.000 651.600 568.650 ;
        RECT 643.950 559.950 646.050 564.750 ;
        RECT 649.950 562.950 652.050 567.000 ;
        RECT 646.950 556.950 649.050 559.050 ;
        RECT 647.400 535.050 648.450 556.950 ;
        RECT 659.400 541.050 660.450 604.800 ;
        RECT 662.400 600.450 663.450 640.950 ;
        RECT 667.950 631.950 670.050 634.050 ;
        RECT 668.400 606.600 669.450 631.950 ;
        RECT 671.400 613.050 672.450 658.950 ;
        RECT 680.400 655.050 681.450 664.950 ;
        RECT 679.950 652.950 682.050 655.050 ;
        RECT 676.950 650.100 679.050 652.200 ;
        RECT 682.950 650.100 685.050 652.200 ;
        RECT 677.400 649.350 678.600 650.100 ;
        RECT 683.400 649.350 684.600 650.100 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 679.950 646.950 682.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 685.950 646.950 688.050 649.050 ;
        RECT 673.950 643.950 676.050 646.050 ;
        RECT 680.400 645.000 681.600 646.650 ;
        RECT 686.400 645.900 687.600 646.650 ;
        RECT 674.400 613.050 675.450 643.950 ;
        RECT 679.950 640.950 682.050 645.000 ;
        RECT 685.950 643.800 688.050 645.900 ;
        RECT 692.400 643.050 693.450 676.800 ;
        RECT 695.400 673.050 696.450 679.950 ;
        RECT 694.950 670.950 697.050 673.050 ;
        RECT 698.400 654.450 699.450 682.950 ;
        RECT 701.400 682.350 702.600 683.100 ;
        RECT 710.400 682.350 711.600 684.000 ;
        RECT 712.950 682.950 715.050 685.050 ;
        RECT 718.950 682.950 721.050 688.050 ;
        RECT 701.400 679.950 703.500 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 716.100 679.950 718.200 682.050 ;
        RECT 707.400 678.000 708.600 679.650 ;
        RECT 716.400 678.900 717.600 679.650 ;
        RECT 706.950 673.950 709.050 678.000 ;
        RECT 715.950 676.800 718.050 678.900 ;
        RECT 722.400 676.050 723.450 715.950 ;
        RECT 725.400 688.050 726.450 724.800 ;
        RECT 731.400 722.400 732.600 724.650 ;
        RECT 731.400 718.050 732.450 722.400 ;
        RECT 730.950 715.950 733.050 718.050 ;
        RECT 733.950 712.950 736.050 715.050 ;
        RECT 730.950 706.950 733.050 709.050 ;
        RECT 724.950 685.950 727.050 688.050 ;
        RECT 731.400 685.200 732.450 706.950 ;
        RECT 734.400 691.050 735.450 712.950 ;
        RECT 736.950 694.950 739.050 697.050 ;
        RECT 733.950 688.950 736.050 691.050 ;
        RECT 724.950 682.800 727.050 684.900 ;
        RECT 730.950 683.100 733.050 685.200 ;
        RECT 737.400 684.600 738.450 694.950 ;
        RECT 740.400 688.050 741.450 754.950 ;
        RECT 743.400 751.050 744.450 772.950 ;
        RECT 746.400 766.050 747.450 796.950 ;
        RECT 749.400 778.050 750.450 805.950 ;
        RECT 758.400 805.350 759.600 807.000 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 757.950 802.950 760.050 805.050 ;
        RECT 760.950 802.950 763.050 805.050 ;
        RECT 755.400 800.400 756.600 802.650 ;
        RECT 761.400 801.450 762.600 802.650 ;
        RECT 761.400 800.400 765.450 801.450 ;
        RECT 755.400 796.050 756.450 800.400 ;
        RECT 754.950 793.950 757.050 796.050 ;
        RECT 748.950 775.950 751.050 778.050 ;
        RECT 755.400 766.050 756.450 793.950 ;
        RECT 764.400 793.050 765.450 800.400 ;
        RECT 763.950 790.950 766.050 793.050 ;
        RECT 757.950 778.950 760.050 781.050 ;
        RECT 745.950 763.950 748.050 766.050 ;
        RECT 754.950 763.950 757.050 766.050 ;
        RECT 758.400 762.600 759.450 778.950 ;
        RECT 749.400 762.450 750.600 762.600 ;
        RECT 746.400 761.400 750.600 762.450 ;
        RECT 742.950 748.950 745.050 751.050 ;
        RECT 746.400 747.450 747.450 761.400 ;
        RECT 749.400 760.350 750.600 761.400 ;
        RECT 758.400 760.350 759.600 762.600 ;
        RECT 749.100 757.950 751.200 760.050 ;
        RECT 754.500 757.950 756.600 760.050 ;
        RECT 757.800 757.950 759.900 760.050 ;
        RECT 755.400 756.900 756.600 757.650 ;
        RECT 754.950 754.800 757.050 756.900 ;
        RECT 760.950 754.950 763.050 757.050 ;
        RECT 743.400 746.400 747.450 747.450 ;
        RECT 743.400 709.050 744.450 746.400 ;
        RECT 761.400 745.050 762.450 754.950 ;
        RECT 764.400 748.050 765.450 790.950 ;
        RECT 767.400 775.050 768.450 817.950 ;
        RECT 770.400 793.050 771.450 835.950 ;
        RECT 779.400 833.400 780.600 835.650 ;
        RECT 785.400 833.400 786.600 835.650 ;
        RECT 779.400 826.050 780.450 833.400 ;
        RECT 785.400 829.050 786.450 833.400 ;
        RECT 785.400 827.400 790.050 829.050 ;
        RECT 786.000 826.950 790.050 827.400 ;
        RECT 778.950 823.950 781.050 826.050 ;
        RECT 784.950 823.950 787.050 826.050 ;
        RECT 785.400 817.050 786.450 823.950 ;
        RECT 784.950 814.950 787.050 817.050 ;
        RECT 778.950 806.100 781.050 808.200 ;
        RECT 785.400 807.600 786.450 814.950 ;
        RECT 779.400 805.350 780.600 806.100 ;
        RECT 785.400 805.350 786.600 807.600 ;
        RECT 791.400 805.050 792.450 854.400 ;
        RECT 796.950 839.100 799.050 841.200 ;
        RECT 803.400 840.600 804.450 856.950 ;
        RECT 797.400 838.350 798.600 839.100 ;
        RECT 803.400 838.350 804.600 840.600 ;
        RECT 796.950 835.950 799.050 838.050 ;
        RECT 799.950 835.950 802.050 838.050 ;
        RECT 802.950 835.950 805.050 838.050 ;
        RECT 800.400 834.900 801.600 835.650 ;
        RECT 809.400 834.900 810.450 862.950 ;
        RECT 842.400 862.050 843.450 910.800 ;
        RECT 847.950 907.950 850.050 912.900 ;
        RECT 854.400 911.400 855.600 913.650 ;
        RECT 854.400 898.050 855.450 911.400 ;
        RECT 863.400 901.050 864.450 925.950 ;
        RECT 868.950 922.950 871.050 925.050 ;
        RECT 928.950 922.950 931.050 925.050 ;
        RECT 869.400 918.600 870.450 922.950 ;
        RECT 869.400 916.350 870.600 918.600 ;
        RECT 874.950 917.100 877.050 919.200 ;
        RECT 875.400 916.350 876.600 917.100 ;
        RECT 883.950 916.950 886.050 919.050 ;
        RECT 892.950 917.100 895.050 919.200 ;
        RECT 898.950 917.100 901.050 919.200 ;
        RECT 868.950 913.950 871.050 916.050 ;
        RECT 871.950 913.950 874.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 872.400 912.900 873.600 913.650 ;
        RECT 878.400 912.900 879.600 913.650 ;
        RECT 871.950 910.800 874.050 912.900 ;
        RECT 877.950 910.800 880.050 912.900 ;
        RECT 884.400 904.050 885.450 916.950 ;
        RECT 893.400 916.350 894.600 917.100 ;
        RECT 899.400 916.350 900.600 917.100 ;
        RECT 907.950 916.950 910.050 919.050 ;
        RECT 916.950 917.100 919.050 919.200 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 892.950 913.950 895.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 898.950 913.950 901.050 916.050 ;
        RECT 890.400 912.900 891.600 913.650 ;
        RECT 889.950 910.800 892.050 912.900 ;
        RECT 896.400 911.400 897.600 913.650 ;
        RECT 883.950 901.950 886.050 904.050 ;
        RECT 862.950 898.950 865.050 901.050 ;
        RECT 892.950 898.950 895.050 901.050 ;
        RECT 853.950 895.950 856.050 898.050 ;
        RECT 862.950 895.800 865.050 897.900 ;
        RECT 850.950 889.950 853.050 892.050 ;
        RECT 851.400 885.600 852.450 889.950 ;
        RECT 851.400 883.350 852.600 885.600 ;
        RECT 856.950 884.100 859.050 886.200 ;
        RECT 857.400 883.350 858.600 884.100 ;
        RECT 847.950 880.950 850.050 883.050 ;
        RECT 850.950 880.950 853.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 848.400 879.900 849.600 880.650 ;
        RECT 847.950 877.800 850.050 879.900 ;
        RECT 854.400 878.400 855.600 880.650 ;
        RECT 854.400 868.050 855.450 878.400 ;
        RECT 859.950 877.950 862.050 880.050 ;
        RECT 853.950 865.950 856.050 868.050 ;
        RECT 841.950 859.950 844.050 862.050 ;
        RECT 832.950 853.950 835.050 856.050 ;
        RECT 817.950 850.950 820.050 853.050 ;
        RECT 811.950 847.950 814.050 850.050 ;
        RECT 799.950 832.800 802.050 834.900 ;
        RECT 808.950 832.800 811.050 834.900 ;
        RECT 812.400 834.450 813.450 847.950 ;
        RECT 818.400 843.450 819.450 850.950 ;
        RECT 826.950 847.950 829.050 850.050 ;
        RECT 818.400 842.400 822.450 843.450 ;
        RECT 821.400 840.600 822.450 842.400 ;
        RECT 827.400 840.600 828.450 847.950 ;
        RECT 821.400 838.350 822.600 840.600 ;
        RECT 827.400 838.350 828.600 840.600 ;
        RECT 817.950 835.950 820.050 838.050 ;
        RECT 820.950 835.950 823.050 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 826.950 835.950 829.050 838.050 ;
        RECT 818.400 834.450 819.600 835.650 ;
        RECT 824.400 834.900 825.600 835.650 ;
        RECT 833.400 834.900 834.450 853.950 ;
        RECT 860.400 844.050 861.450 877.950 ;
        RECT 863.400 867.450 864.450 895.800 ;
        RECT 865.950 883.950 868.050 886.050 ;
        RECT 871.950 884.100 874.050 886.200 ;
        RECT 877.950 884.100 880.050 886.200 ;
        RECT 866.400 871.050 867.450 883.950 ;
        RECT 872.400 883.350 873.600 884.100 ;
        RECT 878.400 883.350 879.600 884.100 ;
        RECT 886.800 883.950 888.900 886.050 ;
        RECT 889.950 883.950 892.050 889.050 ;
        RECT 893.400 885.600 894.450 898.950 ;
        RECT 896.400 892.050 897.450 911.400 ;
        RECT 904.950 910.950 907.050 913.050 ;
        RECT 898.950 895.950 901.050 898.050 ;
        RECT 895.950 889.950 898.050 892.050 ;
        RECT 899.400 886.200 900.450 895.950 ;
        RECT 871.950 880.950 874.050 883.050 ;
        RECT 874.950 880.950 877.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 880.950 880.950 883.050 883.050 ;
        RECT 868.950 877.950 871.050 880.050 ;
        RECT 875.400 878.400 876.600 880.650 ;
        RECT 881.400 878.400 882.600 880.650 ;
        RECT 887.400 879.900 888.450 883.950 ;
        RECT 893.400 883.350 894.600 885.600 ;
        RECT 898.950 884.100 901.050 886.200 ;
        RECT 905.400 886.050 906.450 910.950 ;
        RECT 908.400 898.050 909.450 916.950 ;
        RECT 917.400 916.350 918.600 917.100 ;
        RECT 913.950 913.950 916.050 916.050 ;
        RECT 916.950 913.950 919.050 916.050 ;
        RECT 914.400 912.900 915.600 913.650 ;
        RECT 929.400 912.900 930.450 922.950 ;
        RECT 913.950 910.800 916.050 912.900 ;
        RECT 928.950 910.800 931.050 912.900 ;
        RECT 907.950 895.950 910.050 898.050 ;
        RECT 907.950 886.950 910.050 889.050 ;
        RECT 899.400 883.350 900.600 884.100 ;
        RECT 904.950 883.950 907.050 886.050 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 901.950 880.950 904.050 883.050 ;
        RECT 865.950 868.950 868.050 871.050 ;
        RECT 869.400 868.050 870.450 877.950 ;
        RECT 863.400 866.400 867.450 867.450 ;
        RECT 853.950 841.950 856.050 844.050 ;
        RECT 859.950 841.950 862.050 844.050 ;
        RECT 841.950 839.100 844.050 841.200 ;
        RECT 849.000 840.600 853.050 841.050 ;
        RECT 842.400 838.350 843.600 839.100 ;
        RECT 848.400 838.950 853.050 840.600 ;
        RECT 848.400 838.350 849.600 838.950 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 841.950 835.950 844.050 838.050 ;
        RECT 844.950 835.950 847.050 838.050 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 812.400 833.400 819.600 834.450 ;
        RECT 823.950 832.800 826.050 834.900 ;
        RECT 832.950 832.800 835.050 834.900 ;
        RECT 839.400 833.400 840.600 835.650 ;
        RECT 845.400 833.400 846.600 835.650 ;
        RECT 839.400 829.050 840.450 833.400 ;
        RECT 811.950 826.950 814.050 829.050 ;
        RECT 838.950 826.950 841.050 829.050 ;
        RECT 805.950 820.950 808.050 823.050 ;
        RECT 796.950 814.950 799.050 817.050 ;
        RECT 797.400 808.050 798.450 814.950 ;
        RECT 793.950 805.950 796.050 808.050 ;
        RECT 796.950 805.950 799.050 808.050 ;
        RECT 799.950 806.100 802.050 808.200 ;
        RECT 806.400 807.600 807.450 820.950 ;
        RECT 812.400 808.200 813.450 826.950 ;
        RECT 814.950 823.950 817.050 826.050 ;
        RECT 832.950 823.950 835.050 826.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 776.400 801.000 777.600 802.650 ;
        RECT 775.950 796.950 778.050 801.000 ;
        RECT 782.400 800.400 783.600 802.650 ;
        RECT 782.400 793.050 783.450 800.400 ;
        RECT 787.950 799.950 790.050 802.050 ;
        RECT 769.950 790.950 772.050 793.050 ;
        RECT 781.950 790.950 784.050 793.050 ;
        RECT 772.950 784.950 775.050 787.050 ;
        RECT 766.950 772.950 769.050 775.050 ;
        RECT 773.400 772.050 774.450 784.950 ;
        RECT 772.800 769.950 774.900 772.050 ;
        RECT 775.950 769.950 778.050 772.050 ;
        RECT 766.950 763.950 769.050 766.050 ;
        RECT 767.400 751.050 768.450 763.950 ;
        RECT 776.400 762.600 777.450 769.950 ;
        RECT 781.950 766.950 784.050 769.050 ;
        RECT 782.400 762.600 783.450 766.950 ;
        RECT 776.400 760.350 777.600 762.600 ;
        RECT 782.400 760.350 783.600 762.600 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 773.400 756.900 774.600 757.650 ;
        RECT 779.400 756.900 780.600 757.650 ;
        RECT 772.950 754.800 775.050 756.900 ;
        RECT 778.950 754.800 781.050 756.900 ;
        RECT 784.950 754.950 787.050 757.050 ;
        RECT 788.400 756.450 789.450 799.950 ;
        RECT 794.400 799.050 795.450 805.950 ;
        RECT 800.400 805.350 801.600 806.100 ;
        RECT 806.400 805.350 807.600 807.600 ;
        RECT 811.950 806.100 814.050 808.200 ;
        RECT 815.400 805.050 816.450 823.950 ;
        RECT 817.950 820.950 820.050 823.050 ;
        RECT 826.950 820.950 829.050 823.050 ;
        RECT 818.400 808.050 819.450 820.950 ;
        RECT 827.400 811.050 828.450 820.950 ;
        RECT 826.950 808.950 829.050 811.050 ;
        RECT 817.950 805.950 820.050 808.050 ;
        RECT 820.950 806.100 823.050 808.200 ;
        RECT 821.400 805.350 822.600 806.100 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 802.950 805.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 820.950 802.950 823.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 796.950 799.950 799.050 802.050 ;
        RECT 803.400 801.900 804.600 802.650 ;
        RECT 809.400 801.900 810.600 802.650 ;
        RECT 793.950 796.950 796.050 799.050 ;
        RECT 797.400 780.450 798.450 799.950 ;
        RECT 802.950 799.800 805.050 801.900 ;
        RECT 808.950 799.800 811.050 801.900 ;
        RECT 811.950 799.950 814.050 802.050 ;
        RECT 824.400 800.400 825.600 802.650 ;
        RECT 809.400 787.050 810.450 799.800 ;
        RECT 808.950 784.950 811.050 787.050 ;
        RECT 794.400 779.400 798.450 780.450 ;
        RECT 790.950 772.950 793.050 775.050 ;
        RECT 791.400 760.050 792.450 772.950 ;
        RECT 794.400 763.050 795.450 779.400 ;
        RECT 796.950 775.950 799.050 778.050 ;
        RECT 793.950 760.950 796.050 763.050 ;
        RECT 797.400 762.600 798.450 775.950 ;
        RECT 812.400 772.050 813.450 799.950 ;
        RECT 824.400 793.050 825.450 800.400 ;
        RECT 829.950 799.950 832.050 802.050 ;
        RECT 823.800 790.950 825.900 793.050 ;
        RECT 826.950 790.950 829.050 793.050 ;
        RECT 817.950 784.950 820.050 787.050 ;
        RECT 818.400 781.050 819.450 784.950 ;
        RECT 817.950 778.950 820.050 781.050 ;
        RECT 827.400 778.050 828.450 790.950 ;
        RECT 826.950 775.950 829.050 778.050 ;
        RECT 811.950 769.950 814.050 772.050 ;
        RECT 830.400 769.050 831.450 799.950 ;
        RECT 833.400 771.450 834.450 823.950 ;
        RECT 845.400 811.050 846.450 833.400 ;
        RECT 854.400 829.050 855.450 841.950 ;
        RECT 866.400 841.200 867.450 866.400 ;
        RECT 868.950 865.950 871.050 868.050 ;
        RECT 871.950 859.950 874.050 862.050 ;
        RECT 872.400 841.200 873.450 859.950 ;
        RECT 875.400 847.050 876.450 878.400 ;
        RECT 877.950 868.950 880.050 871.050 ;
        RECT 874.950 844.950 877.050 847.050 ;
        RECT 856.950 838.950 859.050 841.050 ;
        RECT 865.950 839.100 868.050 841.200 ;
        RECT 871.950 839.100 874.050 841.200 ;
        RECT 857.400 834.900 858.450 838.950 ;
        RECT 866.400 838.350 867.600 839.100 ;
        RECT 872.400 838.350 873.600 839.100 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 865.950 835.950 868.050 838.050 ;
        RECT 868.950 835.950 871.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 863.400 834.900 864.600 835.650 ;
        RECT 856.950 832.800 859.050 834.900 ;
        RECT 862.950 832.800 865.050 834.900 ;
        RECT 869.400 833.400 870.600 835.650 ;
        RECT 853.950 828.450 856.050 829.050 ;
        RECT 851.400 827.400 856.050 828.450 ;
        RECT 847.950 814.950 850.050 817.050 ;
        RECT 841.800 810.000 843.900 811.050 ;
        RECT 841.800 808.950 844.050 810.000 ;
        RECT 844.950 808.950 847.050 811.050 ;
        RECT 841.950 807.000 844.050 808.950 ;
        RECT 848.400 807.600 849.450 814.950 ;
        RECT 851.400 808.050 852.450 827.400 ;
        RECT 853.950 826.950 856.050 827.400 ;
        RECT 857.400 820.050 858.450 832.800 ;
        RECT 869.400 826.050 870.450 833.400 ;
        RECT 874.950 832.950 877.050 835.050 ;
        RECT 868.950 823.950 871.050 826.050 ;
        RECT 856.950 817.950 859.050 820.050 ;
        RECT 842.400 805.350 843.600 807.000 ;
        RECT 848.400 805.350 849.600 807.600 ;
        RECT 850.950 805.950 853.050 808.050 ;
        RECT 856.950 805.950 859.050 808.050 ;
        RECT 862.950 806.100 865.050 808.200 ;
        RECT 868.950 806.100 871.050 808.200 ;
        RECT 875.400 808.050 876.450 832.950 ;
        RECT 878.400 808.050 879.450 868.950 ;
        RECT 881.400 865.050 882.450 878.400 ;
        RECT 886.950 877.800 889.050 879.900 ;
        RECT 889.950 877.950 892.050 880.050 ;
        RECT 896.400 878.400 897.600 880.650 ;
        RECT 902.400 879.900 903.600 880.650 ;
        RECT 880.950 862.950 883.050 865.050 ;
        RECT 887.400 856.050 888.450 877.800 ;
        RECT 890.400 874.050 891.450 877.950 ;
        RECT 889.950 871.950 892.050 874.050 ;
        RECT 886.950 853.950 889.050 856.050 ;
        RECT 896.400 847.050 897.450 878.400 ;
        RECT 901.950 877.800 904.050 879.900 ;
        RECT 901.950 874.650 904.050 876.750 ;
        RECT 892.950 844.950 895.050 847.050 ;
        RECT 895.950 844.950 898.050 847.050 ;
        RECT 886.950 840.000 889.050 844.050 ;
        RECT 893.400 840.600 894.450 844.950 ;
        RECT 887.400 838.350 888.600 840.000 ;
        RECT 893.400 838.350 894.600 840.600 ;
        RECT 883.950 835.950 886.050 838.050 ;
        RECT 886.950 835.950 889.050 838.050 ;
        RECT 889.950 835.950 892.050 838.050 ;
        RECT 892.950 835.950 895.050 838.050 ;
        RECT 884.400 833.400 885.600 835.650 ;
        RECT 890.400 834.900 891.600 835.650 ;
        RECT 884.400 829.050 885.450 833.400 ;
        RECT 889.950 832.800 892.050 834.900 ;
        RECT 898.950 832.800 901.050 834.900 ;
        RECT 883.950 826.950 886.050 829.050 ;
        RECT 880.950 820.950 883.050 823.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 841.950 802.950 844.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 839.400 800.400 840.600 802.650 ;
        RECT 845.400 801.900 846.600 802.650 ;
        RECT 839.400 781.050 840.450 800.400 ;
        RECT 844.950 799.800 847.050 801.900 ;
        RECT 850.950 799.950 853.050 802.050 ;
        RECT 857.400 801.450 858.450 805.950 ;
        RECT 863.400 805.350 864.600 806.100 ;
        RECT 869.400 805.350 870.600 806.100 ;
        RECT 874.950 805.950 877.050 808.050 ;
        RECT 877.950 805.950 880.050 808.050 ;
        RECT 862.950 802.950 865.050 805.050 ;
        RECT 865.950 802.950 868.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 866.400 801.900 867.600 802.650 ;
        RECT 857.400 800.400 861.450 801.450 ;
        RECT 841.950 793.950 844.050 796.050 ;
        RECT 838.950 780.450 841.050 781.050 ;
        RECT 836.400 779.400 841.050 780.450 ;
        RECT 836.400 775.050 837.450 779.400 ;
        RECT 838.950 778.950 841.050 779.400 ;
        RECT 835.950 772.950 838.050 775.050 ;
        RECT 833.400 770.400 837.450 771.450 ;
        RECT 823.950 766.950 826.050 769.050 ;
        RECT 829.950 766.950 832.050 769.050 ;
        RECT 797.400 760.350 798.600 762.600 ;
        RECT 802.950 761.100 805.050 763.200 ;
        RECT 808.950 761.100 811.050 763.200 ;
        RECT 803.400 760.350 804.600 761.100 ;
        RECT 809.400 760.350 810.600 761.100 ;
        RECT 814.950 760.950 817.050 763.050 ;
        RECT 824.400 762.600 825.450 766.950 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 805.950 757.950 808.050 760.050 ;
        RECT 808.950 757.950 811.050 760.050 ;
        RECT 800.400 756.900 801.600 757.650 ;
        RECT 788.400 755.400 792.450 756.450 ;
        RECT 766.950 748.950 769.050 751.050 ;
        RECT 763.950 745.950 766.050 748.050 ;
        RECT 760.950 742.950 763.050 745.050 ;
        RECT 785.400 742.050 786.450 754.950 ;
        RECT 787.950 745.950 790.050 748.050 ;
        RECT 748.950 739.950 751.050 742.050 ;
        RECT 763.950 739.950 766.050 742.050 ;
        RECT 784.950 739.950 787.050 742.050 ;
        RECT 749.400 729.600 750.450 739.950 ;
        RECT 764.400 736.050 765.450 739.950 ;
        RECT 766.950 736.950 769.050 739.050 ;
        RECT 781.950 738.900 786.000 739.050 ;
        RECT 781.950 736.950 787.050 738.900 ;
        RECT 763.950 733.950 766.050 736.050 ;
        RECT 749.400 727.350 750.600 729.600 ;
        RECT 754.950 728.100 757.050 730.200 ;
        RECT 755.400 727.350 756.600 728.100 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 754.950 724.950 757.050 727.050 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 752.400 723.000 753.600 724.650 ;
        RECT 758.400 723.900 759.600 724.650 ;
        RECT 764.400 723.900 765.450 733.950 ;
        RECT 767.400 730.050 768.450 736.950 ;
        RECT 784.950 736.800 787.050 736.950 ;
        RECT 784.950 733.800 787.050 735.900 ;
        RECT 766.950 727.950 769.050 730.050 ;
        RECT 772.950 729.000 775.050 733.050 ;
        RECT 773.400 727.350 774.600 729.000 ;
        RECT 778.950 728.100 781.050 730.200 ;
        RECT 779.400 727.350 780.600 728.100 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 772.950 724.950 775.050 727.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 751.950 718.950 754.050 723.000 ;
        RECT 757.950 721.800 760.050 723.900 ;
        RECT 763.950 721.800 766.050 723.900 ;
        RECT 770.400 722.400 771.600 724.650 ;
        RECT 776.400 723.900 777.600 724.650 ;
        RECT 785.400 723.900 786.450 733.800 ;
        RECT 770.400 709.050 771.450 722.400 ;
        RECT 775.950 721.800 778.050 723.900 ;
        RECT 784.950 721.800 787.050 723.900 ;
        RECT 772.950 715.950 775.050 718.050 ;
        RECT 742.950 706.950 745.050 709.050 ;
        RECT 769.950 706.950 772.050 709.050 ;
        RECT 763.950 700.950 766.050 703.050 ;
        RECT 748.950 691.950 751.050 694.050 ;
        RECT 739.950 685.950 742.050 688.050 ;
        RECT 745.950 685.950 748.050 688.050 ;
        RECT 725.400 679.050 726.450 682.800 ;
        RECT 731.400 682.350 732.600 683.100 ;
        RECT 737.400 682.350 738.600 684.600 ;
        RECT 730.950 679.950 733.050 682.050 ;
        RECT 733.950 679.950 736.050 682.050 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 724.950 676.950 727.050 679.050 ;
        RECT 734.400 677.400 735.600 679.650 ;
        RECT 740.400 677.400 741.600 679.650 ;
        RECT 721.950 673.950 724.050 676.050 ;
        RECT 725.400 667.050 726.450 676.950 ;
        RECT 727.950 673.950 730.050 676.050 ;
        RECT 724.950 664.950 727.050 667.050 ;
        RECT 698.400 653.400 702.450 654.450 ;
        RECT 701.400 652.200 702.450 653.400 ;
        RECT 712.950 652.950 715.050 655.050 ;
        RECT 700.950 650.100 703.050 652.200 ;
        RECT 706.950 650.100 709.050 652.200 ;
        RECT 701.400 649.350 702.600 650.100 ;
        RECT 707.400 649.350 708.600 650.100 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 706.950 646.950 709.050 649.050 ;
        RECT 698.400 645.900 699.600 646.650 ;
        RECT 697.950 643.800 700.050 645.900 ;
        RECT 704.400 645.000 705.600 646.650 ;
        RECT 691.950 640.950 694.050 643.050 ;
        RECT 703.950 640.950 706.050 645.000 ;
        RECT 682.950 637.950 685.050 640.050 ;
        RECT 697.950 637.950 700.050 640.050 ;
        RECT 670.950 610.950 673.050 613.050 ;
        RECT 673.950 610.950 676.050 613.050 ;
        RECT 679.950 610.950 682.050 613.050 ;
        RECT 668.400 604.350 669.600 606.600 ;
        RECT 673.950 605.100 676.050 607.200 ;
        RECT 674.400 604.350 675.600 605.100 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 671.400 600.900 672.600 601.650 ;
        RECT 680.400 600.900 681.450 610.950 ;
        RECT 664.950 600.450 667.050 600.900 ;
        RECT 662.400 599.400 667.050 600.450 ;
        RECT 664.950 598.800 667.050 599.400 ;
        RECT 670.950 598.800 673.050 600.900 ;
        RECT 679.950 598.800 682.050 600.900 ;
        RECT 661.950 595.800 664.050 597.900 ;
        RECT 662.400 559.050 663.450 595.800 ;
        RECT 665.400 574.050 666.450 598.800 ;
        RECT 676.950 592.950 679.050 595.050 ;
        RECT 664.950 571.950 667.050 574.050 ;
        RECT 670.950 573.000 673.050 577.050 ;
        RECT 677.400 574.200 678.450 592.950 ;
        RECT 671.400 571.350 672.600 573.000 ;
        RECT 676.950 572.100 679.050 574.200 ;
        RECT 677.400 571.350 678.600 572.100 ;
        RECT 683.400 571.050 684.450 637.950 ;
        RECT 688.950 634.950 691.050 637.050 ;
        RECT 685.950 610.950 688.050 613.050 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 676.950 568.950 679.050 571.050 ;
        RECT 682.950 568.950 685.050 571.050 ;
        RECT 668.400 566.400 669.600 568.650 ;
        RECT 674.400 567.000 675.600 568.650 ;
        RECT 668.400 559.050 669.450 566.400 ;
        RECT 670.950 562.950 673.050 565.050 ;
        RECT 673.950 562.950 676.050 567.000 ;
        RECT 679.950 562.950 682.050 565.050 ;
        RECT 661.950 556.950 664.050 559.050 ;
        RECT 667.950 556.950 670.050 559.050 ;
        RECT 658.950 538.950 661.050 541.050 ;
        RECT 646.950 532.950 649.050 535.050 ;
        RECT 655.950 532.950 658.050 535.050 ;
        RECT 640.950 527.100 643.050 529.200 ;
        RECT 647.400 528.600 648.450 532.950 ;
        RECT 652.950 529.950 655.050 532.050 ;
        RECT 641.400 526.350 642.600 527.100 ;
        RECT 647.400 526.350 648.600 528.600 ;
        RECT 640.950 523.950 643.050 526.050 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 644.400 522.900 645.600 523.650 ;
        RECT 643.950 520.800 646.050 522.900 ;
        RECT 649.950 505.950 652.050 508.050 ;
        RECT 625.950 493.950 628.050 496.050 ;
        RECT 628.950 495.000 631.050 499.050 ;
        RECT 634.950 496.950 637.050 499.050 ;
        RECT 650.400 495.600 651.450 505.950 ;
        RECT 653.400 505.050 654.450 529.950 ;
        RECT 656.400 511.050 657.450 532.950 ;
        RECT 664.950 527.100 667.050 529.200 ;
        RECT 671.400 528.600 672.450 562.950 ;
        RECT 673.950 559.800 676.050 561.900 ;
        RECT 674.400 529.050 675.450 559.800 ;
        RECT 676.950 547.950 679.050 550.050 ;
        RECT 665.400 526.350 666.600 527.100 ;
        RECT 671.400 526.350 672.600 528.600 ;
        RECT 673.950 526.950 676.050 529.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 662.400 521.400 663.600 523.650 ;
        RECT 668.400 521.400 669.600 523.650 ;
        RECT 659.400 511.050 660.450 520.950 ;
        RECT 662.400 520.050 663.450 521.400 ;
        RECT 661.950 517.950 664.050 520.050 ;
        RECT 655.800 508.950 657.900 511.050 ;
        RECT 658.950 508.950 661.050 511.050 ;
        RECT 652.950 502.950 655.050 505.050 ;
        RECT 635.400 495.450 636.600 495.600 ;
        RECT 629.400 493.350 630.600 495.000 ;
        RECT 635.400 494.400 642.450 495.450 ;
        RECT 635.400 493.350 636.600 494.400 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 631.950 490.950 634.050 493.050 ;
        RECT 634.950 490.950 637.050 493.050 ;
        RECT 632.400 488.400 633.600 490.650 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 619.950 466.950 622.050 469.050 ;
        RECT 632.400 466.050 633.450 488.400 ;
        RECT 631.950 463.950 634.050 466.050 ;
        RECT 616.950 460.950 619.050 463.050 ;
        RECT 641.400 460.050 642.450 494.400 ;
        RECT 650.400 493.350 651.600 495.600 ;
        RECT 658.950 493.950 661.050 496.050 ;
        RECT 646.950 490.950 649.050 493.050 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 652.950 490.950 655.050 493.050 ;
        RECT 647.400 489.900 648.600 490.650 ;
        RECT 646.950 487.800 649.050 489.900 ;
        RECT 653.400 488.400 654.600 490.650 ;
        RECT 659.400 489.900 660.450 493.950 ;
        RECT 653.400 486.450 654.450 488.400 ;
        RECT 658.950 487.800 661.050 489.900 ;
        RECT 650.400 485.400 654.450 486.450 ;
        RECT 650.400 472.050 651.450 485.400 ;
        RECT 662.400 481.050 663.450 517.950 ;
        RECT 668.400 505.050 669.450 521.400 ;
        RECT 673.950 517.950 676.050 523.050 ;
        RECT 677.400 514.050 678.450 547.950 ;
        RECT 680.400 529.050 681.450 562.950 ;
        RECT 686.400 535.050 687.450 610.950 ;
        RECT 689.400 606.600 690.450 634.950 ;
        RECT 698.400 628.050 699.450 637.950 ;
        RECT 697.950 625.950 700.050 628.050 ;
        RECT 700.950 619.950 703.050 622.050 ;
        RECT 697.950 610.950 700.050 613.050 ;
        RECT 689.400 604.350 690.600 606.600 ;
        RECT 689.100 601.950 691.200 604.050 ;
        RECT 694.500 601.950 696.600 604.050 ;
        RECT 695.400 600.900 696.600 601.650 ;
        RECT 694.950 598.800 697.050 600.900 ;
        RECT 695.400 577.050 696.450 598.800 ;
        RECT 688.950 573.000 691.050 577.050 ;
        RECT 694.950 574.950 697.050 577.050 ;
        RECT 689.400 571.350 690.600 573.000 ;
        RECT 689.400 568.950 691.500 571.050 ;
        RECT 694.800 568.950 696.900 571.050 ;
        RECT 695.400 566.400 696.600 568.650 ;
        RECT 695.400 553.050 696.450 566.400 ;
        RECT 694.950 550.950 697.050 553.050 ;
        RECT 694.950 541.950 697.050 544.050 ;
        RECT 685.950 532.950 688.050 535.050 ;
        RECT 679.950 526.950 682.050 529.050 ;
        RECT 685.950 528.000 688.050 531.900 ;
        RECT 691.950 528.000 694.050 532.050 ;
        RECT 695.400 529.050 696.450 541.950 ;
        RECT 686.400 526.350 687.600 528.000 ;
        RECT 692.400 526.350 693.600 528.000 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 679.950 520.950 682.050 523.050 ;
        RECT 683.400 521.400 684.600 523.650 ;
        RECT 689.400 522.900 690.600 523.650 ;
        RECT 676.950 511.950 679.050 514.050 ;
        RECT 667.950 502.950 670.050 505.050 ;
        RECT 664.950 499.950 667.050 502.050 ;
        RECT 665.400 496.050 666.450 499.950 ;
        RECT 664.950 493.950 667.050 496.050 ;
        RECT 670.950 494.100 673.050 496.200 ;
        RECT 671.400 493.350 672.600 494.100 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 664.950 487.950 667.050 490.050 ;
        RECT 668.400 489.900 669.600 490.650 ;
        RECT 652.950 478.950 655.050 481.050 ;
        RECT 661.950 478.950 664.050 481.050 ;
        RECT 649.950 469.950 652.050 472.050 ;
        RECT 640.950 457.950 643.050 460.050 ;
        RECT 649.950 457.950 652.050 460.050 ;
        RECT 613.950 454.950 616.050 457.050 ;
        RECT 637.950 454.950 640.050 457.050 ;
        RECT 608.400 452.400 612.450 453.450 ;
        RECT 604.950 448.950 607.050 451.050 ;
        RECT 608.400 450.600 609.450 452.400 ;
        RECT 608.400 448.350 609.600 450.600 ;
        RECT 613.950 449.100 616.050 451.200 ;
        RECT 619.950 449.100 622.050 451.200 ;
        RECT 631.950 449.100 634.050 451.200 ;
        RECT 638.400 450.600 639.450 454.950 ;
        RECT 614.400 448.350 615.600 449.100 ;
        RECT 620.400 448.350 621.600 449.100 ;
        RECT 632.400 448.350 633.600 449.100 ;
        RECT 638.400 448.350 639.600 450.600 ;
        RECT 646.950 449.100 649.050 451.200 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 604.950 442.950 607.050 445.050 ;
        RECT 611.400 444.000 612.600 445.650 ;
        RECT 601.950 439.950 604.050 442.050 ;
        RECT 598.950 433.950 601.050 436.050 ;
        RECT 589.950 424.950 592.050 427.050 ;
        RECT 595.950 424.950 598.050 427.050 ;
        RECT 601.950 424.950 604.050 427.050 ;
        RECT 586.950 406.950 589.050 409.050 ;
        RECT 590.400 403.050 591.450 424.950 ;
        RECT 592.950 418.950 595.050 421.050 ;
        RECT 580.950 400.950 583.050 403.050 ;
        RECT 589.950 400.950 592.050 403.050 ;
        RECT 577.950 388.950 580.050 391.050 ;
        RECT 581.400 388.050 582.450 400.950 ;
        RECT 580.950 385.950 583.050 388.050 ;
        RECT 586.950 379.950 589.050 382.050 ;
        RECT 574.950 373.950 577.050 376.050 ;
        RECT 587.400 372.600 588.450 379.950 ;
        RECT 578.400 372.450 579.600 372.600 ;
        RECT 575.400 372.000 579.600 372.450 ;
        RECT 574.950 371.400 579.600 372.000 ;
        RECT 574.950 367.950 577.050 371.400 ;
        RECT 578.400 370.350 579.600 371.400 ;
        RECT 587.400 370.350 588.600 372.600 ;
        RECT 589.950 370.950 592.050 373.050 ;
        RECT 578.100 367.950 580.200 370.050 ;
        RECT 583.500 367.950 585.600 370.050 ;
        RECT 586.800 367.950 588.900 370.050 ;
        RECT 584.400 365.400 585.600 367.650 ;
        RECT 571.950 355.950 574.050 358.050 ;
        RECT 556.950 352.950 559.050 355.050 ;
        RECT 562.950 352.950 565.050 355.050 ;
        RECT 553.950 346.950 556.050 349.050 ;
        RECT 557.400 345.450 558.450 352.950 ;
        RECT 562.950 346.950 565.050 349.050 ;
        RECT 554.400 345.000 558.450 345.450 ;
        RECT 553.950 344.400 558.450 345.000 ;
        RECT 553.950 340.950 556.050 344.400 ;
        RECT 545.400 338.400 549.450 339.450 ;
        RECT 532.950 334.950 535.050 337.050 ;
        RECT 535.950 334.950 538.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 536.400 333.900 537.600 334.650 ;
        RECT 535.950 331.800 538.050 333.900 ;
        RECT 542.400 332.400 543.600 334.650 ;
        RECT 532.950 328.950 535.050 331.050 ;
        RECT 529.950 316.950 532.050 319.050 ;
        RECT 530.400 313.050 531.450 316.950 ;
        RECT 529.950 310.950 532.050 313.050 ;
        RECT 526.950 292.950 529.050 295.050 ;
        RECT 530.400 294.600 531.450 310.950 ;
        RECT 533.400 301.050 534.450 328.950 ;
        RECT 535.950 322.950 538.050 325.050 ;
        RECT 532.950 298.950 535.050 301.050 ;
        RECT 536.400 295.200 537.450 322.950 ;
        RECT 530.400 292.350 531.600 294.600 ;
        RECT 535.950 293.100 538.050 295.200 ;
        RECT 536.400 292.350 537.600 293.100 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 535.950 289.950 538.050 292.050 ;
        RECT 533.400 288.900 534.600 289.650 ;
        RECT 542.400 289.050 543.450 332.400 ;
        RECT 544.950 331.950 547.050 334.050 ;
        RECT 545.400 295.050 546.450 331.950 ;
        RECT 548.400 316.050 549.450 338.400 ;
        RECT 550.950 337.950 553.050 340.050 ;
        RECT 556.950 338.100 559.050 343.050 ;
        RECT 563.400 340.200 564.450 346.950 ;
        RECT 562.950 338.100 565.050 340.200 ;
        RECT 557.400 337.350 558.600 338.100 ;
        RECT 563.400 337.350 564.600 338.100 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 554.400 333.900 555.600 334.650 ;
        RECT 553.950 331.800 556.050 333.900 ;
        RECT 560.400 332.400 561.600 334.650 ;
        RECT 566.400 332.400 567.600 334.650 ;
        RECT 550.950 322.950 553.050 325.050 ;
        RECT 547.950 313.950 550.050 316.050 ;
        RECT 551.400 298.050 552.450 322.950 ;
        RECT 554.400 319.050 555.450 331.800 ;
        RECT 560.400 325.050 561.450 332.400 ;
        RECT 566.400 330.450 567.450 332.400 ;
        RECT 568.950 331.950 571.050 334.050 ;
        RECT 563.400 329.400 567.450 330.450 ;
        RECT 563.400 325.050 564.450 329.400 ;
        RECT 569.400 327.450 570.450 331.950 ;
        RECT 566.400 326.400 570.450 327.450 ;
        RECT 559.800 322.950 561.900 325.050 ;
        RECT 562.950 322.950 565.050 325.050 ;
        RECT 553.950 316.950 556.050 319.050 ;
        RECT 563.400 316.050 564.450 322.950 ;
        RECT 562.950 313.950 565.050 316.050 ;
        RECT 556.950 307.950 559.050 310.050 ;
        RECT 550.950 295.950 553.050 298.050 ;
        RECT 544.950 292.950 547.050 295.050 ;
        RECT 551.400 294.600 552.450 295.950 ;
        RECT 557.400 294.600 558.450 307.950 ;
        RECT 566.400 307.050 567.450 326.400 ;
        RECT 559.950 304.950 562.050 307.050 ;
        RECT 565.950 304.950 568.050 307.050 ;
        RECT 560.400 298.050 561.450 304.950 ;
        RECT 572.400 304.050 573.450 355.950 ;
        RECT 574.950 343.950 577.050 346.050 ;
        RECT 575.400 313.050 576.450 343.950 ;
        RECT 584.400 343.050 585.450 365.400 ;
        RECT 590.400 358.050 591.450 370.950 ;
        RECT 589.950 355.950 592.050 358.050 ;
        RECT 590.400 346.050 591.450 355.950 ;
        RECT 589.950 343.950 592.050 346.050 ;
        RECT 583.950 339.000 586.050 343.050 ;
        RECT 590.400 339.600 591.450 343.950 ;
        RECT 593.400 343.050 594.450 418.950 ;
        RECT 602.400 417.600 603.450 424.950 ;
        RECT 605.400 421.050 606.450 442.950 ;
        RECT 607.950 439.950 610.050 442.050 ;
        RECT 610.950 439.950 613.050 444.000 ;
        RECT 617.400 443.400 618.600 445.650 ;
        RECT 604.950 418.950 607.050 421.050 ;
        RECT 602.400 415.350 603.600 417.600 ;
        RECT 596.100 412.950 598.200 415.050 ;
        RECT 601.500 412.950 603.600 415.050 ;
        RECT 604.800 412.950 606.900 415.050 ;
        RECT 596.400 411.000 597.600 412.650 ;
        RECT 605.400 411.900 606.600 412.650 ;
        RECT 595.950 406.950 598.050 411.000 ;
        RECT 604.950 409.800 607.050 411.900 ;
        RECT 608.400 409.050 609.450 439.950 ;
        RECT 601.950 406.950 604.050 409.050 ;
        RECT 607.950 406.950 610.050 409.050 ;
        RECT 598.950 397.950 601.050 400.050 ;
        RECT 595.950 394.950 598.050 397.050 ;
        RECT 596.400 367.050 597.450 394.950 ;
        RECT 599.400 373.050 600.450 397.950 ;
        RECT 602.400 385.050 603.450 406.950 ;
        RECT 608.400 396.450 609.450 406.950 ;
        RECT 611.400 400.050 612.450 439.950 ;
        RECT 617.400 430.050 618.450 443.400 ;
        RECT 622.950 439.950 625.050 445.050 ;
        RECT 626.400 439.050 627.450 445.950 ;
        RECT 635.400 443.400 636.600 445.650 ;
        RECT 641.400 443.400 642.600 445.650 ;
        RECT 647.400 445.050 648.450 449.100 ;
        RECT 628.950 441.450 633.000 442.050 ;
        RECT 628.950 439.950 633.450 441.450 ;
        RECT 625.800 436.950 627.900 439.050 ;
        RECT 628.950 436.800 631.050 438.900 ;
        RECT 629.400 433.050 630.450 436.800 ;
        RECT 622.950 430.950 625.050 433.050 ;
        RECT 628.950 430.950 631.050 433.050 ;
        RECT 616.950 427.950 619.050 430.050 ;
        RECT 613.950 421.950 616.050 424.050 ;
        RECT 623.400 423.450 624.450 430.950 ;
        RECT 632.400 426.450 633.450 439.950 ;
        RECT 635.400 430.050 636.450 443.400 ;
        RECT 641.400 433.050 642.450 443.400 ;
        RECT 646.950 442.950 649.050 445.050 ;
        RECT 650.400 436.050 651.450 457.950 ;
        RECT 653.400 451.050 654.450 478.950 ;
        RECT 658.950 472.950 661.050 475.050 ;
        RECT 652.950 448.950 655.050 451.050 ;
        RECT 659.400 450.600 660.450 472.950 ;
        RECT 665.400 454.200 666.450 487.950 ;
        RECT 667.950 487.800 670.050 489.900 ;
        RECT 674.400 488.400 675.600 490.650 ;
        RECT 674.400 486.450 675.450 488.400 ;
        RECT 680.400 487.050 681.450 520.950 ;
        RECT 683.400 514.050 684.450 521.400 ;
        RECT 688.950 520.800 691.050 522.900 ;
        RECT 694.950 520.950 697.050 523.050 ;
        RECT 682.950 511.950 685.050 514.050 ;
        RECT 691.950 508.950 694.050 511.050 ;
        RECT 685.950 495.000 688.050 499.050 ;
        RECT 692.400 495.600 693.450 508.950 ;
        RECT 695.400 508.050 696.450 520.950 ;
        RECT 698.400 511.050 699.450 610.950 ;
        RECT 701.400 601.050 702.450 619.950 ;
        RECT 713.400 613.050 714.450 652.950 ;
        RECT 715.950 649.950 718.050 652.050 ;
        RECT 721.950 650.100 724.050 652.200 ;
        RECT 728.400 651.600 729.450 673.950 ;
        RECT 716.400 622.050 717.450 649.950 ;
        RECT 722.400 649.350 723.600 650.100 ;
        RECT 728.400 649.350 729.600 651.600 ;
        RECT 734.400 651.450 735.450 677.400 ;
        RECT 740.400 673.050 741.450 677.400 ;
        RECT 742.950 676.800 745.050 678.900 ;
        RECT 739.950 670.950 742.050 673.050 ;
        RECT 739.950 664.950 742.050 667.050 ;
        RECT 740.400 652.050 741.450 664.950 ;
        RECT 734.400 650.400 738.450 651.450 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 725.400 645.900 726.600 646.650 ;
        RECT 724.950 643.800 727.050 645.900 ;
        RECT 731.400 644.400 732.600 646.650 ;
        RECT 731.400 634.050 732.450 644.400 ;
        RECT 733.950 643.950 736.050 646.050 ;
        RECT 737.400 645.900 738.450 650.400 ;
        RECT 739.950 649.950 742.050 652.050 ;
        RECT 743.400 651.450 744.450 676.800 ;
        RECT 746.400 655.050 747.450 685.950 ;
        RECT 749.400 667.050 750.450 691.950 ;
        RECT 757.950 683.100 760.050 685.200 ;
        RECT 758.400 682.350 759.600 683.100 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 755.400 678.900 756.600 679.650 ;
        RECT 754.950 676.800 757.050 678.900 ;
        RECT 764.400 670.050 765.450 700.950 ;
        RECT 766.950 694.950 769.050 697.050 ;
        RECT 763.950 667.950 766.050 670.050 ;
        RECT 748.950 664.950 751.050 667.050 ;
        RECT 751.950 655.950 754.050 658.050 ;
        RECT 745.950 652.950 748.050 655.050 ;
        RECT 752.400 651.600 753.450 655.950 ;
        RECT 746.400 651.450 747.600 651.600 ;
        RECT 743.400 650.400 747.600 651.450 ;
        RECT 746.400 649.350 747.600 650.400 ;
        RECT 752.400 649.350 753.600 651.600 ;
        RECT 760.950 649.950 763.050 652.050 ;
        RECT 763.950 650.100 766.050 652.200 ;
        RECT 767.400 652.050 768.450 694.950 ;
        RECT 773.400 685.200 774.450 715.950 ;
        RECT 785.400 685.200 786.450 721.800 ;
        RECT 772.950 683.100 775.050 685.200 ;
        RECT 778.950 683.100 781.050 685.200 ;
        RECT 784.950 683.100 787.050 685.200 ;
        RECT 773.400 682.350 774.600 683.100 ;
        RECT 779.400 682.350 780.600 683.100 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 775.950 679.950 778.050 682.050 ;
        RECT 778.950 679.950 781.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 776.400 678.000 777.600 679.650 ;
        RECT 775.950 673.950 778.050 678.000 ;
        RECT 782.400 677.400 783.600 679.650 ;
        RECT 788.400 679.050 789.450 745.950 ;
        RECT 791.400 745.050 792.450 755.400 ;
        RECT 799.950 754.800 802.050 756.900 ;
        RECT 806.400 756.000 807.600 757.650 ;
        RECT 802.950 751.950 805.050 754.050 ;
        RECT 805.950 751.950 808.050 756.000 ;
        RECT 811.950 754.950 814.050 757.050 ;
        RECT 790.950 742.950 793.050 745.050 ;
        RECT 790.950 736.950 796.050 739.050 ;
        RECT 796.950 736.950 799.050 739.050 ;
        RECT 803.400 738.450 804.450 751.950 ;
        RECT 805.950 742.950 808.050 745.050 ;
        RECT 800.400 738.000 804.450 738.450 ;
        RECT 799.950 737.400 804.450 738.000 ;
        RECT 797.400 729.600 798.450 736.950 ;
        RECT 799.950 736.050 802.050 737.400 ;
        RECT 799.800 735.000 802.050 736.050 ;
        RECT 799.800 733.950 801.900 735.000 ;
        RECT 802.950 733.950 805.050 736.050 ;
        RECT 803.400 730.200 804.450 733.950 ;
        RECT 797.400 727.350 798.600 729.600 ;
        RECT 802.950 728.100 805.050 730.200 ;
        RECT 806.400 730.050 807.450 742.950 ;
        RECT 812.400 736.050 813.450 754.950 ;
        RECT 815.400 754.050 816.450 760.950 ;
        RECT 824.400 760.350 825.600 762.600 ;
        RECT 829.950 761.100 832.050 765.900 ;
        RECT 830.400 760.350 831.600 761.100 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 821.400 756.000 822.600 757.650 ;
        RECT 827.400 756.900 828.600 757.650 ;
        RECT 814.950 751.950 817.050 754.050 ;
        RECT 820.950 751.950 823.050 756.000 ;
        RECT 826.950 754.800 829.050 756.900 ;
        RECT 829.950 742.950 832.050 745.050 ;
        RECT 811.950 733.950 814.050 736.050 ;
        RECT 820.950 733.950 823.050 736.050 ;
        RECT 826.950 733.950 829.050 736.050 ;
        RECT 808.950 730.950 811.050 733.050 ;
        RECT 803.400 727.350 804.600 728.100 ;
        RECT 805.950 727.950 808.050 730.050 ;
        RECT 793.950 724.950 796.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 794.400 722.400 795.600 724.650 ;
        RECT 800.400 723.900 801.600 724.650 ;
        RECT 775.950 667.950 778.050 670.050 ;
        RECT 776.400 652.200 777.450 667.950 ;
        RECT 739.950 646.800 742.050 648.900 ;
        RECT 745.950 646.950 748.050 649.050 ;
        RECT 748.950 646.950 751.050 649.050 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 734.400 640.050 735.450 643.950 ;
        RECT 736.950 643.800 739.050 645.900 ;
        RECT 733.950 637.950 736.050 640.050 ;
        RECT 730.950 631.950 733.050 634.050 ;
        RECT 715.950 619.950 718.050 622.050 ;
        RECT 724.950 619.950 727.050 622.050 ;
        RECT 715.950 613.950 718.050 616.050 ;
        RECT 712.950 610.950 715.050 613.050 ;
        RECT 716.400 606.600 717.450 613.950 ;
        RECT 716.400 604.350 717.600 606.600 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 715.950 601.950 718.050 604.050 ;
        RECT 718.950 601.950 721.050 604.050 ;
        RECT 700.950 598.950 703.050 601.050 ;
        RECT 713.400 600.900 714.600 601.650 ;
        RECT 712.950 598.800 715.050 600.900 ;
        RECT 719.400 600.000 720.600 601.650 ;
        RECT 718.950 595.950 721.050 600.000 ;
        RECT 721.950 598.950 724.050 601.050 ;
        RECT 725.400 600.900 726.450 619.950 ;
        RECT 740.400 610.050 741.450 646.800 ;
        RECT 749.400 645.900 750.600 646.650 ;
        RECT 748.950 643.800 751.050 645.900 ;
        RECT 755.400 645.000 756.600 646.650 ;
        RECT 761.400 645.900 762.450 649.950 ;
        RECT 754.950 640.950 757.050 645.000 ;
        RECT 760.950 643.800 763.050 645.900 ;
        RECT 764.400 622.050 765.450 650.100 ;
        RECT 766.950 649.950 769.050 652.050 ;
        RECT 769.950 650.100 772.050 652.200 ;
        RECT 775.950 650.100 778.050 652.200 ;
        RECT 770.400 649.350 771.600 650.100 ;
        RECT 776.400 649.350 777.600 650.100 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 775.950 646.950 778.050 649.050 ;
        RECT 766.950 643.950 769.050 646.050 ;
        RECT 773.400 644.400 774.600 646.650 ;
        RECT 763.950 619.950 766.050 622.050 ;
        RECT 757.950 613.950 760.050 616.050 ;
        RECT 727.950 605.100 730.050 610.050 ;
        RECT 739.950 607.950 742.050 610.050 ;
        RECT 745.950 607.950 748.050 610.050 ;
        RECT 733.950 605.100 736.050 607.200 ;
        RECT 741.000 606.600 745.050 607.050 ;
        RECT 734.400 604.350 735.600 605.100 ;
        RECT 740.400 604.950 745.050 606.600 ;
        RECT 740.400 604.350 741.600 604.950 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 733.950 601.950 736.050 604.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 718.950 577.950 721.050 580.050 ;
        RECT 709.950 572.100 712.050 574.200 ;
        RECT 710.400 571.350 711.600 572.100 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 701.400 546.450 702.450 568.950 ;
        RECT 713.400 567.900 714.600 568.650 ;
        RECT 712.950 565.800 715.050 567.900 ;
        RECT 701.400 545.400 705.450 546.450 ;
        RECT 700.950 541.950 703.050 544.050 ;
        RECT 701.400 538.050 702.450 541.950 ;
        RECT 704.400 541.050 705.450 545.400 ;
        RECT 703.950 538.950 706.050 541.050 ;
        RECT 700.950 535.950 703.050 538.050 ;
        RECT 701.400 517.050 702.450 535.950 ;
        RECT 703.950 532.950 706.050 535.050 ;
        RECT 704.400 529.050 705.450 532.950 ;
        RECT 713.400 529.200 714.450 565.800 ;
        RECT 715.950 550.950 718.050 553.050 ;
        RECT 716.400 532.050 717.450 550.950 ;
        RECT 719.400 537.450 720.450 577.950 ;
        RECT 722.400 568.050 723.450 598.950 ;
        RECT 724.950 598.800 727.050 600.900 ;
        RECT 731.400 600.000 732.600 601.650 ;
        RECT 725.400 574.200 726.450 598.800 ;
        RECT 730.950 595.950 733.050 600.000 ;
        RECT 737.400 599.400 738.600 601.650 ;
        RECT 737.400 595.050 738.450 599.400 ;
        RECT 746.400 598.050 747.450 607.950 ;
        RECT 748.950 604.950 751.050 607.050 ;
        RECT 758.400 606.600 759.450 613.950 ;
        RECT 745.950 597.450 748.050 598.050 ;
        RECT 743.400 596.400 748.050 597.450 ;
        RECT 736.950 592.950 739.050 595.050 ;
        RECT 733.950 577.950 736.050 580.050 ;
        RECT 724.950 573.450 727.050 574.200 ;
        RECT 734.400 573.600 735.450 577.950 ;
        RECT 739.950 574.950 742.050 580.050 ;
        RECT 728.400 573.450 729.600 573.600 ;
        RECT 724.950 572.400 729.600 573.450 ;
        RECT 724.950 572.100 727.050 572.400 ;
        RECT 728.400 571.350 729.600 572.400 ;
        RECT 734.400 571.350 735.600 573.600 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 733.950 568.950 736.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 721.950 565.950 724.050 568.050 ;
        RECT 731.400 567.900 732.600 568.650 ;
        RECT 737.400 567.900 738.600 568.650 ;
        RECT 730.950 565.800 733.050 567.900 ;
        RECT 736.950 565.800 739.050 567.900 ;
        RECT 724.950 556.950 727.050 559.050 ;
        RECT 725.400 550.050 726.450 556.950 ;
        RECT 727.950 553.950 730.050 556.050 ;
        RECT 724.950 547.950 727.050 550.050 ;
        RECT 719.400 536.400 723.450 537.450 ;
        RECT 718.950 532.950 721.050 535.050 ;
        RECT 715.950 529.950 718.050 532.050 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 712.950 527.100 715.050 529.200 ;
        RECT 719.400 529.050 720.450 532.950 ;
        RECT 713.400 526.350 714.600 527.100 ;
        RECT 718.950 526.950 721.050 529.050 ;
        RECT 722.400 526.050 723.450 536.400 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 715.950 523.950 718.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 703.950 520.950 706.050 523.050 ;
        RECT 710.400 522.900 711.600 523.650 ;
        RECT 700.950 514.950 703.050 517.050 ;
        RECT 704.400 514.050 705.450 520.950 ;
        RECT 709.950 520.800 712.050 522.900 ;
        RECT 716.400 521.400 717.600 523.650 ;
        RECT 718.950 522.900 723.000 523.050 ;
        RECT 709.950 514.950 712.050 517.050 ;
        RECT 703.950 511.950 706.050 514.050 ;
        RECT 697.950 508.950 700.050 511.050 ;
        RECT 694.950 505.950 697.050 508.050 ;
        RECT 697.950 502.950 700.050 505.050 ;
        RECT 703.950 502.950 706.050 505.050 ;
        RECT 686.400 493.350 687.600 495.000 ;
        RECT 692.400 493.350 693.600 495.600 ;
        RECT 698.400 495.450 699.450 502.950 ;
        RECT 704.400 496.200 705.450 502.950 ;
        RECT 710.400 496.200 711.450 514.950 ;
        RECT 716.400 514.050 717.450 521.400 ;
        RECT 718.950 520.950 724.050 522.900 ;
        RECT 721.950 520.800 724.050 520.950 ;
        RECT 718.950 517.800 721.050 519.900 ;
        RECT 715.950 511.950 718.050 514.050 ;
        RECT 719.400 498.450 720.450 517.800 ;
        RECT 721.950 502.950 724.050 505.050 ;
        RECT 716.400 497.400 720.450 498.450 ;
        RECT 698.400 494.400 702.450 495.450 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 694.950 490.950 697.050 493.050 ;
        RECT 689.400 488.400 690.600 490.650 ;
        RECT 695.400 489.900 696.600 490.650 ;
        RECT 671.400 485.400 675.450 486.450 ;
        RECT 667.950 475.950 670.050 478.050 ;
        RECT 668.400 466.050 669.450 475.950 ;
        RECT 667.950 463.950 670.050 466.050 ;
        RECT 667.950 460.800 670.050 462.900 ;
        RECT 668.400 457.050 669.450 460.800 ;
        RECT 667.950 456.450 670.050 457.050 ;
        RECT 671.400 456.450 672.450 485.400 ;
        RECT 679.950 484.950 682.050 487.050 ;
        RECT 682.950 481.950 685.050 484.050 ;
        RECT 679.950 472.950 682.050 475.050 ;
        RECT 680.400 469.050 681.450 472.950 ;
        RECT 679.950 466.950 682.050 469.050 ;
        RECT 667.950 455.400 672.450 456.450 ;
        RECT 667.950 454.950 670.050 455.400 ;
        RECT 676.950 454.950 679.050 457.050 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 664.950 452.100 667.050 454.200 ;
        RECT 670.950 451.800 673.050 453.900 ;
        RECT 659.400 448.350 660.600 450.600 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 665.400 448.350 666.600 448.950 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 656.400 445.050 657.600 445.650 ;
        RECT 652.950 443.400 657.600 445.050 ;
        RECT 662.400 444.900 663.600 445.650 ;
        RECT 652.950 442.950 657.000 443.400 ;
        RECT 653.400 439.050 654.450 442.950 ;
        RECT 661.950 442.800 664.050 444.900 ;
        RECT 667.950 442.950 670.050 445.050 ;
        RECT 664.950 439.950 667.050 442.050 ;
        RECT 652.950 436.950 655.050 439.050 ;
        RECT 643.950 433.950 646.050 436.050 ;
        RECT 649.950 433.950 652.050 436.050 ;
        RECT 658.950 433.950 661.050 436.050 ;
        RECT 640.950 430.950 643.050 433.050 ;
        RECT 634.950 427.950 637.050 430.050 ;
        RECT 644.400 429.450 645.450 433.950 ;
        RECT 641.400 428.400 645.450 429.450 ;
        RECT 632.400 425.400 636.450 426.450 ;
        RECT 620.400 422.400 624.450 423.450 ;
        RECT 614.400 418.050 615.450 421.950 ;
        RECT 620.400 418.050 621.450 422.400 ;
        RECT 631.950 421.950 634.050 424.050 ;
        RECT 613.950 415.950 616.050 418.050 ;
        RECT 616.950 417.600 621.450 418.050 ;
        RECT 616.950 415.950 621.600 417.600 ;
        RECT 625.950 416.100 628.050 418.200 ;
        RECT 632.400 418.050 633.450 421.950 ;
        RECT 620.400 415.350 621.600 415.950 ;
        RECT 626.400 415.350 627.600 416.100 ;
        RECT 631.950 415.950 634.050 418.050 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 623.400 411.000 624.600 412.650 ;
        RECT 629.400 411.900 630.600 412.650 ;
        RECT 617.400 405.450 618.450 409.950 ;
        RECT 622.950 406.950 625.050 411.000 ;
        RECT 628.950 409.800 631.050 411.900 ;
        RECT 617.400 404.400 621.450 405.450 ;
        RECT 610.950 397.950 613.050 400.050 ;
        RECT 605.400 395.400 609.450 396.450 ;
        RECT 601.950 382.950 604.050 385.050 ;
        RECT 605.400 373.200 606.450 395.400 ;
        RECT 607.950 391.950 610.050 394.050 ;
        RECT 608.400 379.050 609.450 391.950 ;
        RECT 610.950 379.950 613.050 382.050 ;
        RECT 607.950 376.950 610.050 379.050 ;
        RECT 598.950 370.950 601.050 373.050 ;
        RECT 604.950 371.100 607.050 373.200 ;
        RECT 611.400 372.600 612.450 379.950 ;
        RECT 620.400 379.050 621.450 404.400 ;
        RECT 631.950 403.950 634.050 406.050 ;
        RECT 625.950 400.950 628.050 403.050 ;
        RECT 622.950 397.950 625.050 400.050 ;
        RECT 619.950 376.950 622.050 379.050 ;
        RECT 623.400 376.050 624.450 397.950 ;
        RECT 626.400 390.450 627.450 400.950 ;
        RECT 626.400 389.400 630.450 390.450 ;
        RECT 625.950 385.950 628.050 388.050 ;
        RECT 622.950 373.950 625.050 376.050 ;
        RECT 605.400 370.350 606.600 371.100 ;
        RECT 611.400 370.350 612.600 372.600 ;
        RECT 616.950 370.950 619.050 373.050 ;
        RECT 626.400 372.600 627.450 385.950 ;
        RECT 629.400 376.050 630.450 389.400 ;
        RECT 632.400 379.050 633.450 403.950 ;
        RECT 631.950 376.950 634.050 379.050 ;
        RECT 629.400 375.900 633.000 376.050 ;
        RECT 629.400 374.400 634.050 375.900 ;
        RECT 630.000 373.950 634.050 374.400 ;
        RECT 631.950 373.800 634.050 373.950 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 610.950 367.950 613.050 370.050 ;
        RECT 595.950 364.950 598.050 367.050 ;
        RECT 602.400 366.900 603.600 367.650 ;
        RECT 601.950 364.800 604.050 366.900 ;
        RECT 608.400 365.400 609.600 367.650 ;
        RECT 595.950 361.800 598.050 363.900 ;
        RECT 604.950 361.950 607.050 364.050 ;
        RECT 596.400 343.050 597.450 361.800 ;
        RECT 605.400 358.050 606.450 361.950 ;
        RECT 604.950 355.950 607.050 358.050 ;
        RECT 608.400 355.050 609.450 365.400 ;
        RECT 607.950 352.950 610.050 355.050 ;
        RECT 613.950 352.950 616.050 355.050 ;
        RECT 610.950 349.950 613.050 352.050 ;
        RECT 598.950 343.950 601.050 346.050 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 584.400 337.350 585.600 339.000 ;
        RECT 590.400 337.350 591.600 339.600 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 581.400 333.900 582.600 334.650 ;
        RECT 580.950 333.450 583.050 333.900 ;
        RECT 578.400 332.400 583.050 333.450 ;
        RECT 574.950 310.950 577.050 313.050 ;
        RECT 562.950 303.900 567.000 304.050 ;
        RECT 562.950 301.950 568.050 303.900 ;
        RECT 571.950 301.950 574.050 304.050 ;
        RECT 565.950 301.800 568.050 301.950 ;
        RECT 568.950 298.950 571.050 301.050 ;
        RECT 559.950 295.950 562.050 298.050 ;
        RECT 569.400 295.050 570.450 298.950 ;
        RECT 551.400 292.350 552.600 294.600 ;
        RECT 557.400 292.350 558.600 294.600 ;
        RECT 565.800 292.950 567.900 295.050 ;
        RECT 568.950 292.950 571.050 295.050 ;
        RECT 571.950 294.000 574.050 298.050 ;
        RECT 578.400 294.600 579.450 332.400 ;
        RECT 580.950 331.800 583.050 332.400 ;
        RECT 587.400 332.400 588.600 334.650 ;
        RECT 593.400 332.400 594.600 334.650 ;
        RECT 583.950 325.950 586.050 328.050 ;
        RECT 584.400 319.050 585.450 325.950 ;
        RECT 583.950 316.950 586.050 319.050 ;
        RECT 587.400 316.050 588.450 332.400 ;
        RECT 593.400 328.050 594.450 332.400 ;
        RECT 592.950 325.950 595.050 328.050 ;
        RECT 589.950 316.950 592.050 319.050 ;
        RECT 586.950 313.950 589.050 316.050 ;
        RECT 580.950 307.950 583.050 310.050 ;
        RECT 581.400 295.050 582.450 307.950 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 559.950 289.950 562.050 292.050 ;
        RECT 532.950 286.800 535.050 288.900 ;
        RECT 541.950 286.950 544.050 289.050 ;
        RECT 548.400 288.900 549.600 289.650 ;
        RECT 547.950 286.800 550.050 288.900 ;
        RECT 554.400 287.400 555.600 289.650 ;
        RECT 560.400 287.400 561.600 289.650 ;
        RECT 523.950 268.950 526.050 271.050 ;
        RECT 533.400 265.050 534.450 286.800 ;
        RECT 547.950 274.950 550.050 277.050 ;
        RECT 541.950 268.950 544.050 271.050 ;
        RECT 515.400 260.400 519.450 261.450 ;
        RECT 523.950 261.000 526.050 265.050 ;
        RECT 529.950 262.950 532.050 265.050 ;
        RECT 532.950 262.950 535.050 265.050 ;
        RECT 497.400 259.350 498.600 260.100 ;
        RECT 503.400 259.350 504.600 260.100 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 499.950 256.950 502.050 259.050 ;
        RECT 502.950 256.950 505.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 493.950 253.950 496.050 256.050 ;
        RECT 500.400 255.000 501.600 256.650 ;
        RECT 506.400 255.900 507.600 256.650 ;
        RECT 490.950 250.950 493.050 253.050 ;
        RECT 481.950 223.950 484.050 226.050 ;
        RECT 490.950 223.950 493.050 226.050 ;
        RECT 478.950 220.950 481.050 223.050 ;
        RECT 472.950 215.100 475.050 220.050 ;
        RECT 479.400 216.600 480.450 220.950 ;
        RECT 479.400 214.350 480.600 216.600 ;
        RECT 484.950 215.100 487.050 217.200 ;
        RECT 485.400 214.350 486.600 215.100 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 481.950 211.950 484.050 214.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 472.950 208.950 475.050 211.050 ;
        RECT 476.400 210.900 477.600 211.650 ;
        RECT 473.400 190.050 474.450 208.950 ;
        RECT 475.950 208.800 478.050 210.900 ;
        RECT 482.400 209.400 483.600 211.650 ;
        RECT 491.400 210.900 492.450 223.950 ;
        RECT 482.400 207.450 483.450 209.400 ;
        RECT 490.950 208.800 493.050 210.900 ;
        RECT 479.400 206.400 483.450 207.450 ;
        RECT 479.400 193.050 480.450 206.400 ;
        RECT 481.950 202.950 484.050 205.050 ;
        RECT 478.950 190.950 481.050 193.050 ;
        RECT 472.950 187.950 475.050 190.050 ;
        RECT 469.950 184.950 472.050 187.050 ;
        RECT 475.950 183.000 478.050 187.050 ;
        RECT 476.400 181.350 477.600 183.000 ;
        RECT 470.100 178.950 472.200 181.050 ;
        RECT 475.500 178.950 477.600 181.050 ;
        RECT 478.800 178.950 480.900 181.050 ;
        RECT 436.950 170.400 441.450 171.450 ;
        RECT 436.950 169.950 439.050 170.400 ;
        RECT 421.950 148.950 424.050 151.050 ;
        RECT 418.950 139.950 421.050 142.050 ;
        RECT 421.950 137.100 424.050 139.200 ;
        RECT 427.950 138.000 430.050 142.050 ;
        RECT 422.400 136.350 423.600 137.100 ;
        RECT 428.400 136.350 429.600 138.000 ;
        RECT 433.950 137.100 436.050 139.200 ;
        RECT 437.400 138.450 438.450 169.950 ;
        RECT 439.950 141.450 444.000 142.050 ;
        RECT 439.950 139.950 444.450 141.450 ;
        RECT 443.400 138.600 444.450 139.950 ;
        RECT 437.400 137.400 441.450 138.450 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 424.950 133.950 427.050 136.050 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 419.400 131.400 420.600 133.650 ;
        RECT 425.400 132.900 426.600 133.650 ;
        RECT 412.950 127.950 415.050 130.050 ;
        RECT 398.100 100.950 400.200 103.050 ;
        RECT 401.400 100.950 403.500 103.050 ;
        RECT 406.800 100.950 408.900 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 398.400 98.400 399.600 100.650 ;
        RECT 407.400 99.450 408.600 100.650 ;
        RECT 410.400 99.450 411.450 100.950 ;
        RECT 407.400 98.400 411.450 99.450 ;
        RECT 398.400 73.050 399.450 98.400 ;
        RECT 413.400 97.050 414.450 127.950 ;
        RECT 419.400 118.050 420.450 131.400 ;
        RECT 424.950 130.800 427.050 132.900 ;
        RECT 434.400 127.050 435.450 137.100 ;
        RECT 436.950 133.950 439.050 136.050 ;
        RECT 433.950 124.950 436.050 127.050 ;
        RECT 437.400 124.050 438.450 133.950 ;
        RECT 436.950 121.950 439.050 124.050 ;
        RECT 418.950 115.950 421.050 118.050 ;
        RECT 436.950 115.950 439.050 118.050 ;
        RECT 427.950 109.950 430.050 112.050 ;
        RECT 421.950 104.100 424.050 106.200 ;
        RECT 428.400 105.600 429.450 109.950 ;
        RECT 422.400 103.350 423.600 104.100 ;
        RECT 428.400 103.350 429.600 105.600 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 421.950 100.950 424.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 419.400 98.400 420.600 100.650 ;
        RECT 425.400 98.400 426.600 100.650 ;
        RECT 431.400 99.900 432.600 100.650 ;
        RECT 412.950 94.950 415.050 97.050 ;
        RECT 419.400 94.050 420.450 98.400 ;
        RECT 418.950 91.950 421.050 94.050 ;
        RECT 415.950 82.950 418.050 85.050 ;
        RECT 400.950 76.950 403.050 79.050 ;
        RECT 397.950 70.950 400.050 73.050 ;
        RECT 394.950 64.950 397.050 67.050 ;
        RECT 391.950 59.100 394.050 61.200 ;
        RECT 401.400 60.600 402.450 76.950 ;
        RECT 412.950 64.950 415.050 67.050 ;
        RECT 392.400 49.050 393.450 59.100 ;
        RECT 401.400 58.350 402.600 60.600 ;
        RECT 406.950 59.100 409.050 61.200 ;
        RECT 407.400 58.350 408.600 59.100 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 400.950 55.950 403.050 58.050 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 398.400 53.400 399.600 55.650 ;
        RECT 404.400 54.900 405.600 55.650 ;
        RECT 391.800 46.950 393.900 49.050 ;
        RECT 385.950 43.950 388.050 46.050 ;
        RECT 388.950 43.950 391.050 46.050 ;
        RECT 394.950 43.950 397.050 49.050 ;
        RECT 386.400 34.050 387.450 43.950 ;
        RECT 398.400 40.050 399.450 53.400 ;
        RECT 403.950 52.800 406.050 54.900 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 404.400 51.450 405.450 52.800 ;
        RECT 406.950 51.450 409.050 52.050 ;
        RECT 404.400 50.400 409.050 51.450 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 400.950 46.950 403.050 49.050 ;
        RECT 397.950 37.950 400.050 40.050 ;
        RECT 401.400 37.050 402.450 46.950 ;
        RECT 400.950 34.950 403.050 37.050 ;
        RECT 385.950 31.950 388.050 34.050 ;
        RECT 400.950 31.800 403.050 33.900 ;
        RECT 370.950 29.400 375.450 31.050 ;
        RECT 370.950 28.950 375.000 29.400 ;
        RECT 368.400 26.400 372.450 27.450 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 325.950 19.800 328.050 21.900 ;
        RECT 334.950 19.800 337.050 21.900 ;
        RECT 341.400 20.400 346.050 22.050 ;
        RECT 342.000 19.950 346.050 20.400 ;
        RECT 349.950 19.800 352.050 22.050 ;
        RECT 356.400 21.900 357.600 22.650 ;
        RECT 362.400 21.900 363.600 22.650 ;
        RECT 371.400 21.900 372.450 26.400 ;
        RECT 373.950 25.950 376.050 28.050 ;
        RECT 382.950 26.100 385.050 28.200 ;
        RECT 388.950 27.000 391.050 31.050 ;
        RECT 401.400 27.600 402.450 31.800 ;
        RECT 407.400 27.600 408.450 49.950 ;
        RECT 410.400 34.050 411.450 52.950 ;
        RECT 409.950 31.950 412.050 34.050 ;
        RECT 413.400 31.050 414.450 64.950 ;
        RECT 416.400 61.050 417.450 82.950 ;
        RECT 425.400 67.050 426.450 98.400 ;
        RECT 430.950 97.800 433.050 99.900 ;
        RECT 427.950 67.950 430.050 70.050 ;
        RECT 424.950 64.950 427.050 67.050 ;
        RECT 428.400 63.450 429.450 67.950 ;
        RECT 433.950 64.950 436.050 67.050 ;
        RECT 425.400 62.400 429.450 63.450 ;
        RECT 415.950 58.950 418.050 61.050 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 425.400 60.600 426.450 62.400 ;
        RECT 419.400 58.350 420.600 59.100 ;
        RECT 425.400 58.350 426.600 60.600 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 422.400 53.400 423.600 55.650 ;
        RECT 428.400 53.400 429.600 55.650 ;
        RECT 416.400 49.050 417.450 52.950 ;
        RECT 422.400 49.050 423.450 53.400 ;
        RECT 415.950 46.950 418.050 49.050 ;
        RECT 421.950 46.950 424.050 49.050 ;
        RECT 428.400 31.050 429.450 53.400 ;
        RECT 430.950 52.950 433.050 55.050 ;
        RECT 412.950 30.450 415.050 31.050 ;
        RECT 412.950 29.400 417.450 30.450 ;
        RECT 412.950 28.950 415.050 29.400 ;
        RECT 355.950 19.800 358.050 21.900 ;
        RECT 361.950 19.800 364.050 21.900 ;
        RECT 370.950 19.800 373.050 21.900 ;
        RECT 374.400 16.050 375.450 25.950 ;
        RECT 383.400 25.350 384.600 26.100 ;
        RECT 389.400 25.350 390.600 27.000 ;
        RECT 401.400 25.350 402.600 27.600 ;
        RECT 407.400 25.350 408.600 27.600 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 382.950 22.950 385.050 25.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 380.400 21.900 381.600 22.650 ;
        RECT 379.950 19.800 382.050 21.900 ;
        RECT 386.400 21.000 387.600 22.650 ;
        RECT 385.950 16.950 388.050 21.000 ;
        RECT 391.950 19.950 394.050 22.050 ;
        RECT 404.400 20.400 405.600 22.650 ;
        RECT 410.400 21.450 411.600 22.650 ;
        RECT 416.400 21.450 417.450 29.400 ;
        RECT 427.950 28.950 430.050 31.050 ;
        RECT 428.400 27.450 429.600 27.600 ;
        RECT 431.400 27.450 432.450 52.950 ;
        RECT 434.400 52.050 435.450 64.950 ;
        RECT 437.400 61.200 438.450 115.950 ;
        RECT 440.400 115.050 441.450 137.400 ;
        RECT 443.400 136.350 444.600 138.600 ;
        RECT 452.400 138.450 453.600 138.600 ;
        RECT 452.400 137.400 456.450 138.450 ;
        RECT 452.400 136.350 453.600 137.400 ;
        RECT 443.100 133.950 445.200 136.050 ;
        RECT 448.500 133.950 450.600 136.050 ;
        RECT 451.800 133.950 453.900 136.050 ;
        RECT 449.400 132.000 450.600 133.650 ;
        RECT 448.950 127.950 451.050 132.000 ;
        RECT 455.400 127.050 456.450 137.400 ;
        RECT 461.400 136.050 462.450 175.950 ;
        RECT 463.950 175.800 466.050 177.900 ;
        RECT 466.950 175.950 469.050 178.050 ;
        RECT 470.400 176.400 471.600 178.650 ;
        RECT 479.400 177.450 480.600 178.650 ;
        RECT 482.400 177.450 483.450 202.950 ;
        RECT 487.950 199.950 490.050 202.050 ;
        RECT 488.400 196.050 489.450 199.950 ;
        RECT 487.950 193.950 490.050 196.050 ;
        RECT 491.400 187.050 492.450 208.800 ;
        RECT 494.400 199.050 495.450 253.950 ;
        RECT 499.950 250.950 502.050 255.000 ;
        RECT 505.950 253.800 508.050 255.900 ;
        RECT 512.400 250.050 513.450 260.100 ;
        RECT 511.950 247.950 514.050 250.050 ;
        RECT 496.950 241.950 499.050 244.050 ;
        RECT 497.400 217.050 498.450 241.950 ;
        RECT 502.950 220.950 505.050 223.050 ;
        RECT 496.950 214.950 499.050 217.050 ;
        RECT 503.400 216.600 504.450 220.950 ;
        RECT 515.400 217.050 516.450 260.400 ;
        RECT 524.400 259.350 525.600 261.000 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 523.950 256.950 526.050 259.050 ;
        RECT 521.400 255.900 522.600 256.650 ;
        RECT 520.950 253.800 523.050 255.900 ;
        RECT 520.950 232.950 523.050 235.050 ;
        RECT 503.400 214.350 504.600 216.600 ;
        RECT 514.950 214.950 517.050 217.050 ;
        RECT 521.400 216.600 522.450 232.950 ;
        RECT 521.400 214.350 522.600 216.600 ;
        RECT 499.950 211.950 502.050 214.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 505.950 211.950 508.050 214.050 ;
        RECT 517.950 211.950 520.050 214.050 ;
        RECT 520.950 211.950 523.050 214.050 ;
        RECT 523.950 211.950 526.050 214.050 ;
        RECT 500.400 210.900 501.600 211.650 ;
        RECT 499.950 208.800 502.050 210.900 ;
        RECT 506.400 209.400 507.600 211.650 ;
        RECT 506.400 205.050 507.450 209.400 ;
        RECT 508.950 208.950 511.050 211.050 ;
        RECT 518.400 210.900 519.600 211.650 ;
        RECT 505.950 202.950 508.050 205.050 ;
        RECT 496.950 199.950 499.050 202.050 ;
        RECT 493.950 196.950 496.050 199.050 ;
        RECT 497.400 196.050 498.450 199.950 ;
        RECT 505.950 199.800 508.050 201.900 ;
        RECT 496.950 193.950 499.050 196.050 ;
        RECT 496.950 187.950 499.050 190.050 ;
        RECT 490.950 186.450 493.050 187.050 ;
        RECT 488.400 185.400 493.050 186.450 ;
        RECT 484.950 181.950 487.050 184.050 ;
        RECT 479.400 176.400 483.450 177.450 ;
        RECT 470.400 175.050 471.450 176.400 ;
        RECT 468.000 174.900 471.450 175.050 ;
        RECT 466.950 173.400 471.450 174.900 ;
        RECT 466.950 172.950 471.000 173.400 ;
        RECT 466.950 172.800 469.050 172.950 ;
        RECT 482.400 172.050 483.450 176.400 ;
        RECT 481.950 169.950 484.050 172.050 ;
        RECT 475.950 163.950 478.050 166.050 ;
        RECT 469.950 137.100 472.050 139.200 ;
        RECT 476.400 138.600 477.450 163.950 ;
        RECT 485.400 163.050 486.450 181.950 ;
        RECT 488.400 177.900 489.450 185.400 ;
        RECT 490.950 184.950 493.050 185.400 ;
        RECT 497.400 183.600 498.450 187.950 ;
        RECT 497.400 181.350 498.600 183.600 ;
        RECT 493.950 178.950 496.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 494.400 177.900 495.600 178.650 ;
        RECT 487.950 175.800 490.050 177.900 ;
        RECT 493.950 175.800 496.050 177.900 ;
        RECT 500.400 176.400 501.600 178.650 ;
        RECT 500.400 172.050 501.450 176.400 ;
        RECT 499.950 169.950 502.050 172.050 ;
        RECT 484.950 160.950 487.050 163.050 ;
        RECT 506.400 157.050 507.450 199.800 ;
        RECT 505.950 154.950 508.050 157.050 ;
        RECT 509.400 151.050 510.450 208.950 ;
        RECT 517.950 208.800 520.050 210.900 ;
        RECT 524.400 209.400 525.600 211.650 ;
        RECT 518.400 202.050 519.450 208.800 ;
        RECT 524.400 205.050 525.450 209.400 ;
        RECT 526.950 205.950 529.050 208.050 ;
        RECT 523.950 202.950 526.050 205.050 ;
        RECT 517.950 199.950 520.050 202.050 ;
        RECT 514.950 190.950 517.050 193.050 ;
        RECT 515.400 183.600 516.450 190.950 ;
        RECT 515.400 181.350 516.600 183.600 ;
        RECT 512.100 178.950 514.200 181.050 ;
        RECT 515.400 178.950 517.500 181.050 ;
        RECT 520.800 178.950 522.900 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 512.400 176.400 513.600 178.650 ;
        RECT 521.400 177.900 522.600 178.650 ;
        RECT 512.400 163.050 513.450 176.400 ;
        RECT 520.950 175.800 523.050 177.900 ;
        RECT 511.950 160.950 514.050 163.050 ;
        RECT 481.950 148.950 484.050 151.050 ;
        RECT 508.950 148.950 511.050 151.050 ;
        RECT 470.400 136.350 471.600 137.100 ;
        RECT 476.400 136.350 477.600 138.600 ;
        RECT 460.950 133.950 463.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 467.400 132.900 468.600 133.650 ;
        RECT 466.950 130.800 469.050 132.900 ;
        RECT 473.400 132.000 474.600 133.650 ;
        RECT 472.950 127.950 475.050 132.000 ;
        RECT 454.950 126.450 457.050 127.050 ;
        RECT 452.400 125.400 457.050 126.450 ;
        RECT 452.400 121.050 453.450 125.400 ;
        RECT 454.950 124.950 457.050 125.400 ;
        RECT 451.950 118.950 454.050 121.050 ;
        RECT 457.950 118.950 460.050 121.050 ;
        RECT 439.950 112.950 442.050 115.050 ;
        RECT 442.950 104.100 445.050 106.200 ;
        RECT 448.950 105.000 451.050 109.050 ;
        RECT 443.400 103.350 444.600 104.100 ;
        RECT 449.400 103.350 450.600 105.000 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 448.950 100.950 451.050 103.050 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 446.400 99.000 447.600 100.650 ;
        RECT 452.400 99.900 453.600 100.650 ;
        RECT 458.400 99.900 459.450 118.950 ;
        RECT 482.400 109.050 483.450 148.950 ;
        RECT 484.950 138.450 487.050 142.050 ;
        RECT 490.500 141.300 492.600 143.400 ;
        RECT 500.100 142.500 502.200 144.600 ;
        RECT 488.400 138.450 489.600 138.600 ;
        RECT 484.950 138.000 489.600 138.450 ;
        RECT 485.400 137.400 489.600 138.000 ;
        RECT 488.400 136.350 489.600 137.400 ;
        RECT 488.100 133.950 490.200 136.050 ;
        RECT 491.400 132.300 492.300 141.300 ;
        RECT 493.800 137.700 495.900 139.800 ;
        RECT 497.400 139.350 498.600 141.600 ;
        RECT 495.000 135.300 495.900 137.700 ;
        RECT 496.800 136.950 498.900 139.050 ;
        RECT 500.700 135.300 501.900 142.500 ;
        RECT 508.950 137.100 511.050 139.200 ;
        RECT 517.950 137.100 520.050 142.050 ;
        RECT 524.400 138.600 525.450 178.950 ;
        RECT 495.000 134.100 501.900 135.300 ;
        RECT 498.000 132.300 500.100 133.200 ;
        RECT 491.400 131.100 500.100 132.300 ;
        RECT 492.900 129.300 495.000 131.100 ;
        RECT 496.800 128.100 498.900 130.200 ;
        RECT 501.000 128.700 501.900 134.100 ;
        RECT 502.800 133.950 504.900 136.050 ;
        RECT 503.400 132.900 504.600 133.650 ;
        RECT 502.950 130.800 505.050 132.900 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 497.400 125.550 498.600 127.800 ;
        RECT 500.100 126.600 502.200 128.700 ;
        RECT 484.950 118.950 487.050 121.050 ;
        RECT 460.950 103.950 463.050 106.050 ;
        RECT 466.950 104.100 469.050 106.200 ;
        RECT 472.950 105.000 475.050 109.050 ;
        RECT 481.950 106.950 484.050 109.050 ;
        RECT 445.950 94.950 448.050 99.000 ;
        RECT 451.950 97.800 454.050 99.900 ;
        RECT 457.950 97.800 460.050 99.900 ;
        RECT 461.400 85.050 462.450 103.950 ;
        RECT 467.400 103.350 468.600 104.100 ;
        RECT 473.400 103.350 474.600 105.000 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 470.400 99.000 471.600 100.650 ;
        RECT 476.400 99.900 477.600 100.650 ;
        RECT 469.950 94.950 472.050 99.000 ;
        RECT 475.950 97.800 478.050 99.900 ;
        RECT 482.400 91.050 483.450 106.950 ;
        RECT 485.400 106.050 486.450 118.950 ;
        RECT 487.950 112.950 490.050 115.050 ;
        RECT 488.400 109.050 489.450 112.950 ;
        RECT 487.950 106.950 490.050 109.050 ;
        RECT 484.950 103.950 487.050 106.050 ;
        RECT 491.400 105.600 492.450 124.950 ;
        RECT 491.400 103.350 492.600 105.600 ;
        RECT 497.400 105.450 498.450 125.550 ;
        RECT 509.400 106.200 510.450 137.100 ;
        RECT 518.400 136.350 519.600 137.100 ;
        RECT 524.400 136.350 525.600 138.600 ;
        RECT 527.400 138.450 528.450 205.950 ;
        RECT 530.400 175.050 531.450 262.950 ;
        RECT 542.400 261.600 543.450 268.950 ;
        RECT 542.400 259.350 543.600 261.600 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 539.400 254.400 540.600 256.650 ;
        RECT 539.400 250.050 540.450 254.400 ;
        RECT 538.950 247.950 541.050 250.050 ;
        RECT 548.400 229.050 549.450 274.950 ;
        RECT 554.400 265.050 555.450 287.400 ;
        RECT 560.400 280.050 561.450 287.400 ;
        RECT 562.950 280.950 565.050 283.050 ;
        RECT 559.950 277.950 562.050 280.050 ;
        RECT 558.000 267.450 562.050 268.050 ;
        RECT 557.400 265.950 562.050 267.450 ;
        RECT 553.950 262.950 556.050 265.050 ;
        RECT 557.400 262.200 558.450 265.950 ;
        RECT 563.400 262.200 564.450 280.950 ;
        RECT 566.400 277.050 567.450 292.950 ;
        RECT 572.400 292.350 573.600 294.000 ;
        RECT 578.400 292.350 579.600 294.600 ;
        RECT 580.950 292.950 583.050 295.050 ;
        RECT 583.950 292.950 586.050 295.050 ;
        RECT 590.400 294.450 591.450 316.950 ;
        RECT 587.400 293.400 591.450 294.450 ;
        RECT 593.400 294.600 594.450 325.950 ;
        RECT 595.950 322.950 598.050 325.050 ;
        RECT 596.400 298.050 597.450 322.950 ;
        RECT 599.400 298.200 600.450 343.950 ;
        RECT 601.950 340.950 604.050 343.050 ;
        RECT 602.400 307.050 603.450 340.950 ;
        RECT 611.400 339.600 612.450 349.950 ;
        RECT 614.400 343.050 615.450 352.950 ;
        RECT 617.400 346.050 618.450 370.950 ;
        RECT 626.400 370.350 627.600 372.600 ;
        RECT 631.950 370.950 634.050 373.050 ;
        RECT 635.400 372.450 636.450 425.400 ;
        RECT 637.950 421.950 640.050 424.050 ;
        RECT 638.400 418.050 639.450 421.950 ;
        RECT 641.400 421.050 642.450 428.400 ;
        RECT 659.400 427.050 660.450 433.950 ;
        RECT 649.950 421.950 652.050 427.050 ;
        RECT 652.950 424.950 655.050 427.050 ;
        RECT 658.950 424.950 661.050 427.050 ;
        RECT 640.950 418.950 643.050 421.050 ;
        RECT 637.950 415.950 640.050 418.050 ;
        RECT 643.950 416.100 646.050 418.200 ;
        RECT 644.400 415.350 645.600 416.100 ;
        RECT 649.950 415.950 652.050 420.900 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 641.400 411.900 642.600 412.650 ;
        RECT 647.400 411.900 648.600 412.650 ;
        RECT 653.400 411.900 654.450 424.950 ;
        RECT 655.950 415.950 661.050 418.050 ;
        RECT 665.400 417.600 666.450 439.950 ;
        RECT 668.400 436.050 669.450 442.950 ;
        RECT 671.400 442.050 672.450 451.800 ;
        RECT 673.950 448.950 676.050 451.050 ;
        RECT 670.950 439.950 673.050 442.050 ;
        RECT 674.400 439.050 675.450 448.950 ;
        RECT 673.950 436.950 676.050 439.050 ;
        RECT 667.950 433.950 670.050 436.050 ;
        RECT 674.400 427.050 675.450 436.950 ;
        RECT 673.950 424.950 676.050 427.050 ;
        RECT 665.400 415.350 666.600 417.600 ;
        RECT 670.950 417.000 673.050 421.050 ;
        RECT 677.400 418.050 678.450 454.950 ;
        RECT 680.400 450.600 681.450 454.950 ;
        RECT 683.400 454.050 684.450 481.950 ;
        RECT 689.400 472.050 690.450 488.400 ;
        RECT 694.950 487.800 697.050 489.900 ;
        RECT 701.400 484.050 702.450 494.400 ;
        RECT 703.950 494.100 706.050 496.200 ;
        RECT 709.950 494.100 712.050 496.200 ;
        RECT 710.400 493.350 711.600 494.100 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 707.400 488.400 708.600 490.650 ;
        RECT 703.950 484.950 706.050 487.050 ;
        RECT 700.950 481.950 703.050 484.050 ;
        RECT 688.950 469.950 691.050 472.050 ;
        RECT 694.950 469.950 697.050 472.050 ;
        RECT 691.950 457.950 694.050 460.050 ;
        RECT 682.950 451.950 685.050 454.050 ;
        RECT 680.400 448.350 681.600 450.600 ;
        RECT 688.950 449.100 691.050 451.200 ;
        RECT 689.400 448.350 690.600 449.100 ;
        RECT 692.400 448.050 693.450 457.950 ;
        RECT 695.400 457.050 696.450 469.950 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 697.950 454.950 700.050 457.050 ;
        RECT 694.950 451.800 697.050 453.900 ;
        RECT 680.100 445.950 682.200 448.050 ;
        RECT 685.500 445.950 687.600 448.050 ;
        RECT 688.800 445.950 690.900 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 686.400 443.400 687.600 445.650 ;
        RECT 682.950 439.950 685.050 442.050 ;
        RECT 683.400 430.050 684.450 439.950 ;
        RECT 682.950 427.950 685.050 430.050 ;
        RECT 686.400 427.050 687.450 443.400 ;
        RECT 691.950 439.950 694.050 444.900 ;
        RECT 695.400 436.050 696.450 451.800 ;
        RECT 698.400 451.050 699.450 454.950 ;
        RECT 704.400 451.200 705.450 484.950 ;
        RECT 707.400 457.050 708.450 488.400 ;
        RECT 712.950 487.950 715.050 490.050 ;
        RECT 713.400 478.050 714.450 487.950 ;
        RECT 712.950 475.950 715.050 478.050 ;
        RECT 716.400 472.050 717.450 497.400 ;
        RECT 722.400 495.600 723.450 502.950 ;
        RECT 725.400 499.050 726.450 547.950 ;
        RECT 728.400 538.050 729.450 553.950 ;
        RECT 727.950 535.950 730.050 538.050 ;
        RECT 733.950 528.000 736.050 532.050 ;
        RECT 743.400 529.200 744.450 596.400 ;
        RECT 745.950 595.950 748.050 596.400 ;
        RECT 745.950 589.950 748.050 592.050 ;
        RECT 746.400 574.050 747.450 589.950 ;
        RECT 749.400 577.050 750.450 604.950 ;
        RECT 758.400 604.350 759.600 606.600 ;
        RECT 763.950 604.950 766.050 610.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 757.950 601.950 760.050 604.050 ;
        RECT 760.950 601.950 763.050 604.050 ;
        RECT 755.400 600.900 756.600 601.650 ;
        RECT 754.950 598.800 757.050 600.900 ;
        RECT 761.400 599.400 762.600 601.650 ;
        RECT 761.400 586.050 762.450 599.400 ;
        RECT 763.950 598.950 766.050 601.050 ;
        RECT 764.400 595.050 765.450 598.950 ;
        RECT 763.950 592.950 766.050 595.050 ;
        RECT 760.950 583.950 763.050 586.050 ;
        RECT 748.800 574.950 750.900 577.050 ;
        RECT 745.950 571.950 748.050 574.050 ;
        RECT 751.950 573.000 754.050 577.050 ;
        RECT 754.950 576.450 759.000 577.050 ;
        RECT 754.950 574.950 759.450 576.450 ;
        RECT 758.400 573.600 759.450 574.950 ;
        RECT 752.400 571.350 753.600 573.000 ;
        RECT 758.400 571.350 759.600 573.600 ;
        RECT 748.950 568.950 751.050 571.050 ;
        RECT 751.950 568.950 754.050 571.050 ;
        RECT 754.950 568.950 757.050 571.050 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 749.400 568.050 750.600 568.650 ;
        RECT 745.950 566.400 750.600 568.050 ;
        RECT 755.400 567.900 756.600 568.650 ;
        RECT 745.950 565.950 750.450 566.400 ;
        RECT 749.400 553.050 750.450 565.950 ;
        RECT 754.950 565.800 757.050 567.900 ;
        RECT 764.400 565.050 765.450 592.950 ;
        RECT 754.950 562.650 757.050 564.750 ;
        RECT 763.950 562.950 766.050 565.050 ;
        RECT 748.950 550.950 751.050 553.050 ;
        RECT 751.950 538.950 754.050 541.050 ;
        RECT 734.400 526.350 735.600 528.000 ;
        RECT 739.800 527.100 741.900 529.200 ;
        RECT 742.950 528.450 745.050 529.200 ;
        RECT 742.950 527.400 747.450 528.450 ;
        RECT 742.950 527.100 745.050 527.400 ;
        RECT 740.400 526.350 741.600 527.100 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 733.950 523.950 736.050 526.050 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 731.400 521.400 732.600 523.650 ;
        RECT 737.400 522.000 738.600 523.650 ;
        RECT 731.400 508.050 732.450 521.400 ;
        RECT 733.950 517.950 736.050 520.050 ;
        RECT 736.950 517.950 739.050 522.000 ;
        RECT 746.400 520.050 747.450 527.400 ;
        RECT 745.950 517.950 748.050 520.050 ;
        RECT 730.950 505.950 733.050 508.050 ;
        RECT 727.950 502.950 730.050 505.050 ;
        RECT 724.950 496.950 727.050 499.050 ;
        RECT 728.400 495.600 729.450 502.950 ;
        RECT 734.400 496.050 735.450 517.950 ;
        RECT 745.950 508.950 748.050 511.050 ;
        RECT 739.950 505.950 742.050 508.050 ;
        RECT 736.950 496.950 739.050 499.050 ;
        RECT 722.400 493.350 723.600 495.600 ;
        RECT 728.400 493.350 729.600 495.600 ;
        RECT 733.950 493.950 736.050 496.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 724.950 490.950 727.050 493.050 ;
        RECT 727.950 490.950 730.050 493.050 ;
        RECT 730.950 490.950 733.050 493.050 ;
        RECT 725.400 488.400 726.600 490.650 ;
        RECT 731.400 489.900 732.600 490.650 ;
        RECT 725.400 484.050 726.450 488.400 ;
        RECT 730.950 487.800 733.050 489.900 ;
        RECT 733.950 487.950 736.050 490.050 ;
        RECT 737.400 489.900 738.450 496.950 ;
        RECT 740.400 496.050 741.450 505.950 ;
        RECT 746.400 496.200 747.450 508.950 ;
        RECT 752.400 499.050 753.450 538.950 ;
        RECT 755.400 526.050 756.450 562.650 ;
        RECT 767.400 541.050 768.450 643.950 ;
        RECT 773.400 628.050 774.450 644.400 ;
        RECT 782.400 634.050 783.450 677.400 ;
        RECT 787.950 676.950 790.050 679.050 ;
        RECT 791.400 673.050 792.450 721.950 ;
        RECT 794.400 718.050 795.450 722.400 ;
        RECT 799.950 721.800 802.050 723.900 ;
        RECT 805.950 721.950 808.050 724.050 ;
        RECT 793.950 715.950 796.050 718.050 ;
        RECT 796.950 703.950 799.050 706.050 ;
        RECT 797.400 694.050 798.450 703.950 ;
        RECT 800.400 697.050 801.450 721.800 ;
        RECT 802.950 712.950 805.050 715.050 ;
        RECT 799.950 694.950 802.050 697.050 ;
        RECT 796.950 691.950 799.050 694.050 ;
        RECT 797.400 684.600 798.450 691.950 ;
        RECT 803.400 684.600 804.450 712.950 ;
        RECT 806.400 706.050 807.450 721.950 ;
        RECT 805.950 703.950 808.050 706.050 ;
        RECT 797.400 682.350 798.600 684.600 ;
        RECT 803.400 682.350 804.600 684.600 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 800.400 677.400 801.600 679.650 ;
        RECT 790.950 670.950 793.050 673.050 ;
        RECT 800.400 667.050 801.450 677.400 ;
        RECT 809.400 676.050 810.450 730.950 ;
        RECT 814.950 728.100 817.050 730.200 ;
        RECT 821.400 729.600 822.450 733.950 ;
        RECT 827.400 730.050 828.450 733.950 ;
        RECT 815.400 727.350 816.600 728.100 ;
        RECT 821.400 727.350 822.600 729.600 ;
        RECT 826.950 727.950 829.050 730.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 818.400 723.000 819.600 724.650 ;
        RECT 824.400 723.900 825.600 724.650 ;
        RECT 830.400 723.900 831.450 742.950 ;
        RECT 836.400 735.450 837.450 770.400 ;
        RECT 842.400 769.050 843.450 793.950 ;
        RECT 851.400 793.050 852.450 799.950 ;
        RECT 856.950 796.950 859.050 799.050 ;
        RECT 850.950 790.950 853.050 793.050 ;
        RECT 841.950 766.950 844.050 769.050 ;
        RECT 847.950 766.950 850.050 769.050 ;
        RECT 841.950 763.950 847.050 766.050 ;
        RECT 841.950 760.950 844.050 763.050 ;
        RECT 848.400 762.600 849.450 766.950 ;
        RECT 842.400 760.350 843.600 760.950 ;
        RECT 848.400 760.350 849.600 762.600 ;
        RECT 841.950 757.950 844.050 760.050 ;
        RECT 844.950 757.950 847.050 760.050 ;
        RECT 847.950 757.950 850.050 760.050 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 845.400 756.900 846.600 757.650 ;
        RECT 844.950 754.800 847.050 756.900 ;
        RECT 851.400 755.400 852.600 757.650 ;
        RECT 857.400 756.450 858.450 796.950 ;
        RECT 860.400 781.050 861.450 800.400 ;
        RECT 865.950 799.800 868.050 801.900 ;
        RECT 872.400 800.400 873.600 802.650 ;
        RECT 866.400 790.050 867.450 799.800 ;
        RECT 865.950 787.950 868.050 790.050 ;
        RECT 872.400 787.050 873.450 800.400 ;
        RECT 877.950 799.950 880.050 804.900 ;
        RECT 881.400 799.050 882.450 820.950 ;
        RECT 889.950 806.100 892.050 808.200 ;
        RECT 895.950 807.000 898.050 811.050 ;
        RECT 899.400 808.050 900.450 832.800 ;
        RECT 890.400 805.350 891.600 806.100 ;
        RECT 896.400 805.350 897.600 807.000 ;
        RECT 898.950 805.950 901.050 808.050 ;
        RECT 886.950 802.950 889.050 805.050 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 895.950 802.950 898.050 805.050 ;
        RECT 887.400 800.400 888.600 802.650 ;
        RECT 893.400 800.400 894.600 802.650 ;
        RECT 880.950 796.950 883.050 799.050 ;
        RECT 887.400 787.050 888.450 800.400 ;
        RECT 893.400 793.050 894.450 800.400 ;
        RECT 898.800 799.950 900.900 802.050 ;
        RECT 902.400 801.900 903.450 874.650 ;
        RECT 908.400 871.050 909.450 886.950 ;
        RECT 916.950 884.100 919.050 886.200 ;
        RECT 922.950 885.000 925.050 889.050 ;
        RECT 917.400 883.350 918.600 884.100 ;
        RECT 923.400 883.350 924.600 885.000 ;
        RECT 913.950 880.950 916.050 883.050 ;
        RECT 916.950 880.950 919.050 883.050 ;
        RECT 919.950 880.950 922.050 883.050 ;
        RECT 922.950 880.950 925.050 883.050 ;
        RECT 914.400 878.400 915.600 880.650 ;
        RECT 920.400 879.000 921.600 880.650 ;
        RECT 914.400 874.050 915.450 878.400 ;
        RECT 919.950 874.950 922.050 879.000 ;
        RECT 913.950 871.950 916.050 874.050 ;
        RECT 907.950 868.950 910.050 871.050 ;
        RECT 919.950 868.950 922.050 871.050 ;
        RECT 913.950 847.950 916.050 850.050 ;
        RECT 904.950 844.950 907.050 847.050 ;
        RECT 905.400 840.600 906.450 844.950 ;
        RECT 914.400 840.600 915.450 847.950 ;
        RECT 905.400 838.350 906.600 840.600 ;
        RECT 914.400 840.450 915.600 840.600 ;
        RECT 914.400 839.400 918.450 840.450 ;
        RECT 914.400 838.350 915.600 839.400 ;
        RECT 905.100 835.950 907.200 838.050 ;
        RECT 910.500 835.950 912.600 838.050 ;
        RECT 913.800 835.950 915.900 838.050 ;
        RECT 911.400 833.400 912.600 835.650 ;
        RECT 911.400 811.050 912.450 833.400 ;
        RECT 917.400 811.050 918.450 839.400 ;
        RECT 920.400 823.050 921.450 868.950 ;
        RECT 929.400 865.050 930.450 910.800 ;
        RECT 931.950 901.950 934.050 904.050 ;
        RECT 928.950 862.950 931.050 865.050 ;
        RECT 929.400 829.050 930.450 862.950 ;
        RECT 932.400 844.050 933.450 901.950 ;
        RECT 931.950 841.950 934.050 844.050 ;
        RECT 928.950 826.950 931.050 829.050 ;
        RECT 919.950 820.950 922.050 823.050 ;
        RECT 904.950 808.950 907.050 811.050 ;
        RECT 892.950 790.950 895.050 793.050 ;
        RECT 871.950 784.950 874.050 787.050 ;
        RECT 886.950 784.950 889.050 787.050 ;
        RECT 859.950 778.950 862.050 781.050 ;
        RECT 874.950 775.950 877.050 778.050 ;
        RECT 859.950 761.100 862.050 763.200 ;
        RECT 868.950 761.100 871.050 763.200 ;
        RECT 875.400 762.600 876.450 775.950 ;
        RECT 899.400 775.050 900.450 799.950 ;
        RECT 901.950 799.800 904.050 801.900 ;
        RECT 905.400 796.050 906.450 808.950 ;
        RECT 910.950 807.000 913.050 811.050 ;
        RECT 916.950 807.000 919.050 811.050 ;
        RECT 922.950 808.950 925.050 811.050 ;
        RECT 928.950 808.950 931.050 811.050 ;
        RECT 911.400 805.350 912.600 807.000 ;
        RECT 917.400 805.350 918.600 807.000 ;
        RECT 910.950 802.950 913.050 805.050 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 916.950 802.950 919.050 805.050 ;
        RECT 914.400 801.900 915.600 802.650 ;
        RECT 913.950 799.800 916.050 801.900 ;
        RECT 904.950 793.950 907.050 796.050 ;
        RECT 916.950 775.950 919.050 778.050 ;
        RECT 889.950 772.950 892.050 775.050 ;
        RECT 898.950 772.950 901.050 775.050 ;
        RECT 913.950 772.950 916.050 775.050 ;
        RECT 890.400 762.600 891.450 772.950 ;
        RECT 901.950 766.950 904.050 769.050 ;
        RECT 854.400 755.400 858.450 756.450 ;
        RECT 841.950 747.450 844.050 751.050 ;
        RECT 851.400 748.050 852.450 755.400 ;
        RECT 841.950 747.000 846.450 747.450 ;
        RECT 842.400 746.400 846.450 747.000 ;
        RECT 841.950 742.950 844.050 745.050 ;
        RECT 833.400 734.400 837.450 735.450 ;
        RECT 817.950 718.950 820.050 723.000 ;
        RECT 823.950 721.800 826.050 723.900 ;
        RECT 829.950 721.800 832.050 723.900 ;
        RECT 833.400 721.050 834.450 734.400 ;
        RECT 842.400 729.600 843.450 742.950 ;
        RECT 845.400 742.050 846.450 746.400 ;
        RECT 850.950 745.950 853.050 748.050 ;
        RECT 844.950 739.950 847.050 742.050 ;
        RECT 842.400 727.350 843.600 729.600 ;
        RECT 847.950 729.000 850.050 733.050 ;
        RECT 850.950 730.950 853.050 736.050 ;
        RECT 848.400 727.350 849.600 729.000 ;
        RECT 838.950 724.950 841.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 839.400 724.050 840.600 724.650 ;
        RECT 835.950 722.400 840.600 724.050 ;
        RECT 845.400 723.000 846.600 724.650 ;
        RECT 835.950 721.950 840.000 722.400 ;
        RECT 832.950 718.950 835.050 721.050 ;
        RECT 838.950 718.950 841.050 721.050 ;
        RECT 844.950 718.950 847.050 723.000 ;
        RECT 854.400 721.050 855.450 755.400 ;
        RECT 856.950 739.950 859.050 742.050 ;
        RECT 857.400 736.050 858.450 739.950 ;
        RECT 856.950 733.950 859.050 736.050 ;
        RECT 860.400 733.050 861.450 761.100 ;
        RECT 869.400 760.350 870.600 761.100 ;
        RECT 875.400 760.350 876.600 762.600 ;
        RECT 890.400 760.350 891.600 762.600 ;
        RECT 895.950 761.100 898.050 763.200 ;
        RECT 896.400 760.350 897.600 761.100 ;
        RECT 865.950 757.950 868.050 760.050 ;
        RECT 868.950 757.950 871.050 760.050 ;
        RECT 871.950 757.950 874.050 760.050 ;
        RECT 874.950 757.950 877.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 889.950 757.950 892.050 760.050 ;
        RECT 892.950 757.950 895.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 866.400 756.900 867.600 757.650 ;
        RECT 872.400 756.900 873.600 757.650 ;
        RECT 865.950 754.800 868.050 756.900 ;
        RECT 871.950 754.800 874.050 756.900 ;
        RECT 887.400 755.400 888.600 757.650 ;
        RECT 893.400 755.400 894.600 757.650 ;
        RECT 862.950 748.950 865.050 751.050 ;
        RECT 863.400 739.050 864.450 748.950 ;
        RECT 862.950 736.950 865.050 739.050 ;
        RECT 856.950 729.450 859.050 732.900 ;
        RECT 859.950 730.950 862.050 733.050 ;
        RECT 860.400 729.450 861.600 729.600 ;
        RECT 856.950 729.000 861.600 729.450 ;
        RECT 857.400 728.400 861.600 729.000 ;
        RECT 860.400 727.350 861.600 728.400 ;
        RECT 865.950 728.100 868.050 733.050 ;
        RECT 872.400 730.050 873.450 754.800 ;
        RECT 874.800 748.950 876.900 751.050 ;
        RECT 877.950 748.950 880.050 751.050 ;
        RECT 866.400 727.350 867.600 728.100 ;
        RECT 871.950 727.950 874.050 730.050 ;
        RECT 859.950 724.950 862.050 727.050 ;
        RECT 862.950 724.950 865.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 856.950 721.950 859.050 724.050 ;
        RECT 863.400 723.000 864.600 724.650 ;
        RECT 869.400 724.050 870.600 724.650 ;
        RECT 853.950 718.950 856.050 721.050 ;
        RECT 814.950 697.950 817.050 700.050 ;
        RECT 815.400 685.050 816.450 697.950 ;
        RECT 835.950 691.950 838.050 694.050 ;
        RECT 811.950 682.950 814.050 685.050 ;
        RECT 814.950 682.950 817.050 685.050 ;
        RECT 817.950 683.100 820.050 685.200 ;
        RECT 823.950 683.100 826.050 685.200 ;
        RECT 802.950 673.950 805.050 676.050 ;
        RECT 808.950 675.450 811.050 676.050 ;
        RECT 806.400 674.400 811.050 675.450 ;
        RECT 799.950 664.950 802.050 667.050 ;
        RECT 784.950 655.950 787.050 658.050 ;
        RECT 781.950 631.950 784.050 634.050 ;
        RECT 772.950 625.950 775.050 628.050 ;
        RECT 781.950 619.950 784.050 622.050 ;
        RECT 769.950 604.950 772.050 610.050 ;
        RECT 772.950 606.000 775.050 610.050 ;
        RECT 778.950 606.000 781.050 610.050 ;
        RECT 782.400 607.050 783.450 619.950 ;
        RECT 773.400 604.350 774.600 606.000 ;
        RECT 779.400 604.350 780.600 606.000 ;
        RECT 781.950 604.950 784.050 607.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 769.950 598.950 772.050 601.050 ;
        RECT 776.400 599.400 777.600 601.650 ;
        RECT 770.400 574.050 771.450 598.950 ;
        RECT 776.400 586.050 777.450 599.400 ;
        RECT 781.950 598.950 784.050 601.050 ;
        RECT 775.950 583.950 778.050 586.050 ;
        RECT 782.400 576.450 783.450 598.950 ;
        RECT 779.400 575.400 783.450 576.450 ;
        RECT 779.400 574.200 780.450 575.400 ;
        RECT 769.950 571.950 772.050 574.050 ;
        RECT 772.950 572.100 775.050 574.200 ;
        RECT 778.950 572.100 781.050 574.200 ;
        RECT 785.400 574.050 786.450 655.950 ;
        RECT 793.950 650.100 796.050 652.200 ;
        RECT 794.400 649.350 795.600 650.100 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 793.950 646.950 796.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 791.400 644.400 792.600 646.650 ;
        RECT 797.400 644.400 798.600 646.650 ;
        RECT 791.400 637.050 792.450 644.400 ;
        RECT 797.400 640.050 798.450 644.400 ;
        RECT 796.950 637.950 799.050 640.050 ;
        RECT 803.400 637.050 804.450 673.950 ;
        RECT 806.400 643.050 807.450 674.400 ;
        RECT 808.950 673.950 811.050 674.400 ;
        RECT 812.400 673.050 813.450 682.950 ;
        RECT 818.400 682.350 819.600 683.100 ;
        RECT 824.400 682.350 825.600 683.100 ;
        RECT 829.950 682.950 832.050 688.050 ;
        RECT 836.400 684.450 837.450 691.950 ;
        RECT 839.400 688.200 840.450 718.950 ;
        RECT 853.950 715.800 856.050 717.900 ;
        RECT 838.950 686.100 841.050 688.200 ;
        RECT 833.400 683.400 837.450 684.450 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 823.950 679.950 826.050 682.050 ;
        RECT 826.950 679.950 829.050 682.050 ;
        RECT 821.400 677.400 822.600 679.650 ;
        RECT 827.400 678.900 828.600 679.650 ;
        RECT 811.950 670.950 814.050 673.050 ;
        RECT 812.400 655.200 813.450 670.950 ;
        RECT 821.400 658.050 822.450 677.400 ;
        RECT 826.950 676.800 829.050 678.900 ;
        RECT 829.950 667.950 832.050 670.050 ;
        RECT 830.400 663.450 831.450 667.950 ;
        RECT 833.400 667.050 834.450 683.400 ;
        RECT 838.950 682.950 841.050 685.050 ;
        RECT 844.950 684.000 847.050 688.050 ;
        RECT 839.400 682.350 840.600 682.950 ;
        RECT 845.400 682.350 846.600 684.000 ;
        RECT 838.950 679.950 841.050 682.050 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 844.950 679.950 847.050 682.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 842.400 677.400 843.600 679.650 ;
        RECT 848.400 677.400 849.600 679.650 ;
        RECT 838.950 673.950 841.050 676.050 ;
        RECT 832.950 664.950 835.050 667.050 ;
        RECT 830.400 662.400 834.450 663.450 ;
        RECT 820.950 655.950 823.050 658.050 ;
        RECT 811.950 653.100 814.050 655.200 ;
        RECT 811.950 649.950 814.050 652.050 ;
        RECT 817.950 651.000 820.050 655.050 ;
        RECT 833.400 654.450 834.450 662.400 ;
        RECT 835.950 661.950 838.050 664.050 ;
        RECT 836.400 654.450 837.450 661.950 ;
        RECT 839.400 658.050 840.450 673.950 ;
        RECT 842.400 673.050 843.450 677.400 ;
        RECT 848.400 673.050 849.450 677.400 ;
        RECT 850.950 676.950 853.050 679.050 ;
        RECT 841.950 670.950 844.050 673.050 ;
        RECT 847.950 670.950 850.050 673.050 ;
        RECT 838.950 655.950 841.050 658.050 ;
        RECT 851.400 655.050 852.450 676.950 ;
        RECT 854.400 670.050 855.450 715.800 ;
        RECT 857.400 684.450 858.450 721.950 ;
        RECT 862.950 718.950 865.050 723.000 ;
        RECT 869.400 721.950 874.050 724.050 ;
        RECT 865.950 718.950 868.050 721.050 ;
        RECT 862.950 703.950 865.050 706.050 ;
        RECT 863.400 687.450 864.450 703.950 ;
        RECT 866.400 697.050 867.450 718.950 ;
        RECT 869.400 715.050 870.450 721.950 ;
        RECT 871.950 720.450 874.050 720.900 ;
        RECT 875.400 720.450 876.450 748.950 ;
        RECT 878.400 739.050 879.450 748.950 ;
        RECT 883.950 742.950 886.050 745.050 ;
        RECT 880.950 739.950 883.050 742.050 ;
        RECT 877.950 736.950 880.050 739.050 ;
        RECT 881.400 735.450 882.450 739.950 ;
        RECT 878.400 734.400 882.450 735.450 ;
        RECT 878.400 730.050 879.450 734.400 ;
        RECT 877.950 727.950 880.050 730.050 ;
        RECT 884.400 729.600 885.450 742.950 ;
        RECT 887.400 733.050 888.450 755.400 ;
        RECT 889.950 748.950 892.050 751.050 ;
        RECT 890.400 733.050 891.450 748.950 ;
        RECT 893.400 745.050 894.450 755.400 ;
        RECT 892.950 742.950 895.050 745.050 ;
        RECT 898.950 736.950 901.050 739.050 ;
        RECT 886.800 730.950 888.900 733.050 ;
        RECT 889.950 730.950 892.050 733.050 ;
        RECT 895.950 730.950 898.050 733.050 ;
        RECT 890.400 729.600 891.450 730.950 ;
        RECT 884.400 727.350 885.600 729.600 ;
        RECT 890.400 727.350 891.600 729.600 ;
        RECT 880.950 724.950 883.050 727.050 ;
        RECT 883.950 724.950 886.050 727.050 ;
        RECT 886.950 724.950 889.050 727.050 ;
        RECT 889.950 724.950 892.050 727.050 ;
        RECT 877.950 721.950 880.050 724.050 ;
        RECT 881.400 723.000 882.600 724.650 ;
        RECT 887.400 723.900 888.600 724.650 ;
        RECT 871.950 719.400 876.450 720.450 ;
        RECT 871.950 718.800 874.050 719.400 ;
        RECT 868.950 712.950 871.050 715.050 ;
        RECT 872.400 712.050 873.450 718.800 ;
        RECT 871.950 709.950 874.050 712.050 ;
        RECT 870.000 702.450 874.050 703.050 ;
        RECT 869.400 700.950 874.050 702.450 ;
        RECT 865.950 694.950 868.050 697.050 ;
        RECT 869.400 688.050 870.450 700.950 ;
        RECT 878.400 694.050 879.450 721.950 ;
        RECT 880.950 720.450 883.050 723.000 ;
        RECT 886.950 721.800 889.050 723.900 ;
        RECT 880.950 720.000 885.450 720.450 ;
        RECT 880.950 719.400 886.050 720.000 ;
        RECT 880.950 718.950 883.050 719.400 ;
        RECT 880.800 715.800 882.900 717.900 ;
        RECT 883.950 715.950 886.050 719.400 ;
        RECT 881.400 709.050 882.450 715.800 ;
        RECT 880.950 706.950 883.050 709.050 ;
        RECT 887.400 699.450 888.450 721.800 ;
        RECT 892.950 712.950 895.050 715.050 ;
        RECT 889.950 709.950 892.050 712.050 ;
        RECT 884.400 698.400 888.450 699.450 ;
        RECT 877.950 691.950 880.050 694.050 ;
        RECT 874.950 688.950 877.050 691.050 ;
        RECT 863.400 686.400 867.450 687.450 ;
        RECT 866.400 684.600 867.450 686.400 ;
        RECT 868.950 685.950 871.050 688.050 ;
        RECT 860.400 684.450 861.600 684.600 ;
        RECT 857.400 683.400 861.600 684.450 ;
        RECT 860.400 682.350 861.600 683.400 ;
        RECT 866.400 682.350 867.600 684.600 ;
        RECT 871.950 683.100 874.050 685.200 ;
        RECT 875.400 685.050 876.450 688.950 ;
        RECT 884.400 688.050 885.450 698.400 ;
        RECT 886.950 688.950 889.050 691.050 ;
        RECT 883.950 685.950 886.050 688.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 679.950 865.050 682.050 ;
        RECT 865.950 679.950 868.050 682.050 ;
        RECT 863.400 678.900 864.600 679.650 ;
        RECT 862.950 676.800 865.050 678.900 ;
        RECT 868.950 676.950 871.050 679.050 ;
        RECT 869.400 673.050 870.450 676.950 ;
        RECT 868.950 670.950 871.050 673.050 ;
        RECT 872.400 670.050 873.450 683.100 ;
        RECT 874.950 682.950 877.050 685.050 ;
        RECT 880.950 683.100 883.050 685.200 ;
        RECT 887.400 684.600 888.450 688.950 ;
        RECT 890.400 685.050 891.450 709.950 ;
        RECT 881.400 682.350 882.600 683.100 ;
        RECT 887.400 682.350 888.600 684.600 ;
        RECT 889.950 682.950 892.050 685.050 ;
        RECT 877.950 679.950 880.050 682.050 ;
        RECT 880.950 679.950 883.050 682.050 ;
        RECT 883.950 679.950 886.050 682.050 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 878.400 677.400 879.600 679.650 ;
        RECT 884.400 677.400 885.600 679.650 ;
        RECT 853.950 667.950 856.050 670.050 ;
        RECT 862.950 667.950 865.050 670.050 ;
        RECT 871.950 667.950 874.050 670.050 ;
        RECT 853.950 664.800 856.050 666.900 ;
        RECT 833.400 653.400 837.450 654.450 ;
        RECT 833.400 651.600 834.450 653.400 ;
        RECT 812.400 649.350 813.600 649.950 ;
        RECT 818.400 649.350 819.600 651.000 ;
        RECT 833.400 649.350 834.600 651.600 ;
        RECT 841.950 650.100 844.050 652.200 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 832.950 646.950 835.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 815.400 644.400 816.600 646.650 ;
        RECT 821.400 645.900 822.600 646.650 ;
        RECT 805.950 640.950 808.050 643.050 ;
        RECT 815.400 642.450 816.450 644.400 ;
        RECT 820.950 643.800 823.050 645.900 ;
        RECT 812.400 641.400 816.450 642.450 ;
        RECT 805.950 637.800 808.050 639.900 ;
        RECT 790.950 634.950 793.050 637.050 ;
        RECT 796.950 634.800 799.050 636.900 ;
        RECT 802.950 634.950 805.050 637.050 ;
        RECT 790.950 605.100 793.050 607.200 ;
        RECT 797.400 607.050 798.450 634.800 ;
        RECT 799.950 631.950 802.050 634.050 ;
        RECT 791.400 604.350 792.600 605.100 ;
        RECT 796.950 604.950 799.050 607.050 ;
        RECT 800.400 604.050 801.450 631.950 ;
        RECT 802.950 607.950 805.050 610.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 794.400 600.000 795.600 601.650 ;
        RECT 793.950 595.950 796.050 600.000 ;
        RECT 799.950 598.800 802.050 600.900 ;
        RECT 800.400 595.050 801.450 598.800 ;
        RECT 799.950 592.950 802.050 595.050 ;
        RECT 803.400 580.050 804.450 607.950 ;
        RECT 806.400 607.050 807.450 637.800 ;
        RECT 808.950 634.950 811.050 637.050 ;
        RECT 805.950 604.950 808.050 607.050 ;
        RECT 809.400 606.600 810.450 634.950 ;
        RECT 812.400 631.050 813.450 641.400 ;
        RECT 817.950 640.950 820.050 643.050 ;
        RECT 814.950 631.950 817.050 634.050 ;
        RECT 811.950 628.950 814.050 631.050 ;
        RECT 815.400 606.600 816.450 631.950 ;
        RECT 818.400 616.050 819.450 640.950 ;
        RECT 827.400 634.050 828.450 646.950 ;
        RECT 836.400 645.900 837.600 646.650 ;
        RECT 835.950 643.800 838.050 645.900 ;
        RECT 842.400 634.050 843.450 650.100 ;
        RECT 844.950 649.950 847.050 655.050 ;
        RECT 850.950 652.950 853.050 655.050 ;
        RECT 847.950 650.100 850.050 652.200 ;
        RECT 854.400 651.600 855.450 664.800 ;
        RECT 863.400 652.050 864.450 667.950 ;
        RECT 878.400 658.050 879.450 677.400 ;
        RECT 880.950 673.950 883.050 676.050 ;
        RECT 877.950 655.950 880.050 658.050 ;
        RECT 848.400 649.350 849.600 650.100 ;
        RECT 854.400 649.350 855.600 651.600 ;
        RECT 862.950 649.950 865.050 652.050 ;
        RECT 865.950 651.600 870.000 652.050 ;
        RECT 865.950 649.950 870.600 651.600 ;
        RECT 874.950 650.100 877.050 652.200 ;
        RECT 881.400 652.050 882.450 673.950 ;
        RECT 884.400 664.050 885.450 677.400 ;
        RECT 889.950 676.950 892.050 679.050 ;
        RECT 883.950 661.950 886.050 664.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 850.950 646.950 853.050 649.050 ;
        RECT 853.950 646.950 856.050 649.050 ;
        RECT 856.950 646.950 859.050 649.050 ;
        RECT 844.950 643.950 847.050 646.050 ;
        RECT 851.400 644.400 852.600 646.650 ;
        RECT 857.400 645.000 858.600 646.650 ;
        RECT 826.950 631.950 829.050 634.050 ;
        RECT 841.950 631.950 844.050 634.050 ;
        RECT 817.950 613.950 820.050 616.050 ;
        RECT 841.950 613.950 844.050 616.050 ;
        RECT 842.400 610.050 843.450 613.950 ;
        RECT 841.950 607.950 844.050 610.050 ;
        RECT 809.400 604.350 810.600 606.600 ;
        RECT 815.400 604.350 816.600 606.600 ;
        RECT 820.950 605.100 823.050 607.200 ;
        RECT 826.950 605.100 829.050 607.200 ;
        RECT 835.950 605.100 838.050 607.200 ;
        RECT 842.400 606.600 843.450 607.950 ;
        RECT 821.400 604.350 822.600 605.100 ;
        RECT 808.950 601.950 811.050 604.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 812.400 599.400 813.600 601.650 ;
        RECT 818.400 600.900 819.600 601.650 ;
        RECT 790.950 577.950 793.050 580.050 ;
        RECT 802.950 577.950 805.050 580.050 ;
        RECT 787.950 574.950 790.050 577.050 ;
        RECT 773.400 571.350 774.600 572.100 ;
        RECT 779.400 571.350 780.600 572.100 ;
        RECT 784.950 571.950 787.050 574.050 ;
        RECT 772.950 568.950 775.050 571.050 ;
        RECT 775.950 568.950 778.050 571.050 ;
        RECT 778.950 568.950 781.050 571.050 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 769.950 565.950 772.050 568.050 ;
        RECT 776.400 566.400 777.600 568.650 ;
        RECT 782.400 567.900 783.600 568.650 ;
        RECT 788.400 567.900 789.450 574.950 ;
        RECT 770.400 556.050 771.450 565.950 ;
        RECT 769.950 553.950 772.050 556.050 ;
        RECT 776.400 553.050 777.450 566.400 ;
        RECT 781.950 565.800 784.050 567.900 ;
        RECT 787.950 565.800 790.050 567.900 ;
        RECT 778.950 553.950 781.050 556.050 ;
        RECT 775.950 550.950 778.050 553.050 ;
        RECT 766.950 538.950 769.050 541.050 ;
        RECT 757.950 528.000 760.050 532.050 ;
        RECT 766.950 528.000 769.050 532.050 ;
        RECT 758.400 526.350 759.600 528.000 ;
        RECT 767.400 526.350 768.600 528.000 ;
        RECT 754.950 523.950 757.050 526.050 ;
        RECT 758.400 523.950 760.500 526.050 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 773.100 523.950 775.200 526.050 ;
        RECT 755.400 520.050 756.450 523.950 ;
        RECT 764.400 522.900 765.600 523.650 ;
        RECT 763.950 520.800 766.050 522.900 ;
        RECT 769.950 520.800 772.050 522.900 ;
        RECT 773.400 522.000 774.600 523.650 ;
        RECT 754.950 517.950 757.050 520.050 ;
        RECT 760.950 517.950 763.050 520.050 ;
        RECT 761.400 511.050 762.450 517.950 ;
        RECT 770.400 517.050 771.450 520.800 ;
        RECT 772.950 517.950 775.050 522.000 ;
        RECT 769.950 514.950 772.050 517.050 ;
        RECT 760.950 508.950 763.050 511.050 ;
        RECT 760.950 499.950 763.050 502.050 ;
        RECT 751.950 496.950 754.050 499.050 ;
        RECT 757.950 496.950 760.050 499.050 ;
        RECT 739.950 493.950 742.050 496.050 ;
        RECT 745.950 494.100 748.050 496.200 ;
        RECT 753.000 495.600 757.050 496.050 ;
        RECT 746.400 493.350 747.600 494.100 ;
        RECT 752.400 493.950 757.050 495.600 ;
        RECT 752.400 493.350 753.600 493.950 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 745.950 490.950 748.050 493.050 ;
        RECT 748.950 490.950 751.050 493.050 ;
        RECT 751.950 490.950 754.050 493.050 ;
        RECT 724.950 481.950 727.050 484.050 ;
        RECT 715.950 469.950 718.050 472.050 ;
        RECT 721.950 457.950 724.050 460.050 ;
        RECT 706.950 454.950 709.050 457.050 ;
        RECT 697.950 448.950 700.050 451.050 ;
        RECT 703.950 449.100 706.050 451.200 ;
        RECT 709.950 449.100 712.050 451.200 ;
        RECT 715.950 449.100 718.050 451.200 ;
        RECT 722.400 450.600 723.450 457.950 ;
        RECT 704.400 448.350 705.600 449.100 ;
        RECT 710.400 448.350 711.600 449.100 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 697.950 442.950 700.050 445.050 ;
        RECT 701.400 444.900 702.600 445.650 ;
        RECT 694.950 433.950 697.050 436.050 ;
        RECT 694.950 427.950 697.050 430.050 ;
        RECT 679.950 424.950 682.050 427.050 ;
        RECT 685.950 424.950 688.050 427.050 ;
        RECT 671.400 415.350 672.600 417.000 ;
        RECT 676.950 415.950 679.050 418.050 ;
        RECT 655.950 412.800 658.050 414.900 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 664.950 412.950 667.050 415.050 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 638.400 388.050 639.450 409.950 ;
        RECT 640.950 409.800 643.050 411.900 ;
        RECT 646.950 409.800 649.050 411.900 ;
        RECT 652.950 409.800 655.050 411.900 ;
        RECT 646.950 400.950 649.050 403.050 ;
        RECT 647.400 394.050 648.450 400.950 ;
        RECT 646.950 391.950 649.050 394.050 ;
        RECT 637.950 385.950 640.050 388.050 ;
        RECT 643.950 379.950 646.050 382.050 ;
        RECT 644.400 372.600 645.450 379.950 ;
        RECT 635.400 371.400 639.450 372.450 ;
        RECT 632.400 370.350 633.600 370.950 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 623.400 367.050 624.600 367.650 ;
        RECT 619.950 365.400 624.600 367.050 ;
        RECT 629.400 365.400 630.600 367.650 ;
        RECT 619.950 364.950 624.000 365.400 ;
        RECT 622.950 352.950 625.050 355.050 ;
        RECT 616.800 343.950 618.900 346.050 ;
        RECT 619.950 343.950 622.050 346.050 ;
        RECT 613.950 340.950 616.050 343.050 ;
        RECT 611.400 337.350 612.600 339.600 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 608.400 333.450 609.600 334.650 ;
        RECT 605.400 332.400 609.600 333.450 ;
        RECT 614.400 332.400 615.600 334.650 ;
        RECT 605.400 325.050 606.450 332.400 ;
        RECT 614.400 328.050 615.450 332.400 ;
        RECT 616.950 331.950 619.050 334.050 ;
        RECT 613.950 325.950 616.050 328.050 ;
        RECT 604.950 322.950 607.050 325.050 ;
        RECT 613.950 322.800 616.050 324.900 ;
        RECT 614.400 316.050 615.450 322.800 ;
        RECT 617.400 319.050 618.450 331.950 ;
        RECT 620.400 319.050 621.450 343.950 ;
        RECT 623.400 340.050 624.450 352.950 ;
        RECT 622.950 337.950 625.050 340.050 ;
        RECT 629.400 339.600 630.450 365.400 ;
        RECT 634.950 343.950 637.050 346.050 ;
        RECT 635.400 339.600 636.450 343.950 ;
        RECT 638.400 340.050 639.450 371.400 ;
        RECT 644.400 370.350 645.600 372.600 ;
        RECT 649.950 371.100 652.050 373.200 ;
        RECT 650.400 370.350 651.600 371.100 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 640.950 364.950 643.050 367.050 ;
        RECT 647.400 365.400 648.600 367.650 ;
        RECT 656.400 366.450 657.450 412.800 ;
        RECT 662.400 410.400 663.600 412.650 ;
        RECT 668.400 410.400 669.600 412.650 ;
        RECT 674.400 411.000 675.600 412.650 ;
        RECT 662.400 391.050 663.450 410.400 ;
        RECT 668.400 406.050 669.450 410.400 ;
        RECT 670.950 406.950 673.050 409.050 ;
        RECT 673.950 406.950 676.050 411.000 ;
        RECT 680.400 409.050 681.450 424.950 ;
        RECT 688.950 421.950 691.050 424.050 ;
        RECT 682.950 415.950 685.050 421.050 ;
        RECT 689.400 417.600 690.450 421.950 ;
        RECT 695.400 418.050 696.450 427.950 ;
        RECT 698.400 421.050 699.450 442.950 ;
        RECT 700.950 442.800 703.050 444.900 ;
        RECT 707.400 443.400 708.600 445.650 ;
        RECT 697.950 418.950 700.050 421.050 ;
        RECT 689.400 415.350 690.600 417.600 ;
        RECT 694.950 415.950 697.050 418.050 ;
        RECT 701.400 417.450 702.450 442.800 ;
        RECT 707.400 436.050 708.450 443.400 ;
        RECT 716.400 439.050 717.450 449.100 ;
        RECT 722.400 448.350 723.600 450.600 ;
        RECT 727.950 450.000 730.050 454.050 ;
        RECT 734.400 451.050 735.450 487.950 ;
        RECT 736.800 487.800 738.900 489.900 ;
        RECT 739.950 487.950 742.050 490.050 ;
        RECT 743.400 488.400 744.600 490.650 ;
        RECT 749.400 488.400 750.600 490.650 ;
        RECT 736.950 460.950 739.050 463.050 ;
        RECT 728.400 448.350 729.600 450.000 ;
        RECT 733.950 448.950 736.050 451.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 718.950 442.950 721.050 445.050 ;
        RECT 725.400 443.400 726.600 445.650 ;
        RECT 731.400 444.900 732.600 445.650 ;
        RECT 737.400 445.050 738.450 460.950 ;
        RECT 740.400 459.450 741.450 487.950 ;
        RECT 743.400 478.050 744.450 488.400 ;
        RECT 742.950 475.950 745.050 478.050 ;
        RECT 745.950 469.950 748.050 472.050 ;
        RECT 740.400 458.400 744.450 459.450 ;
        RECT 739.950 454.950 742.050 457.050 ;
        RECT 715.950 436.950 718.050 439.050 ;
        RECT 706.950 433.950 709.050 436.050 ;
        RECT 715.950 433.800 718.050 435.900 ;
        RECT 716.400 427.050 717.450 433.800 ;
        RECT 719.400 430.050 720.450 442.950 ;
        RECT 721.950 439.950 724.050 442.050 ;
        RECT 718.950 427.950 721.050 430.050 ;
        RECT 715.950 424.950 718.050 427.050 ;
        RECT 718.950 421.950 721.050 424.050 ;
        RECT 698.400 416.400 702.450 417.450 ;
        RECT 703.950 417.000 706.050 421.050 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 686.400 411.900 687.600 412.650 ;
        RECT 692.400 411.900 693.600 412.650 ;
        RECT 685.950 409.800 688.050 411.900 ;
        RECT 691.950 409.800 694.050 411.900 ;
        RECT 679.950 406.950 682.050 409.050 ;
        RECT 667.950 403.950 670.050 406.050 ;
        RECT 661.950 388.950 664.050 391.050 ;
        RECT 667.950 388.950 670.050 391.050 ;
        RECT 661.950 385.800 664.050 387.900 ;
        RECT 662.400 373.200 663.450 385.800 ;
        RECT 668.400 373.200 669.450 388.950 ;
        RECT 661.950 371.100 664.050 373.200 ;
        RECT 667.950 371.100 670.050 373.200 ;
        RECT 671.400 373.050 672.450 406.950 ;
        RECT 686.400 406.050 687.450 409.800 ;
        RECT 692.400 409.050 693.450 409.800 ;
        RECT 688.950 407.400 693.450 409.050 ;
        RECT 688.950 406.950 693.000 407.400 ;
        RECT 694.950 406.950 697.050 409.050 ;
        RECT 675.000 405.450 679.050 406.050 ;
        RECT 674.400 403.950 679.050 405.450 ;
        RECT 685.950 403.950 688.050 406.050 ;
        RECT 674.400 379.050 675.450 403.950 ;
        RECT 676.950 394.950 679.050 397.050 ;
        RECT 673.950 376.950 676.050 379.050 ;
        RECT 662.400 370.350 663.600 371.100 ;
        RECT 668.400 370.350 669.600 371.100 ;
        RECT 670.950 370.950 673.050 373.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 653.400 365.400 657.450 366.450 ;
        RECT 665.400 365.400 666.600 367.650 ;
        RECT 641.400 355.050 642.450 364.950 ;
        RECT 640.950 352.950 643.050 355.050 ;
        RECT 647.400 349.050 648.450 365.400 ;
        RECT 649.950 352.950 652.050 355.050 ;
        RECT 646.950 346.950 649.050 349.050 ;
        RECT 646.950 343.800 649.050 345.900 ;
        RECT 640.950 340.950 643.050 343.050 ;
        RECT 629.400 337.350 630.600 339.600 ;
        RECT 635.400 337.350 636.600 339.600 ;
        RECT 637.950 337.950 640.050 340.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 628.950 334.950 631.050 337.050 ;
        RECT 631.950 334.950 634.050 337.050 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 626.400 333.450 627.600 334.650 ;
        RECT 623.400 332.400 627.600 333.450 ;
        RECT 632.400 333.000 633.600 334.650 ;
        RECT 616.800 316.950 618.900 319.050 ;
        RECT 619.950 316.950 622.050 319.050 ;
        RECT 613.950 313.950 616.050 316.050 ;
        RECT 601.950 306.450 604.050 307.050 ;
        RECT 601.950 305.400 606.450 306.450 ;
        RECT 601.950 304.950 604.050 305.400 ;
        RECT 595.950 295.950 598.050 298.050 ;
        RECT 598.950 296.100 601.050 298.200 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 575.400 287.400 576.600 289.650 ;
        RECT 575.400 280.050 576.450 287.400 ;
        RECT 580.950 283.950 583.050 286.050 ;
        RECT 581.400 280.050 582.450 283.950 ;
        RECT 574.950 277.950 577.050 280.050 ;
        RECT 580.950 277.950 583.050 280.050 ;
        RECT 565.950 274.950 568.050 277.050 ;
        RECT 568.950 268.950 571.050 271.050 ;
        RECT 550.950 259.950 553.050 262.050 ;
        RECT 556.950 260.100 559.050 262.200 ;
        RECT 562.950 260.100 565.050 262.200 ;
        RECT 547.950 226.950 550.050 229.050 ;
        RECT 551.400 220.050 552.450 259.950 ;
        RECT 557.400 259.350 558.600 260.100 ;
        RECT 563.400 259.350 564.600 260.100 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 560.400 254.400 561.600 256.650 ;
        RECT 560.400 238.050 561.450 254.400 ;
        RECT 569.400 249.450 570.450 268.950 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 575.400 261.600 576.450 265.950 ;
        RECT 584.400 265.050 585.450 292.950 ;
        RECT 587.400 271.050 588.450 293.400 ;
        RECT 593.400 292.350 594.600 294.600 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 599.400 292.350 600.600 292.950 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 589.950 283.950 592.050 289.050 ;
        RECT 596.400 288.000 597.600 289.650 ;
        RECT 595.950 283.950 598.050 288.000 ;
        RECT 601.950 286.950 604.050 289.050 ;
        RECT 602.400 280.050 603.450 286.950 ;
        RECT 605.400 283.050 606.450 305.400 ;
        RECT 607.950 295.950 610.050 298.050 ;
        RECT 617.400 297.450 618.450 316.950 ;
        RECT 623.400 304.050 624.450 332.400 ;
        RECT 631.950 328.950 634.050 333.000 ;
        RECT 637.950 331.950 640.050 334.050 ;
        RECT 628.950 325.950 631.050 328.050 ;
        RECT 629.400 316.050 630.450 325.950 ;
        RECT 628.950 313.950 631.050 316.050 ;
        RECT 628.950 310.800 631.050 312.900 ;
        RECT 622.950 301.950 625.050 304.050 ;
        RECT 614.400 296.400 618.450 297.450 ;
        RECT 604.950 280.950 607.050 283.050 ;
        RECT 601.950 277.950 604.050 280.050 ;
        RECT 586.950 268.950 589.050 271.050 ;
        RECT 598.950 268.950 601.050 271.050 ;
        RECT 583.950 262.950 586.050 265.050 ;
        RECT 575.400 259.350 576.600 261.600 ;
        RECT 580.950 260.100 583.050 262.200 ;
        RECT 581.400 259.350 582.600 260.100 ;
        RECT 586.950 259.950 589.050 265.050 ;
        RECT 589.950 262.950 592.050 265.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 583.950 256.950 586.050 259.050 ;
        RECT 578.400 255.900 579.600 256.650 ;
        RECT 584.400 255.900 585.600 256.650 ;
        RECT 577.950 253.800 580.050 255.900 ;
        RECT 583.950 253.800 586.050 255.900 ;
        RECT 566.400 248.400 570.450 249.450 ;
        RECT 562.950 238.950 565.050 241.050 ;
        RECT 559.950 235.950 562.050 238.050 ;
        RECT 563.400 235.050 564.450 238.950 ;
        RECT 562.950 232.950 565.050 235.050 ;
        RECT 550.950 217.950 553.050 220.050 ;
        RECT 532.950 216.600 537.000 217.050 ;
        RECT 532.950 214.950 537.600 216.600 ;
        RECT 541.950 215.100 544.050 217.200 ;
        RECT 536.400 214.350 537.600 214.950 ;
        RECT 542.400 214.350 543.600 215.100 ;
        RECT 550.950 214.800 553.050 216.900 ;
        RECT 556.950 215.100 559.050 217.200 ;
        RECT 563.400 216.600 564.450 232.950 ;
        RECT 566.400 217.200 567.450 248.400 ;
        RECT 590.400 241.050 591.450 262.950 ;
        RECT 599.400 261.600 600.450 268.950 ;
        RECT 604.950 265.950 607.050 268.050 ;
        RECT 599.400 259.350 600.600 261.600 ;
        RECT 595.950 256.950 598.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 592.950 253.950 595.050 256.050 ;
        RECT 596.400 255.900 597.600 256.650 ;
        RECT 593.400 244.050 594.450 253.950 ;
        RECT 595.950 253.800 598.050 255.900 ;
        RECT 601.950 250.950 604.050 256.050 ;
        RECT 605.400 247.050 606.450 265.950 ;
        RECT 608.400 262.050 609.450 295.950 ;
        RECT 614.400 294.600 615.450 296.400 ;
        RECT 614.400 292.350 615.600 294.600 ;
        RECT 619.950 294.000 622.050 298.050 ;
        RECT 623.400 295.050 624.450 301.950 ;
        RECT 625.950 295.950 628.050 298.050 ;
        RECT 620.400 292.350 621.600 294.000 ;
        RECT 622.950 292.950 625.050 295.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 617.400 288.900 618.600 289.650 ;
        RECT 616.950 286.800 619.050 288.900 ;
        RECT 626.400 280.050 627.450 295.950 ;
        RECT 610.950 277.950 613.050 280.050 ;
        RECT 625.950 277.950 628.050 280.050 ;
        RECT 611.400 271.050 612.450 277.950 ;
        RECT 622.950 274.950 625.050 277.050 ;
        RECT 610.950 268.950 613.050 271.050 ;
        RECT 613.950 265.950 616.050 268.050 ;
        RECT 607.950 259.950 610.050 262.050 ;
        RECT 614.400 261.600 615.450 265.950 ;
        RECT 614.400 259.350 615.600 261.600 ;
        RECT 623.400 259.050 624.450 274.950 ;
        RECT 626.400 262.050 627.450 277.950 ;
        RECT 629.400 265.050 630.450 310.800 ;
        RECT 634.950 297.450 637.050 298.050 ;
        RECT 638.400 297.450 639.450 331.950 ;
        RECT 641.400 313.050 642.450 340.950 ;
        RECT 647.400 339.600 648.450 343.800 ;
        RECT 650.400 343.050 651.450 352.950 ;
        RECT 649.950 340.950 652.050 343.050 ;
        RECT 653.400 340.050 654.450 365.400 ;
        RECT 665.400 355.050 666.450 365.400 ;
        RECT 670.950 361.950 673.050 367.050 ;
        RECT 674.400 366.900 675.450 376.950 ;
        RECT 673.950 364.800 676.050 366.900 ;
        RECT 664.950 352.950 667.050 355.050 ;
        RECT 658.950 346.950 661.050 349.050 ;
        RECT 673.950 346.950 676.050 349.050 ;
        RECT 655.950 343.950 658.050 346.050 ;
        RECT 647.400 337.350 648.600 339.600 ;
        RECT 652.950 337.950 655.050 340.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 649.950 334.950 652.050 337.050 ;
        RECT 650.400 333.900 651.600 334.650 ;
        RECT 649.950 331.800 652.050 333.900 ;
        RECT 652.950 331.950 655.050 334.050 ;
        RECT 653.400 328.050 654.450 331.950 ;
        RECT 646.950 325.950 649.050 328.050 ;
        RECT 652.950 325.950 655.050 328.050 ;
        RECT 640.950 310.950 643.050 313.050 ;
        RECT 640.950 304.950 643.050 307.050 ;
        RECT 634.950 296.400 639.450 297.450 ;
        RECT 634.950 295.950 637.050 296.400 ;
        RECT 635.400 294.600 636.450 295.950 ;
        RECT 641.400 294.600 642.450 304.950 ;
        RECT 647.400 295.050 648.450 325.950 ;
        RECT 656.400 325.050 657.450 343.950 ;
        RECT 659.400 331.050 660.450 346.950 ;
        RECT 667.950 338.100 670.050 340.200 ;
        RECT 674.400 339.600 675.450 346.950 ;
        RECT 677.400 340.050 678.450 394.950 ;
        RECT 689.400 382.050 690.450 406.950 ;
        RECT 691.950 403.950 694.050 406.050 ;
        RECT 692.400 391.050 693.450 403.950 ;
        RECT 695.400 403.050 696.450 406.950 ;
        RECT 694.950 400.950 697.050 403.050 ;
        RECT 698.400 400.050 699.450 416.400 ;
        RECT 704.400 415.350 705.600 417.000 ;
        RECT 709.950 416.100 712.050 418.200 ;
        RECT 710.400 415.350 711.600 416.100 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 707.400 411.900 708.600 412.650 ;
        RECT 713.400 411.900 714.600 412.650 ;
        RECT 719.400 411.900 720.450 421.950 ;
        RECT 706.950 409.800 709.050 411.900 ;
        RECT 712.950 409.800 715.050 411.900 ;
        RECT 718.950 409.800 721.050 411.900 ;
        RECT 713.400 403.050 714.450 409.800 ;
        RECT 722.400 409.050 723.450 439.950 ;
        RECT 725.400 436.050 726.450 443.400 ;
        RECT 730.950 442.800 733.050 444.900 ;
        RECT 736.950 442.950 739.050 445.050 ;
        RECT 731.400 439.050 732.450 442.800 ;
        RECT 736.950 439.800 739.050 441.900 ;
        RECT 730.950 436.950 733.050 439.050 ;
        RECT 724.950 433.950 727.050 436.050 ;
        RECT 730.950 416.100 733.050 418.200 ;
        RECT 737.400 418.050 738.450 439.800 ;
        RECT 731.400 415.350 732.600 416.100 ;
        RECT 736.950 415.950 739.050 418.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 728.400 410.400 729.600 412.650 ;
        RECT 734.400 411.000 735.600 412.650 ;
        RECT 715.950 406.950 718.050 409.050 ;
        RECT 721.950 406.950 724.050 409.050 ;
        RECT 712.950 400.950 715.050 403.050 ;
        RECT 697.950 397.950 700.050 400.050 ;
        RECT 716.400 397.050 717.450 406.950 ;
        RECT 718.950 397.950 721.050 400.050 ;
        RECT 715.950 394.950 718.050 397.050 ;
        RECT 719.400 391.050 720.450 397.950 ;
        RECT 725.400 397.050 726.450 409.950 ;
        RECT 724.950 394.950 727.050 397.050 ;
        RECT 691.950 388.950 694.050 391.050 ;
        RECT 718.950 388.950 721.050 391.050 ;
        RECT 697.950 385.950 700.050 388.050 ;
        RECT 715.950 387.900 720.000 388.050 ;
        RECT 715.950 385.950 721.050 387.900 ;
        RECT 721.950 385.950 724.050 388.050 ;
        RECT 724.950 385.950 727.050 391.050 ;
        RECT 688.950 379.950 691.050 382.050 ;
        RECT 694.950 379.950 697.050 382.050 ;
        RECT 682.950 371.100 685.050 373.200 ;
        RECT 688.950 372.000 691.050 376.050 ;
        RECT 695.400 372.600 696.450 379.950 ;
        RECT 698.400 373.050 699.450 385.950 ;
        RECT 718.950 385.800 721.050 385.950 ;
        RECT 712.950 382.950 715.050 385.050 ;
        RECT 706.950 379.950 709.050 382.050 ;
        RECT 700.950 373.950 703.050 376.050 ;
        RECT 683.400 370.350 684.600 371.100 ;
        RECT 689.400 370.350 690.600 372.000 ;
        RECT 695.400 370.350 696.600 372.600 ;
        RECT 697.950 370.950 700.050 373.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 679.950 364.950 682.050 367.050 ;
        RECT 686.400 366.900 687.600 367.650 ;
        RECT 692.400 366.900 693.600 367.650 ;
        RECT 668.400 337.350 669.600 338.100 ;
        RECT 674.400 337.350 675.600 339.600 ;
        RECT 676.950 337.950 679.050 340.050 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 665.400 332.400 666.600 334.650 ;
        RECT 671.400 333.000 672.600 334.650 ;
        RECT 680.400 333.900 681.450 364.950 ;
        RECT 685.950 364.800 688.050 366.900 ;
        RECT 691.950 364.800 694.050 366.900 ;
        RECT 701.400 364.050 702.450 373.950 ;
        RECT 707.400 372.600 708.450 379.950 ;
        RECT 713.400 372.600 714.450 382.950 ;
        RECT 707.400 370.350 708.600 372.600 ;
        RECT 713.400 370.350 714.600 372.600 ;
        RECT 706.950 367.950 709.050 370.050 ;
        RECT 709.950 367.950 712.050 370.050 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 703.950 364.950 706.050 367.050 ;
        RECT 710.400 366.900 711.600 367.650 ;
        RECT 700.950 361.950 703.050 364.050 ;
        RECT 704.400 361.050 705.450 364.950 ;
        RECT 709.950 364.800 712.050 366.900 ;
        RECT 716.400 366.450 717.600 367.650 ;
        RECT 722.400 366.450 723.450 385.950 ;
        RECT 728.400 385.050 729.450 410.400 ;
        RECT 733.950 406.950 736.050 411.000 ;
        RECT 740.400 409.050 741.450 454.950 ;
        RECT 743.400 427.050 744.450 458.400 ;
        RECT 746.400 451.200 747.450 469.950 ;
        RECT 749.400 457.050 750.450 488.400 ;
        RECT 754.950 484.950 757.050 490.050 ;
        RECT 758.400 469.050 759.450 496.950 ;
        RECT 761.400 496.050 762.450 499.950 ;
        RECT 760.950 493.950 763.050 496.050 ;
        RECT 766.950 494.100 769.050 496.200 ;
        RECT 775.950 495.450 778.050 496.200 ;
        RECT 779.400 495.450 780.450 553.950 ;
        RECT 782.400 499.050 783.450 565.800 ;
        RECT 784.950 547.950 787.050 550.050 ;
        RECT 785.400 538.050 786.450 547.950 ;
        RECT 784.950 535.950 787.050 538.050 ;
        RECT 785.400 529.050 786.450 535.950 ;
        RECT 791.400 532.050 792.450 577.950 ;
        RECT 793.950 571.950 796.050 577.050 ;
        RECT 796.950 573.000 799.050 577.050 ;
        RECT 797.400 571.350 798.600 573.000 ;
        RECT 802.950 572.100 805.050 574.200 ;
        RECT 803.400 571.350 804.600 572.100 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 805.950 568.950 808.050 571.050 ;
        RECT 800.400 567.900 801.600 568.650 ;
        RECT 799.950 565.800 802.050 567.900 ;
        RECT 806.400 566.400 807.600 568.650 ;
        RECT 790.950 529.950 793.050 532.050 ;
        RECT 784.950 526.950 787.050 529.050 ;
        RECT 787.950 527.100 790.050 529.200 ;
        RECT 793.950 527.100 796.050 529.200 ;
        RECT 800.400 529.050 801.450 565.800 ;
        RECT 806.400 553.050 807.450 566.400 ;
        RECT 808.950 562.950 811.050 568.050 ;
        RECT 805.950 550.950 808.050 553.050 ;
        RECT 812.400 532.200 813.450 599.400 ;
        RECT 817.950 598.800 820.050 600.900 ;
        RECT 823.950 598.950 826.050 601.050 ;
        RECT 827.400 600.450 828.450 605.100 ;
        RECT 836.400 604.350 837.600 605.100 ;
        RECT 842.400 604.350 843.600 606.600 ;
        RECT 845.400 606.450 846.450 643.950 ;
        RECT 851.400 631.050 852.450 644.400 ;
        RECT 856.950 640.950 859.050 645.000 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 863.400 645.900 864.450 649.950 ;
        RECT 869.400 649.350 870.600 649.950 ;
        RECT 875.400 649.350 876.600 650.100 ;
        RECT 880.950 649.950 883.050 652.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 874.950 646.950 877.050 649.050 ;
        RECT 877.950 646.950 880.050 649.050 ;
        RECT 850.950 628.950 853.050 631.050 ;
        RECT 851.400 616.050 852.450 628.950 ;
        RECT 850.950 613.950 853.050 616.050 ;
        RECT 860.400 615.450 861.450 643.950 ;
        RECT 862.950 643.800 865.050 645.900 ;
        RECT 872.400 644.400 873.600 646.650 ;
        RECT 878.400 644.400 879.600 646.650 ;
        RECT 865.950 640.950 868.050 643.050 ;
        RECT 866.400 637.050 867.450 640.950 ;
        RECT 865.950 634.950 868.050 637.050 ;
        RECT 872.400 616.050 873.450 644.400 ;
        RECT 878.400 634.050 879.450 644.400 ;
        RECT 880.950 643.950 883.050 646.050 ;
        RECT 877.950 631.950 880.050 634.050 ;
        RECT 874.950 616.950 877.050 619.050 ;
        RECT 860.400 614.400 864.450 615.450 ;
        RECT 859.950 610.950 862.050 613.050 ;
        RECT 845.400 605.400 849.450 606.450 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 838.950 601.950 841.050 604.050 ;
        RECT 841.950 601.950 844.050 604.050 ;
        RECT 827.400 599.400 831.450 600.450 ;
        RECT 814.950 592.950 817.050 595.050 ;
        RECT 815.400 559.050 816.450 592.950 ;
        RECT 818.400 574.050 819.450 598.800 ;
        RECT 817.950 571.950 820.050 574.050 ;
        RECT 824.400 573.600 825.450 598.950 ;
        RECT 830.400 574.050 831.450 599.400 ;
        RECT 833.400 599.400 834.600 601.650 ;
        RECT 839.400 600.000 840.600 601.650 ;
        RECT 833.400 592.050 834.450 599.400 ;
        RECT 838.950 595.950 841.050 600.000 ;
        RECT 844.950 598.950 847.050 601.050 ;
        RECT 832.950 589.950 835.050 592.050 ;
        RECT 824.400 571.350 825.600 573.600 ;
        RECT 829.950 571.950 832.050 574.050 ;
        RECT 832.950 572.100 835.050 574.200 ;
        RECT 838.950 572.100 841.050 574.200 ;
        RECT 845.400 573.600 846.450 598.950 ;
        RECT 848.400 580.050 849.450 605.400 ;
        RECT 853.950 605.100 856.050 607.200 ;
        RECT 860.400 606.600 861.450 610.950 ;
        RECT 863.400 610.050 864.450 614.400 ;
        RECT 871.950 613.950 874.050 616.050 ;
        RECT 862.950 607.950 865.050 610.050 ;
        RECT 854.400 604.350 855.600 605.100 ;
        RECT 860.400 604.350 861.600 606.600 ;
        RECT 865.950 606.000 868.050 610.050 ;
        RECT 866.400 604.350 867.600 606.000 ;
        RECT 871.950 605.100 874.050 607.200 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 856.950 601.950 859.050 604.050 ;
        RECT 859.950 601.950 862.050 604.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 857.400 599.400 858.600 601.650 ;
        RECT 863.400 600.000 864.600 601.650 ;
        RECT 857.400 595.050 858.450 599.400 ;
        RECT 862.950 595.950 865.050 600.000 ;
        RECT 856.950 592.950 859.050 595.050 ;
        RECT 862.950 592.800 865.050 594.900 ;
        RECT 847.950 577.950 850.050 580.050 ;
        RECT 853.950 577.950 856.050 580.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 826.950 568.950 829.050 571.050 ;
        RECT 817.950 565.950 820.050 568.050 ;
        RECT 821.400 566.400 822.600 568.650 ;
        RECT 827.400 566.400 828.600 568.650 ;
        RECT 814.950 556.950 817.050 559.050 ;
        RECT 818.400 550.050 819.450 565.950 ;
        RECT 821.400 565.050 822.450 566.400 ;
        RECT 820.950 562.950 823.050 565.050 ;
        RECT 817.950 547.950 820.050 550.050 ;
        RECT 802.950 529.950 805.050 532.050 ;
        RECT 811.950 530.100 814.050 532.200 ;
        RECT 788.400 526.350 789.600 527.100 ;
        RECT 794.400 526.350 795.600 527.100 ;
        RECT 799.950 526.950 802.050 529.050 ;
        RECT 787.950 523.950 790.050 526.050 ;
        RECT 790.950 523.950 793.050 526.050 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 791.400 522.900 792.600 523.650 ;
        RECT 790.950 520.800 793.050 522.900 ;
        RECT 797.400 522.450 798.600 523.650 ;
        RECT 803.400 522.450 804.450 529.950 ;
        RECT 821.400 529.050 822.450 562.950 ;
        RECT 827.400 553.050 828.450 566.400 ;
        RECT 826.950 550.950 829.050 553.050 ;
        RECT 823.950 538.950 826.050 541.050 ;
        RECT 811.950 526.950 814.050 529.050 ;
        RECT 819.000 528.600 823.050 529.050 ;
        RECT 818.400 526.950 823.050 528.600 ;
        RECT 812.400 526.350 813.600 526.950 ;
        RECT 818.400 526.350 819.600 526.950 ;
        RECT 808.950 523.950 811.050 526.050 ;
        RECT 811.950 523.950 814.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 797.400 521.400 804.450 522.450 ;
        RECT 796.950 505.950 799.050 508.050 ;
        RECT 781.950 496.950 784.050 499.050 ;
        RECT 793.950 496.950 796.050 499.050 ;
        RECT 775.950 494.400 780.450 495.450 ;
        RECT 775.950 494.100 778.050 494.400 ;
        RECT 784.950 494.100 787.050 496.200 ;
        RECT 767.400 493.350 768.600 494.100 ;
        RECT 763.950 490.950 766.050 493.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 769.950 490.950 772.050 493.050 ;
        RECT 760.950 487.950 763.050 490.050 ;
        RECT 764.400 489.900 765.600 490.650 ;
        RECT 761.400 469.050 762.450 487.950 ;
        RECT 763.950 487.800 766.050 489.900 ;
        RECT 770.400 488.400 771.600 490.650 ;
        RECT 763.950 486.450 768.000 487.050 ;
        RECT 763.950 484.950 768.450 486.450 ;
        RECT 763.950 481.800 766.050 483.900 ;
        RECT 757.800 466.950 759.900 469.050 ;
        RECT 760.950 466.950 763.050 469.050 ;
        RECT 748.950 456.450 751.050 457.050 ;
        RECT 748.950 455.400 753.450 456.450 ;
        RECT 748.950 454.950 751.050 455.400 ;
        RECT 752.400 453.450 753.450 455.400 ;
        RECT 760.950 454.950 763.050 457.050 ;
        RECT 752.400 452.400 756.450 453.450 ;
        RECT 745.950 449.100 748.050 451.200 ;
        RECT 755.400 450.600 756.450 452.400 ;
        RECT 757.950 451.950 760.050 454.050 ;
        RECT 746.400 448.350 747.600 449.100 ;
        RECT 755.400 448.350 756.600 450.600 ;
        RECT 746.100 445.950 748.200 448.050 ;
        RECT 751.500 445.950 753.600 448.050 ;
        RECT 754.800 445.950 756.900 448.050 ;
        RECT 752.400 444.900 753.600 445.650 ;
        RECT 758.400 444.900 759.450 451.950 ;
        RECT 751.950 442.800 754.050 444.900 ;
        RECT 757.950 442.800 760.050 444.900 ;
        RECT 761.400 433.050 762.450 454.950 ;
        RECT 760.950 430.950 763.050 433.050 ;
        RECT 742.950 424.950 745.050 427.050 ;
        RECT 757.800 424.950 759.900 427.050 ;
        RECT 760.950 424.950 763.050 427.050 ;
        RECT 745.950 421.950 748.050 424.050 ;
        RECT 751.950 421.950 754.050 424.050 ;
        RECT 754.950 421.950 757.050 424.050 ;
        RECT 746.400 417.600 747.450 421.950 ;
        RECT 752.400 417.600 753.450 421.950 ;
        RECT 755.400 418.050 756.450 421.950 ;
        RECT 746.400 415.350 747.600 417.600 ;
        RECT 752.400 415.350 753.600 417.600 ;
        RECT 754.950 415.950 757.050 418.050 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 748.950 412.950 751.050 415.050 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 742.950 409.950 745.050 412.050 ;
        RECT 749.400 410.400 750.600 412.650 ;
        RECT 739.950 406.950 742.050 409.050 ;
        RECT 739.950 400.950 742.050 403.050 ;
        RECT 727.950 382.950 730.050 385.050 ;
        RECT 724.950 376.950 727.050 379.050 ;
        RECT 733.950 376.950 736.050 379.050 ;
        RECT 716.400 365.400 723.450 366.450 ;
        RECT 703.950 358.950 706.050 361.050 ;
        RECT 700.950 352.950 703.050 355.050 ;
        RECT 682.950 337.950 685.050 340.050 ;
        RECT 691.950 338.100 694.050 340.200 ;
        RECT 658.950 328.950 661.050 331.050 ;
        RECT 665.400 328.050 666.450 332.400 ;
        RECT 670.950 328.950 673.050 333.000 ;
        RECT 679.950 331.800 682.050 333.900 ;
        RECT 658.950 325.800 661.050 327.900 ;
        RECT 664.950 325.950 667.050 328.050 ;
        RECT 655.950 322.950 658.050 325.050 ;
        RECT 649.950 304.950 652.050 307.050 ;
        RECT 635.400 292.350 636.600 294.600 ;
        RECT 641.400 292.350 642.600 294.600 ;
        RECT 646.950 292.950 649.050 295.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 638.400 287.400 639.600 289.650 ;
        RECT 644.400 288.900 645.600 289.650 ;
        RECT 631.950 268.950 634.050 271.050 ;
        RECT 628.950 262.950 631.050 265.050 ;
        RECT 625.950 259.950 628.050 262.050 ;
        RECT 632.400 261.600 633.450 268.950 ;
        RECT 638.400 262.200 639.450 287.400 ;
        RECT 643.950 286.800 646.050 288.900 ;
        RECT 644.400 283.050 645.450 286.800 ;
        RECT 643.950 280.950 646.050 283.050 ;
        RECT 640.950 271.950 643.050 274.050 ;
        RECT 632.400 259.350 633.600 261.600 ;
        RECT 637.950 259.950 640.050 262.200 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 622.950 256.950 625.050 259.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 611.400 255.000 612.600 256.650 ;
        RECT 610.950 250.950 613.050 255.000 ;
        RECT 617.400 254.400 618.600 256.650 ;
        RECT 613.950 250.950 616.050 253.050 ;
        RECT 604.950 244.950 607.050 247.050 ;
        RECT 592.950 241.950 595.050 244.050 ;
        RECT 589.950 238.950 592.050 241.050 ;
        RECT 610.950 238.950 613.050 241.050 ;
        RECT 568.950 226.950 571.050 229.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 532.950 208.950 535.050 211.050 ;
        RECT 539.400 210.900 540.600 211.650 ;
        RECT 533.400 193.050 534.450 208.950 ;
        RECT 538.950 208.800 541.050 210.900 ;
        RECT 545.400 209.400 546.600 211.650 ;
        RECT 545.400 205.050 546.450 209.400 ;
        RECT 544.950 202.950 547.050 205.050 ;
        RECT 551.400 202.050 552.450 214.800 ;
        RECT 557.400 214.350 558.600 215.100 ;
        RECT 563.400 214.350 564.600 216.600 ;
        RECT 565.950 215.100 568.050 217.200 ;
        RECT 556.950 211.950 559.050 214.050 ;
        RECT 559.950 211.950 562.050 214.050 ;
        RECT 562.950 211.950 565.050 214.050 ;
        RECT 560.400 210.000 561.600 211.650 ;
        RECT 559.950 205.950 562.050 210.000 ;
        RECT 550.950 199.950 553.050 202.050 ;
        RECT 565.950 199.950 568.050 202.050 ;
        RECT 551.400 196.050 552.450 199.950 ;
        RECT 566.400 196.050 567.450 199.950 ;
        RECT 550.800 193.950 552.900 196.050 ;
        RECT 532.950 190.950 535.050 193.050 ;
        RECT 547.950 190.950 550.050 193.050 ;
        RECT 553.950 192.450 556.050 196.050 ;
        RECT 565.950 193.950 568.050 196.050 ;
        RECT 569.400 193.050 570.450 226.950 ;
        RECT 604.950 223.950 607.050 226.050 ;
        RECT 571.950 220.950 574.050 223.050 ;
        RECT 577.950 220.950 580.050 223.050 ;
        RECT 592.950 220.950 595.050 223.050 ;
        RECT 572.400 202.050 573.450 220.950 ;
        RECT 578.400 216.600 579.450 220.950 ;
        RECT 589.950 217.950 592.050 220.050 ;
        RECT 578.400 214.350 579.600 216.600 ;
        RECT 583.950 215.100 586.050 217.200 ;
        RECT 584.400 214.350 585.600 215.100 ;
        RECT 577.950 211.950 580.050 214.050 ;
        RECT 580.950 211.950 583.050 214.050 ;
        RECT 583.950 211.950 586.050 214.050 ;
        RECT 581.400 209.400 582.600 211.650 ;
        RECT 581.400 205.050 582.450 209.400 ;
        RECT 580.950 202.950 583.050 205.050 ;
        RECT 571.950 199.950 574.050 202.050 ;
        RECT 551.400 192.000 556.050 192.450 ;
        RECT 551.400 191.400 555.450 192.000 ;
        RECT 538.950 182.100 541.050 184.200 ;
        RECT 539.400 181.350 540.600 182.100 ;
        RECT 535.950 178.950 538.050 181.050 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 536.400 177.000 537.600 178.650 ;
        RECT 529.950 172.950 532.050 175.050 ;
        RECT 535.950 172.950 538.050 177.000 ;
        RECT 542.400 176.400 543.600 178.650 ;
        RECT 542.400 163.050 543.450 176.400 ;
        RECT 548.400 166.050 549.450 190.950 ;
        RECT 551.400 177.900 552.450 191.400 ;
        RECT 568.950 190.950 571.050 193.050 ;
        RECT 574.950 190.950 577.050 193.050 ;
        RECT 553.950 187.950 556.050 190.050 ;
        RECT 565.950 187.950 568.050 190.050 ;
        RECT 550.950 175.800 553.050 177.900 ;
        RECT 547.950 163.950 550.050 166.050 ;
        RECT 541.950 160.950 544.050 163.050 ;
        RECT 532.950 154.950 535.050 157.050 ;
        RECT 527.400 137.400 531.450 138.450 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 523.950 133.950 526.050 136.050 ;
        RECT 515.400 132.900 516.600 133.650 ;
        RECT 514.950 130.800 517.050 132.900 ;
        RECT 521.400 131.400 522.600 133.650 ;
        RECT 530.400 132.900 531.450 137.400 ;
        RECT 521.400 129.450 522.450 131.400 ;
        RECT 529.950 130.800 532.050 132.900 ;
        RECT 518.400 128.400 522.450 129.450 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 497.400 104.400 501.450 105.450 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 488.400 99.900 489.600 100.650 ;
        RECT 487.950 97.800 490.050 99.900 ;
        RECT 494.400 98.400 495.600 100.650 ;
        RECT 494.400 91.050 495.450 98.400 ;
        RECT 481.950 88.950 484.050 91.050 ;
        RECT 493.950 88.950 496.050 91.050 ;
        RECT 460.950 82.950 463.050 85.050 ;
        RECT 439.950 76.950 442.050 79.050 ;
        RECT 436.950 59.100 439.050 61.200 ;
        RECT 440.400 60.600 441.450 76.950 ;
        RECT 500.400 70.050 501.450 104.400 ;
        RECT 502.950 104.100 505.050 106.200 ;
        RECT 508.950 104.100 511.050 106.200 ;
        RECT 515.400 105.600 516.450 121.950 ;
        RECT 518.400 106.050 519.450 128.400 ;
        RECT 520.950 124.950 523.050 127.050 ;
        RECT 469.950 67.950 472.050 70.050 ;
        RECT 499.950 67.950 502.050 70.050 ;
        RECT 440.400 58.350 441.600 60.600 ;
        RECT 445.950 59.100 448.050 64.050 ;
        RECT 463.950 60.000 466.050 64.050 ;
        RECT 470.400 61.200 471.450 67.950 ;
        RECT 478.950 61.950 481.050 64.050 ;
        RECT 446.400 58.350 447.600 59.100 ;
        RECT 464.400 58.350 465.600 60.000 ;
        RECT 469.950 59.100 472.050 61.200 ;
        RECT 475.950 59.100 478.050 61.200 ;
        RECT 470.400 58.350 471.600 59.100 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 448.950 55.950 451.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 443.400 53.400 444.600 55.650 ;
        RECT 449.400 54.000 450.600 55.650 ;
        RECT 461.400 54.000 462.600 55.650 ;
        RECT 467.400 54.900 468.600 55.650 ;
        RECT 433.950 49.950 436.050 52.050 ;
        RECT 433.950 28.950 436.050 31.050 ;
        RECT 428.400 26.400 432.450 27.450 ;
        RECT 428.400 25.350 429.600 26.400 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 410.400 20.400 417.450 21.450 ;
        RECT 425.400 20.400 426.600 22.650 ;
        RECT 373.950 13.950 376.050 16.050 ;
        RECT 392.400 13.050 393.450 19.950 ;
        RECT 404.400 16.050 405.450 20.400 ;
        RECT 425.400 16.050 426.450 20.400 ;
        RECT 430.950 19.950 433.050 22.050 ;
        RECT 403.950 13.950 406.050 16.050 ;
        RECT 424.950 13.950 427.050 16.050 ;
        RECT 431.400 13.050 432.450 19.950 ;
        RECT 434.400 19.050 435.450 28.950 ;
        RECT 443.400 27.600 444.450 53.400 ;
        RECT 448.950 49.950 451.050 54.000 ;
        RECT 460.950 49.950 463.050 54.000 ;
        RECT 466.950 52.800 469.050 54.900 ;
        RECT 476.400 49.050 477.450 59.100 ;
        RECT 479.400 55.050 480.450 61.950 ;
        RECT 487.950 60.000 490.050 64.050 ;
        RECT 499.950 61.950 502.050 64.050 ;
        RECT 488.400 58.350 489.600 60.000 ;
        RECT 493.950 59.100 496.050 61.200 ;
        RECT 494.400 58.350 495.600 59.100 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 490.950 55.950 493.050 58.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 478.950 52.950 481.050 55.050 ;
        RECT 485.400 53.400 486.600 55.650 ;
        RECT 491.400 53.400 492.600 55.650 ;
        RECT 475.950 46.950 478.050 49.050 ;
        RECT 460.950 43.950 463.050 46.050 ;
        RECT 454.950 34.950 457.050 37.050 ;
        RECT 443.400 25.350 444.600 27.600 ;
        RECT 448.950 26.100 451.050 28.200 ;
        RECT 449.400 25.350 450.600 26.100 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 445.950 22.950 448.050 25.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 440.400 21.900 441.600 22.650 ;
        RECT 439.950 19.800 442.050 21.900 ;
        RECT 446.400 21.000 447.600 22.650 ;
        RECT 455.400 21.900 456.450 34.950 ;
        RECT 461.400 27.600 462.450 43.950 ;
        RECT 466.950 40.950 469.050 43.050 ;
        RECT 467.400 34.050 468.450 40.950 ;
        RECT 485.400 34.050 486.450 53.400 ;
        RECT 491.400 40.050 492.450 53.400 ;
        RECT 490.950 37.950 493.050 40.050 ;
        RECT 500.400 37.050 501.450 61.950 ;
        RECT 503.400 43.050 504.450 104.100 ;
        RECT 509.400 103.350 510.600 104.100 ;
        RECT 515.400 103.350 516.600 105.600 ;
        RECT 517.950 103.950 520.050 106.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 512.400 99.900 513.600 100.650 ;
        RECT 511.950 97.800 514.050 99.900 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 508.950 60.000 511.050 64.050 ;
        RECT 518.400 61.200 519.450 97.950 ;
        RECT 521.400 94.050 522.450 124.950 ;
        RECT 533.400 105.600 534.450 154.950 ;
        RECT 538.800 142.200 540.900 144.300 ;
        RECT 547.800 142.500 549.900 144.600 ;
        RECT 535.950 137.100 538.050 139.200 ;
        RECT 536.400 136.350 537.600 137.100 ;
        RECT 536.100 133.950 538.200 136.050 ;
        RECT 539.100 129.600 540.000 142.200 ;
        RECT 545.400 139.350 546.600 141.600 ;
        RECT 545.100 136.950 547.200 139.050 ;
        RECT 540.900 135.900 543.000 136.200 ;
        RECT 549.000 135.900 549.900 142.500 ;
        RECT 554.400 139.200 555.450 187.950 ;
        RECT 559.500 185.400 561.600 187.500 ;
        RECT 566.400 187.200 567.600 187.950 ;
        RECT 557.100 178.950 559.200 181.050 ;
        RECT 557.400 177.900 558.600 178.650 ;
        RECT 556.950 175.800 559.050 177.900 ;
        RECT 560.100 172.800 561.000 185.400 ;
        RECT 566.100 184.800 568.200 186.900 ;
        RECT 569.400 185.100 571.500 187.200 ;
        RECT 561.900 183.000 564.000 183.900 ;
        RECT 561.900 181.800 569.100 183.000 ;
        RECT 567.000 180.900 569.100 181.800 ;
        RECT 561.900 180.000 564.000 180.900 ;
        RECT 570.000 180.000 570.900 185.100 ;
        RECT 571.950 182.100 574.050 184.200 ;
        RECT 572.400 181.350 573.600 182.100 ;
        RECT 561.900 179.100 570.900 180.000 ;
        RECT 561.900 178.800 564.000 179.100 ;
        RECT 566.100 175.950 568.200 178.050 ;
        RECT 566.400 173.400 567.600 175.650 ;
        RECT 559.800 170.700 561.900 172.800 ;
        RECT 570.000 172.500 570.900 179.100 ;
        RECT 571.800 178.950 573.900 181.050 ;
        RECT 568.800 170.400 570.900 172.500 ;
        RECT 575.400 172.050 576.450 190.950 ;
        RECT 590.400 187.050 591.450 217.950 ;
        RECT 593.400 202.050 594.450 220.950 ;
        RECT 605.400 220.050 606.450 223.950 ;
        RECT 598.950 219.450 603.000 220.050 ;
        RECT 598.950 217.950 603.450 219.450 ;
        RECT 604.950 217.950 607.050 220.050 ;
        RECT 602.400 216.600 603.450 217.950 ;
        RECT 602.400 214.350 603.600 216.600 ;
        RECT 598.950 211.950 601.050 214.050 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 599.400 210.900 600.600 211.650 ;
        RECT 605.400 210.900 606.600 211.650 ;
        RECT 598.950 208.800 601.050 210.900 ;
        RECT 604.950 208.800 607.050 210.900 ;
        RECT 595.950 205.950 598.050 208.050 ;
        RECT 592.950 199.950 595.050 202.050 ;
        RECT 596.400 196.050 597.450 205.950 ;
        RECT 595.950 193.950 598.050 196.050 ;
        RECT 611.400 187.050 612.450 238.950 ;
        RECT 614.400 210.900 615.450 250.950 ;
        RECT 617.400 238.050 618.450 254.400 ;
        RECT 625.950 253.950 628.050 256.050 ;
        RECT 629.400 254.400 630.600 256.650 ;
        RECT 635.400 255.900 636.600 256.650 ;
        RECT 616.950 235.950 619.050 238.050 ;
        RECT 619.950 232.950 622.050 235.050 ;
        RECT 620.400 216.600 621.450 232.950 ;
        RECT 626.400 216.600 627.450 253.950 ;
        RECT 629.400 238.050 630.450 254.400 ;
        RECT 634.950 253.800 637.050 255.900 ;
        RECT 628.950 235.950 631.050 238.050 ;
        RECT 641.400 229.050 642.450 271.950 ;
        RECT 650.400 268.050 651.450 304.950 ;
        RECT 652.950 301.950 655.050 304.050 ;
        RECT 653.400 295.050 654.450 301.950 ;
        RECT 652.950 292.950 655.050 295.050 ;
        RECT 659.400 294.600 660.450 325.800 ;
        RECT 664.950 295.950 667.050 298.050 ;
        RECT 659.400 292.350 660.600 294.600 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 656.400 288.900 657.600 289.650 ;
        RECT 655.950 286.800 658.050 288.900 ;
        RECT 658.950 280.950 661.050 283.050 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 649.950 260.100 652.050 262.200 ;
        RECT 655.950 260.100 658.050 262.200 ;
        RECT 659.400 262.050 660.450 280.950 ;
        RECT 665.400 274.050 666.450 295.950 ;
        RECT 671.400 294.600 672.450 328.950 ;
        RECT 676.950 322.950 679.050 325.050 ;
        RECT 679.950 322.950 682.050 325.050 ;
        RECT 677.400 294.600 678.450 322.950 ;
        RECT 680.400 316.050 681.450 322.950 ;
        RECT 679.950 313.950 682.050 316.050 ;
        RECT 683.400 307.050 684.450 337.950 ;
        RECT 692.400 337.350 693.600 338.100 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 689.400 333.900 690.600 334.650 ;
        RECT 695.400 333.900 696.600 334.650 ;
        RECT 686.400 325.050 687.450 331.950 ;
        RECT 688.950 331.800 691.050 333.900 ;
        RECT 694.950 331.800 697.050 333.900 ;
        RECT 695.400 328.050 696.450 331.800 ;
        RECT 685.950 322.950 688.050 325.050 ;
        RECT 688.950 322.950 691.050 328.050 ;
        RECT 694.950 325.950 697.050 328.050 ;
        RECT 682.950 304.950 685.050 307.050 ;
        RECT 671.400 292.350 672.600 294.600 ;
        RECT 677.400 292.350 678.600 294.600 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 673.950 289.950 676.050 292.050 ;
        RECT 676.950 289.950 679.050 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 674.400 287.400 675.600 289.650 ;
        RECT 680.400 288.900 681.600 289.650 ;
        RECT 674.400 280.050 675.450 287.400 ;
        RECT 679.800 286.800 681.900 288.900 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 673.950 277.950 676.050 280.050 ;
        RECT 664.950 271.950 667.050 274.050 ;
        RECT 676.950 268.950 679.050 271.050 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 650.400 259.350 651.600 260.100 ;
        RECT 656.400 259.350 657.600 260.100 ;
        RECT 658.950 259.950 661.050 262.050 ;
        RECT 646.950 256.950 649.050 259.050 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 643.950 253.950 646.050 256.050 ;
        RECT 647.400 255.900 648.600 256.650 ;
        RECT 644.400 238.050 645.450 253.950 ;
        RECT 646.950 253.800 649.050 255.900 ;
        RECT 653.400 254.400 654.600 256.650 ;
        RECT 649.950 250.950 652.050 253.050 ;
        RECT 650.400 244.050 651.450 250.950 ;
        RECT 653.400 247.050 654.450 254.400 ;
        RECT 658.950 253.950 661.050 256.050 ;
        RECT 652.950 244.950 655.050 247.050 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 643.950 235.950 646.050 238.050 ;
        RECT 640.950 226.950 643.050 229.050 ;
        RECT 646.950 226.950 649.050 229.050 ;
        RECT 647.400 217.200 648.450 226.950 ;
        RECT 652.950 217.950 655.050 220.050 ;
        RECT 620.400 214.350 621.600 216.600 ;
        RECT 626.400 214.350 627.600 216.600 ;
        RECT 638.400 216.450 639.600 216.600 ;
        RECT 635.400 215.400 639.600 216.450 ;
        RECT 619.950 211.950 622.050 214.050 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 625.950 211.950 628.050 214.050 ;
        RECT 613.950 208.800 616.050 210.900 ;
        RECT 623.400 209.400 624.600 211.650 ;
        RECT 613.950 196.950 616.050 199.050 ;
        RECT 580.950 184.950 583.050 187.050 ;
        RECT 589.950 184.950 592.050 187.050 ;
        RECT 604.950 184.950 607.050 187.050 ;
        RECT 610.950 184.950 613.050 187.050 ;
        RECT 577.950 178.950 580.050 181.050 ;
        RECT 574.950 171.450 577.050 172.050 ;
        RECT 572.400 170.400 577.050 171.450 ;
        RECT 565.950 154.950 568.050 157.050 ;
        RECT 556.950 145.950 559.050 148.050 ;
        RECT 553.950 137.100 556.050 139.200 ;
        RECT 540.900 135.000 549.900 135.900 ;
        RECT 540.900 134.100 543.000 135.000 ;
        RECT 546.000 133.200 548.100 134.100 ;
        RECT 540.900 132.000 548.100 133.200 ;
        RECT 540.900 131.100 543.000 132.000 ;
        RECT 538.500 127.500 540.600 129.600 ;
        RECT 545.100 128.100 547.200 130.200 ;
        RECT 549.000 129.900 549.900 135.000 ;
        RECT 550.800 133.950 552.900 136.050 ;
        RECT 551.400 132.900 552.600 133.650 ;
        RECT 550.950 130.800 553.050 132.900 ;
        RECT 548.400 127.800 550.500 129.900 ;
        RECT 545.400 125.550 546.600 127.800 ;
        RECT 541.950 115.950 544.050 118.050 ;
        RECT 533.400 103.350 534.600 105.600 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 530.400 98.400 531.600 100.650 ;
        RECT 536.400 99.900 537.600 100.650 ;
        RECT 542.400 99.900 543.450 115.950 ;
        RECT 545.400 109.050 546.450 125.550 ;
        RECT 557.400 115.050 558.450 145.950 ;
        RECT 566.400 138.600 567.450 154.950 ;
        RECT 572.400 139.200 573.450 170.400 ;
        RECT 574.950 169.950 577.050 170.400 ;
        RECT 578.400 153.450 579.450 178.950 ;
        RECT 581.400 163.050 582.450 184.950 ;
        RECT 586.950 182.100 589.050 184.200 ;
        RECT 592.950 182.100 595.050 184.200 ;
        RECT 601.950 182.100 604.050 184.200 ;
        RECT 587.400 181.350 588.600 182.100 ;
        RECT 593.400 181.350 594.600 182.100 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 590.400 176.400 591.600 178.650 ;
        RECT 596.400 176.400 597.600 178.650 ;
        RECT 590.400 163.050 591.450 176.400 ;
        RECT 596.400 172.050 597.450 176.400 ;
        RECT 595.950 169.950 598.050 172.050 ;
        RECT 580.950 160.950 583.050 163.050 ;
        RECT 589.950 160.950 592.050 163.050 ;
        RECT 590.400 157.050 591.450 160.950 ;
        RECT 595.950 157.950 598.050 160.050 ;
        RECT 589.950 154.950 592.050 157.050 ;
        RECT 575.400 152.400 579.450 153.450 ;
        RECT 575.400 148.050 576.450 152.400 ;
        RECT 577.950 148.950 580.050 151.050 ;
        RECT 583.950 148.950 586.050 151.050 ;
        RECT 574.950 145.950 577.050 148.050 ;
        RECT 566.400 136.350 567.600 138.600 ;
        RECT 571.950 137.100 574.050 139.200 ;
        RECT 572.400 136.350 573.600 137.100 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 563.400 131.400 564.600 133.650 ;
        RECT 569.400 132.900 570.600 133.650 ;
        RECT 578.400 132.900 579.450 148.950 ;
        RECT 584.400 138.600 585.450 148.950 ;
        RECT 584.400 136.350 585.600 138.600 ;
        RECT 589.950 137.100 592.050 139.200 ;
        RECT 590.400 136.350 591.600 137.100 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 556.950 112.950 559.050 115.050 ;
        RECT 544.950 106.950 547.050 109.050 ;
        RECT 544.950 103.800 547.050 105.900 ;
        RECT 553.950 104.100 556.050 106.200 ;
        RECT 559.950 105.000 562.050 109.050 ;
        RECT 563.400 106.200 564.450 131.400 ;
        RECT 568.950 130.800 571.050 132.900 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 587.400 131.400 588.600 133.650 ;
        RECT 565.950 112.950 568.050 115.050 ;
        RECT 530.400 94.050 531.450 98.400 ;
        RECT 535.950 97.800 538.050 99.900 ;
        RECT 541.950 97.800 544.050 99.900 ;
        RECT 520.950 91.950 523.050 94.050 ;
        RECT 529.950 91.950 532.050 94.050 ;
        RECT 541.950 91.950 544.050 94.050 ;
        RECT 526.950 85.950 529.050 88.050 ;
        RECT 509.400 58.350 510.600 60.000 ;
        RECT 517.950 59.100 520.050 61.200 ;
        RECT 527.400 60.600 528.450 85.950 ;
        RECT 532.950 67.950 535.050 70.050 ;
        RECT 533.400 60.600 534.450 67.950 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 512.400 54.450 513.600 55.650 ;
        RECT 518.400 54.450 519.450 59.100 ;
        RECT 527.400 58.350 528.600 60.600 ;
        RECT 533.400 58.350 534.600 60.600 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 512.400 53.400 519.450 54.450 ;
        RECT 524.400 53.400 525.600 55.650 ;
        RECT 530.400 54.000 531.600 55.650 ;
        RECT 524.400 49.050 525.450 53.400 ;
        RECT 529.950 49.950 532.050 54.000 ;
        RECT 523.950 46.950 526.050 49.050 ;
        RECT 542.400 46.050 543.450 91.950 ;
        RECT 545.400 79.050 546.450 103.800 ;
        RECT 554.400 103.350 555.600 104.100 ;
        RECT 560.400 103.350 561.600 105.000 ;
        RECT 562.950 104.100 565.050 106.200 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 551.400 99.000 552.600 100.650 ;
        RECT 557.400 99.000 558.600 100.650 ;
        RECT 550.950 96.450 553.050 99.000 ;
        RECT 548.400 95.400 553.050 96.450 ;
        RECT 544.950 76.950 547.050 79.050 ;
        RECT 548.400 61.200 549.450 95.400 ;
        RECT 550.950 94.950 553.050 95.400 ;
        RECT 556.950 94.950 559.050 99.000 ;
        RECT 566.400 97.050 567.450 112.950 ;
        RECT 587.400 112.050 588.450 131.400 ;
        RECT 589.950 121.950 592.050 124.050 ;
        RECT 586.950 109.950 589.050 112.050 ;
        RECT 568.950 103.950 571.050 106.050 ;
        RECT 574.950 104.100 577.050 106.200 ;
        RECT 580.950 104.100 583.050 106.200 ;
        RECT 587.400 106.050 588.450 109.950 ;
        RECT 569.400 97.050 570.450 103.950 ;
        RECT 575.400 103.350 576.600 104.100 ;
        RECT 581.400 103.350 582.600 104.100 ;
        RECT 586.950 103.950 589.050 106.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 583.950 100.950 586.050 103.050 ;
        RECT 578.400 98.400 579.600 100.650 ;
        RECT 584.400 99.900 585.600 100.650 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 568.950 94.950 571.050 97.050 ;
        RECT 578.400 88.050 579.450 98.400 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 577.950 85.950 580.050 88.050 ;
        RECT 590.400 82.050 591.450 121.950 ;
        RECT 596.400 121.050 597.450 157.950 ;
        RECT 602.400 151.050 603.450 182.100 ;
        RECT 605.400 177.450 606.450 184.950 ;
        RECT 614.400 183.600 615.450 196.950 ;
        RECT 619.950 193.950 622.050 196.050 ;
        RECT 614.400 181.350 615.600 183.600 ;
        RECT 608.100 178.950 610.200 181.050 ;
        RECT 613.500 178.950 615.600 181.050 ;
        RECT 616.800 178.950 618.900 181.050 ;
        RECT 608.400 177.450 609.600 178.650 ;
        RECT 605.400 177.000 609.600 177.450 ;
        RECT 605.400 176.400 610.050 177.000 ;
        RECT 607.950 172.950 610.050 176.400 ;
        RECT 617.400 176.400 618.600 178.650 ;
        RECT 601.950 148.950 604.050 151.050 ;
        RECT 617.400 142.050 618.450 176.400 ;
        RECT 620.400 166.050 621.450 193.950 ;
        RECT 623.400 169.050 624.450 209.400 ;
        RECT 635.400 190.050 636.450 215.400 ;
        RECT 638.400 214.350 639.600 215.400 ;
        RECT 646.950 215.100 649.050 217.200 ;
        RECT 647.400 214.350 648.600 215.100 ;
        RECT 638.100 211.950 640.200 214.050 ;
        RECT 643.500 211.950 645.600 214.050 ;
        RECT 646.800 211.950 648.900 214.050 ;
        RECT 644.400 210.900 645.600 211.650 ;
        RECT 653.400 210.900 654.450 217.950 ;
        RECT 659.400 216.450 660.450 253.950 ;
        RECT 662.400 220.050 663.450 265.950 ;
        RECT 664.950 259.950 667.050 262.050 ;
        RECT 670.950 260.100 673.050 262.200 ;
        RECT 677.400 261.600 678.450 268.950 ;
        RECT 683.400 262.050 684.450 286.950 ;
        RECT 661.950 217.950 664.050 220.050 ;
        RECT 665.400 219.450 666.450 259.950 ;
        RECT 671.400 259.350 672.600 260.100 ;
        RECT 677.400 259.350 678.600 261.600 ;
        RECT 682.950 259.950 685.050 262.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 667.950 253.950 670.050 256.050 ;
        RECT 674.400 255.000 675.600 256.650 ;
        RECT 680.400 255.900 681.600 256.650 ;
        RECT 668.400 226.050 669.450 253.950 ;
        RECT 673.950 250.950 676.050 255.000 ;
        RECT 679.950 253.800 682.050 255.900 ;
        RECT 680.400 235.050 681.450 253.800 ;
        RECT 679.950 232.950 682.050 235.050 ;
        RECT 686.400 226.050 687.450 322.950 ;
        RECT 701.400 322.050 702.450 352.950 ;
        RECT 704.400 340.050 705.450 358.950 ;
        RECT 712.950 346.950 715.050 349.050 ;
        RECT 703.950 337.950 706.050 340.050 ;
        RECT 706.950 339.000 709.050 343.050 ;
        RECT 713.400 340.050 714.450 346.950 ;
        RECT 707.400 337.350 708.600 339.000 ;
        RECT 712.950 337.950 715.050 340.050 ;
        RECT 706.950 334.950 709.050 337.050 ;
        RECT 709.950 334.950 712.050 337.050 ;
        RECT 710.400 332.400 711.600 334.650 ;
        RECT 710.400 325.050 711.450 332.400 ;
        RECT 712.950 331.950 715.050 334.050 ;
        RECT 709.950 322.950 712.050 325.050 ;
        RECT 688.800 319.800 690.900 321.900 ;
        RECT 691.950 319.950 694.050 322.050 ;
        RECT 700.950 319.950 703.050 322.050 ;
        RECT 689.400 295.050 690.450 319.800 ;
        RECT 692.400 298.050 693.450 319.950 ;
        RECT 694.950 316.950 700.050 319.050 ;
        RECT 702.000 318.900 706.050 319.050 ;
        RECT 700.950 316.950 706.050 318.900 ;
        RECT 700.950 316.800 703.050 316.950 ;
        RECT 700.950 310.950 703.050 313.050 ;
        RECT 691.950 295.950 694.050 298.050 ;
        RECT 688.950 292.950 691.050 295.050 ;
        RECT 694.950 293.100 697.050 295.200 ;
        RECT 695.400 292.350 696.600 293.100 ;
        RECT 691.950 289.950 694.050 292.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 688.950 286.950 691.050 289.050 ;
        RECT 692.400 287.400 693.600 289.650 ;
        RECT 689.400 283.050 690.450 286.950 ;
        RECT 688.950 280.950 691.050 283.050 ;
        RECT 692.400 277.050 693.450 287.400 ;
        RECT 691.950 276.450 694.050 277.050 ;
        RECT 689.400 275.400 694.050 276.450 ;
        RECT 689.400 262.050 690.450 275.400 ;
        RECT 691.950 274.950 694.050 275.400 ;
        RECT 694.950 268.950 697.050 271.050 ;
        RECT 688.950 259.950 691.050 262.050 ;
        RECT 695.400 261.600 696.450 268.950 ;
        RECT 701.400 265.050 702.450 310.950 ;
        RECT 703.950 301.950 706.050 304.050 ;
        RECT 713.400 303.450 714.450 331.950 ;
        RECT 716.400 328.050 717.450 365.400 ;
        RECT 718.950 361.950 721.050 364.050 ;
        RECT 721.950 361.950 724.050 364.050 ;
        RECT 719.400 355.050 720.450 361.950 ;
        RECT 722.400 355.050 723.450 361.950 ;
        RECT 718.800 352.950 720.900 355.050 ;
        RECT 721.950 352.950 724.050 355.050 ;
        RECT 718.950 349.800 721.050 351.900 ;
        RECT 719.400 340.050 720.450 349.800 ;
        RECT 718.950 337.950 721.050 340.050 ;
        RECT 722.400 339.600 723.450 352.950 ;
        RECT 725.400 343.050 726.450 376.950 ;
        RECT 734.400 372.600 735.450 376.950 ;
        RECT 740.400 373.050 741.450 400.950 ;
        RECT 734.400 370.350 735.600 372.600 ;
        RECT 739.950 370.950 742.050 373.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 731.400 366.000 732.600 367.650 ;
        RECT 737.400 366.900 738.600 367.650 ;
        RECT 730.950 361.950 733.050 366.000 ;
        RECT 736.950 364.800 739.050 366.900 ;
        RECT 727.950 346.950 730.050 349.050 ;
        RECT 724.950 340.950 727.050 343.050 ;
        RECT 728.400 339.600 729.450 346.950 ;
        RECT 743.400 345.450 744.450 409.950 ;
        RECT 749.400 406.050 750.450 410.400 ;
        RECT 754.950 409.950 757.050 412.050 ;
        RECT 748.950 403.950 751.050 406.050 ;
        RECT 755.400 391.050 756.450 409.950 ;
        RECT 754.950 388.950 757.050 391.050 ;
        RECT 748.950 371.100 751.050 373.200 ;
        RECT 749.400 370.350 750.600 371.100 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 752.400 365.400 753.600 367.650 ;
        RECT 748.950 361.950 751.050 364.050 ;
        RECT 749.400 358.050 750.450 361.950 ;
        RECT 748.950 355.950 751.050 358.050 ;
        RECT 740.400 344.400 744.450 345.450 ;
        RECT 736.950 340.950 739.050 343.050 ;
        RECT 722.400 337.350 723.600 339.600 ;
        RECT 728.400 337.350 729.600 339.600 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 727.950 334.950 730.050 337.050 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 718.950 331.950 721.050 334.050 ;
        RECT 725.400 333.900 726.600 334.650 ;
        RECT 715.950 325.950 718.050 328.050 ;
        RECT 719.400 322.050 720.450 331.950 ;
        RECT 724.950 331.800 727.050 333.900 ;
        RECT 731.400 332.400 732.600 334.650 ;
        RECT 731.400 328.050 732.450 332.400 ;
        RECT 733.950 331.950 736.050 334.050 ;
        RECT 737.400 333.900 738.450 340.950 ;
        RECT 740.400 340.050 741.450 344.400 ;
        RECT 739.950 337.950 742.050 340.050 ;
        RECT 742.950 338.100 745.050 340.200 ;
        RECT 749.400 339.600 750.450 355.950 ;
        RECT 752.400 352.050 753.450 365.400 ;
        RECT 751.950 349.950 754.050 352.050 ;
        RECT 743.400 337.350 744.600 338.100 ;
        RECT 749.400 337.350 750.600 339.600 ;
        RECT 754.950 337.950 757.050 343.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 746.400 333.900 747.600 334.650 ;
        RECT 752.400 333.900 753.600 334.650 ;
        RECT 730.950 325.950 733.050 328.050 ;
        RECT 718.950 319.950 721.050 322.050 ;
        RECT 734.400 304.050 735.450 331.950 ;
        RECT 736.950 331.800 739.050 333.900 ;
        RECT 745.950 331.800 748.050 333.900 ;
        RECT 751.950 331.800 754.050 333.900 ;
        RECT 754.950 331.950 757.050 334.050 ;
        RECT 755.400 316.050 756.450 331.950 ;
        RECT 754.950 313.950 757.050 316.050 ;
        RECT 713.400 302.400 717.450 303.450 ;
        RECT 704.400 288.450 705.450 301.950 ;
        RECT 710.100 298.500 712.200 300.600 ;
        RECT 707.100 289.950 709.200 292.050 ;
        RECT 710.100 291.900 711.000 298.500 ;
        RECT 716.400 298.050 717.450 302.400 ;
        RECT 727.950 301.950 730.050 304.050 ;
        RECT 733.950 301.950 736.050 304.050 ;
        RECT 719.100 298.200 721.200 300.300 ;
        RECT 724.950 298.950 727.050 301.050 ;
        RECT 713.400 295.350 714.600 297.600 ;
        RECT 715.950 295.950 718.050 298.050 ;
        RECT 712.800 292.950 714.900 295.050 ;
        RECT 717.000 291.900 719.100 292.200 ;
        RECT 710.100 291.000 719.100 291.900 ;
        RECT 707.400 288.450 708.600 289.650 ;
        RECT 704.400 287.400 708.600 288.450 ;
        RECT 710.100 285.900 711.000 291.000 ;
        RECT 717.000 290.100 719.100 291.000 ;
        RECT 711.900 289.200 714.000 290.100 ;
        RECT 711.900 288.000 719.100 289.200 ;
        RECT 717.000 287.100 719.100 288.000 ;
        RECT 709.500 283.800 711.600 285.900 ;
        RECT 712.800 284.100 714.900 286.200 ;
        RECT 720.000 285.600 720.900 298.200 ;
        RECT 722.400 294.450 723.600 294.600 ;
        RECT 725.400 294.450 726.450 298.950 ;
        RECT 722.400 293.400 726.450 294.450 ;
        RECT 722.400 292.350 723.600 293.400 ;
        RECT 721.800 289.950 723.900 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 713.400 283.050 714.600 283.800 ;
        RECT 719.400 283.500 721.500 285.600 ;
        RECT 712.950 280.950 715.050 283.050 ;
        RECT 706.950 277.950 709.050 280.050 ;
        RECT 700.950 262.950 703.050 265.050 ;
        RECT 702.000 261.600 706.050 262.050 ;
        RECT 695.400 259.350 696.600 261.600 ;
        RECT 701.400 259.950 706.050 261.600 ;
        RECT 701.400 259.350 702.600 259.950 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 692.400 255.900 693.600 256.650 ;
        RECT 691.950 253.800 694.050 255.900 ;
        RECT 698.400 255.000 699.600 256.650 ;
        RECT 697.950 250.950 700.050 255.000 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 700.950 250.950 703.050 253.050 ;
        RECT 667.950 223.950 670.050 226.050 ;
        RECT 679.950 223.950 682.050 226.050 ;
        RECT 685.950 223.950 688.050 226.050 ;
        RECT 676.950 220.950 679.050 223.050 ;
        RECT 665.400 218.400 669.450 219.450 ;
        RECT 668.400 216.600 669.450 218.400 ;
        RECT 662.400 216.450 663.600 216.600 ;
        RECT 659.400 215.400 663.600 216.450 ;
        RECT 662.400 214.350 663.600 215.400 ;
        RECT 668.400 214.350 669.600 216.600 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 643.950 208.800 646.050 210.900 ;
        RECT 652.950 208.800 655.050 210.900 ;
        RECT 665.400 209.400 666.600 211.650 ;
        RECT 646.950 205.950 649.050 208.050 ;
        RECT 661.950 205.950 664.050 208.050 ;
        RECT 647.400 202.050 648.450 205.950 ;
        RECT 658.950 202.950 661.050 205.050 ;
        RECT 646.950 199.950 649.050 202.050 ;
        RECT 659.400 199.050 660.450 202.950 ;
        RECT 662.400 202.050 663.450 205.950 ;
        RECT 661.950 199.950 664.050 202.050 ;
        RECT 652.950 196.950 655.050 199.050 ;
        RECT 658.950 196.950 661.050 199.050 ;
        RECT 625.950 187.950 628.050 190.050 ;
        RECT 634.950 187.950 637.050 190.050 ;
        RECT 622.950 166.950 625.050 169.050 ;
        RECT 619.950 163.950 622.050 166.050 ;
        RECT 626.400 160.050 627.450 187.950 ;
        RECT 653.400 184.200 654.450 196.950 ;
        RECT 665.400 193.050 666.450 209.400 ;
        RECT 664.950 190.950 667.050 193.050 ;
        RECT 634.950 182.100 637.050 184.200 ;
        RECT 652.950 182.100 655.050 184.200 ;
        RECT 658.950 183.000 661.050 187.050 ;
        RECT 667.950 184.950 670.050 187.050 ;
        RECT 635.400 181.350 636.600 182.100 ;
        RECT 653.400 181.350 654.600 182.100 ;
        RECT 659.400 181.350 660.600 183.000 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 628.950 175.950 631.050 178.050 ;
        RECT 632.400 177.000 633.600 178.650 ;
        RECT 638.400 177.900 639.600 178.650 ;
        RECT 625.950 157.950 628.050 160.050 ;
        RECT 629.400 151.050 630.450 175.950 ;
        RECT 631.950 172.950 634.050 177.000 ;
        RECT 637.950 175.800 640.050 177.900 ;
        RECT 650.400 177.000 651.600 178.650 ;
        RECT 649.950 172.950 652.050 177.000 ;
        RECT 656.400 176.400 657.600 178.650 ;
        RECT 662.400 176.400 663.600 178.650 ;
        RECT 637.950 157.950 640.050 160.050 ;
        RECT 656.400 159.450 657.450 176.400 ;
        RECT 662.400 172.050 663.450 176.400 ;
        RECT 661.950 169.950 664.050 172.050 ;
        RECT 662.400 160.050 663.450 169.950 ;
        RECT 656.400 158.400 660.450 159.450 ;
        RECT 628.950 148.950 631.050 151.050 ;
        RECT 616.950 139.950 619.050 142.050 ;
        RECT 601.950 137.100 604.050 139.200 ;
        RECT 607.950 137.100 610.050 139.200 ;
        RECT 625.950 138.000 628.050 142.050 ;
        RECT 602.400 136.350 603.600 137.100 ;
        RECT 608.400 136.350 609.600 137.100 ;
        RECT 626.400 136.350 627.600 138.000 ;
        RECT 631.950 137.100 634.050 142.050 ;
        RECT 634.950 139.950 637.050 145.050 ;
        RECT 632.400 136.350 633.600 137.100 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 610.950 133.950 613.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 631.950 133.950 634.050 136.050 ;
        RECT 605.400 132.000 606.600 133.650 ;
        RECT 604.950 127.950 607.050 132.000 ;
        RECT 611.400 131.400 612.600 133.650 ;
        RECT 611.400 121.050 612.450 131.400 ;
        RECT 595.950 118.950 598.050 121.050 ;
        RECT 610.950 118.950 613.050 121.050 ;
        RECT 617.400 115.050 618.450 133.950 ;
        RECT 623.400 131.400 624.600 133.650 ;
        RECT 629.400 132.900 630.600 133.650 ;
        RECT 638.400 132.900 639.450 157.950 ;
        RECT 655.950 154.950 658.050 157.050 ;
        RECT 649.950 137.100 652.050 139.200 ;
        RECT 656.400 138.600 657.450 154.950 ;
        RECT 650.400 136.350 651.600 137.100 ;
        RECT 656.400 136.350 657.600 138.600 ;
        RECT 659.400 138.450 660.450 158.400 ;
        RECT 661.950 157.950 664.050 160.050 ;
        RECT 668.400 157.050 669.450 184.950 ;
        RECT 670.950 181.950 673.050 184.050 ;
        RECT 677.400 183.600 678.450 220.950 ;
        RECT 680.400 186.450 681.450 223.950 ;
        RECT 686.100 220.500 688.200 222.600 ;
        RECT 683.100 211.950 685.200 214.050 ;
        RECT 686.100 213.900 687.000 220.500 ;
        RECT 695.100 220.200 697.200 222.300 ;
        RECT 689.400 217.350 690.600 219.600 ;
        RECT 688.800 214.950 690.900 217.050 ;
        RECT 693.000 213.900 695.100 214.200 ;
        RECT 686.100 213.000 695.100 213.900 ;
        RECT 683.400 210.900 684.600 211.650 ;
        RECT 682.950 208.800 685.050 210.900 ;
        RECT 686.100 207.900 687.000 213.000 ;
        RECT 693.000 212.100 695.100 213.000 ;
        RECT 687.900 211.200 690.000 212.100 ;
        RECT 687.900 210.000 695.100 211.200 ;
        RECT 693.000 209.100 695.100 210.000 ;
        RECT 685.500 205.800 687.600 207.900 ;
        RECT 688.800 206.100 690.900 208.200 ;
        RECT 696.000 207.600 696.900 220.200 ;
        RECT 697.950 215.100 700.050 217.200 ;
        RECT 698.400 214.350 699.600 215.100 ;
        RECT 697.800 211.950 699.900 214.050 ;
        RECT 689.400 203.550 690.600 205.800 ;
        RECT 695.400 205.500 697.500 207.600 ;
        RECT 680.400 185.400 684.450 186.450 ;
        RECT 683.400 183.600 684.450 185.400 ;
        RECT 671.400 163.050 672.450 181.950 ;
        RECT 677.400 181.350 678.600 183.600 ;
        RECT 683.400 181.350 684.600 183.600 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 682.950 178.950 685.050 181.050 ;
        RECT 680.400 177.000 681.600 178.650 ;
        RECT 679.950 172.950 682.050 177.000 ;
        RECT 682.950 169.950 685.050 172.050 ;
        RECT 670.950 160.950 673.050 163.050 ;
        RECT 667.950 154.950 670.050 157.050 ;
        RECT 664.950 139.950 667.050 142.050 ;
        RECT 659.400 137.400 663.450 138.450 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 655.950 133.950 658.050 136.050 ;
        RECT 623.400 115.050 624.450 131.400 ;
        RECT 628.950 130.800 631.050 132.900 ;
        RECT 637.950 130.800 640.050 132.900 ;
        RECT 647.400 131.400 648.600 133.650 ;
        RECT 653.400 132.900 654.600 133.650 ;
        RECT 647.400 124.050 648.450 131.400 ;
        RECT 652.950 130.800 655.050 132.900 ;
        RECT 662.400 127.050 663.450 137.400 ;
        RECT 661.950 124.950 664.050 127.050 ;
        RECT 646.950 121.950 649.050 124.050 ;
        RECT 625.950 118.950 628.050 121.050 ;
        RECT 610.950 112.950 613.050 115.050 ;
        RECT 616.950 112.950 619.050 115.050 ;
        RECT 622.950 112.950 625.050 115.050 ;
        RECT 598.950 104.100 601.050 106.200 ;
        RECT 599.400 103.350 600.600 104.100 ;
        RECT 607.950 103.950 610.050 106.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 596.400 99.900 597.600 100.650 ;
        RECT 602.400 99.900 603.600 100.650 ;
        RECT 595.950 97.800 598.050 99.900 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 601.950 91.950 604.050 94.050 ;
        RECT 589.950 79.950 592.050 82.050 ;
        RECT 586.950 73.950 589.050 76.050 ;
        RECT 553.950 67.950 556.050 70.050 ;
        RECT 571.950 67.950 574.050 70.050 ;
        RECT 547.950 59.100 550.050 61.200 ;
        RECT 554.400 60.600 555.450 67.950 ;
        RECT 572.400 60.600 573.450 67.950 ;
        RECT 548.400 58.350 549.600 59.100 ;
        RECT 554.400 58.350 555.600 60.600 ;
        RECT 572.400 58.350 573.600 60.600 ;
        RECT 577.950 59.100 580.050 61.200 ;
        RECT 578.400 58.350 579.600 59.100 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 580.950 55.950 583.050 58.050 ;
        RECT 551.400 54.900 552.600 55.650 ;
        RECT 550.950 49.950 553.050 54.900 ;
        RECT 557.400 53.400 558.600 55.650 ;
        RECT 575.400 54.000 576.600 55.650 ;
        RECT 581.400 54.000 582.600 55.650 ;
        RECT 587.400 55.050 588.450 73.950 ;
        RECT 602.400 70.050 603.450 91.950 ;
        RECT 608.400 76.050 609.450 103.950 ;
        RECT 611.400 99.900 612.450 112.950 ;
        RECT 617.400 105.600 618.450 112.950 ;
        RECT 622.950 109.800 625.050 111.900 ;
        RECT 623.400 105.600 624.450 109.800 ;
        RECT 626.400 106.050 627.450 118.950 ;
        RECT 628.950 115.950 631.050 118.050 ;
        RECT 617.400 103.350 618.600 105.600 ;
        RECT 623.400 103.350 624.600 105.600 ;
        RECT 625.950 103.950 628.050 106.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 622.950 100.950 625.050 103.050 ;
        RECT 610.950 97.800 613.050 99.900 ;
        RECT 620.400 98.400 621.600 100.650 ;
        RECT 620.400 88.050 621.450 98.400 ;
        RECT 629.400 94.050 630.450 115.950 ;
        RECT 640.950 112.950 643.050 115.050 ;
        RECT 652.950 114.450 655.050 115.050 ;
        RECT 652.950 113.400 663.450 114.450 ;
        RECT 652.950 112.950 655.050 113.400 ;
        RECT 631.950 106.950 634.050 109.050 ;
        RECT 632.400 99.900 633.450 106.950 ;
        RECT 641.400 105.600 642.450 112.950 ;
        RECT 655.950 109.950 658.050 112.050 ;
        RECT 641.400 103.350 642.600 105.600 ;
        RECT 646.950 105.000 649.050 109.050 ;
        RECT 652.950 106.950 655.050 109.050 ;
        RECT 647.400 103.350 648.600 105.000 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 640.950 100.950 643.050 103.050 ;
        RECT 643.950 100.950 646.050 103.050 ;
        RECT 646.950 100.950 649.050 103.050 ;
        RECT 638.400 100.050 639.600 100.650 ;
        RECT 631.950 97.800 634.050 99.900 ;
        RECT 634.950 98.400 639.600 100.050 ;
        RECT 644.400 99.900 645.600 100.650 ;
        RECT 634.950 97.950 639.000 98.400 ;
        RECT 643.950 97.800 646.050 99.900 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 619.950 85.950 622.050 88.050 ;
        RECT 607.950 73.950 610.050 76.050 ;
        RECT 640.950 73.950 643.050 76.050 ;
        RECT 601.950 67.950 604.050 70.050 ;
        RECT 607.950 67.950 610.050 70.050 ;
        RECT 634.950 67.950 637.050 70.050 ;
        RECT 595.950 60.000 598.050 64.050 ;
        RECT 602.400 60.600 603.450 67.950 ;
        RECT 596.400 58.350 597.600 60.000 ;
        RECT 602.400 58.350 603.600 60.600 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 557.400 49.050 558.450 53.400 ;
        RECT 574.950 49.950 577.050 54.000 ;
        RECT 580.950 49.950 583.050 54.000 ;
        RECT 586.950 52.950 589.050 55.050 ;
        RECT 593.400 53.400 594.600 55.650 ;
        RECT 599.400 54.900 600.600 55.650 ;
        RECT 608.400 54.900 609.450 67.950 ;
        RECT 628.950 64.950 631.050 67.050 ;
        RECT 613.950 59.100 616.050 61.200 ;
        RECT 619.950 60.000 622.050 64.050 ;
        RECT 614.400 58.350 615.600 59.100 ;
        RECT 620.400 58.350 621.600 60.000 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 617.400 54.900 618.600 55.650 ;
        RECT 556.950 46.950 559.050 49.050 ;
        RECT 571.950 48.450 574.050 49.050 ;
        RECT 577.950 48.450 580.050 49.050 ;
        RECT 571.950 47.400 580.050 48.450 ;
        RECT 571.950 46.950 574.050 47.400 ;
        RECT 577.950 46.950 580.050 47.400 ;
        RECT 593.400 46.050 594.450 53.400 ;
        RECT 595.950 49.050 598.050 52.050 ;
        RECT 598.950 49.950 601.050 54.900 ;
        RECT 607.950 52.800 610.050 54.900 ;
        RECT 616.950 52.800 619.050 54.900 ;
        RECT 623.400 53.400 624.600 55.650 ;
        RECT 610.950 51.450 613.050 52.050 ;
        RECT 619.950 51.450 622.050 52.050 ;
        RECT 610.950 50.400 622.050 51.450 ;
        RECT 610.950 49.950 613.050 50.400 ;
        RECT 619.950 49.950 622.050 50.400 ;
        RECT 595.800 48.000 598.050 49.050 ;
        RECT 595.800 46.950 597.900 48.000 ;
        RECT 541.950 43.950 544.050 46.050 ;
        RECT 547.950 43.950 550.050 46.050 ;
        RECT 592.950 43.950 595.050 46.050 ;
        RECT 610.950 43.950 613.050 46.050 ;
        RECT 502.950 40.950 505.050 43.050 ;
        RECT 526.950 40.950 529.050 43.050 ;
        RECT 499.950 34.950 502.050 37.050 ;
        RECT 466.950 31.950 469.050 34.050 ;
        RECT 484.950 31.950 487.050 34.050 ;
        RECT 496.950 31.950 499.050 34.050 ;
        RECT 508.950 31.950 511.050 34.050 ;
        RECT 467.400 27.600 468.450 31.950 ;
        RECT 461.400 25.350 462.600 27.600 ;
        RECT 467.400 25.350 468.600 27.600 ;
        RECT 475.950 25.950 478.050 28.050 ;
        RECT 484.950 26.100 487.050 28.200 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 469.950 22.950 472.050 25.050 ;
        RECT 433.950 16.950 436.050 19.050 ;
        RECT 445.950 16.950 448.050 21.000 ;
        RECT 454.950 19.800 457.050 21.900 ;
        RECT 464.400 20.400 465.600 22.650 ;
        RECT 470.400 21.900 471.600 22.650 ;
        RECT 464.400 16.050 465.450 20.400 ;
        RECT 469.950 19.800 472.050 21.900 ;
        RECT 463.950 13.950 466.050 16.050 ;
        RECT 238.950 11.400 246.450 12.450 ;
        RECT 238.950 10.950 241.050 11.400 ;
        RECT 322.950 10.950 325.050 13.050 ;
        RECT 391.950 10.950 394.050 13.050 ;
        RECT 430.950 10.950 433.050 13.050 ;
        RECT 476.400 7.050 477.450 25.950 ;
        RECT 485.400 25.350 486.600 26.100 ;
        RECT 493.950 25.950 496.050 28.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 482.400 21.900 483.600 22.650 ;
        RECT 488.400 22.050 489.600 22.650 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 488.400 20.400 493.050 22.050 ;
        RECT 489.000 19.950 493.050 20.400 ;
        RECT 494.400 13.050 495.450 25.950 ;
        RECT 497.400 22.050 498.450 31.950 ;
        RECT 502.950 26.100 505.050 28.200 ;
        RECT 509.400 27.600 510.450 31.950 ;
        RECT 517.950 28.950 520.050 31.050 ;
        RECT 503.400 25.350 504.600 26.100 ;
        RECT 509.400 25.350 510.600 27.600 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 496.950 19.950 499.050 22.050 ;
        RECT 506.400 20.400 507.600 22.650 ;
        RECT 512.400 21.450 513.600 22.650 ;
        RECT 518.400 21.450 519.450 28.950 ;
        RECT 527.400 27.600 528.450 40.950 ;
        RECT 527.400 25.350 528.600 27.600 ;
        RECT 532.950 26.100 535.050 28.200 ;
        RECT 548.400 27.600 549.450 43.950 ;
        RECT 565.950 40.950 568.050 43.050 ;
        RECT 562.950 31.950 565.050 34.050 ;
        RECT 533.400 25.350 534.600 26.100 ;
        RECT 548.400 25.350 549.600 27.600 ;
        RECT 553.950 26.100 556.050 28.200 ;
        RECT 554.400 25.350 555.600 26.100 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 550.950 22.950 553.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 512.400 20.400 519.450 21.450 ;
        RECT 530.400 21.000 531.600 22.650 ;
        RECT 536.400 21.900 537.600 22.650 ;
        RECT 493.950 10.950 496.050 13.050 ;
        RECT 506.400 7.050 507.450 20.400 ;
        RECT 529.950 16.950 532.050 21.000 ;
        RECT 535.950 19.800 538.050 21.900 ;
        RECT 551.400 21.000 552.600 22.650 ;
        RECT 557.400 21.900 558.600 22.650 ;
        RECT 563.400 21.900 564.450 31.950 ;
        RECT 538.950 16.950 544.050 19.050 ;
        RECT 550.950 16.950 553.050 21.000 ;
        RECT 556.950 19.800 559.050 21.900 ;
        RECT 562.950 19.800 565.050 21.900 ;
        RECT 566.400 19.050 567.450 40.950 ;
        RECT 592.950 37.950 595.050 40.050 ;
        RECT 596.400 38.400 606.450 39.450 ;
        RECT 568.950 34.950 571.050 37.050 ;
        RECT 586.950 34.950 589.050 37.050 ;
        RECT 569.400 28.200 570.450 34.950 ;
        RECT 568.950 26.100 571.050 28.200 ;
        RECT 574.950 26.100 577.050 28.200 ;
        RECT 580.950 26.100 583.050 28.200 ;
        RECT 575.400 25.350 576.600 26.100 ;
        RECT 581.400 25.350 582.600 26.100 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 572.400 21.900 573.600 22.650 ;
        RECT 571.950 19.800 574.050 21.900 ;
        RECT 578.400 20.400 579.600 22.650 ;
        RECT 587.400 22.050 588.450 34.950 ;
        RECT 593.400 28.050 594.450 37.950 ;
        RECT 592.950 25.950 595.050 28.050 ;
        RECT 596.400 27.600 597.450 38.400 ;
        RECT 601.950 34.950 604.050 37.050 ;
        RECT 602.400 27.600 603.450 34.950 ;
        RECT 605.400 30.450 606.450 38.400 ;
        RECT 605.400 30.000 609.450 30.450 ;
        RECT 605.400 29.400 610.050 30.000 ;
        RECT 596.400 25.350 597.600 27.600 ;
        RECT 602.400 25.350 603.600 27.600 ;
        RECT 607.950 25.950 610.050 29.400 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 565.950 16.950 568.050 19.050 ;
        RECT 574.950 16.950 577.050 19.050 ;
        RECT 575.400 13.050 576.450 16.950 ;
        RECT 574.950 10.950 577.050 13.050 ;
        RECT 578.400 10.050 579.450 20.400 ;
        RECT 586.950 19.950 589.050 22.050 ;
        RECT 590.400 19.050 591.450 22.950 ;
        RECT 592.950 19.950 595.050 22.050 ;
        RECT 599.400 21.900 600.600 22.650 ;
        RECT 589.950 16.950 592.050 19.050 ;
        RECT 593.400 16.050 594.450 19.950 ;
        RECT 598.950 19.800 601.050 21.900 ;
        RECT 605.400 20.400 606.600 22.650 ;
        RECT 605.400 16.050 606.450 20.400 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 608.400 16.050 609.450 19.950 ;
        RECT 592.950 13.950 595.050 16.050 ;
        RECT 598.950 13.950 604.050 16.050 ;
        RECT 604.950 13.950 607.050 16.050 ;
        RECT 607.950 13.950 610.050 16.050 ;
        RECT 611.400 10.050 612.450 43.950 ;
        RECT 616.950 31.950 619.050 34.050 ;
        RECT 617.400 27.600 618.450 31.950 ;
        RECT 623.400 31.050 624.450 53.400 ;
        RECT 629.400 43.050 630.450 64.950 ;
        RECT 635.400 60.600 636.450 67.950 ;
        RECT 641.400 60.600 642.450 73.950 ;
        RECT 653.400 61.200 654.450 106.950 ;
        RECT 656.400 106.050 657.450 109.950 ;
        RECT 655.950 103.950 658.050 106.050 ;
        RECT 662.400 105.600 663.450 113.400 ;
        RECT 665.400 108.450 666.450 139.950 ;
        RECT 673.950 138.000 676.050 142.050 ;
        RECT 674.400 136.350 675.600 138.000 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 671.400 132.900 672.600 133.650 ;
        RECT 677.400 133.050 678.600 133.650 ;
        RECT 683.400 133.050 684.450 169.950 ;
        RECT 689.400 148.050 690.450 203.550 ;
        RECT 701.400 190.050 702.450 250.950 ;
        RECT 704.400 223.050 705.450 253.950 ;
        RECT 703.950 220.950 706.050 223.050 ;
        RECT 691.950 187.950 694.050 190.050 ;
        RECT 700.950 187.950 703.050 190.050 ;
        RECT 692.400 163.050 693.450 187.950 ;
        RECT 707.400 187.050 708.450 277.950 ;
        RECT 709.950 268.950 712.050 271.050 ;
        RECT 710.400 262.050 711.450 268.950 ;
        RECT 715.950 265.950 718.050 268.050 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 716.400 261.600 717.450 265.950 ;
        RECT 716.400 259.350 717.600 261.600 ;
        RECT 721.950 260.100 724.050 262.200 ;
        RECT 725.400 262.050 726.450 289.950 ;
        RECT 722.400 259.350 723.600 260.100 ;
        RECT 724.950 259.950 727.050 262.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 721.950 256.950 724.050 259.050 ;
        RECT 713.400 256.050 714.600 256.650 ;
        RECT 709.950 254.400 714.600 256.050 ;
        RECT 719.400 255.900 720.600 256.650 ;
        RECT 728.400 256.050 729.450 301.950 ;
        RECT 748.950 298.950 751.050 301.050 ;
        RECT 730.950 293.100 733.050 295.200 ;
        RECT 736.950 293.100 739.050 295.200 ;
        RECT 742.950 293.100 745.050 295.200 ;
        RECT 731.400 286.050 732.450 293.100 ;
        RECT 737.400 292.350 738.600 293.100 ;
        RECT 743.400 292.350 744.600 293.100 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 740.400 287.400 741.600 289.650 ;
        RECT 730.950 283.950 733.050 286.050 ;
        RECT 731.400 271.050 732.450 283.950 ;
        RECT 740.400 283.050 741.450 287.400 ;
        RECT 749.400 283.050 750.450 298.950 ;
        RECT 758.400 297.450 759.450 424.950 ;
        RECT 761.400 412.050 762.450 424.950 ;
        RECT 764.400 424.050 765.450 481.800 ;
        RECT 767.400 472.050 768.450 484.950 ;
        RECT 770.400 478.050 771.450 488.400 ;
        RECT 772.950 487.950 775.050 490.050 ;
        RECT 769.950 475.950 772.050 478.050 ;
        RECT 766.950 469.950 769.050 472.050 ;
        RECT 769.950 460.950 772.050 463.050 ;
        RECT 770.400 450.600 771.450 460.950 ;
        RECT 773.400 454.050 774.450 487.950 ;
        RECT 776.400 484.050 777.450 494.100 ;
        RECT 785.400 493.350 786.600 494.100 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 782.400 488.400 783.600 490.650 ;
        RECT 788.400 489.900 789.600 490.650 ;
        RECT 775.950 481.950 778.050 484.050 ;
        RECT 782.400 481.050 783.450 488.400 ;
        RECT 787.950 487.800 790.050 489.900 ;
        RECT 790.950 487.950 793.050 490.050 ;
        RECT 781.950 478.950 784.050 481.050 ;
        RECT 782.400 475.050 783.450 478.950 ;
        RECT 781.950 472.950 784.050 475.050 ;
        RECT 778.950 460.950 781.050 463.050 ;
        RECT 775.950 454.950 778.050 457.050 ;
        RECT 772.950 451.950 775.050 454.050 ;
        RECT 776.400 450.600 777.450 454.950 ;
        RECT 779.400 451.050 780.450 460.950 ;
        RECT 791.400 460.050 792.450 487.950 ;
        RECT 790.950 457.950 793.050 460.050 ;
        RECT 794.400 457.050 795.450 496.950 ;
        RECT 797.400 489.900 798.450 505.950 ;
        RECT 800.400 496.050 801.450 521.400 ;
        RECT 805.950 520.950 808.050 523.050 ;
        RECT 809.400 521.400 810.600 523.650 ;
        RECT 815.400 522.900 816.600 523.650 ;
        RECT 806.400 505.050 807.450 520.950 ;
        RECT 809.400 517.050 810.450 521.400 ;
        RECT 814.950 520.800 817.050 522.900 ;
        RECT 808.950 514.950 811.050 517.050 ;
        RECT 815.400 514.050 816.450 520.800 ;
        RECT 814.950 511.950 817.050 514.050 ;
        RECT 824.400 510.450 825.450 538.950 ;
        RECT 827.400 529.050 828.450 550.950 ;
        RECT 829.950 547.950 832.050 550.050 ;
        RECT 826.950 526.950 829.050 529.050 ;
        RECT 830.400 528.600 831.450 547.950 ;
        RECT 833.400 547.050 834.450 572.100 ;
        RECT 839.400 571.350 840.600 572.100 ;
        RECT 845.400 571.350 846.600 573.600 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 835.950 565.950 838.050 568.050 ;
        RECT 842.400 566.400 843.600 568.650 ;
        RECT 848.400 566.400 849.600 568.650 ;
        RECT 832.950 544.950 835.050 547.050 ;
        RECT 836.400 544.050 837.450 565.950 ;
        RECT 835.950 541.950 838.050 544.050 ;
        RECT 830.400 526.350 831.600 528.600 ;
        RECT 835.950 527.100 838.050 529.200 ;
        RECT 842.400 529.050 843.450 566.400 ;
        RECT 844.950 559.950 847.050 562.050 ;
        RECT 845.400 556.050 846.450 559.950 ;
        RECT 848.400 556.050 849.450 566.400 ;
        RECT 844.800 553.950 846.900 556.050 ;
        RECT 847.950 553.950 850.050 556.050 ;
        RECT 850.950 544.950 853.050 547.050 ;
        RECT 847.950 532.950 850.050 535.050 ;
        RECT 836.400 526.350 837.600 527.100 ;
        RECT 841.950 526.950 844.050 529.050 ;
        RECT 844.950 527.100 847.050 529.200 ;
        RECT 829.950 523.950 832.050 526.050 ;
        RECT 832.950 523.950 835.050 526.050 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 826.950 517.950 829.050 523.050 ;
        RECT 833.400 522.000 834.600 523.650 ;
        RECT 839.400 523.050 840.600 523.650 ;
        RECT 832.950 517.950 835.050 522.000 ;
        RECT 839.400 521.400 844.050 523.050 ;
        RECT 840.000 520.950 844.050 521.400 ;
        RECT 845.400 514.050 846.450 527.100 ;
        RECT 844.950 511.950 847.050 514.050 ;
        RECT 824.400 509.400 828.450 510.450 ;
        RECT 823.950 505.950 826.050 508.050 ;
        RECT 805.950 502.950 808.050 505.050 ;
        RECT 811.950 499.950 814.050 502.050 ;
        RECT 805.500 497.400 807.600 499.500 ;
        RECT 812.400 499.200 813.600 499.950 ;
        RECT 799.950 493.950 802.050 496.050 ;
        RECT 799.950 490.800 802.050 492.900 ;
        RECT 803.100 490.950 805.200 493.050 ;
        RECT 796.950 487.800 799.050 489.900 ;
        RECT 781.950 454.950 784.050 457.050 ;
        RECT 793.950 454.950 796.050 457.050 ;
        RECT 770.400 448.350 771.600 450.600 ;
        RECT 776.400 448.350 777.600 450.600 ;
        RECT 778.950 448.950 781.050 451.050 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 773.400 444.900 774.600 445.650 ;
        RECT 772.950 442.800 775.050 444.900 ;
        RECT 775.950 427.950 778.050 430.050 ;
        RECT 763.950 421.950 766.050 424.050 ;
        RECT 769.950 417.000 772.050 421.050 ;
        RECT 776.400 417.600 777.450 427.950 ;
        RECT 770.400 415.350 771.600 417.000 ;
        RECT 776.400 415.350 777.600 417.600 ;
        RECT 766.950 412.950 769.050 415.050 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 760.950 409.950 763.050 412.050 ;
        RECT 767.400 411.900 768.600 412.650 ;
        RECT 766.950 409.800 769.050 411.900 ;
        RECT 773.400 411.000 774.600 412.650 ;
        RECT 767.400 397.050 768.450 409.800 ;
        RECT 772.950 406.950 775.050 411.000 ;
        RECT 778.950 409.950 781.050 412.050 ;
        RECT 769.950 405.450 772.050 406.050 ;
        RECT 775.950 405.450 778.050 406.050 ;
        RECT 769.950 404.400 778.050 405.450 ;
        RECT 769.950 403.950 772.050 404.400 ;
        RECT 775.950 403.950 778.050 404.400 ;
        RECT 779.400 400.050 780.450 409.950 ;
        RECT 778.950 397.950 781.050 400.050 ;
        RECT 766.950 394.950 769.050 397.050 ;
        RECT 778.950 391.950 781.050 394.050 ;
        RECT 772.950 385.950 775.050 388.050 ;
        RECT 760.950 371.100 763.050 373.200 ;
        RECT 766.950 371.100 769.050 373.200 ;
        RECT 773.400 372.600 774.450 385.950 ;
        RECT 779.400 373.050 780.450 391.950 ;
        RECT 761.400 364.050 762.450 371.100 ;
        RECT 767.400 370.350 768.600 371.100 ;
        RECT 773.400 370.350 774.600 372.600 ;
        RECT 778.950 370.950 781.050 373.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 769.950 367.950 772.050 370.050 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 770.400 365.400 771.600 367.650 ;
        RECT 776.400 366.900 777.600 367.650 ;
        RECT 760.950 361.950 763.050 364.050 ;
        RECT 766.950 352.950 769.050 355.050 ;
        RECT 767.400 339.600 768.450 352.950 ;
        RECT 770.400 352.050 771.450 365.400 ;
        RECT 775.950 364.800 778.050 366.900 ;
        RECT 772.950 361.950 775.050 364.050 ;
        RECT 769.950 349.950 772.050 352.050 ;
        RECT 767.400 337.350 768.600 339.600 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 764.400 333.900 765.600 334.650 ;
        RECT 773.400 334.050 774.450 361.950 ;
        RECT 782.400 343.050 783.450 454.950 ;
        RECT 787.950 451.950 790.050 454.050 ;
        RECT 800.400 453.450 801.450 490.800 ;
        RECT 803.400 489.900 804.600 490.650 ;
        RECT 802.950 487.800 805.050 489.900 ;
        RECT 806.100 484.800 807.000 497.400 ;
        RECT 812.100 496.800 814.200 498.900 ;
        RECT 815.400 497.100 817.500 499.200 ;
        RECT 807.900 495.000 810.000 495.900 ;
        RECT 807.900 493.800 815.100 495.000 ;
        RECT 813.000 492.900 815.100 493.800 ;
        RECT 807.900 492.000 810.000 492.900 ;
        RECT 816.000 492.000 816.900 497.100 ;
        RECT 818.400 495.450 819.600 495.600 ;
        RECT 818.400 494.400 822.450 495.450 ;
        RECT 818.400 493.350 819.600 494.400 ;
        RECT 807.900 491.100 816.900 492.000 ;
        RECT 807.900 490.800 810.000 491.100 ;
        RECT 812.100 487.950 814.200 490.050 ;
        RECT 812.400 485.400 813.600 487.650 ;
        RECT 805.800 482.700 807.900 484.800 ;
        RECT 816.000 484.500 816.900 491.100 ;
        RECT 817.800 490.950 819.900 493.050 ;
        RECT 814.800 482.400 816.900 484.500 ;
        RECT 821.400 481.050 822.450 494.400 ;
        RECT 824.400 487.050 825.450 505.950 ;
        RECT 827.400 505.050 828.450 509.400 ;
        RECT 826.950 502.950 829.050 505.050 ;
        RECT 832.950 499.950 835.050 502.050 ;
        RECT 826.950 493.950 829.050 496.050 ;
        RECT 833.400 495.600 834.450 499.950 ;
        RECT 823.950 484.950 826.050 487.050 ;
        RECT 820.950 478.950 823.050 481.050 ;
        RECT 827.400 478.050 828.450 493.950 ;
        RECT 833.400 493.350 834.600 495.600 ;
        RECT 838.950 494.100 841.050 496.200 ;
        RECT 845.400 496.050 846.450 511.950 ;
        RECT 839.400 493.350 840.600 494.100 ;
        RECT 844.950 493.950 847.050 496.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 835.950 490.950 838.050 493.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 836.400 489.900 837.600 490.650 ;
        RECT 835.950 487.800 838.050 489.900 ;
        RECT 842.400 488.400 843.600 490.650 ;
        RECT 842.400 484.050 843.450 488.400 ;
        RECT 844.950 487.950 847.050 490.050 ;
        RECT 841.950 481.950 844.050 484.050 ;
        RECT 826.950 475.950 829.050 478.050 ;
        RECT 820.950 472.950 823.050 475.050 ;
        RECT 811.950 469.950 814.050 472.050 ;
        RECT 808.950 463.950 811.050 466.050 ;
        RECT 805.950 457.950 808.050 460.050 ;
        RECT 800.400 452.400 804.450 453.450 ;
        RECT 784.950 449.100 787.050 451.200 ;
        RECT 785.400 439.050 786.450 449.100 ;
        RECT 784.950 436.950 787.050 439.050 ;
        RECT 788.400 435.450 789.450 451.950 ;
        RECT 790.950 449.100 793.050 451.200 ;
        RECT 799.950 449.100 802.050 451.200 ;
        RECT 791.400 448.350 792.600 449.100 ;
        RECT 800.400 448.350 801.600 449.100 ;
        RECT 791.100 445.950 793.200 448.050 ;
        RECT 796.500 445.950 798.600 448.050 ;
        RECT 799.800 445.950 801.900 448.050 ;
        RECT 797.400 443.400 798.600 445.650 ;
        RECT 797.400 436.050 798.450 443.400 ;
        RECT 799.950 439.950 802.050 442.050 ;
        RECT 788.400 434.400 792.450 435.450 ;
        RECT 787.950 430.950 790.050 433.050 ;
        RECT 784.950 427.950 787.050 430.050 ;
        RECT 785.400 400.050 786.450 427.950 ;
        RECT 788.400 418.050 789.450 430.950 ;
        RECT 791.400 424.050 792.450 434.400 ;
        RECT 796.950 433.950 799.050 436.050 ;
        RECT 790.950 421.950 793.050 424.050 ;
        RECT 787.950 415.950 790.050 418.050 ;
        RECT 793.950 417.000 796.050 421.050 ;
        RECT 800.400 417.600 801.450 439.950 ;
        RECT 803.400 418.050 804.450 452.400 ;
        RECT 806.400 436.050 807.450 457.950 ;
        RECT 805.950 433.950 808.050 436.050 ;
        RECT 805.950 418.950 808.050 421.050 ;
        RECT 794.400 415.350 795.600 417.000 ;
        RECT 800.400 415.350 801.600 417.600 ;
        RECT 802.950 415.950 805.050 418.050 ;
        RECT 806.400 415.050 807.450 418.950 ;
        RECT 809.400 418.050 810.450 463.950 ;
        RECT 812.400 451.050 813.450 469.950 ;
        RECT 811.950 448.950 814.050 451.050 ;
        RECT 814.950 450.000 817.050 454.050 ;
        RECT 821.400 450.600 822.450 472.950 ;
        RECT 845.400 469.050 846.450 487.950 ;
        RECT 848.400 477.450 849.450 532.950 ;
        RECT 851.400 529.050 852.450 544.950 ;
        RECT 854.400 535.050 855.450 577.950 ;
        RECT 863.400 573.600 864.450 592.800 ;
        RECT 872.400 586.050 873.450 605.100 ;
        RECT 871.950 583.950 874.050 586.050 ;
        RECT 875.400 574.200 876.450 616.950 ;
        RECT 877.950 607.950 880.050 610.050 ;
        RECT 878.400 585.450 879.450 607.950 ;
        RECT 881.400 606.600 882.450 643.950 ;
        RECT 884.400 640.050 885.450 661.950 ;
        RECT 890.400 655.050 891.450 676.950 ;
        RECT 893.400 658.050 894.450 712.950 ;
        RECT 896.400 706.050 897.450 730.950 ;
        RECT 895.950 703.950 898.050 706.050 ;
        RECT 895.950 694.950 898.050 697.050 ;
        RECT 896.400 691.050 897.450 694.950 ;
        RECT 899.400 691.050 900.450 736.950 ;
        RECT 902.400 730.050 903.450 766.950 ;
        RECT 904.950 760.950 907.050 763.050 ;
        RECT 914.400 762.600 915.450 772.950 ;
        RECT 917.400 766.050 918.450 775.950 ;
        RECT 923.400 766.050 924.450 808.950 ;
        RECT 916.950 763.950 919.050 766.050 ;
        RECT 922.950 763.950 925.050 766.050 ;
        RECT 905.400 751.050 906.450 760.950 ;
        RECT 914.400 760.350 915.600 762.600 ;
        RECT 919.950 761.100 922.050 763.200 ;
        RECT 925.950 761.100 928.050 763.200 ;
        RECT 920.400 760.350 921.600 761.100 ;
        RECT 910.950 757.950 913.050 760.050 ;
        RECT 913.950 757.950 916.050 760.050 ;
        RECT 916.950 757.950 919.050 760.050 ;
        RECT 919.950 757.950 922.050 760.050 ;
        RECT 911.400 756.900 912.600 757.650 ;
        RECT 910.950 754.800 913.050 756.900 ;
        RECT 917.400 755.400 918.600 757.650 ;
        RECT 917.400 751.050 918.450 755.400 ;
        RECT 922.950 754.950 925.050 757.050 ;
        RECT 904.950 748.950 907.050 751.050 ;
        RECT 916.950 748.950 919.050 751.050 ;
        RECT 905.400 736.050 906.450 748.950 ;
        RECT 913.950 742.950 916.050 745.050 ;
        RECT 904.950 733.950 907.050 736.050 ;
        RECT 901.950 727.950 904.050 730.050 ;
        RECT 907.950 728.100 910.050 730.200 ;
        RECT 914.400 729.600 915.450 742.950 ;
        RECT 908.400 727.350 909.600 728.100 ;
        RECT 914.400 727.350 915.600 729.600 ;
        RECT 919.950 728.100 922.050 730.200 ;
        RECT 904.950 724.950 907.050 727.050 ;
        RECT 907.950 724.950 910.050 727.050 ;
        RECT 910.950 724.950 913.050 727.050 ;
        RECT 913.950 724.950 916.050 727.050 ;
        RECT 905.400 722.400 906.600 724.650 ;
        RECT 911.400 723.000 912.600 724.650 ;
        RECT 901.950 718.950 904.050 721.050 ;
        RECT 902.400 715.050 903.450 718.950 ;
        RECT 901.950 712.950 904.050 715.050 ;
        RECT 901.950 703.950 904.050 706.050 ;
        RECT 895.950 688.950 898.050 691.050 ;
        RECT 898.950 688.950 901.050 691.050 ;
        RECT 896.400 685.050 897.450 688.950 ;
        RECT 895.950 682.950 898.050 685.050 ;
        RECT 899.400 684.600 900.450 688.950 ;
        RECT 902.400 687.450 903.450 703.950 ;
        RECT 905.400 697.050 906.450 722.400 ;
        RECT 910.950 718.950 913.050 723.000 ;
        RECT 916.950 718.950 919.050 721.050 ;
        RECT 904.950 694.950 907.050 697.050 ;
        RECT 902.400 686.400 906.450 687.450 ;
        RECT 905.400 684.600 906.450 686.400 ;
        RECT 899.400 682.350 900.600 684.600 ;
        RECT 905.400 682.350 906.600 684.600 ;
        RECT 913.950 683.100 916.050 685.200 ;
        RECT 898.950 679.950 901.050 682.050 ;
        RECT 901.950 679.950 904.050 682.050 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 895.950 675.450 898.050 679.050 ;
        RECT 902.400 678.000 903.600 679.650 ;
        RECT 908.400 678.900 909.600 679.650 ;
        RECT 895.950 675.000 900.450 675.450 ;
        RECT 896.400 674.400 900.450 675.000 ;
        RECT 892.950 655.950 895.050 658.050 ;
        RECT 890.400 653.550 895.050 655.050 ;
        RECT 891.000 652.950 895.050 653.550 ;
        RECT 892.950 649.950 895.050 652.050 ;
        RECT 893.400 649.350 894.600 649.950 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 890.400 644.400 891.600 646.650 ;
        RECT 883.950 637.950 886.050 640.050 ;
        RECT 890.400 634.050 891.450 644.400 ;
        RECT 895.950 643.950 898.050 646.050 ;
        RECT 892.950 637.950 895.050 643.050 ;
        RECT 889.950 631.950 892.050 634.050 ;
        RECT 896.400 628.050 897.450 643.950 ;
        RECT 899.400 634.050 900.450 674.400 ;
        RECT 901.950 673.950 904.050 678.000 ;
        RECT 907.950 676.800 910.050 678.900 ;
        RECT 914.400 670.050 915.450 683.100 ;
        RECT 910.800 667.950 912.900 670.050 ;
        RECT 913.950 667.950 916.050 670.050 ;
        RECT 901.950 655.950 904.050 658.050 ;
        RECT 898.950 631.950 901.050 634.050 ;
        RECT 895.950 625.950 898.050 628.050 ;
        RECT 898.950 622.950 901.050 625.050 ;
        RECT 892.950 619.950 895.050 622.050 ;
        RECT 881.400 604.350 882.600 606.600 ;
        RECT 889.950 605.100 892.050 607.200 ;
        RECT 890.400 604.350 891.600 605.100 ;
        RECT 881.100 601.950 883.200 604.050 ;
        RECT 884.400 601.950 886.500 604.050 ;
        RECT 889.800 601.950 891.900 604.050 ;
        RECT 884.400 599.400 885.600 601.650 ;
        RECT 878.400 584.400 882.450 585.450 ;
        RECT 877.950 580.950 880.050 583.050 ;
        RECT 863.400 571.350 864.600 573.600 ;
        RECT 868.950 572.100 871.050 574.200 ;
        RECT 869.400 571.350 870.600 572.100 ;
        RECT 874.950 571.950 877.050 574.200 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 871.950 568.950 874.050 571.050 ;
        RECT 866.400 566.400 867.600 568.650 ;
        RECT 872.400 567.900 873.600 568.650 ;
        RECT 856.950 553.950 859.050 556.050 ;
        RECT 853.950 532.950 856.050 535.050 ;
        RECT 850.950 526.950 853.050 529.050 ;
        RECT 857.400 528.600 858.450 553.950 ;
        RECT 866.400 552.450 867.450 566.400 ;
        RECT 871.950 565.800 874.050 567.900 ;
        RECT 874.950 565.950 877.050 568.050 ;
        RECT 866.400 551.400 870.450 552.450 ;
        RECT 865.950 538.950 868.050 541.050 ;
        RECT 857.400 526.350 858.600 528.600 ;
        RECT 862.950 527.100 865.050 529.200 ;
        RECT 866.400 529.050 867.450 538.950 ;
        RECT 863.400 526.350 864.600 527.100 ;
        RECT 865.950 526.950 868.050 529.050 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 850.950 520.950 853.050 523.050 ;
        RECT 854.400 521.400 855.600 523.650 ;
        RECT 860.400 521.400 861.600 523.650 ;
        RECT 851.400 502.050 852.450 520.950 ;
        RECT 854.400 511.050 855.450 521.400 ;
        RECT 860.400 517.050 861.450 521.400 ;
        RECT 865.950 520.950 868.050 523.050 ;
        RECT 862.950 517.950 865.050 520.050 ;
        RECT 859.950 514.950 862.050 517.050 ;
        RECT 853.950 508.950 856.050 511.050 ;
        RECT 860.400 508.050 861.450 514.950 ;
        RECT 859.950 505.950 862.050 508.050 ;
        RECT 850.800 499.950 852.900 502.050 ;
        RECT 853.950 498.450 856.050 502.050 ;
        RECT 851.400 498.000 856.050 498.450 ;
        RECT 850.950 497.400 855.450 498.000 ;
        RECT 850.950 493.950 853.050 497.400 ;
        RECT 856.950 494.100 859.050 496.200 ;
        RECT 863.400 495.600 864.450 517.950 ;
        RECT 866.400 502.050 867.450 520.950 ;
        RECT 869.400 517.050 870.450 551.400 ;
        RECT 872.400 550.050 873.450 565.800 ;
        RECT 871.950 547.950 874.050 550.050 ;
        RECT 872.400 532.050 873.450 547.950 ;
        RECT 875.400 532.050 876.450 565.950 ;
        RECT 878.400 562.050 879.450 580.950 ;
        RECT 881.400 574.050 882.450 584.400 ;
        RECT 884.400 583.050 885.450 599.400 ;
        RECT 883.950 580.950 886.050 583.050 ;
        RECT 880.950 571.950 883.050 574.050 ;
        RECT 883.950 573.000 886.050 577.050 ;
        RECT 884.400 571.350 885.600 573.000 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 880.950 565.950 883.050 568.050 ;
        RECT 887.400 566.400 888.600 568.650 ;
        RECT 877.950 559.950 880.050 562.050 ;
        RECT 877.950 544.950 880.050 547.050 ;
        RECT 871.800 529.950 873.900 532.050 ;
        RECT 874.950 529.950 877.050 532.050 ;
        RECT 878.400 528.600 879.450 544.950 ;
        RECT 881.400 532.050 882.450 565.950 ;
        RECT 887.400 556.050 888.450 566.400 ;
        RECT 886.950 555.450 889.050 556.050 ;
        RECT 886.950 554.400 891.450 555.450 ;
        RECT 886.950 553.950 889.050 554.400 ;
        RECT 883.950 547.950 886.050 550.050 ;
        RECT 884.400 541.050 885.450 547.950 ;
        RECT 883.950 538.950 886.050 541.050 ;
        RECT 880.950 529.950 883.050 532.050 ;
        RECT 878.400 526.350 879.600 528.600 ;
        RECT 883.950 527.100 886.050 532.050 ;
        RECT 884.400 526.350 885.600 527.100 ;
        RECT 874.950 523.950 877.050 526.050 ;
        RECT 877.950 523.950 880.050 526.050 ;
        RECT 880.950 523.950 883.050 526.050 ;
        RECT 883.950 523.950 886.050 526.050 ;
        RECT 875.400 521.400 876.600 523.650 ;
        RECT 881.400 522.900 882.600 523.650 ;
        RECT 890.400 522.900 891.450 554.400 ;
        RECT 893.400 550.050 894.450 619.950 ;
        RECT 899.400 607.050 900.450 622.950 ;
        RECT 902.400 610.050 903.450 655.950 ;
        RECT 911.400 655.050 912.450 667.950 ;
        RECT 913.950 655.950 916.050 658.050 ;
        RECT 910.950 652.950 913.050 655.050 ;
        RECT 907.950 650.100 910.050 652.200 ;
        RECT 914.400 651.600 915.450 655.950 ;
        RECT 917.400 655.050 918.450 718.950 ;
        RECT 920.400 709.050 921.450 728.100 ;
        RECT 923.400 715.050 924.450 754.950 ;
        RECT 926.400 745.050 927.450 761.100 ;
        RECT 925.950 742.950 928.050 745.050 ;
        RECT 922.950 712.950 925.050 715.050 ;
        RECT 919.950 706.950 922.050 709.050 ;
        RECT 929.400 703.050 930.450 808.950 ;
        RECT 928.950 700.950 931.050 703.050 ;
        RECT 932.400 691.050 933.450 841.950 ;
        RECT 934.950 763.950 937.050 766.050 ;
        RECT 935.400 700.050 936.450 763.950 ;
        RECT 934.950 697.950 937.050 700.050 ;
        RECT 919.950 688.950 922.050 691.050 ;
        RECT 931.950 688.950 934.050 691.050 ;
        RECT 920.400 685.050 921.450 688.950 ;
        RECT 919.950 682.950 922.050 685.050 ;
        RECT 925.950 683.100 928.050 685.200 ;
        RECT 931.950 683.100 934.050 685.200 ;
        RECT 926.400 682.350 927.600 683.100 ;
        RECT 932.400 682.350 933.600 683.100 ;
        RECT 922.950 679.950 925.050 682.050 ;
        RECT 925.950 679.950 928.050 682.050 ;
        RECT 928.950 679.950 931.050 682.050 ;
        RECT 931.950 679.950 934.050 682.050 ;
        RECT 919.950 676.950 922.050 679.050 ;
        RECT 923.400 677.400 924.600 679.650 ;
        RECT 929.400 678.900 930.600 679.650 ;
        RECT 916.950 652.950 919.050 655.050 ;
        RECT 920.400 652.050 921.450 676.950 ;
        RECT 923.400 661.050 924.450 677.400 ;
        RECT 928.950 676.800 931.050 678.900 ;
        RECT 934.950 676.950 937.050 679.050 ;
        RECT 925.950 670.950 928.050 673.050 ;
        RECT 922.950 658.950 925.050 661.050 ;
        RECT 922.950 655.800 925.050 657.900 ;
        RECT 908.400 649.350 909.600 650.100 ;
        RECT 914.400 649.350 915.600 651.600 ;
        RECT 919.950 649.950 922.050 652.050 ;
        RECT 907.950 646.950 910.050 649.050 ;
        RECT 910.950 646.950 913.050 649.050 ;
        RECT 913.950 646.950 916.050 649.050 ;
        RECT 916.950 646.950 919.050 649.050 ;
        RECT 904.950 643.950 907.050 646.050 ;
        RECT 911.400 645.000 912.600 646.650 ;
        RECT 917.400 645.900 918.600 646.650 ;
        RECT 901.950 607.950 904.050 610.050 ;
        RECT 895.800 604.950 897.900 607.050 ;
        RECT 898.950 604.950 901.050 607.050 ;
        RECT 905.400 606.600 906.450 643.950 ;
        RECT 910.950 640.950 913.050 645.000 ;
        RECT 916.950 643.800 919.050 645.900 ;
        RECT 919.950 643.950 922.050 646.050 ;
        RECT 913.950 634.950 916.050 637.050 ;
        RECT 896.400 592.050 897.450 604.950 ;
        RECT 905.400 604.350 906.600 606.600 ;
        RECT 910.950 606.000 913.050 610.050 ;
        RECT 914.400 606.450 915.450 634.950 ;
        RECT 917.400 622.050 918.450 643.800 ;
        RECT 920.400 637.050 921.450 643.950 ;
        RECT 919.950 634.950 922.050 637.050 ;
        RECT 919.950 625.950 922.050 628.050 ;
        RECT 916.950 619.950 919.050 622.050 ;
        RECT 916.950 610.950 919.050 616.050 ;
        RECT 911.400 604.350 912.600 606.000 ;
        RECT 914.400 605.400 918.450 606.450 ;
        RECT 901.950 601.950 904.050 604.050 ;
        RECT 904.950 601.950 907.050 604.050 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 898.950 598.950 901.050 601.050 ;
        RECT 902.400 599.400 903.600 601.650 ;
        RECT 908.400 599.400 909.600 601.650 ;
        RECT 895.950 589.950 898.050 592.050 ;
        RECT 899.400 589.050 900.450 598.950 ;
        RECT 898.950 586.950 901.050 589.050 ;
        RECT 902.400 577.050 903.450 599.400 ;
        RECT 908.400 577.200 909.450 599.400 ;
        RECT 913.950 598.950 916.050 601.050 ;
        RECT 910.950 595.950 913.050 598.050 ;
        RECT 911.400 586.050 912.450 595.950 ;
        RECT 910.950 583.950 913.050 586.050 ;
        RECT 901.950 574.950 904.050 577.050 ;
        RECT 907.950 575.100 910.050 577.200 ;
        RECT 914.400 574.050 915.450 598.950 ;
        RECT 902.400 573.450 903.600 573.600 ;
        RECT 896.400 572.400 903.600 573.450 ;
        RECT 892.950 547.950 895.050 550.050 ;
        RECT 896.400 547.050 897.450 572.400 ;
        RECT 902.400 571.350 903.600 572.400 ;
        RECT 907.950 571.950 910.050 574.050 ;
        RECT 913.950 571.950 916.050 574.050 ;
        RECT 908.400 571.350 909.600 571.950 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 907.950 568.950 910.050 571.050 ;
        RECT 910.950 568.950 913.050 571.050 ;
        RECT 898.950 565.950 901.050 568.050 ;
        RECT 905.400 567.000 906.600 568.650 ;
        RECT 899.400 559.050 900.450 565.950 ;
        RECT 904.950 562.950 907.050 567.000 ;
        RECT 911.400 566.400 912.600 568.650 ;
        RECT 898.950 556.950 901.050 559.050 ;
        RECT 911.400 553.050 912.450 566.400 ;
        RECT 913.950 565.950 916.050 568.050 ;
        RECT 910.950 550.950 913.050 553.050 ;
        RECT 895.950 544.950 898.050 547.050 ;
        RECT 898.950 532.950 901.050 535.050 ;
        RECT 899.400 528.600 900.450 532.950 ;
        RECT 911.400 532.050 912.450 550.950 ;
        RECT 910.950 529.950 913.050 532.050 ;
        RECT 899.400 526.350 900.600 528.600 ;
        RECT 904.950 527.100 907.050 529.200 ;
        RECT 905.400 526.350 906.600 527.100 ;
        RECT 910.950 526.800 913.050 528.900 ;
        RECT 895.950 523.950 898.050 526.050 ;
        RECT 898.950 523.950 901.050 526.050 ;
        RECT 901.950 523.950 904.050 526.050 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 868.950 514.950 871.050 517.050 ;
        RECT 865.950 499.950 868.050 502.050 ;
        RECT 868.950 501.450 871.050 505.050 ;
        RECT 868.950 501.000 873.450 501.450 ;
        RECT 869.400 500.400 873.450 501.000 ;
        RECT 857.400 493.350 858.600 494.100 ;
        RECT 863.400 493.350 864.600 495.600 ;
        RECT 868.950 493.950 871.050 496.050 ;
        RECT 853.950 490.950 856.050 493.050 ;
        RECT 856.950 490.950 859.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 854.400 488.400 855.600 490.650 ;
        RECT 860.400 489.900 861.600 490.650 ;
        RECT 848.400 476.400 852.450 477.450 ;
        RECT 847.950 472.950 850.050 475.050 ;
        RECT 844.950 466.950 847.050 469.050 ;
        RECT 832.950 463.950 835.050 466.050 ;
        RECT 833.400 450.600 834.450 463.950 ;
        RECT 815.400 448.350 816.600 450.000 ;
        RECT 821.400 448.350 822.600 450.600 ;
        RECT 833.400 448.350 834.600 450.600 ;
        RECT 838.950 449.100 841.050 451.200 ;
        RECT 839.400 448.350 840.600 449.100 ;
        RECT 814.950 445.950 817.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 838.950 445.950 841.050 448.050 ;
        RECT 841.950 445.950 844.050 448.050 ;
        RECT 818.400 443.400 819.600 445.650 ;
        RECT 836.400 444.900 837.600 445.650 ;
        RECT 818.400 442.050 819.450 443.400 ;
        RECT 826.950 442.800 829.050 444.900 ;
        RECT 835.950 442.800 838.050 444.900 ;
        RECT 842.400 443.400 843.600 445.650 ;
        RECT 817.950 439.950 820.050 442.050 ;
        RECT 818.400 421.050 819.450 439.950 ;
        RECT 823.950 436.950 826.050 439.050 ;
        RECT 820.950 427.950 823.050 430.050 ;
        RECT 821.400 421.050 822.450 427.950 ;
        RECT 808.950 415.950 811.050 418.050 ;
        RECT 811.950 417.000 814.050 421.050 ;
        RECT 817.950 418.950 820.050 421.050 ;
        RECT 820.950 418.950 823.050 421.050 ;
        RECT 812.400 415.350 813.600 417.000 ;
        RECT 820.950 415.800 823.050 417.900 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 796.950 412.950 799.050 415.050 ;
        RECT 799.950 412.950 802.050 415.050 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 791.400 411.900 792.600 412.650 ;
        RECT 790.950 409.800 793.050 411.900 ;
        RECT 797.400 410.400 798.600 412.650 ;
        RECT 797.400 406.050 798.450 410.400 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 815.400 411.900 816.600 412.650 ;
        RECT 796.950 403.950 799.050 406.050 ;
        RECT 784.950 397.950 787.050 400.050 ;
        RECT 793.950 376.950 796.050 379.050 ;
        RECT 787.950 371.100 790.050 373.200 ;
        RECT 794.400 372.600 795.450 376.950 ;
        RECT 788.400 370.350 789.600 371.100 ;
        RECT 794.400 370.350 795.600 372.600 ;
        RECT 787.950 367.950 790.050 370.050 ;
        RECT 790.950 367.950 793.050 370.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 784.950 364.950 787.050 367.050 ;
        RECT 791.400 366.000 792.600 367.650 ;
        RECT 785.400 352.050 786.450 364.950 ;
        RECT 790.950 361.950 793.050 366.000 ;
        RECT 797.400 365.400 798.600 367.650 ;
        RECT 787.950 355.950 790.050 358.050 ;
        RECT 784.950 349.950 787.050 352.050 ;
        RECT 788.400 349.050 789.450 355.950 ;
        RECT 797.400 355.050 798.450 365.400 ;
        RECT 796.950 352.950 799.050 355.050 ;
        RECT 787.950 346.950 790.050 349.050 ;
        RECT 775.950 340.950 778.050 343.050 ;
        RECT 781.950 340.950 784.050 343.050 ;
        RECT 788.400 342.450 789.450 346.950 ;
        RECT 803.400 343.050 804.450 409.950 ;
        RECT 805.950 409.800 808.050 411.900 ;
        RECT 814.950 409.800 817.050 411.900 ;
        RECT 817.950 409.950 820.050 412.050 ;
        RECT 806.400 397.050 807.450 409.800 ;
        RECT 818.400 403.050 819.450 409.950 ;
        RECT 814.800 400.950 816.900 403.050 ;
        RECT 817.950 400.950 820.050 403.050 ;
        RECT 805.950 394.950 808.050 397.050 ;
        RECT 805.950 388.950 808.050 391.050 ;
        RECT 806.400 373.050 807.450 388.950 ;
        RECT 815.400 388.050 816.450 400.950 ;
        RECT 821.400 397.050 822.450 415.800 ;
        RECT 817.800 394.950 819.900 397.050 ;
        RECT 820.950 394.950 823.050 397.050 ;
        RECT 814.950 385.950 817.050 388.050 ;
        RECT 808.950 382.950 811.050 385.050 ;
        RECT 809.400 376.050 810.450 382.950 ;
        RECT 811.950 376.950 814.050 379.050 ;
        RECT 808.950 373.950 811.050 376.050 ;
        RECT 805.950 370.950 808.050 373.050 ;
        RECT 812.400 372.600 813.450 376.950 ;
        RECT 818.400 376.200 819.450 394.950 ;
        RECT 817.950 374.100 820.050 376.200 ;
        RECT 812.400 370.350 813.600 372.600 ;
        RECT 817.950 370.950 820.050 373.050 ;
        RECT 818.400 370.350 819.600 370.950 ;
        RECT 808.950 367.950 811.050 370.050 ;
        RECT 811.950 367.950 814.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 805.950 361.950 808.050 367.050 ;
        RECT 809.400 365.400 810.600 367.650 ;
        RECT 815.400 366.900 816.600 367.650 ;
        RECT 809.400 355.050 810.450 365.400 ;
        RECT 814.950 364.800 817.050 366.900 ;
        RECT 820.950 364.950 823.050 367.050 ;
        RECT 808.950 352.950 811.050 355.050 ;
        RECT 814.950 352.950 817.050 355.050 ;
        RECT 785.400 341.400 789.450 342.450 ;
        RECT 763.950 331.800 766.050 333.900 ;
        RECT 772.950 331.950 775.050 334.050 ;
        RECT 776.400 313.050 777.450 340.950 ;
        RECT 785.400 339.600 786.450 341.400 ;
        RECT 796.950 340.950 799.050 343.050 ;
        RECT 802.950 340.950 805.050 343.050 ;
        RECT 785.400 337.350 786.600 339.600 ;
        RECT 790.950 338.100 793.050 340.200 ;
        RECT 791.400 337.350 792.600 338.100 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 782.400 333.900 783.600 334.650 ;
        RECT 781.950 331.800 784.050 333.900 ;
        RECT 788.400 332.400 789.600 334.650 ;
        RECT 788.400 328.050 789.450 332.400 ;
        RECT 787.950 325.950 790.050 328.050 ;
        RECT 775.950 310.950 778.050 313.050 ;
        RECT 769.950 301.950 772.050 304.050 ;
        RECT 755.400 296.400 759.450 297.450 ;
        RECT 755.400 294.600 756.450 296.400 ;
        RECT 755.400 292.350 756.600 294.600 ;
        RECT 760.950 293.100 763.050 295.200 ;
        RECT 761.400 292.350 762.600 293.100 ;
        RECT 754.950 289.950 757.050 292.050 ;
        RECT 757.950 289.950 760.050 292.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 758.400 288.900 759.600 289.650 ;
        RECT 757.950 286.800 760.050 288.900 ;
        RECT 764.400 287.400 765.600 289.650 ;
        RECT 739.950 280.950 742.050 283.050 ;
        RECT 748.950 280.950 751.050 283.050 ;
        RECT 758.400 280.050 759.450 286.800 ;
        RECT 757.950 277.950 760.050 280.050 ;
        RECT 764.400 274.050 765.450 287.400 ;
        RECT 766.950 283.950 769.050 289.050 ;
        RECT 763.950 271.950 766.050 274.050 ;
        RECT 730.950 268.950 733.050 271.050 ;
        RECT 748.950 265.950 751.050 268.050 ;
        RECT 754.950 265.950 757.050 268.050 ;
        RECT 733.950 260.100 736.050 262.200 ;
        RECT 739.950 260.100 742.050 262.200 ;
        RECT 734.400 259.350 735.600 260.100 ;
        RECT 740.400 259.350 741.600 260.100 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 736.950 256.950 739.050 259.050 ;
        RECT 739.950 256.950 742.050 259.050 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 709.950 253.950 714.000 254.400 ;
        RECT 718.950 253.800 721.050 255.900 ;
        RECT 727.950 253.950 730.050 256.050 ;
        RECT 737.400 255.000 738.600 256.650 ;
        RECT 743.400 255.900 744.600 256.650 ;
        RECT 727.950 250.800 730.050 252.900 ;
        RECT 736.950 250.950 739.050 255.000 ;
        RECT 742.950 253.800 745.050 255.900 ;
        RECT 712.800 220.500 714.900 222.600 ;
        RECT 710.100 211.950 712.200 214.050 ;
        RECT 713.100 213.300 714.300 220.500 ;
        RECT 716.400 217.350 717.600 219.600 ;
        RECT 722.400 219.300 724.500 221.400 ;
        RECT 716.100 214.950 718.200 217.050 ;
        RECT 719.100 215.700 721.200 217.800 ;
        RECT 719.100 213.300 720.000 215.700 ;
        RECT 713.100 212.100 720.000 213.300 ;
        RECT 710.400 210.900 711.600 211.650 ;
        RECT 709.950 208.800 712.050 210.900 ;
        RECT 713.100 206.700 714.000 212.100 ;
        RECT 714.900 210.300 717.000 211.200 ;
        RECT 722.700 210.300 723.600 219.300 ;
        RECT 724.950 215.100 727.050 217.200 ;
        RECT 725.400 214.350 726.600 215.100 ;
        RECT 724.800 211.950 726.900 214.050 ;
        RECT 714.900 209.100 723.600 210.300 ;
        RECT 712.800 204.600 714.900 206.700 ;
        RECT 716.100 206.100 718.200 208.200 ;
        RECT 720.000 207.300 722.100 209.100 ;
        RECT 716.400 203.550 717.600 205.800 ;
        RECT 716.400 190.050 717.450 203.550 ;
        RECT 715.950 187.950 718.050 190.050 ;
        RECT 706.950 184.950 709.050 187.050 ;
        RECT 712.950 184.950 715.050 187.050 ;
        RECT 700.950 182.100 703.050 184.200 ;
        RECT 708.000 183.600 712.050 184.050 ;
        RECT 701.400 181.350 702.600 182.100 ;
        RECT 707.400 181.950 712.050 183.600 ;
        RECT 707.400 181.350 708.600 181.950 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 698.400 176.400 699.600 178.650 ;
        RECT 704.400 177.000 705.600 178.650 ;
        RECT 691.950 160.950 694.050 163.050 ;
        RECT 688.950 145.950 691.050 148.050 ;
        RECT 692.400 141.450 693.450 160.950 ;
        RECT 698.400 157.050 699.450 176.400 ;
        RECT 703.950 172.950 706.050 177.000 ;
        RECT 709.950 175.950 712.050 178.050 ;
        RECT 700.950 166.950 703.050 169.050 ;
        RECT 706.950 166.950 709.050 169.050 ;
        RECT 697.950 154.950 700.050 157.050 ;
        RECT 694.950 145.950 697.050 148.050 ;
        RECT 689.400 140.400 693.450 141.450 ;
        RECT 689.400 139.050 690.450 140.400 ;
        RECT 695.400 139.200 696.450 145.950 ;
        RECT 685.950 138.600 690.450 139.050 ;
        RECT 685.950 136.950 690.600 138.600 ;
        RECT 694.950 137.100 697.050 139.200 ;
        RECT 689.400 136.350 690.600 136.950 ;
        RECT 695.400 136.350 696.600 137.100 ;
        RECT 688.950 133.950 691.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 670.950 130.800 673.050 132.900 ;
        RECT 677.400 131.400 682.050 133.050 ;
        RECT 678.000 130.950 682.050 131.400 ;
        RECT 682.950 130.950 685.050 133.050 ;
        RECT 692.400 132.900 693.600 133.650 ;
        RECT 691.950 130.800 694.050 132.900 ;
        RECT 676.950 112.950 679.050 115.050 ;
        RECT 665.400 107.400 669.450 108.450 ;
        RECT 668.400 105.600 669.450 107.400 ;
        RECT 662.400 103.350 663.600 105.600 ;
        RECT 668.400 103.350 669.600 105.600 ;
        RECT 673.950 103.950 676.050 106.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 664.950 100.950 667.050 103.050 ;
        RECT 667.950 100.950 670.050 103.050 ;
        RECT 659.400 99.900 660.600 100.650 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 665.400 98.400 666.600 100.650 ;
        RECT 665.400 91.050 666.450 98.400 ;
        RECT 674.400 94.050 675.450 103.950 ;
        RECT 677.400 99.900 678.450 112.950 ;
        RECT 701.400 112.050 702.450 166.950 ;
        RECT 707.400 163.050 708.450 166.950 ;
        RECT 706.950 160.950 709.050 163.050 ;
        RECT 710.400 151.050 711.450 175.950 ;
        RECT 709.950 148.950 712.050 151.050 ;
        RECT 706.950 145.950 709.050 148.050 ;
        RECT 707.400 138.600 708.450 145.950 ;
        RECT 713.400 142.200 714.450 184.950 ;
        RECT 716.400 183.450 717.450 187.950 ;
        RECT 719.400 183.450 720.600 183.600 ;
        RECT 716.400 182.400 720.600 183.450 ;
        RECT 719.400 181.350 720.600 182.400 ;
        RECT 725.400 183.450 726.600 183.600 ;
        RECT 728.400 183.450 729.450 250.800 ;
        RECT 745.950 244.950 748.050 247.050 ;
        RECT 733.950 235.950 736.050 238.050 ;
        RECT 734.400 210.900 735.450 235.950 ;
        RECT 739.950 232.950 742.050 235.050 ;
        RECT 740.400 216.600 741.450 232.950 ;
        RECT 746.400 217.200 747.450 244.950 ;
        RECT 749.400 232.050 750.450 265.950 ;
        RECT 755.400 261.450 756.450 265.950 ;
        RECT 752.400 260.400 756.450 261.450 ;
        RECT 752.400 255.900 753.450 260.400 ;
        RECT 757.950 260.100 760.050 262.200 ;
        RECT 763.950 260.100 766.050 262.200 ;
        RECT 770.400 262.050 771.450 301.950 ;
        RECT 797.400 301.050 798.450 340.950 ;
        RECT 805.950 338.100 808.050 340.200 ;
        RECT 806.400 337.350 807.600 338.100 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 803.400 332.400 804.600 334.650 ;
        RECT 809.400 332.400 810.600 334.650 ;
        RECT 803.400 322.050 804.450 332.400 ;
        RECT 809.400 331.050 810.450 332.400 ;
        RECT 808.950 328.950 811.050 331.050 ;
        RECT 802.950 319.950 805.050 322.050 ;
        RECT 809.400 319.050 810.450 328.950 ;
        RECT 808.950 316.950 811.050 319.050 ;
        RECT 784.950 298.950 787.050 301.050 ;
        RECT 796.950 298.950 799.050 301.050 ;
        RECT 772.950 294.600 777.000 295.050 ;
        RECT 772.950 292.950 777.600 294.600 ;
        RECT 776.400 292.350 777.600 292.950 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 779.400 288.900 780.600 289.650 ;
        RECT 778.950 286.800 781.050 288.900 ;
        RECT 775.950 277.950 778.050 280.050 ;
        RECT 772.950 271.950 775.050 274.050 ;
        RECT 758.400 259.350 759.600 260.100 ;
        RECT 764.400 259.350 765.600 260.100 ;
        RECT 769.950 259.950 772.050 262.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 751.950 253.800 754.050 255.900 ;
        RECT 761.400 255.000 762.600 256.650 ;
        RECT 760.950 250.950 763.050 255.000 ;
        RECT 767.400 254.400 768.600 256.650 ;
        RECT 748.950 229.950 751.050 232.050 ;
        RECT 767.400 226.050 768.450 254.400 ;
        RECT 769.950 250.950 772.050 256.050 ;
        RECT 766.950 223.950 769.050 226.050 ;
        RECT 740.400 214.350 741.600 216.600 ;
        RECT 745.950 215.100 748.050 217.200 ;
        RECT 760.950 215.100 763.050 217.200 ;
        RECT 766.950 215.100 769.050 217.200 ;
        RECT 746.400 214.350 747.600 215.100 ;
        RECT 761.400 214.350 762.600 215.100 ;
        RECT 767.400 214.350 768.600 215.100 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 742.950 211.950 745.050 214.050 ;
        RECT 745.950 211.950 748.050 214.050 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 743.400 210.900 744.600 211.650 ;
        RECT 733.950 208.800 736.050 210.900 ;
        RECT 742.950 208.800 745.050 210.900 ;
        RECT 749.400 209.400 750.600 211.650 ;
        RECT 764.400 210.000 765.600 211.650 ;
        RECT 749.400 205.050 750.450 209.400 ;
        RECT 763.950 205.950 766.050 210.000 ;
        RECT 769.950 205.950 772.050 208.050 ;
        RECT 748.950 202.950 751.050 205.050 ;
        RECT 760.950 204.450 763.050 205.050 ;
        RECT 766.950 204.450 769.050 205.050 ;
        RECT 760.950 203.400 769.050 204.450 ;
        RECT 760.950 202.950 763.050 203.400 ;
        RECT 766.950 202.950 769.050 203.400 ;
        RECT 770.400 202.050 771.450 205.950 ;
        RECT 769.950 199.950 772.050 202.050 ;
        RECT 773.400 199.050 774.450 271.950 ;
        RECT 776.400 271.050 777.450 277.950 ;
        RECT 779.400 277.050 780.450 286.800 ;
        RECT 778.950 274.950 781.050 277.050 ;
        RECT 775.950 268.950 778.050 271.050 ;
        RECT 785.400 265.050 786.450 298.950 ;
        RECT 796.950 294.000 799.050 297.900 ;
        RECT 797.400 292.350 798.600 294.000 ;
        RECT 802.950 293.100 805.050 295.200 ;
        RECT 815.400 294.450 816.450 352.950 ;
        RECT 821.400 349.050 822.450 364.950 ;
        RECT 820.950 346.950 823.050 349.050 ;
        RECT 824.400 343.050 825.450 436.950 ;
        RECT 827.400 418.050 828.450 442.800 ;
        RECT 838.950 433.950 841.050 436.050 ;
        RECT 839.400 418.200 840.450 433.950 ;
        RECT 842.400 430.050 843.450 443.400 ;
        RECT 841.950 427.950 844.050 430.050 ;
        RECT 841.950 421.950 844.050 424.050 ;
        RECT 826.950 415.950 829.050 418.050 ;
        RECT 832.950 416.100 835.050 418.200 ;
        RECT 838.950 416.100 841.050 418.200 ;
        RECT 842.400 418.050 843.450 421.950 ;
        RECT 833.400 415.350 834.600 416.100 ;
        RECT 839.400 415.350 840.600 416.100 ;
        RECT 841.950 415.950 844.050 418.050 ;
        RECT 848.400 417.450 849.450 472.950 ;
        RECT 851.400 451.050 852.450 476.400 ;
        RECT 854.400 463.050 855.450 488.400 ;
        RECT 859.950 487.800 862.050 489.900 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 857.400 466.050 858.450 484.950 ;
        RECT 860.400 481.050 861.450 487.800 ;
        RECT 859.950 478.950 862.050 481.050 ;
        RECT 869.400 475.050 870.450 493.950 ;
        RECT 872.400 480.450 873.450 500.400 ;
        RECT 875.400 496.050 876.450 521.400 ;
        RECT 880.950 520.800 883.050 522.900 ;
        RECT 889.950 520.800 892.050 522.900 ;
        RECT 892.950 520.950 895.050 523.050 ;
        RECT 896.400 521.400 897.600 523.650 ;
        RECT 902.400 521.400 903.600 523.650 ;
        RECT 886.950 502.950 889.050 505.050 ;
        RECT 874.950 493.950 877.050 496.050 ;
        RECT 880.950 494.100 883.050 496.200 ;
        RECT 887.400 495.600 888.450 502.950 ;
        RECT 881.400 493.350 882.600 494.100 ;
        RECT 887.400 493.350 888.600 495.600 ;
        RECT 877.950 490.950 880.050 493.050 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 878.400 488.400 879.600 490.650 ;
        RECT 884.400 488.400 885.600 490.650 ;
        RECT 872.400 479.400 876.450 480.450 ;
        RECT 871.950 475.950 874.050 478.050 ;
        RECT 868.950 472.950 871.050 475.050 ;
        RECT 856.950 463.950 859.050 466.050 ;
        RECT 865.950 463.950 868.050 466.050 ;
        RECT 853.950 460.950 856.050 463.050 ;
        RECT 854.400 457.050 855.450 460.950 ;
        RECT 859.950 457.950 862.050 460.050 ;
        RECT 853.950 454.950 856.050 457.050 ;
        RECT 850.950 448.950 853.050 451.050 ;
        RECT 853.950 450.000 856.050 453.900 ;
        RECT 860.400 450.600 861.450 457.950 ;
        RECT 866.400 451.050 867.450 463.950 ;
        RECT 868.950 457.950 871.050 460.050 ;
        RECT 869.400 454.050 870.450 457.950 ;
        RECT 868.950 451.950 871.050 454.050 ;
        RECT 854.400 448.350 855.600 450.000 ;
        RECT 860.400 448.350 861.600 450.600 ;
        RECT 865.950 448.950 868.050 451.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 850.950 442.950 853.050 445.050 ;
        RECT 857.400 443.400 858.600 445.650 ;
        RECT 863.400 444.900 864.600 445.650 ;
        RECT 851.400 424.050 852.450 442.950 ;
        RECT 857.400 439.050 858.450 443.400 ;
        RECT 862.950 442.800 865.050 444.900 ;
        RECT 856.950 436.950 859.050 439.050 ;
        RECT 857.400 433.050 858.450 436.950 ;
        RECT 856.950 430.950 859.050 433.050 ;
        RECT 869.400 430.050 870.450 451.950 ;
        RECT 856.950 427.800 859.050 429.900 ;
        RECT 868.950 427.950 871.050 430.050 ;
        RECT 850.950 421.950 853.050 424.050 ;
        RECT 845.400 416.400 849.450 417.450 ;
        RECT 829.950 412.950 832.050 415.050 ;
        RECT 832.950 412.950 835.050 415.050 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 826.950 409.950 829.050 412.050 ;
        RECT 830.400 411.900 831.600 412.650 ;
        RECT 827.400 384.450 828.450 409.950 ;
        RECT 829.950 409.800 832.050 411.900 ;
        RECT 836.400 410.400 837.600 412.650 ;
        RECT 836.400 409.050 837.450 410.400 ;
        RECT 835.950 403.950 838.050 409.050 ;
        RECT 841.950 406.950 844.050 409.050 ;
        RECT 835.950 400.800 838.050 402.900 ;
        RECT 829.950 384.450 832.050 385.050 ;
        RECT 827.400 383.400 832.050 384.450 ;
        RECT 829.950 382.950 832.050 383.400 ;
        RECT 830.400 372.600 831.450 382.950 ;
        RECT 836.400 379.050 837.450 400.800 ;
        RECT 838.950 397.950 841.050 400.050 ;
        RECT 835.950 376.950 838.050 379.050 ;
        RECT 839.400 376.050 840.450 397.950 ;
        RECT 838.950 373.950 841.050 376.050 ;
        RECT 830.400 370.350 831.600 372.600 ;
        RECT 835.950 371.100 838.050 373.200 ;
        RECT 842.400 372.600 843.450 406.950 ;
        RECT 836.400 370.350 837.600 371.100 ;
        RECT 842.400 370.350 843.600 372.600 ;
        RECT 845.400 372.450 846.450 416.400 ;
        RECT 850.950 416.100 853.050 418.200 ;
        RECT 857.400 417.600 858.450 427.800 ;
        RECT 862.950 421.950 865.050 424.050 ;
        RECT 851.400 415.350 852.600 416.100 ;
        RECT 857.400 415.350 858.600 417.600 ;
        RECT 863.400 417.450 864.450 421.950 ;
        RECT 872.400 420.450 873.450 475.950 ;
        RECT 875.400 451.050 876.450 479.400 ;
        RECT 878.400 466.050 879.450 488.400 ;
        RECT 884.400 478.050 885.450 488.400 ;
        RECT 883.950 475.950 886.050 478.050 ;
        RECT 884.400 472.050 885.450 475.950 ;
        RECT 883.950 469.950 886.050 472.050 ;
        RECT 886.950 466.950 889.050 469.050 ;
        RECT 877.950 463.950 880.050 466.050 ;
        RECT 874.950 448.950 877.050 451.050 ;
        RECT 877.950 450.000 880.050 454.050 ;
        RECT 883.950 453.450 886.050 454.050 ;
        RECT 887.400 453.450 888.450 466.950 ;
        RECT 883.950 452.400 888.450 453.450 ;
        RECT 883.950 451.950 886.050 452.400 ;
        RECT 884.400 450.600 885.450 451.950 ;
        RECT 878.400 448.350 879.600 450.000 ;
        RECT 884.400 448.350 885.600 450.600 ;
        RECT 877.950 445.950 880.050 448.050 ;
        RECT 880.950 445.950 883.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 881.400 443.400 882.600 445.650 ;
        RECT 887.400 444.900 888.600 445.650 ;
        RECT 874.950 439.950 877.050 442.050 ;
        RECT 869.400 420.000 873.450 420.450 ;
        RECT 868.950 419.400 873.450 420.000 ;
        RECT 863.400 416.400 867.450 417.450 ;
        RECT 850.950 412.950 853.050 415.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 847.950 409.950 850.050 412.050 ;
        RECT 854.400 411.000 855.600 412.650 ;
        RECT 860.400 411.900 861.600 412.650 ;
        RECT 848.400 406.050 849.450 409.950 ;
        RECT 853.950 406.950 856.050 411.000 ;
        RECT 859.950 409.800 862.050 411.900 ;
        RECT 862.950 409.950 865.050 412.050 ;
        RECT 866.400 411.450 867.450 416.400 ;
        RECT 868.950 415.950 871.050 419.400 ;
        RECT 875.400 418.200 876.450 439.950 ;
        RECT 881.400 439.050 882.450 443.400 ;
        RECT 886.950 442.800 889.050 444.900 ;
        RECT 883.950 439.950 886.050 442.050 ;
        RECT 880.950 436.950 883.050 439.050 ;
        RECT 874.950 416.100 877.050 418.200 ;
        RECT 880.950 417.000 883.050 421.050 ;
        RECT 884.400 418.050 885.450 439.950 ;
        RECT 886.950 430.950 889.050 433.050 ;
        RECT 887.400 421.050 888.450 430.950 ;
        RECT 886.950 418.950 889.050 421.050 ;
        RECT 875.400 415.350 876.600 416.100 ;
        RECT 881.400 415.350 882.600 417.000 ;
        RECT 883.950 415.950 886.050 418.050 ;
        RECT 871.950 412.950 874.050 415.050 ;
        RECT 874.950 412.950 877.050 415.050 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 866.400 410.400 870.450 411.450 ;
        RECT 847.950 403.950 850.050 406.050 ;
        RECT 847.950 397.950 850.050 400.050 ;
        RECT 848.400 376.050 849.450 397.950 ;
        RECT 853.950 385.950 856.050 388.050 ;
        RECT 850.950 376.950 853.050 379.050 ;
        RECT 847.950 373.950 850.050 376.050 ;
        RECT 845.400 371.400 849.450 372.450 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 835.950 367.950 838.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 833.400 366.000 834.600 367.650 ;
        RECT 839.400 366.900 840.600 367.650 ;
        RECT 832.950 361.950 835.050 366.000 ;
        RECT 838.950 364.800 841.050 366.900 ;
        RECT 844.950 364.950 847.050 367.050 ;
        RECT 835.950 361.950 838.050 364.050 ;
        RECT 817.950 340.950 820.050 343.050 ;
        RECT 823.950 340.950 826.050 343.050 ;
        RECT 818.400 315.450 819.450 340.950 ;
        RECT 829.950 338.100 832.050 340.200 ;
        RECT 830.400 337.350 831.600 338.100 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 824.100 334.950 826.200 337.050 ;
        RECT 829.500 334.950 831.600 337.050 ;
        RECT 832.800 334.950 834.900 337.050 ;
        RECT 821.400 322.050 822.450 334.950 ;
        RECT 824.400 333.000 825.600 334.650 ;
        RECT 823.950 328.950 826.050 333.000 ;
        RECT 833.400 332.400 834.600 334.650 ;
        RECT 820.950 319.950 823.050 322.050 ;
        RECT 818.400 314.400 822.450 315.450 ;
        RECT 817.950 310.950 820.050 313.050 ;
        RECT 818.400 298.050 819.450 310.950 ;
        RECT 821.400 304.050 822.450 314.400 ;
        RECT 829.950 304.950 832.050 307.050 ;
        RECT 820.950 301.950 823.050 304.050 ;
        RECT 817.950 295.950 820.050 298.050 ;
        RECT 812.400 293.400 816.450 294.450 ;
        RECT 818.400 294.600 819.450 295.950 ;
        RECT 803.400 292.350 804.600 293.100 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 794.400 287.400 795.600 289.650 ;
        RECT 800.400 287.400 801.600 289.650 ;
        RECT 787.950 280.950 790.050 283.050 ;
        RECT 784.950 262.950 787.050 265.050 ;
        RECT 781.950 260.100 784.050 262.200 ;
        RECT 788.400 261.600 789.450 280.950 ;
        RECT 794.400 277.050 795.450 287.400 ;
        RECT 800.400 283.050 801.450 287.400 ;
        RECT 799.950 280.950 802.050 283.050 ;
        RECT 793.950 274.950 796.050 277.050 ;
        RECT 808.950 271.950 811.050 274.050 ;
        RECT 802.950 265.950 805.050 268.050 ;
        RECT 793.950 262.950 796.050 265.050 ;
        RECT 782.400 259.350 783.600 260.100 ;
        RECT 788.400 259.350 789.600 261.600 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 775.950 253.950 778.050 256.050 ;
        RECT 779.400 255.000 780.600 256.650 ;
        RECT 776.400 244.050 777.450 253.950 ;
        RECT 778.950 250.950 781.050 255.000 ;
        RECT 785.400 254.400 786.600 256.650 ;
        RECT 794.400 255.900 795.450 262.950 ;
        RECT 803.400 261.600 804.450 265.950 ;
        RECT 809.400 261.600 810.450 271.950 ;
        RECT 812.400 262.050 813.450 293.400 ;
        RECT 818.400 292.350 819.600 294.600 ;
        RECT 823.950 293.100 826.050 295.200 ;
        RECT 830.400 294.450 831.450 304.950 ;
        RECT 833.400 301.050 834.450 332.400 ;
        RECT 836.400 325.050 837.450 361.950 ;
        RECT 838.950 355.950 841.050 358.050 ;
        RECT 835.950 322.950 838.050 325.050 ;
        RECT 832.950 298.950 835.050 301.050 ;
        RECT 836.400 295.200 837.450 322.950 ;
        RECT 839.400 313.050 840.450 355.950 ;
        RECT 841.950 346.950 844.050 349.050 ;
        RECT 842.400 343.050 843.450 346.950 ;
        RECT 841.950 340.950 844.050 343.050 ;
        RECT 845.400 339.450 846.450 364.950 ;
        RECT 848.400 352.050 849.450 371.400 ;
        RECT 847.950 349.950 850.050 352.050 ;
        RECT 847.950 346.800 850.050 348.900 ;
        RECT 842.400 338.400 846.450 339.450 ;
        RECT 848.400 339.600 849.450 346.800 ;
        RECT 851.400 346.050 852.450 376.950 ;
        RECT 854.400 373.050 855.450 385.950 ;
        RECT 853.950 370.950 856.050 373.050 ;
        RECT 860.400 372.600 861.450 409.800 ;
        RECT 863.400 376.050 864.450 409.950 ;
        RECT 865.950 406.950 868.050 409.050 ;
        RECT 862.950 373.950 865.050 376.050 ;
        RECT 866.400 372.600 867.450 406.950 ;
        RECT 869.400 373.050 870.450 410.400 ;
        RECT 872.400 410.400 873.600 412.650 ;
        RECT 878.400 411.000 879.600 412.650 ;
        RECT 872.400 406.050 873.450 410.400 ;
        RECT 877.950 406.950 880.050 411.000 ;
        RECT 883.950 409.950 886.050 412.050 ;
        RECT 871.950 403.950 874.050 406.050 ;
        RECT 884.400 400.050 885.450 409.950 ;
        RECT 887.400 409.050 888.450 418.950 ;
        RECT 893.400 417.450 894.450 520.950 ;
        RECT 896.400 514.050 897.450 521.400 ;
        RECT 895.950 511.950 898.050 514.050 ;
        RECT 902.400 511.050 903.450 521.400 ;
        RECT 911.400 520.050 912.450 526.800 ;
        RECT 904.950 517.950 907.050 520.050 ;
        RECT 910.950 517.950 913.050 520.050 ;
        RECT 901.950 508.950 904.050 511.050 ;
        RECT 902.400 505.050 903.450 508.950 ;
        RECT 901.950 502.950 904.050 505.050 ;
        RECT 905.400 501.450 906.450 517.950 ;
        RECT 911.400 508.050 912.450 517.950 ;
        RECT 910.950 505.950 913.050 508.050 ;
        RECT 902.400 500.400 906.450 501.450 ;
        RECT 902.400 495.600 903.450 500.400 ;
        RECT 902.400 493.350 903.600 495.600 ;
        RECT 907.950 494.100 910.050 496.200 ;
        RECT 908.400 493.350 909.600 494.100 ;
        RECT 898.950 490.950 901.050 493.050 ;
        RECT 901.950 490.950 904.050 493.050 ;
        RECT 904.950 490.950 907.050 493.050 ;
        RECT 907.950 490.950 910.050 493.050 ;
        RECT 899.400 488.400 900.600 490.650 ;
        RECT 905.400 489.000 906.600 490.650 ;
        RECT 895.950 478.950 898.050 481.050 ;
        RECT 896.400 457.050 897.450 478.950 ;
        RECT 899.400 460.050 900.450 488.400 ;
        RECT 904.950 484.950 907.050 489.000 ;
        RECT 904.950 481.800 907.050 483.900 ;
        RECT 898.950 457.950 901.050 460.050 ;
        RECT 895.950 454.950 898.050 457.050 ;
        RECT 890.400 416.400 894.450 417.450 ;
        RECT 896.400 417.600 897.450 454.950 ;
        RECT 899.400 451.050 900.450 457.950 ;
        RECT 905.400 451.200 906.450 481.800 ;
        RECT 914.400 469.050 915.450 565.950 ;
        RECT 917.400 565.050 918.450 605.400 ;
        RECT 920.400 595.050 921.450 625.950 ;
        RECT 923.400 625.050 924.450 655.800 ;
        RECT 922.950 622.950 925.050 625.050 ;
        RECT 926.400 618.450 927.450 670.950 ;
        RECT 929.400 655.050 930.450 676.800 ;
        RECT 935.400 673.050 936.450 676.950 ;
        RECT 934.950 670.950 937.050 673.050 ;
        RECT 934.950 667.800 937.050 669.900 ;
        RECT 931.950 658.950 934.050 661.050 ;
        RECT 928.950 652.950 931.050 655.050 ;
        RECT 928.950 649.800 931.050 651.900 ;
        RECT 929.400 628.050 930.450 649.800 ;
        RECT 928.950 625.950 931.050 628.050 ;
        RECT 923.400 617.400 927.450 618.450 ;
        RECT 923.400 607.050 924.450 617.400 ;
        RECT 932.400 616.050 933.450 658.950 ;
        RECT 925.950 613.950 931.050 616.050 ;
        RECT 931.950 613.950 934.050 616.050 ;
        RECT 935.400 610.050 936.450 667.800 ;
        RECT 934.950 607.950 937.050 610.050 ;
        RECT 922.950 604.950 925.050 607.050 ;
        RECT 925.950 605.100 928.050 607.200 ;
        RECT 931.950 605.100 934.050 607.200 ;
        RECT 926.400 604.350 927.600 605.100 ;
        RECT 932.400 604.350 933.600 605.100 ;
        RECT 925.950 601.950 928.050 604.050 ;
        RECT 928.950 601.950 931.050 604.050 ;
        RECT 931.950 601.950 934.050 604.050 ;
        RECT 929.400 599.400 930.600 601.650 ;
        RECT 919.950 592.950 922.050 595.050 ;
        RECT 922.950 586.950 925.050 589.050 ;
        RECT 919.950 571.950 922.050 574.050 ;
        RECT 916.950 562.950 919.050 565.050 ;
        RECT 920.400 561.450 921.450 571.950 ;
        RECT 923.400 571.050 924.450 586.950 ;
        RECT 922.950 568.950 925.050 571.050 ;
        RECT 922.950 565.800 925.050 567.900 ;
        RECT 917.400 560.400 921.450 561.450 ;
        RECT 917.400 529.050 918.450 560.400 ;
        RECT 923.400 535.050 924.450 565.800 ;
        RECT 929.400 559.050 930.450 599.400 ;
        RECT 934.950 598.950 937.050 601.050 ;
        RECT 931.950 592.950 934.050 595.050 ;
        RECT 928.950 556.950 931.050 559.050 ;
        RECT 922.950 532.950 925.050 535.050 ;
        RECT 916.950 526.950 919.050 529.050 ;
        RECT 923.400 528.600 924.450 532.950 ;
        RECT 923.400 526.350 924.600 528.600 ;
        RECT 928.950 527.100 931.050 529.200 ;
        RECT 932.400 528.450 933.450 592.950 ;
        RECT 935.400 592.050 936.450 598.950 ;
        RECT 934.950 589.950 937.050 592.050 ;
        RECT 934.950 586.800 937.050 588.900 ;
        RECT 935.400 553.050 936.450 586.800 ;
        RECT 934.950 550.950 937.050 553.050 ;
        RECT 932.400 527.400 936.450 528.450 ;
        RECT 929.400 526.350 930.600 527.100 ;
        RECT 919.950 523.950 922.050 526.050 ;
        RECT 922.950 523.950 925.050 526.050 ;
        RECT 925.950 523.950 928.050 526.050 ;
        RECT 928.950 523.950 931.050 526.050 ;
        RECT 916.950 520.950 919.050 523.050 ;
        RECT 920.400 521.400 921.600 523.650 ;
        RECT 926.400 521.400 927.600 523.650 ;
        RECT 917.400 514.050 918.450 520.950 ;
        RECT 920.400 517.050 921.450 521.400 ;
        RECT 926.400 519.450 927.450 521.400 ;
        RECT 923.400 518.400 927.450 519.450 ;
        RECT 919.950 514.950 922.050 517.050 ;
        RECT 916.950 511.950 919.050 514.050 ;
        RECT 923.400 508.050 924.450 518.400 ;
        RECT 928.950 517.950 931.050 520.050 ;
        RECT 925.950 511.950 928.050 514.050 ;
        RECT 922.950 505.950 925.050 508.050 ;
        RECT 919.950 494.100 922.050 496.200 ;
        RECT 926.400 495.600 927.450 511.950 ;
        RECT 929.400 511.050 930.450 517.950 ;
        RECT 928.950 508.950 931.050 511.050 ;
        RECT 935.400 502.050 936.450 527.400 ;
        RECT 934.950 499.950 937.050 502.050 ;
        RECT 920.400 493.350 921.600 494.100 ;
        RECT 926.400 493.350 927.600 495.600 ;
        RECT 934.950 494.100 937.050 496.200 ;
        RECT 919.950 490.950 922.050 493.050 ;
        RECT 922.950 490.950 925.050 493.050 ;
        RECT 925.950 490.950 928.050 493.050 ;
        RECT 928.950 490.950 931.050 493.050 ;
        RECT 923.400 488.400 924.600 490.650 ;
        RECT 929.400 488.400 930.600 490.650 ;
        RECT 923.400 487.050 924.450 488.400 ;
        RECT 922.950 484.950 925.050 487.050 ;
        RECT 913.950 466.950 916.050 469.050 ;
        RECT 910.950 463.950 913.050 466.050 ;
        RECT 898.950 448.950 901.050 451.050 ;
        RECT 904.950 449.100 907.050 451.200 ;
        RECT 911.400 450.600 912.450 463.950 ;
        RECT 923.400 454.200 924.450 484.950 ;
        RECT 929.400 478.050 930.450 488.400 ;
        RECT 931.950 487.950 934.050 490.050 ;
        RECT 928.950 477.450 931.050 478.050 ;
        RECT 926.400 476.400 931.050 477.450 ;
        RECT 926.400 457.050 927.450 476.400 ;
        RECT 928.950 475.950 931.050 476.400 ;
        RECT 925.950 454.950 928.050 457.050 ;
        RECT 932.400 456.450 933.450 487.950 ;
        RECT 935.400 484.050 936.450 494.100 ;
        RECT 934.950 481.950 937.050 484.050 ;
        RECT 932.400 455.400 936.450 456.450 ;
        RECT 916.950 451.950 919.050 454.050 ;
        RECT 922.950 452.100 925.050 454.200 ;
        RECT 905.400 448.350 906.600 449.100 ;
        RECT 911.400 448.350 912.600 450.600 ;
        RECT 901.950 445.950 904.050 448.050 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 907.950 445.950 910.050 448.050 ;
        RECT 910.950 445.950 913.050 448.050 ;
        RECT 902.400 445.050 903.600 445.650 ;
        RECT 898.950 443.400 903.600 445.050 ;
        RECT 908.400 443.400 909.600 445.650 ;
        RECT 898.950 442.950 903.000 443.400 ;
        RECT 908.400 427.050 909.450 443.400 ;
        RECT 913.950 433.950 916.050 436.050 ;
        RECT 907.950 424.950 910.050 427.050 ;
        RECT 890.400 411.900 891.450 416.400 ;
        RECT 896.400 415.350 897.600 417.600 ;
        RECT 901.950 416.100 904.050 418.200 ;
        RECT 910.950 416.100 913.050 418.200 ;
        RECT 902.400 415.350 903.600 416.100 ;
        RECT 895.950 412.950 898.050 415.050 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 904.950 412.950 907.050 415.050 ;
        RECT 899.400 411.900 900.600 412.650 ;
        RECT 889.950 409.800 892.050 411.900 ;
        RECT 886.950 406.950 889.050 409.050 ;
        RECT 898.950 406.950 901.050 411.900 ;
        RECT 905.400 411.000 906.600 412.650 ;
        RECT 904.950 406.950 907.050 411.000 ;
        RECT 883.950 397.950 886.050 400.050 ;
        RECT 911.400 397.050 912.450 416.100 ;
        RECT 910.950 394.950 913.050 397.050 ;
        RECT 883.950 391.950 886.050 394.050 ;
        RECT 871.950 373.950 874.050 376.050 ;
        RECT 860.400 370.350 861.600 372.600 ;
        RECT 866.400 370.350 867.600 372.600 ;
        RECT 868.950 370.950 871.050 373.050 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 857.400 366.900 858.600 367.650 ;
        RECT 863.400 366.900 864.600 367.650 ;
        RECT 856.950 364.800 859.050 366.900 ;
        RECT 862.950 364.800 865.050 366.900 ;
        RECT 872.400 358.050 873.450 373.950 ;
        RECT 884.400 373.200 885.450 391.950 ;
        RECT 914.400 379.050 915.450 433.950 ;
        RECT 917.400 430.050 918.450 451.950 ;
        RECT 922.950 448.950 925.050 451.050 ;
        RECT 928.950 450.000 931.050 454.050 ;
        RECT 935.400 451.050 936.450 455.400 ;
        RECT 923.400 448.350 924.600 448.950 ;
        RECT 929.400 448.350 930.600 450.000 ;
        RECT 934.950 448.950 937.050 451.050 ;
        RECT 922.950 445.950 925.050 448.050 ;
        RECT 925.950 445.950 928.050 448.050 ;
        RECT 928.950 445.950 931.050 448.050 ;
        RECT 931.950 445.950 934.050 448.050 ;
        RECT 926.400 444.900 927.600 445.650 ;
        RECT 925.950 442.800 928.050 444.900 ;
        RECT 932.400 443.400 933.600 445.650 ;
        RECT 932.400 436.050 933.450 443.400 ;
        RECT 934.950 442.950 937.050 445.050 ;
        RECT 931.950 433.950 934.050 436.050 ;
        RECT 922.950 430.950 925.050 433.050 ;
        RECT 916.950 427.950 919.050 430.050 ;
        RECT 923.400 417.600 924.450 430.950 ;
        RECT 928.950 427.950 931.050 430.050 ;
        RECT 935.400 429.450 936.450 442.950 ;
        RECT 932.400 428.400 936.450 429.450 ;
        RECT 929.400 417.600 930.450 427.950 ;
        RECT 932.400 418.050 933.450 428.400 ;
        RECT 934.950 424.950 937.050 427.050 ;
        RECT 923.400 415.350 924.600 417.600 ;
        RECT 929.400 415.350 930.600 417.600 ;
        RECT 931.950 415.950 934.050 418.050 ;
        RECT 919.950 412.950 922.050 415.050 ;
        RECT 922.950 412.950 925.050 415.050 ;
        RECT 925.950 412.950 928.050 415.050 ;
        RECT 928.950 412.950 931.050 415.050 ;
        RECT 920.400 410.400 921.600 412.650 ;
        RECT 926.400 411.000 927.600 412.650 ;
        RECT 920.400 397.050 921.450 410.400 ;
        RECT 925.950 406.950 928.050 411.000 ;
        RECT 931.950 409.950 934.050 412.050 ;
        RECT 919.950 394.950 922.050 397.050 ;
        RECT 898.950 376.950 901.050 379.050 ;
        RECT 913.950 376.950 916.050 379.050 ;
        RECT 874.950 370.950 877.050 373.050 ;
        RECT 883.950 371.100 886.050 373.200 ;
        RECT 889.950 372.000 892.050 376.050 ;
        RECT 895.950 373.950 898.050 376.050 ;
        RECT 875.400 364.050 876.450 370.950 ;
        RECT 884.400 370.350 885.600 371.100 ;
        RECT 890.400 370.350 891.600 372.000 ;
        RECT 880.950 367.950 883.050 370.050 ;
        RECT 883.950 367.950 886.050 370.050 ;
        RECT 886.950 367.950 889.050 370.050 ;
        RECT 889.950 367.950 892.050 370.050 ;
        RECT 881.400 365.400 882.600 367.650 ;
        RECT 887.400 365.400 888.600 367.650 ;
        RECT 896.400 367.050 897.450 373.950 ;
        RECT 874.950 361.950 877.050 364.050 ;
        RECT 871.950 355.950 874.050 358.050 ;
        RECT 853.950 352.950 856.050 355.050 ;
        RECT 865.950 352.950 868.050 355.050 ;
        RECT 850.950 343.950 853.050 346.050 ;
        RECT 854.400 339.600 855.450 352.950 ;
        RECT 862.950 349.950 865.050 352.050 ;
        RECT 859.950 343.950 862.050 346.050 ;
        RECT 860.400 340.050 861.450 343.950 ;
        RECT 838.950 310.950 841.050 313.050 ;
        RECT 842.400 307.050 843.450 338.400 ;
        RECT 848.400 337.350 849.600 339.600 ;
        RECT 854.400 337.350 855.600 339.600 ;
        RECT 859.950 337.950 862.050 340.050 ;
        RECT 847.950 334.950 850.050 337.050 ;
        RECT 850.950 334.950 853.050 337.050 ;
        RECT 853.950 334.950 856.050 337.050 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 844.950 331.950 847.050 334.050 ;
        RECT 851.400 333.900 852.600 334.650 ;
        RECT 857.400 334.050 858.600 334.650 ;
        RECT 845.400 328.050 846.450 331.950 ;
        RECT 850.950 331.800 853.050 333.900 ;
        RECT 857.400 332.400 862.050 334.050 ;
        RECT 858.000 331.950 862.050 332.400 ;
        RECT 844.950 325.950 847.050 328.050 ;
        RECT 841.950 304.950 844.050 307.050 ;
        RECT 847.950 295.950 850.050 301.050 ;
        RECT 853.950 295.950 856.050 298.050 ;
        RECT 830.400 293.400 834.450 294.450 ;
        RECT 824.400 292.350 825.600 293.100 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 821.400 287.400 822.600 289.650 ;
        RECT 827.400 287.400 828.600 289.650 ;
        RECT 821.400 283.050 822.450 287.400 ;
        RECT 823.950 283.950 826.050 286.050 ;
        RECT 820.950 280.950 823.050 283.050 ;
        RECT 814.950 271.950 817.050 274.050 ;
        RECT 803.400 259.350 804.600 261.600 ;
        RECT 809.400 259.350 810.600 261.600 ;
        RECT 811.950 259.950 814.050 262.050 ;
        RECT 799.950 256.950 802.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 800.400 255.900 801.600 256.650 ;
        RECT 785.400 253.050 786.450 254.400 ;
        RECT 793.950 253.800 796.050 255.900 ;
        RECT 799.950 253.800 802.050 255.900 ;
        RECT 806.400 254.400 807.600 256.650 ;
        RECT 784.950 250.950 787.050 253.050 ;
        RECT 775.950 241.950 778.050 244.050 ;
        RECT 785.400 238.050 786.450 250.950 ;
        RECT 784.950 235.950 787.050 238.050 ;
        RECT 787.950 220.950 790.050 223.050 ;
        RECT 775.950 215.100 778.050 217.200 ;
        RECT 781.950 215.100 784.050 217.200 ;
        RECT 788.400 216.600 789.450 220.950 ;
        RECT 776.400 205.050 777.450 215.100 ;
        RECT 782.400 214.350 783.600 215.100 ;
        RECT 788.400 214.350 789.600 216.600 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 787.950 211.950 790.050 214.050 ;
        RECT 785.400 209.400 786.600 211.650 ;
        RECT 778.950 205.950 781.050 208.050 ;
        RECT 781.950 205.950 784.050 208.050 ;
        RECT 775.950 202.950 778.050 205.050 ;
        RECT 772.950 196.950 775.050 199.050 ;
        RECT 754.950 187.950 757.050 190.050 ;
        RECT 725.400 182.400 732.450 183.450 ;
        RECT 725.400 181.350 726.600 182.400 ;
        RECT 718.950 178.950 721.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 715.950 172.950 718.050 178.050 ;
        RECT 722.400 177.900 723.600 178.650 ;
        RECT 721.950 175.800 724.050 177.900 ;
        RECT 731.400 175.050 732.450 182.400 ;
        RECT 733.950 181.950 736.050 184.050 ;
        RECT 742.950 182.100 745.050 184.200 ;
        RECT 718.950 172.950 721.050 175.050 ;
        RECT 730.950 172.950 733.050 175.050 ;
        RECT 712.950 140.100 715.050 142.200 ;
        RECT 707.400 136.350 708.600 138.600 ;
        RECT 712.950 136.950 715.050 139.050 ;
        RECT 713.400 136.350 714.600 136.950 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 709.950 133.950 712.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 710.400 132.000 711.600 133.650 ;
        RECT 709.950 127.950 712.050 132.000 ;
        RECT 712.950 118.950 715.050 121.050 ;
        RECT 700.950 109.950 703.050 112.050 ;
        RECT 682.950 104.100 685.050 106.200 ;
        RECT 688.950 104.100 691.050 106.200 ;
        RECT 697.950 104.100 700.050 106.200 ;
        RECT 706.950 104.100 709.050 106.200 ;
        RECT 713.400 105.600 714.450 118.950 ;
        RECT 719.400 106.050 720.450 172.950 ;
        RECT 734.400 157.050 735.450 181.950 ;
        RECT 743.400 181.350 744.600 182.100 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 739.950 178.950 742.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 740.400 177.000 741.600 178.650 ;
        RECT 746.400 177.900 747.600 178.650 ;
        RECT 739.950 172.950 742.050 177.000 ;
        RECT 745.950 175.800 748.050 177.900 ;
        RECT 733.950 154.950 736.050 157.050 ;
        RECT 730.950 148.950 733.050 151.050 ;
        RECT 721.950 139.950 724.050 142.050 ;
        RECT 683.400 103.350 684.600 104.100 ;
        RECT 689.400 103.350 690.600 104.100 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 685.950 100.950 688.050 103.050 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 686.400 99.900 687.600 100.650 ;
        RECT 692.400 99.900 693.600 100.650 ;
        RECT 676.950 97.800 679.050 99.900 ;
        RECT 685.950 97.800 688.050 99.900 ;
        RECT 691.950 97.800 694.050 99.900 ;
        RECT 673.950 91.950 676.050 94.050 ;
        RECT 679.950 91.950 682.050 94.050 ;
        RECT 664.950 88.950 667.050 91.050 ;
        RECT 673.950 85.950 676.050 88.050 ;
        RECT 655.950 73.950 658.050 76.050 ;
        RECT 635.400 58.350 636.600 60.600 ;
        RECT 641.400 58.350 642.600 60.600 ;
        RECT 652.950 59.100 655.050 61.200 ;
        RECT 656.400 60.600 657.450 73.950 ;
        RECT 656.400 58.350 657.600 60.600 ;
        RECT 661.950 59.100 664.050 61.200 ;
        RECT 662.400 58.350 663.600 59.100 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 638.400 53.400 639.600 55.650 ;
        RECT 644.400 53.400 645.600 55.650 ;
        RECT 659.400 53.400 660.600 55.650 ;
        RECT 665.400 54.000 666.600 55.650 ;
        RECT 638.400 49.050 639.450 53.400 ;
        RECT 637.950 46.950 640.050 49.050 ;
        RECT 644.400 43.050 645.450 53.400 ;
        RECT 646.950 43.950 649.050 46.050 ;
        RECT 628.950 40.950 631.050 43.050 ;
        RECT 643.950 40.950 646.050 43.050 ;
        RECT 647.400 37.050 648.450 43.950 ;
        RECT 659.400 37.050 660.450 53.400 ;
        RECT 664.950 49.950 667.050 54.000 ;
        RECT 646.950 34.950 649.050 37.050 ;
        RECT 658.950 34.950 661.050 37.050 ;
        RECT 670.950 34.950 673.050 37.050 ;
        RECT 664.950 31.950 667.050 34.050 ;
        RECT 622.950 28.950 625.050 31.050 ;
        RECT 623.400 27.600 624.450 28.950 ;
        RECT 617.400 25.350 618.600 27.600 ;
        RECT 623.400 25.350 624.600 27.600 ;
        RECT 637.950 26.100 640.050 28.200 ;
        RECT 658.950 27.000 661.050 31.050 ;
        RECT 665.400 27.600 666.450 31.950 ;
        RECT 638.400 25.350 639.600 26.100 ;
        RECT 659.400 25.350 660.600 27.000 ;
        RECT 665.400 25.350 666.600 27.600 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 620.400 20.400 621.600 22.650 ;
        RECT 626.400 21.900 627.600 22.650 ;
        RECT 641.400 21.900 642.600 22.650 ;
        RECT 656.400 21.900 657.600 22.650 ;
        RECT 662.400 21.900 663.600 22.650 ;
        RECT 671.400 21.900 672.450 34.950 ;
        RECT 674.400 34.050 675.450 85.950 ;
        RECT 680.400 82.050 681.450 91.950 ;
        RECT 692.400 88.050 693.450 97.800 ;
        RECT 691.950 85.950 694.050 88.050 ;
        RECT 698.400 85.050 699.450 104.100 ;
        RECT 707.400 103.350 708.600 104.100 ;
        RECT 713.400 103.350 714.600 105.600 ;
        RECT 718.950 103.950 721.050 106.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 709.950 100.950 712.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 704.400 98.400 705.600 100.650 ;
        RECT 710.400 98.400 711.600 100.650 ;
        RECT 716.400 99.000 717.600 100.650 ;
        RECT 704.400 85.050 705.450 98.400 ;
        RECT 710.400 94.050 711.450 98.400 ;
        RECT 715.950 94.950 718.050 99.000 ;
        RECT 718.950 97.950 721.050 100.050 ;
        RECT 709.950 91.950 712.050 94.050 ;
        RECT 697.950 82.950 700.050 85.050 ;
        RECT 703.950 82.950 706.050 85.050 ;
        RECT 679.950 79.950 682.050 82.050 ;
        RECT 688.950 76.950 691.050 79.050 ;
        RECT 689.400 64.050 690.450 76.950 ;
        RECT 694.950 67.950 697.050 70.050 ;
        RECT 688.950 61.950 691.050 64.050 ;
        RECT 682.950 59.100 685.050 61.200 ;
        RECT 689.400 60.600 690.450 61.950 ;
        RECT 683.400 58.350 684.600 59.100 ;
        RECT 689.400 58.350 690.600 60.600 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 680.400 54.000 681.600 55.650 ;
        RECT 679.950 49.950 682.050 54.000 ;
        RECT 686.400 53.400 687.600 55.650 ;
        RECT 686.400 46.050 687.450 53.400 ;
        RECT 688.950 46.950 691.050 49.050 ;
        RECT 685.950 43.950 688.050 46.050 ;
        RECT 686.400 34.050 687.450 43.950 ;
        RECT 673.950 31.950 676.050 34.050 ;
        RECT 679.950 31.950 682.050 34.050 ;
        RECT 685.950 31.950 688.050 34.050 ;
        RECT 680.400 27.600 681.450 31.950 ;
        RECT 689.400 30.450 690.450 46.950 ;
        RECT 695.400 46.050 696.450 67.950 ;
        RECT 698.400 49.050 699.450 82.950 ;
        RECT 706.950 60.000 709.050 64.050 ;
        RECT 707.400 58.350 708.600 60.000 ;
        RECT 715.950 58.950 718.050 61.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 704.400 54.000 705.600 55.650 ;
        RECT 710.400 54.000 711.600 55.650 ;
        RECT 703.950 49.950 706.050 54.000 ;
        RECT 709.950 49.950 712.050 54.000 ;
        RECT 716.400 52.050 717.450 58.950 ;
        RECT 719.400 54.900 720.450 97.950 ;
        RECT 722.400 61.200 723.450 139.950 ;
        RECT 731.400 138.600 732.450 148.950 ;
        RECT 731.400 136.350 732.600 138.600 ;
        RECT 736.950 138.000 739.050 142.050 ;
        RECT 740.400 139.050 741.450 172.950 ;
        RECT 742.950 148.950 745.050 151.050 ;
        RECT 737.400 136.350 738.600 138.000 ;
        RECT 739.950 136.950 742.050 139.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 728.400 131.400 729.600 133.650 ;
        RECT 734.400 132.000 735.600 133.650 ;
        RECT 743.400 133.050 744.450 148.950 ;
        RECT 752.400 142.200 753.450 181.950 ;
        RECT 755.400 177.900 756.450 187.950 ;
        RECT 779.400 187.050 780.450 205.950 ;
        RECT 782.400 202.050 783.450 205.950 ;
        RECT 781.950 199.950 784.050 202.050 ;
        RECT 785.400 196.050 786.450 209.400 ;
        RECT 794.400 208.050 795.450 253.800 ;
        RECT 806.400 241.050 807.450 254.400 ;
        RECT 811.950 253.950 814.050 256.050 ;
        RECT 805.950 238.950 808.050 241.050 ;
        RECT 799.950 235.950 802.050 238.050 ;
        RECT 800.400 216.600 801.450 235.950 ;
        RECT 806.400 216.600 807.450 238.950 ;
        RECT 800.400 214.350 801.600 216.600 ;
        RECT 806.400 214.350 807.600 216.600 ;
        RECT 812.400 216.450 813.450 253.950 ;
        RECT 815.400 235.050 816.450 271.950 ;
        RECT 824.400 261.600 825.450 283.950 ;
        RECT 827.400 271.050 828.450 287.400 ;
        RECT 829.950 271.950 832.050 274.050 ;
        RECT 826.950 268.950 829.050 271.050 ;
        RECT 830.400 261.600 831.450 271.950 ;
        RECT 833.400 262.050 834.450 293.400 ;
        RECT 835.950 293.100 838.050 295.200 ;
        RECT 841.950 293.100 844.050 295.200 ;
        RECT 848.400 294.600 849.450 295.950 ;
        RECT 842.400 292.350 843.600 293.100 ;
        RECT 848.400 292.350 849.600 294.600 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 841.950 289.950 844.050 292.050 ;
        RECT 844.950 289.950 847.050 292.050 ;
        RECT 847.950 289.950 850.050 292.050 ;
        RECT 839.400 287.400 840.600 289.650 ;
        RECT 845.400 288.900 846.600 289.650 ;
        RECT 839.400 264.450 840.450 287.400 ;
        RECT 844.950 286.800 847.050 288.900 ;
        RECT 854.400 265.050 855.450 295.950 ;
        RECT 860.400 294.600 861.450 331.950 ;
        RECT 863.400 298.050 864.450 349.950 ;
        RECT 866.400 328.050 867.450 352.950 ;
        RECT 881.400 352.050 882.450 365.400 ;
        RECT 883.950 361.950 886.050 364.050 ;
        RECT 868.950 349.950 871.050 352.050 ;
        RECT 874.950 349.950 877.050 352.050 ;
        RECT 880.950 349.950 883.050 352.050 ;
        RECT 884.400 351.450 885.450 361.950 ;
        RECT 887.400 355.050 888.450 365.400 ;
        RECT 895.950 364.950 898.050 367.050 ;
        RECT 886.950 352.950 889.050 355.050 ;
        RECT 884.400 350.400 888.450 351.450 ;
        RECT 869.400 340.050 870.450 349.950 ;
        RECT 868.950 337.950 871.050 340.050 ;
        RECT 875.400 339.600 876.450 349.950 ;
        RECT 882.000 348.600 886.050 349.050 ;
        RECT 881.400 346.950 886.050 348.600 ;
        RECT 881.400 339.600 882.450 346.950 ;
        RECT 883.950 343.800 886.050 345.900 ;
        RECT 884.400 340.050 885.450 343.800 ;
        RECT 875.400 337.350 876.600 339.600 ;
        RECT 881.400 337.350 882.600 339.600 ;
        RECT 883.950 337.950 886.050 340.050 ;
        RECT 871.950 334.950 874.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 880.950 334.950 883.050 337.050 ;
        RECT 872.400 333.900 873.600 334.650 ;
        RECT 871.950 331.800 874.050 333.900 ;
        RECT 878.400 333.000 879.600 334.650 ;
        RECT 877.950 328.950 880.050 333.000 ;
        RECT 865.950 325.950 868.050 328.050 ;
        RECT 874.950 310.950 877.050 313.050 ;
        RECT 865.950 304.950 868.050 307.050 ;
        RECT 866.400 298.050 867.450 304.950 ;
        RECT 862.950 295.950 865.050 298.050 ;
        RECT 860.400 292.350 861.600 294.600 ;
        RECT 865.950 294.000 868.050 298.050 ;
        RECT 866.400 292.350 867.600 294.000 ;
        RECT 859.950 289.950 862.050 292.050 ;
        RECT 862.950 289.950 865.050 292.050 ;
        RECT 865.950 289.950 868.050 292.050 ;
        RECT 868.950 289.950 871.050 292.050 ;
        RECT 863.400 288.900 864.600 289.650 ;
        RECT 862.950 286.800 865.050 288.900 ;
        RECT 869.400 287.400 870.600 289.650 ;
        RECT 869.400 280.050 870.450 287.400 ;
        RECT 868.950 277.950 871.050 280.050 ;
        RECT 868.950 271.950 871.050 274.050 ;
        RECT 862.950 265.950 865.050 268.050 ;
        RECT 836.400 263.400 840.450 264.450 ;
        RECT 824.400 259.350 825.600 261.600 ;
        RECT 830.400 259.350 831.600 261.600 ;
        RECT 832.950 259.950 835.050 262.050 ;
        RECT 820.950 256.950 823.050 259.050 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 821.400 254.400 822.600 256.650 ;
        RECT 827.400 254.400 828.600 256.650 ;
        RECT 821.400 252.450 822.450 254.400 ;
        RECT 821.400 251.400 825.450 252.450 ;
        RECT 814.950 232.950 817.050 235.050 ;
        RECT 824.400 226.050 825.450 251.400 ;
        RECT 827.400 241.050 828.450 254.400 ;
        RECT 832.950 253.950 835.050 256.050 ;
        RECT 826.950 238.950 829.050 241.050 ;
        RECT 823.950 223.950 826.050 226.050 ;
        RECT 824.400 216.600 825.450 223.950 ;
        RECT 833.400 219.450 834.450 253.950 ;
        RECT 830.400 218.400 834.450 219.450 ;
        RECT 812.400 215.400 816.450 216.450 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 803.400 209.400 804.600 211.650 ;
        RECT 809.400 210.000 810.600 211.650 ;
        RECT 793.950 205.950 796.050 208.050 ;
        RECT 784.950 193.950 787.050 196.050 ;
        RECT 778.950 186.450 781.050 187.050 ;
        RECT 776.400 185.400 781.050 186.450 ;
        RECT 763.950 182.100 766.050 184.200 ;
        RECT 764.400 181.350 765.600 182.100 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 761.400 177.900 762.600 178.650 ;
        RECT 754.950 175.800 757.050 177.900 ;
        RECT 760.950 175.800 763.050 177.900 ;
        RECT 767.400 176.400 768.600 178.650 ;
        RECT 767.400 169.050 768.450 176.400 ;
        RECT 766.950 166.950 769.050 169.050 ;
        RECT 773.400 166.050 774.450 178.950 ;
        RECT 772.950 163.950 775.050 166.050 ;
        RECT 751.950 140.100 754.050 142.200 ;
        RECT 776.400 142.050 777.450 185.400 ;
        RECT 778.950 184.950 781.050 185.400 ;
        RECT 781.950 182.100 784.050 184.200 ;
        RECT 787.950 182.100 790.050 184.200 ;
        RECT 796.950 182.100 799.050 184.200 ;
        RECT 803.400 184.050 804.450 209.400 ;
        RECT 808.950 205.950 811.050 210.000 ;
        RECT 782.400 181.350 783.600 182.100 ;
        RECT 788.400 181.350 789.600 182.100 ;
        RECT 781.950 178.950 784.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 785.400 176.400 786.600 178.650 ;
        RECT 791.400 177.900 792.600 178.650 ;
        RECT 785.400 172.050 786.450 176.400 ;
        RECT 790.950 175.800 793.050 177.900 ;
        RECT 790.950 172.650 793.050 174.750 ;
        RECT 784.950 169.950 787.050 172.050 ;
        RECT 787.950 166.950 790.050 169.050 ;
        RECT 778.950 142.950 781.050 145.050 ;
        RECT 745.950 136.950 748.050 139.050 ;
        RECT 751.950 136.950 754.050 139.050 ;
        RECT 757.950 138.000 760.050 142.050 ;
        RECT 766.950 139.950 769.050 142.050 ;
        RECT 775.950 139.950 778.050 142.050 ;
        RECT 728.400 105.450 729.450 131.400 ;
        RECT 733.950 127.950 736.050 132.000 ;
        RECT 742.950 130.950 745.050 133.050 ;
        RECT 746.400 130.050 747.450 136.950 ;
        RECT 752.400 136.350 753.600 136.950 ;
        RECT 758.400 136.350 759.600 138.000 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 760.950 133.950 763.050 136.050 ;
        RECT 755.400 132.900 756.600 133.650 ;
        RECT 761.400 132.900 762.600 133.650 ;
        RECT 745.950 127.950 748.050 130.050 ;
        RECT 748.950 127.950 751.050 132.900 ;
        RECT 754.950 130.800 757.050 132.900 ;
        RECT 760.950 130.800 763.050 132.900 ;
        RECT 745.950 112.950 748.050 115.050 ;
        RECT 739.950 109.950 742.050 112.050 ;
        RECT 725.400 104.400 729.450 105.450 ;
        RECT 725.400 91.050 726.450 104.400 ;
        RECT 730.950 104.100 733.050 106.200 ;
        RECT 731.400 103.350 732.600 104.100 ;
        RECT 730.950 100.950 733.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 734.400 99.900 735.600 100.650 ;
        RECT 733.950 97.800 736.050 99.900 ;
        RECT 724.950 88.950 727.050 91.050 ;
        RECT 740.400 73.050 741.450 109.950 ;
        RECT 746.400 105.600 747.450 112.950 ;
        RECT 767.400 109.050 768.450 139.950 ;
        RECT 772.950 137.100 775.050 139.200 ;
        RECT 779.400 138.600 780.450 142.950 ;
        RECT 773.400 136.350 774.600 137.100 ;
        RECT 779.400 136.350 780.600 138.600 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 781.950 133.950 784.050 136.050 ;
        RECT 776.400 131.400 777.600 133.650 ;
        RECT 782.400 131.400 783.600 133.650 ;
        RECT 776.400 124.050 777.450 131.400 ;
        RECT 778.950 127.950 781.050 130.050 ;
        RECT 775.950 121.950 778.050 124.050 ;
        RECT 779.400 121.050 780.450 127.950 ;
        RECT 778.950 118.950 781.050 121.050 ;
        RECT 775.950 115.950 778.050 118.050 ;
        RECT 760.950 106.950 763.050 109.050 ;
        RECT 766.950 106.950 769.050 109.050 ;
        RECT 746.400 103.350 747.600 105.600 ;
        RECT 751.950 104.100 754.050 106.200 ;
        RECT 752.400 103.350 753.600 104.100 ;
        RECT 745.950 100.950 748.050 103.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 751.950 100.950 754.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 749.400 99.900 750.600 100.650 ;
        RECT 755.400 99.900 756.600 100.650 ;
        RECT 761.400 99.900 762.450 106.950 ;
        RECT 769.950 104.100 772.050 106.200 ;
        RECT 776.400 105.600 777.450 115.950 ;
        RECT 770.400 103.350 771.600 104.100 ;
        RECT 776.400 103.350 777.600 105.600 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 767.400 99.900 768.600 100.650 ;
        RECT 748.950 97.800 751.050 99.900 ;
        RECT 754.950 97.800 757.050 99.900 ;
        RECT 760.950 97.800 763.050 99.900 ;
        RECT 766.950 97.800 769.050 99.900 ;
        RECT 773.400 99.000 774.600 100.650 ;
        RECT 772.950 94.950 775.050 99.000 ;
        RECT 739.950 70.950 742.050 73.050 ;
        RECT 751.950 70.950 754.050 73.050 ;
        RECT 757.950 70.950 760.050 73.050 ;
        RECT 775.950 70.950 778.050 73.050 ;
        RECT 736.950 64.950 739.050 67.050 ;
        RECT 721.950 59.100 724.050 61.200 ;
        RECT 730.950 59.100 733.050 61.200 ;
        RECT 722.400 58.350 723.600 59.100 ;
        RECT 731.400 58.350 732.600 59.100 ;
        RECT 722.100 55.950 724.200 58.050 ;
        RECT 727.500 55.950 729.600 58.050 ;
        RECT 730.800 55.950 732.900 58.050 ;
        RECT 728.400 54.900 729.600 55.650 ;
        RECT 737.400 54.900 738.450 64.950 ;
        RECT 745.950 59.100 748.050 61.200 ;
        RECT 752.400 60.600 753.450 70.950 ;
        RECT 746.400 58.350 747.600 59.100 ;
        RECT 752.400 58.350 753.600 60.600 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 745.950 55.950 748.050 58.050 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 743.400 54.900 744.600 55.650 ;
        RECT 718.950 52.800 721.050 54.900 ;
        RECT 727.950 52.800 730.050 54.900 ;
        RECT 736.950 52.800 739.050 54.900 ;
        RECT 742.950 52.800 745.050 54.900 ;
        RECT 749.400 53.400 750.600 55.650 ;
        RECT 758.400 54.900 759.450 70.950 ;
        RECT 767.400 60.450 768.600 60.600 ;
        RECT 767.400 59.400 774.450 60.450 ;
        RECT 767.400 58.350 768.600 59.400 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 764.400 54.900 765.600 55.650 ;
        RECT 715.950 49.950 718.050 52.050 ;
        RECT 697.950 46.950 700.050 49.050 ;
        RECT 706.950 46.950 709.050 49.050 ;
        RECT 694.950 43.950 697.050 46.050 ;
        RECT 691.950 40.950 694.050 43.050 ;
        RECT 686.400 29.400 690.450 30.450 ;
        RECT 686.400 27.600 687.450 29.400 ;
        RECT 680.400 25.350 681.600 27.600 ;
        RECT 686.400 25.350 687.600 27.600 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 677.400 21.900 678.600 22.650 ;
        RECT 683.400 21.900 684.600 22.650 ;
        RECT 692.400 21.900 693.450 40.950 ;
        RECT 707.400 37.050 708.450 46.950 ;
        RECT 712.950 37.950 715.050 40.050 ;
        RECT 700.950 34.950 703.050 37.050 ;
        RECT 706.950 34.950 709.050 37.050 ;
        RECT 701.400 27.600 702.450 34.950 ;
        RECT 701.400 25.350 702.600 27.600 ;
        RECT 706.950 26.100 709.050 28.200 ;
        RECT 713.400 28.050 714.450 37.950 ;
        RECT 707.400 25.350 708.600 26.100 ;
        RECT 712.950 25.950 715.050 28.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 620.400 13.050 621.450 20.400 ;
        RECT 625.950 19.800 628.050 21.900 ;
        RECT 640.950 19.800 643.050 21.900 ;
        RECT 655.950 19.800 658.050 21.900 ;
        RECT 661.950 19.800 664.050 21.900 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 676.950 19.800 679.050 21.900 ;
        RECT 682.950 19.800 685.050 21.900 ;
        RECT 691.950 19.800 694.050 21.900 ;
        RECT 704.400 20.400 705.600 22.650 ;
        RECT 710.400 21.900 711.600 22.650 ;
        RECT 641.400 16.050 642.450 19.800 ;
        RECT 640.950 13.950 643.050 16.050 ;
        RECT 671.400 13.050 672.450 19.800 ;
        RECT 619.950 10.950 622.050 13.050 ;
        RECT 670.950 10.950 673.050 13.050 ;
        RECT 704.400 10.050 705.450 20.400 ;
        RECT 709.950 19.800 712.050 21.900 ;
        RECT 716.400 16.050 717.450 49.950 ;
        RECT 719.400 31.050 720.450 52.800 ;
        RECT 727.950 37.950 730.050 40.050 ;
        RECT 718.950 28.950 721.050 31.050 ;
        RECT 719.400 21.900 720.450 28.950 ;
        RECT 728.400 27.600 729.450 37.950 ;
        RECT 728.400 25.350 729.600 27.600 ;
        RECT 724.950 22.950 727.050 25.050 ;
        RECT 727.950 22.950 730.050 25.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 725.400 21.900 726.600 22.650 ;
        RECT 718.950 19.800 721.050 21.900 ;
        RECT 724.950 19.800 727.050 21.900 ;
        RECT 731.400 20.400 732.600 22.650 ;
        RECT 731.400 16.050 732.450 20.400 ;
        RECT 715.950 13.950 718.050 16.050 ;
        RECT 730.950 13.950 733.050 16.050 ;
        RECT 737.400 10.050 738.450 52.800 ;
        RECT 749.400 34.050 750.450 53.400 ;
        RECT 757.950 52.800 760.050 54.900 ;
        RECT 763.950 52.800 766.050 54.900 ;
        RECT 758.400 49.050 759.450 52.800 ;
        RECT 757.950 46.950 760.050 49.050 ;
        RECT 769.950 37.950 772.050 40.050 ;
        RECT 748.950 31.950 751.050 34.050 ;
        RECT 745.950 27.000 748.050 31.050 ;
        RECT 760.950 28.950 763.050 31.050 ;
        RECT 746.400 25.350 747.600 27.000 ;
        RECT 743.100 22.950 745.200 25.050 ;
        RECT 746.400 22.950 748.500 25.050 ;
        RECT 751.800 22.950 753.900 25.050 ;
        RECT 743.400 20.400 744.600 22.650 ;
        RECT 752.400 20.400 753.600 22.650 ;
        RECT 761.400 21.900 762.450 28.950 ;
        RECT 770.400 27.600 771.450 37.950 ;
        RECT 773.400 31.050 774.450 59.400 ;
        RECT 776.400 43.050 777.450 70.950 ;
        RECT 782.400 63.450 783.450 131.400 ;
        RECT 788.400 118.050 789.450 166.950 ;
        RECT 791.400 139.050 792.450 172.650 ;
        RECT 797.400 169.050 798.450 182.100 ;
        RECT 802.950 181.950 805.050 184.050 ;
        RECT 805.950 183.000 808.050 187.050 ;
        RECT 806.400 181.350 807.600 183.000 ;
        RECT 799.950 178.950 802.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 800.400 175.050 801.450 178.950 ;
        RECT 809.400 176.400 810.600 178.650 ;
        RECT 799.950 172.950 802.050 175.050 ;
        RECT 802.950 172.950 805.050 175.050 ;
        RECT 796.950 166.950 799.050 169.050 ;
        RECT 803.400 163.050 804.450 172.950 ;
        RECT 802.950 160.950 805.050 163.050 ;
        RECT 809.400 145.050 810.450 176.400 ;
        RECT 790.950 136.950 793.050 139.050 ;
        RECT 796.950 138.000 799.050 145.050 ;
        RECT 808.950 142.950 811.050 145.050 ;
        RECT 815.400 142.200 816.450 215.400 ;
        RECT 824.400 214.350 825.600 216.600 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 821.400 210.000 822.600 211.650 ;
        RECT 820.950 205.950 823.050 210.000 ;
        RECT 830.400 205.050 831.450 218.400 ;
        RECT 836.400 216.450 837.450 263.400 ;
        RECT 853.950 262.950 856.050 265.050 ;
        RECT 859.950 262.950 862.050 265.050 ;
        RECT 838.950 259.950 841.050 262.050 ;
        RECT 844.950 260.100 847.050 262.200 ;
        RECT 850.950 260.100 853.050 262.200 ;
        RECT 839.400 244.050 840.450 259.950 ;
        RECT 845.400 259.350 846.600 260.100 ;
        RECT 851.400 259.350 852.600 260.100 ;
        RECT 844.950 256.950 847.050 259.050 ;
        RECT 847.950 256.950 850.050 259.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 848.400 255.000 849.600 256.650 ;
        RECT 854.400 255.000 855.600 256.650 ;
        RECT 847.950 250.950 850.050 255.000 ;
        RECT 853.950 250.950 856.050 255.000 ;
        RECT 856.800 253.950 858.900 256.050 ;
        RECT 860.400 255.900 861.450 262.950 ;
        RECT 853.950 249.450 856.050 249.900 ;
        RECT 857.400 249.450 858.450 253.950 ;
        RECT 859.950 253.800 862.050 255.900 ;
        RECT 853.950 248.400 858.450 249.450 ;
        RECT 853.950 247.800 856.050 248.400 ;
        RECT 838.950 241.950 841.050 244.050 ;
        RECT 839.400 220.050 840.450 241.950 ;
        RECT 850.950 238.950 853.050 241.050 ;
        RECT 841.950 232.950 844.050 235.050 ;
        RECT 838.950 217.950 841.050 220.050 ;
        RECT 833.400 215.400 837.450 216.450 ;
        RECT 842.400 216.600 843.450 232.950 ;
        RECT 847.950 223.950 850.050 226.050 ;
        RECT 848.400 216.600 849.450 223.950 ;
        RECT 851.400 217.050 852.450 238.950 ;
        RECT 829.950 202.950 832.050 205.050 ;
        RECT 829.950 199.800 832.050 201.900 ;
        RECT 817.950 184.950 820.050 187.050 ;
        RECT 797.400 136.350 798.600 138.000 ;
        RECT 802.950 137.100 805.050 142.050 ;
        RECT 808.950 139.800 811.050 141.900 ;
        RECT 814.950 140.100 817.050 142.200 ;
        RECT 818.400 141.450 819.450 184.950 ;
        RECT 823.950 182.100 826.050 184.200 ;
        RECT 830.400 183.600 831.450 199.800 ;
        RECT 833.400 187.050 834.450 215.400 ;
        RECT 842.400 214.350 843.600 216.600 ;
        RECT 848.400 214.350 849.600 216.600 ;
        RECT 850.950 214.950 853.050 217.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 839.400 209.400 840.600 211.650 ;
        RECT 845.400 210.900 846.600 211.650 ;
        RECT 835.950 202.950 838.050 205.050 ;
        RECT 832.950 184.950 835.050 187.050 ;
        RECT 836.400 184.050 837.450 202.950 ;
        RECT 824.400 181.350 825.600 182.100 ;
        RECT 830.400 181.350 831.600 183.600 ;
        RECT 835.950 181.950 838.050 184.050 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 827.400 176.400 828.600 178.650 ;
        RECT 833.400 177.900 834.600 178.650 ;
        RECT 818.400 140.400 822.450 141.450 ;
        RECT 803.400 136.350 804.600 137.100 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 790.950 130.950 793.050 133.050 ;
        RECT 794.400 131.400 795.600 133.650 ;
        RECT 800.400 132.900 801.600 133.650 ;
        RECT 791.400 126.450 792.450 130.950 ;
        RECT 794.400 129.450 795.450 131.400 ;
        RECT 799.950 130.800 802.050 132.900 ;
        RECT 794.400 128.400 798.450 129.450 ;
        RECT 791.400 125.400 795.450 126.450 ;
        RECT 787.950 115.950 790.050 118.050 ;
        RECT 794.400 117.450 795.450 125.400 ;
        RECT 797.400 120.450 798.450 128.400 ;
        RECT 800.400 124.050 801.450 130.800 ;
        RECT 799.950 121.950 802.050 124.050 ;
        RECT 797.400 119.400 801.450 120.450 ;
        RECT 794.400 116.400 798.450 117.450 ;
        RECT 790.950 112.950 793.050 115.050 ;
        RECT 791.400 106.200 792.450 112.950 ;
        RECT 790.950 104.100 793.050 106.200 ;
        RECT 797.400 105.600 798.450 116.400 ;
        RECT 800.400 106.050 801.450 119.400 ;
        RECT 805.950 115.950 808.050 118.050 ;
        RECT 791.400 103.350 792.600 104.100 ;
        RECT 797.400 103.350 798.600 105.600 ;
        RECT 799.950 103.950 802.050 106.050 ;
        RECT 806.400 105.450 807.450 115.950 ;
        RECT 809.400 109.050 810.450 139.800 ;
        RECT 821.400 139.200 822.450 140.400 ;
        RECT 814.950 136.950 817.050 139.050 ;
        RECT 820.950 137.100 823.050 139.200 ;
        RECT 827.400 139.050 828.450 176.400 ;
        RECT 832.950 175.800 835.050 177.900 ;
        RECT 835.950 175.950 838.050 178.050 ;
        RECT 839.400 177.900 840.450 209.400 ;
        RECT 844.950 208.800 847.050 210.900 ;
        RECT 854.400 210.450 855.450 247.800 ;
        RECT 859.950 232.950 862.050 235.050 ;
        RECT 856.950 220.950 859.050 223.050 ;
        RECT 851.400 209.400 855.450 210.450 ;
        RECT 841.950 196.950 844.050 199.050 ;
        RECT 836.400 142.050 837.450 175.950 ;
        RECT 838.950 175.800 841.050 177.900 ;
        RECT 838.950 142.950 841.050 145.050 ;
        RECT 835.950 139.950 838.050 142.050 ;
        RECT 815.400 136.350 816.600 136.950 ;
        RECT 821.400 136.350 822.600 137.100 ;
        RECT 826.950 136.950 829.050 139.050 ;
        RECT 829.950 136.950 832.050 139.050 ;
        RECT 839.400 138.600 840.450 142.950 ;
        RECT 842.400 142.050 843.450 196.950 ;
        RECT 844.950 190.950 847.050 193.050 ;
        RECT 845.400 184.050 846.450 190.950 ;
        RECT 844.950 181.950 847.050 184.050 ;
        RECT 851.400 183.600 852.450 209.400 ;
        RECT 857.400 199.050 858.450 220.950 ;
        RECT 860.400 217.050 861.450 232.950 ;
        RECT 863.400 229.050 864.450 265.950 ;
        RECT 869.400 261.600 870.450 271.950 ;
        RECT 875.400 268.050 876.450 310.950 ;
        RECT 878.400 295.050 879.450 328.950 ;
        RECT 887.400 310.050 888.450 350.400 ;
        RECT 889.950 346.950 892.050 349.050 ;
        RECT 890.400 340.050 891.450 346.950 ;
        RECT 899.400 346.050 900.450 376.950 ;
        RECT 904.950 371.100 907.050 373.200 ;
        RECT 910.950 372.000 913.050 376.050 ;
        RECT 905.400 370.350 906.600 371.100 ;
        RECT 911.400 370.350 912.600 372.000 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 907.950 367.950 910.050 370.050 ;
        RECT 910.950 367.950 913.050 370.050 ;
        RECT 913.950 367.950 916.050 370.050 ;
        RECT 908.400 365.400 909.600 367.650 ;
        RECT 914.400 365.400 915.600 367.650 ;
        RECT 901.950 358.950 904.050 361.050 ;
        RECT 898.950 343.950 901.050 346.050 ;
        RECT 902.400 340.200 903.450 358.950 ;
        RECT 908.400 355.050 909.450 365.400 ;
        RECT 907.950 352.950 910.050 355.050 ;
        RECT 914.400 354.450 915.450 365.400 ;
        RECT 925.950 355.950 928.050 358.050 ;
        RECT 914.400 353.400 918.450 354.450 ;
        RECT 913.950 349.950 916.050 352.050 ;
        RECT 910.950 346.950 913.050 349.050 ;
        RECT 907.950 343.950 910.050 346.050 ;
        RECT 889.950 337.950 892.050 340.050 ;
        RECT 895.950 338.100 898.050 340.200 ;
        RECT 901.950 338.100 904.050 340.200 ;
        RECT 896.400 337.350 897.600 338.100 ;
        RECT 902.400 337.350 903.600 338.100 ;
        RECT 892.950 334.950 895.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 901.950 334.950 904.050 337.050 ;
        RECT 889.950 331.950 892.050 334.050 ;
        RECT 893.400 332.400 894.600 334.650 ;
        RECT 899.400 333.900 900.600 334.650 ;
        RECT 886.950 307.950 889.050 310.050 ;
        RECT 890.400 301.050 891.450 331.950 ;
        RECT 893.400 307.050 894.450 332.400 ;
        RECT 898.950 331.800 901.050 333.900 ;
        RECT 904.950 331.950 907.050 334.050 ;
        RECT 895.950 328.950 898.050 331.050 ;
        RECT 892.950 304.950 895.050 307.050 ;
        RECT 889.950 298.950 892.050 301.050 ;
        RECT 877.950 292.950 880.050 295.050 ;
        RECT 883.950 294.000 886.050 298.050 ;
        RECT 896.400 295.200 897.450 328.950 ;
        RECT 905.400 325.050 906.450 331.950 ;
        RECT 904.950 322.950 907.050 325.050 ;
        RECT 901.950 298.950 904.050 301.050 ;
        RECT 884.400 292.350 885.600 294.000 ;
        RECT 889.950 293.100 892.050 295.200 ;
        RECT 895.950 293.100 898.050 295.200 ;
        RECT 902.400 294.600 903.450 298.950 ;
        RECT 908.400 298.050 909.450 343.950 ;
        RECT 911.400 333.900 912.450 346.950 ;
        RECT 914.400 340.050 915.450 349.950 ;
        RECT 917.400 343.050 918.450 353.400 ;
        RECT 919.950 343.950 922.050 346.050 ;
        RECT 916.950 340.950 919.050 343.050 ;
        RECT 913.950 337.950 916.050 340.050 ;
        RECT 920.400 339.600 921.450 343.950 ;
        RECT 926.400 339.600 927.450 355.950 ;
        RECT 932.400 352.050 933.450 409.950 ;
        RECT 931.950 349.950 934.050 352.050 ;
        RECT 931.950 343.950 934.050 346.050 ;
        RECT 920.400 337.350 921.600 339.600 ;
        RECT 926.400 337.350 927.600 339.600 ;
        RECT 916.950 334.950 919.050 337.050 ;
        RECT 919.950 334.950 922.050 337.050 ;
        RECT 922.950 334.950 925.050 337.050 ;
        RECT 925.950 334.950 928.050 337.050 ;
        RECT 910.950 331.800 913.050 333.900 ;
        RECT 913.950 331.950 916.050 334.050 ;
        RECT 917.400 333.900 918.600 334.650 ;
        RECT 923.400 333.900 924.600 334.650 ;
        RECT 907.950 295.950 910.050 298.050 ;
        RECT 908.400 294.600 909.450 295.950 ;
        RECT 914.400 295.050 915.450 331.950 ;
        RECT 916.950 331.800 919.050 333.900 ;
        RECT 922.950 331.800 925.050 333.900 ;
        RECT 916.950 307.950 919.050 310.050 ;
        RECT 890.400 292.350 891.600 293.100 ;
        RECT 880.950 289.950 883.050 292.050 ;
        RECT 883.950 289.950 886.050 292.050 ;
        RECT 886.950 289.950 889.050 292.050 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 881.400 287.400 882.600 289.650 ;
        RECT 887.400 288.900 888.600 289.650 ;
        RECT 896.400 288.900 897.450 293.100 ;
        RECT 902.400 292.350 903.600 294.600 ;
        RECT 908.400 292.350 909.600 294.600 ;
        RECT 913.950 292.950 916.050 295.050 ;
        RECT 901.950 289.950 904.050 292.050 ;
        RECT 904.950 289.950 907.050 292.050 ;
        RECT 907.950 289.950 910.050 292.050 ;
        RECT 910.950 289.950 913.050 292.050 ;
        RECT 905.400 288.900 906.600 289.650 ;
        RECT 874.950 265.950 877.050 268.050 ;
        RECT 869.400 259.350 870.600 261.600 ;
        RECT 874.950 261.000 877.050 264.900 ;
        RECT 881.400 262.050 882.450 287.400 ;
        RECT 886.950 286.800 889.050 288.900 ;
        RECT 895.950 286.800 898.050 288.900 ;
        RECT 904.950 286.800 907.050 288.900 ;
        RECT 911.400 287.400 912.600 289.650 ;
        RECT 883.950 277.950 886.050 280.050 ;
        RECT 898.950 277.950 901.050 280.050 ;
        RECT 875.400 259.350 876.600 261.000 ;
        RECT 880.950 259.950 883.050 262.050 ;
        RECT 868.950 256.950 871.050 259.050 ;
        RECT 871.950 256.950 874.050 259.050 ;
        RECT 874.950 256.950 877.050 259.050 ;
        RECT 877.950 256.950 880.050 259.050 ;
        RECT 872.400 255.900 873.600 256.650 ;
        RECT 871.950 253.800 874.050 255.900 ;
        RECT 878.400 254.400 879.600 256.650 ;
        RECT 865.950 252.450 868.050 253.050 ;
        RECT 871.950 252.450 874.050 252.750 ;
        RECT 865.950 251.400 874.050 252.450 ;
        RECT 865.950 250.950 868.050 251.400 ;
        RECT 871.950 250.650 874.050 251.400 ;
        RECT 878.400 250.050 879.450 254.400 ;
        RECT 880.950 253.950 883.050 256.050 ;
        RECT 877.950 247.950 880.050 250.050 ;
        RECT 877.950 244.800 880.050 246.900 ;
        RECT 862.950 226.950 865.050 229.050 ;
        RECT 863.400 219.450 864.450 226.950 ;
        RECT 863.400 218.400 867.450 219.450 ;
        RECT 859.950 214.950 862.050 217.050 ;
        RECT 866.400 216.600 867.450 218.400 ;
        RECT 873.000 216.600 877.050 217.050 ;
        RECT 866.400 214.350 867.600 216.600 ;
        RECT 872.400 214.950 877.050 216.600 ;
        RECT 872.400 214.350 873.600 214.950 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 871.950 211.950 874.050 214.050 ;
        RECT 863.400 210.900 864.600 211.650 ;
        RECT 869.400 210.900 870.600 211.650 ;
        RECT 862.950 208.800 865.050 210.900 ;
        RECT 868.950 208.800 871.050 210.900 ;
        RECT 874.950 208.950 877.050 211.050 ;
        RECT 871.950 205.950 874.050 208.050 ;
        RECT 862.950 199.950 865.050 202.050 ;
        RECT 856.950 196.950 859.050 199.050 ;
        RECT 859.950 193.950 862.050 196.050 ;
        RECT 856.950 187.950 859.050 190.050 ;
        RECT 857.400 183.600 858.450 187.950 ;
        RECT 860.400 184.050 861.450 193.950 ;
        RECT 851.400 181.350 852.600 183.600 ;
        RECT 857.400 181.350 858.600 183.600 ;
        RECT 859.950 181.950 862.050 184.050 ;
        RECT 847.950 178.950 850.050 181.050 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 856.950 178.950 859.050 181.050 ;
        RECT 848.400 177.900 849.600 178.650 ;
        RECT 847.950 175.800 850.050 177.900 ;
        RECT 854.400 177.000 855.600 178.650 ;
        RECT 853.950 172.950 856.050 177.000 ;
        RECT 853.950 160.950 856.050 163.050 ;
        RECT 844.950 142.950 847.050 145.050 ;
        RECT 841.950 139.950 844.050 142.050 ;
        RECT 845.400 138.600 846.450 142.950 ;
        RECT 850.950 139.950 853.050 142.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 817.950 133.950 820.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 823.950 133.950 826.050 136.050 ;
        RECT 818.400 132.900 819.600 133.650 ;
        RECT 817.950 130.800 820.050 132.900 ;
        RECT 824.400 131.400 825.600 133.650 ;
        RECT 814.950 115.950 817.050 118.050 ;
        RECT 808.950 106.950 811.050 109.050 ;
        RECT 815.400 105.600 816.450 115.950 ;
        RECT 824.400 111.450 825.450 131.400 ;
        RECT 824.400 110.400 828.450 111.450 ;
        RECT 823.950 106.950 826.050 109.050 ;
        RECT 809.400 105.450 810.600 105.600 ;
        RECT 803.400 104.400 810.600 105.450 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 788.400 99.000 789.600 100.650 ;
        RECT 794.400 99.900 795.600 100.650 ;
        RECT 787.950 94.950 790.050 99.000 ;
        RECT 793.950 97.800 796.050 99.900 ;
        RECT 799.950 97.950 802.050 100.050 ;
        RECT 796.950 76.950 799.050 79.050 ;
        RECT 782.400 62.400 786.450 63.450 ;
        RECT 785.400 60.600 786.450 62.400 ;
        RECT 785.400 58.350 786.600 60.600 ;
        RECT 790.950 60.000 793.050 64.050 ;
        RECT 791.400 58.350 792.600 60.000 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 782.400 53.400 783.600 55.650 ;
        RECT 788.400 54.900 789.600 55.650 ;
        RECT 797.400 55.050 798.450 76.950 ;
        RECT 800.400 64.050 801.450 97.950 ;
        RECT 799.950 61.950 802.050 64.050 ;
        RECT 803.400 60.450 804.450 104.400 ;
        RECT 809.400 103.350 810.600 104.400 ;
        RECT 815.400 103.350 816.600 105.600 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 814.950 100.950 817.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 812.400 98.400 813.600 100.650 ;
        RECT 818.400 99.900 819.600 100.650 ;
        RECT 812.400 91.050 813.450 98.400 ;
        RECT 817.950 97.800 820.050 99.900 ;
        RECT 808.950 88.950 811.050 91.050 ;
        RECT 811.950 88.950 814.050 91.050 ;
        RECT 800.400 59.400 804.450 60.450 ;
        RECT 809.400 60.600 810.450 88.950 ;
        RECT 824.400 64.050 825.450 106.950 ;
        RECT 827.400 106.050 828.450 110.400 ;
        RECT 830.400 109.050 831.450 136.950 ;
        RECT 839.400 136.350 840.600 138.600 ;
        RECT 845.400 136.350 846.600 138.600 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 844.950 133.950 847.050 136.050 ;
        RECT 836.400 133.050 837.600 133.650 ;
        RECT 832.950 131.400 837.600 133.050 ;
        RECT 842.400 131.400 843.600 133.650 ;
        RECT 832.950 130.950 837.000 131.400 ;
        RECT 842.400 127.050 843.450 131.400 ;
        RECT 844.950 127.950 847.050 130.050 ;
        RECT 841.950 124.950 844.050 127.050 ;
        RECT 832.950 115.950 835.050 118.050 ;
        RECT 829.950 106.950 832.050 109.050 ;
        RECT 826.950 103.950 829.050 106.050 ;
        RECT 833.400 105.600 834.450 115.950 ;
        RECT 833.400 103.350 834.600 105.600 ;
        RECT 838.950 104.100 841.050 106.200 ;
        RECT 839.400 103.350 840.600 104.100 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 830.400 99.900 831.600 100.650 ;
        RECT 836.400 99.900 837.600 100.650 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 835.950 97.800 838.050 99.900 ;
        RECT 830.400 88.050 831.450 97.800 ;
        RECT 829.950 85.950 832.050 88.050 ;
        RECT 836.400 73.050 837.450 97.800 ;
        RECT 845.400 94.050 846.450 127.950 ;
        RECT 851.400 105.450 852.450 139.950 ;
        RECT 854.400 133.050 855.450 160.950 ;
        RECT 863.400 157.050 864.450 199.950 ;
        RECT 872.400 199.050 873.450 205.950 ;
        RECT 871.950 196.950 874.050 199.050 ;
        RECT 865.950 193.950 868.050 196.050 ;
        RECT 866.400 190.050 867.450 193.950 ;
        RECT 865.950 187.950 868.050 190.050 ;
        RECT 865.950 181.950 868.050 186.900 ;
        RECT 872.400 183.600 873.450 196.950 ;
        RECT 875.400 187.050 876.450 208.950 ;
        RECT 878.400 196.050 879.450 244.800 ;
        RECT 881.400 217.050 882.450 253.950 ;
        RECT 884.400 220.050 885.450 277.950 ;
        RECT 886.950 265.950 889.050 268.050 ;
        RECT 887.400 223.050 888.450 265.950 ;
        RECT 892.950 260.100 895.050 262.200 ;
        RECT 899.400 261.600 900.450 277.950 ;
        RECT 911.400 262.200 912.450 287.400 ;
        RECT 917.400 268.050 918.450 307.950 ;
        RECT 932.400 298.050 933.450 343.950 ;
        RECT 925.950 295.950 928.050 298.050 ;
        RECT 931.950 295.950 934.050 298.050 ;
        RECT 916.950 265.950 919.050 268.050 ;
        RECT 893.400 259.350 894.600 260.100 ;
        RECT 899.400 259.350 900.600 261.600 ;
        RECT 910.950 261.450 913.050 262.200 ;
        RECT 908.400 260.400 913.050 261.450 ;
        RECT 892.950 256.950 895.050 259.050 ;
        RECT 895.950 256.950 898.050 259.050 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 901.950 256.950 904.050 259.050 ;
        RECT 889.950 253.950 892.050 256.050 ;
        RECT 896.400 254.400 897.600 256.650 ;
        RECT 902.400 255.900 903.600 256.650 ;
        RECT 890.400 250.050 891.450 253.950 ;
        RECT 889.950 247.950 892.050 250.050 ;
        RECT 896.400 244.050 897.450 254.400 ;
        RECT 901.950 253.800 904.050 255.900 ;
        RECT 895.950 241.950 898.050 244.050 ;
        RECT 889.950 235.950 892.050 238.050 ;
        RECT 886.950 220.950 889.050 223.050 ;
        RECT 890.400 220.050 891.450 235.950 ;
        RECT 898.950 232.950 901.050 235.050 ;
        RECT 892.950 226.950 895.050 229.050 ;
        RECT 893.400 220.200 894.450 226.950 ;
        RECT 883.950 217.950 886.050 220.050 ;
        RECT 880.950 214.950 883.050 217.050 ;
        RECT 886.950 216.000 889.050 219.900 ;
        RECT 889.950 217.950 892.050 220.050 ;
        RECT 892.950 218.100 895.050 220.200 ;
        RECT 899.400 217.050 900.450 232.950 ;
        RECT 908.400 232.050 909.450 260.400 ;
        RECT 910.950 260.100 913.050 260.400 ;
        RECT 916.950 260.100 919.050 262.200 ;
        RECT 922.950 260.100 925.050 262.200 ;
        RECT 926.400 262.050 927.450 295.950 ;
        RECT 931.950 292.800 934.050 294.900 ;
        RECT 917.400 259.350 918.600 260.100 ;
        RECT 923.400 259.350 924.600 260.100 ;
        RECT 925.950 259.950 928.050 262.050 ;
        RECT 928.950 259.950 931.050 262.050 ;
        RECT 913.950 256.950 916.050 259.050 ;
        RECT 916.950 256.950 919.050 259.050 ;
        RECT 919.950 256.950 922.050 259.050 ;
        RECT 922.950 256.950 925.050 259.050 ;
        RECT 914.400 254.400 915.600 256.650 ;
        RECT 920.400 254.400 921.600 256.650 ;
        RECT 907.950 229.950 910.050 232.050 ;
        RECT 914.400 229.050 915.450 254.400 ;
        RECT 913.950 226.950 916.050 229.050 ;
        RECT 920.400 217.200 921.450 254.400 ;
        RECT 925.950 250.950 928.050 255.900 ;
        RECT 922.950 226.950 925.050 229.050 ;
        RECT 887.400 214.350 888.600 216.000 ;
        RECT 892.950 214.950 895.050 217.050 ;
        RECT 898.950 214.950 901.050 217.050 ;
        RECT 904.950 215.100 907.050 217.200 ;
        RECT 910.950 215.100 913.050 217.200 ;
        RECT 919.950 215.100 922.050 217.200 ;
        RECT 893.400 214.350 894.600 214.950 ;
        RECT 883.950 211.950 886.050 214.050 ;
        RECT 886.950 211.950 889.050 214.050 ;
        RECT 889.950 211.950 892.050 214.050 ;
        RECT 892.950 211.950 895.050 214.050 ;
        RECT 880.950 208.950 883.050 211.050 ;
        RECT 884.400 210.000 885.600 211.650 ;
        RECT 877.950 193.950 880.050 196.050 ;
        RECT 874.950 184.950 877.050 187.050 ;
        RECT 878.400 183.600 879.450 193.950 ;
        RECT 872.400 181.350 873.600 183.600 ;
        RECT 878.400 181.350 879.600 183.600 ;
        RECT 881.400 183.450 882.450 208.950 ;
        RECT 883.950 205.950 886.050 210.000 ;
        RECT 890.400 209.400 891.600 211.650 ;
        RECT 890.400 207.450 891.450 209.400 ;
        RECT 895.950 208.950 898.050 211.050 ;
        RECT 887.400 206.400 891.450 207.450 ;
        RECT 887.400 199.050 888.450 206.400 ;
        RECT 889.950 199.950 892.050 202.050 ;
        RECT 886.950 196.950 889.050 199.050 ;
        RECT 886.950 193.800 889.050 195.900 ;
        RECT 887.400 184.050 888.450 193.800 ;
        RECT 881.400 182.400 885.450 183.450 ;
        RECT 868.950 178.950 871.050 181.050 ;
        RECT 871.950 178.950 874.050 181.050 ;
        RECT 874.950 178.950 877.050 181.050 ;
        RECT 877.950 178.950 880.050 181.050 ;
        RECT 869.400 177.900 870.600 178.650 ;
        RECT 868.950 175.800 871.050 177.900 ;
        RECT 875.400 177.000 876.600 178.650 ;
        RECT 874.950 172.950 877.050 177.000 ;
        RECT 875.400 169.050 876.450 172.950 ;
        RECT 874.950 166.950 877.050 169.050 ;
        RECT 884.400 160.050 885.450 182.400 ;
        RECT 886.950 181.950 889.050 184.050 ;
        RECT 890.400 183.600 891.450 199.950 ;
        RECT 896.400 193.050 897.450 208.950 ;
        RECT 899.400 205.050 900.450 214.950 ;
        RECT 905.400 214.350 906.600 215.100 ;
        RECT 911.400 214.350 912.600 215.100 ;
        RECT 904.950 211.950 907.050 214.050 ;
        RECT 907.950 211.950 910.050 214.050 ;
        RECT 910.950 211.950 913.050 214.050 ;
        RECT 913.950 211.950 916.050 214.050 ;
        RECT 908.400 210.900 909.600 211.650 ;
        RECT 907.950 208.800 910.050 210.900 ;
        RECT 914.400 209.400 915.600 211.650 ;
        RECT 898.950 202.950 901.050 205.050 ;
        RECT 895.950 190.950 898.050 193.050 ;
        RECT 896.400 183.600 897.450 190.950 ;
        RECT 890.400 181.350 891.600 183.600 ;
        RECT 896.400 181.350 897.600 183.600 ;
        RECT 908.400 183.450 909.450 208.800 ;
        RECT 910.950 205.950 913.050 208.050 ;
        RECT 911.400 187.050 912.450 205.950 ;
        RECT 914.400 205.050 915.450 209.400 ;
        RECT 913.950 202.950 916.050 205.050 ;
        RECT 920.400 187.050 921.450 215.100 ;
        RECT 923.400 208.050 924.450 226.950 ;
        RECT 922.950 205.950 925.050 208.050 ;
        RECT 905.400 182.400 909.450 183.450 ;
        RECT 910.950 183.000 913.050 187.050 ;
        RECT 919.950 184.950 922.050 187.050 ;
        RECT 889.950 178.950 892.050 181.050 ;
        RECT 892.950 178.950 895.050 181.050 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 898.950 178.950 901.050 181.050 ;
        RECT 886.950 175.950 889.050 178.050 ;
        RECT 893.400 176.400 894.600 178.650 ;
        RECT 899.400 177.900 900.600 178.650 ;
        RECT 905.400 177.900 906.450 182.400 ;
        RECT 911.400 181.350 912.600 183.000 ;
        RECT 916.950 182.100 919.050 184.200 ;
        RECT 917.400 181.350 918.600 182.100 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 913.950 178.950 916.050 181.050 ;
        RECT 916.950 178.950 919.050 181.050 ;
        RECT 919.950 178.950 922.050 181.050 ;
        RECT 887.400 172.050 888.450 175.950 ;
        RECT 886.950 169.950 889.050 172.050 ;
        RECT 893.400 169.050 894.450 176.400 ;
        RECT 898.950 175.800 901.050 177.900 ;
        RECT 904.800 175.800 906.900 177.900 ;
        RECT 907.950 175.950 910.050 178.050 ;
        RECT 914.400 176.400 915.600 178.650 ;
        RECT 920.400 177.900 921.600 178.650 ;
        RECT 892.950 166.950 895.050 169.050 ;
        RECT 883.950 157.950 886.050 160.050 ;
        RECT 862.950 154.950 865.050 157.050 ;
        RECT 883.950 154.800 886.050 156.900 ;
        RECT 868.950 145.950 871.050 148.050 ;
        RECT 874.950 145.950 877.050 148.050 ;
        RECT 856.950 142.950 859.050 145.050 ;
        RECT 857.400 139.200 858.450 142.950 ;
        RECT 856.950 137.100 859.050 139.200 ;
        RECT 862.950 137.100 865.050 139.200 ;
        RECT 869.400 138.600 870.450 145.950 ;
        RECT 871.950 142.950 874.050 145.050 ;
        RECT 872.400 139.050 873.450 142.950 ;
        RECT 863.400 136.350 864.600 137.100 ;
        RECT 869.400 136.350 870.600 138.600 ;
        RECT 871.950 136.950 874.050 139.050 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 862.950 133.950 865.050 136.050 ;
        RECT 865.950 133.950 868.050 136.050 ;
        RECT 868.950 133.950 871.050 136.050 ;
        RECT 853.950 130.950 856.050 133.050 ;
        RECT 860.400 132.900 861.600 133.650 ;
        RECT 859.950 130.800 862.050 132.900 ;
        RECT 866.400 131.400 867.600 133.650 ;
        RECT 862.950 127.950 865.050 130.050 ;
        RECT 856.950 115.950 859.050 118.050 ;
        RECT 848.400 104.400 852.450 105.450 ;
        RECT 857.400 105.600 858.450 115.950 ;
        RECT 863.400 105.600 864.450 127.950 ;
        RECT 866.400 127.050 867.450 131.400 ;
        RECT 875.400 130.050 876.450 145.950 ;
        RECT 884.400 139.200 885.450 154.800 ;
        RECT 889.950 145.950 892.050 148.050 ;
        RECT 883.950 137.100 886.050 139.200 ;
        RECT 890.400 138.600 891.450 145.950 ;
        RECT 908.400 141.450 909.450 175.950 ;
        RECT 914.400 172.050 915.450 176.400 ;
        RECT 919.950 175.800 922.050 177.900 ;
        RECT 913.950 169.950 916.050 172.050 ;
        RECT 913.950 157.950 916.050 160.050 ;
        RECT 910.950 145.950 913.050 148.050 ;
        RECT 905.400 140.400 909.450 141.450 ;
        RECT 905.400 139.200 906.450 140.400 ;
        RECT 884.400 136.350 885.600 137.100 ;
        RECT 890.400 136.350 891.600 138.600 ;
        RECT 895.950 136.950 898.050 139.050 ;
        RECT 904.950 137.100 907.050 139.200 ;
        RECT 911.400 138.600 912.450 145.950 ;
        RECT 914.400 139.050 915.450 157.950 ;
        RECT 880.950 133.950 883.050 136.050 ;
        RECT 883.950 133.950 886.050 136.050 ;
        RECT 886.950 133.950 889.050 136.050 ;
        RECT 889.950 133.950 892.050 136.050 ;
        RECT 881.400 133.050 882.600 133.650 ;
        RECT 877.950 131.400 882.600 133.050 ;
        RECT 887.400 131.400 888.600 133.650 ;
        RECT 877.950 130.950 882.000 131.400 ;
        RECT 874.950 129.450 877.050 130.050 ;
        RECT 872.400 128.400 877.050 129.450 ;
        RECT 865.950 124.950 868.050 127.050 ;
        RECT 866.400 112.050 867.450 124.950 ;
        RECT 865.950 109.950 868.050 112.050 ;
        RECT 844.950 91.950 847.050 94.050 ;
        RECT 838.950 88.950 841.050 91.050 ;
        RECT 835.950 70.950 838.050 73.050 ;
        RECT 782.400 43.050 783.450 53.400 ;
        RECT 787.950 52.800 790.050 54.900 ;
        RECT 796.950 52.950 799.050 55.050 ;
        RECT 800.400 52.050 801.450 59.400 ;
        RECT 809.400 58.350 810.600 60.600 ;
        RECT 814.950 60.000 817.050 64.050 ;
        RECT 823.950 61.950 826.050 64.050 ;
        RECT 826.950 61.950 829.050 64.050 ;
        RECT 815.400 58.350 816.600 60.000 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 811.950 55.950 814.050 58.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 806.400 54.000 807.600 55.650 ;
        RECT 799.950 49.950 802.050 52.050 ;
        RECT 805.950 49.950 808.050 54.000 ;
        RECT 812.400 53.400 813.600 55.650 ;
        RECT 775.950 40.950 778.050 43.050 ;
        RECT 781.950 40.950 784.050 43.050 ;
        RECT 793.950 40.950 796.050 43.050 ;
        RECT 772.950 28.950 775.050 31.050 ;
        RECT 770.400 25.350 771.600 27.600 ;
        RECT 775.950 26.100 778.050 28.200 ;
        RECT 776.400 25.350 777.600 26.100 ;
        RECT 784.950 25.950 787.050 28.050 ;
        RECT 794.400 27.600 795.450 40.950 ;
        RECT 812.400 40.050 813.450 53.400 ;
        RECT 824.400 52.050 825.450 61.950 ;
        RECT 817.950 49.950 823.050 52.050 ;
        RECT 823.950 49.950 826.050 52.050 ;
        RECT 811.950 37.950 814.050 40.050 ;
        RECT 802.950 31.950 805.050 34.050 ;
        RECT 814.950 31.950 817.050 34.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 767.400 21.900 768.600 22.650 ;
        RECT 743.400 16.050 744.450 20.400 ;
        RECT 752.400 19.050 753.450 20.400 ;
        RECT 760.950 19.800 763.050 21.900 ;
        RECT 766.950 19.800 769.050 21.900 ;
        RECT 773.400 21.000 774.600 22.650 ;
        RECT 785.400 21.900 786.450 25.950 ;
        RECT 794.400 25.350 795.600 27.600 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 791.400 21.900 792.600 22.650 ;
        RECT 797.400 21.900 798.600 22.650 ;
        RECT 803.400 21.900 804.450 31.950 ;
        RECT 815.400 27.600 816.450 31.950 ;
        RECT 820.950 28.950 823.050 31.050 ;
        RECT 815.400 25.350 816.600 27.600 ;
        RECT 809.100 22.950 811.200 25.050 ;
        RECT 814.500 22.950 816.600 25.050 ;
        RECT 817.800 22.950 819.900 25.050 ;
        RECT 752.400 17.400 757.050 19.050 ;
        RECT 753.000 16.950 757.050 17.400 ;
        RECT 772.950 16.950 775.050 21.000 ;
        RECT 784.950 19.800 787.050 21.900 ;
        RECT 790.950 16.950 793.050 21.900 ;
        RECT 796.950 19.800 799.050 21.900 ;
        RECT 802.950 19.800 805.050 21.900 ;
        RECT 809.400 21.000 810.600 22.650 ;
        RECT 818.400 21.450 819.600 22.650 ;
        RECT 821.400 21.450 822.450 28.950 ;
        RECT 827.400 25.050 828.450 61.950 ;
        RECT 839.400 60.600 840.450 88.950 ;
        RECT 848.400 82.050 849.450 104.400 ;
        RECT 857.400 103.350 858.600 105.600 ;
        RECT 863.400 103.350 864.600 105.600 ;
        RECT 868.950 103.950 871.050 106.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 854.400 99.900 855.600 100.650 ;
        RECT 853.950 97.800 856.050 99.900 ;
        RECT 860.400 98.400 861.600 100.650 ;
        RECT 869.400 99.900 870.450 103.950 ;
        RECT 860.400 88.050 861.450 98.400 ;
        RECT 868.950 97.800 871.050 99.900 ;
        RECT 869.400 88.050 870.450 97.800 ;
        RECT 859.950 85.950 862.050 88.050 ;
        RECT 868.950 85.950 871.050 88.050 ;
        RECT 847.950 79.950 850.050 82.050 ;
        RECT 856.950 79.950 859.050 82.050 ;
        RECT 853.950 73.950 856.050 76.050 ;
        RECT 847.950 70.950 850.050 73.050 ;
        RECT 848.400 60.600 849.450 70.950 ;
        RECT 839.400 58.350 840.600 60.600 ;
        RECT 848.400 58.350 849.600 60.600 ;
        RECT 850.950 59.100 853.050 61.200 ;
        RECT 832.800 55.950 834.900 58.050 ;
        RECT 838.950 55.950 841.050 58.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 847.500 55.950 849.600 58.050 ;
        RECT 833.400 54.000 834.600 55.650 ;
        RECT 842.400 54.000 843.600 55.650 ;
        RECT 832.950 49.950 835.050 54.000 ;
        RECT 841.950 49.950 844.050 54.000 ;
        RECT 851.400 51.450 852.450 59.100 ;
        RECT 854.400 55.050 855.450 73.950 ;
        RECT 853.950 52.950 856.050 55.050 ;
        RECT 848.400 50.400 852.450 51.450 ;
        RECT 841.950 37.950 844.050 40.050 ;
        RECT 835.950 31.950 838.050 34.050 ;
        RECT 836.400 27.600 837.450 31.950 ;
        RECT 842.400 27.600 843.450 37.950 ;
        RECT 848.400 31.050 849.450 50.400 ;
        RECT 853.950 49.800 856.050 51.900 ;
        RECT 854.400 46.050 855.450 49.800 ;
        RECT 857.400 49.050 858.450 79.950 ;
        RECT 872.400 76.050 873.450 128.400 ;
        RECT 874.950 127.950 877.050 128.400 ;
        RECT 880.950 127.950 883.050 130.050 ;
        RECT 877.950 115.950 880.050 118.050 ;
        RECT 878.400 105.600 879.450 115.950 ;
        RECT 881.400 112.050 882.450 127.950 ;
        RECT 887.400 124.050 888.450 131.400 ;
        RECT 886.950 121.950 889.050 124.050 ;
        RECT 892.950 115.950 895.050 118.050 ;
        RECT 883.950 112.950 886.050 115.050 ;
        RECT 880.950 109.950 883.050 112.050 ;
        RECT 884.400 105.600 885.450 112.950 ;
        RECT 889.950 109.950 892.050 112.050 ;
        RECT 890.400 106.050 891.450 109.950 ;
        RECT 893.400 106.200 894.450 115.950 ;
        RECT 896.400 112.050 897.450 136.950 ;
        RECT 905.400 136.350 906.600 137.100 ;
        RECT 911.400 136.350 912.600 138.600 ;
        RECT 913.950 136.950 916.050 139.050 ;
        RECT 901.950 133.950 904.050 136.050 ;
        RECT 904.950 133.950 907.050 136.050 ;
        RECT 907.950 133.950 910.050 136.050 ;
        RECT 910.950 133.950 913.050 136.050 ;
        RECT 902.400 131.400 903.600 133.650 ;
        RECT 908.400 132.000 909.600 133.650 ;
        RECT 898.950 127.950 901.050 130.050 ;
        RECT 899.400 118.050 900.450 127.950 ;
        RECT 898.950 115.950 901.050 118.050 ;
        RECT 895.950 109.950 898.050 112.050 ;
        RECT 902.400 108.450 903.450 131.400 ;
        RECT 904.950 127.950 907.050 130.050 ;
        RECT 907.950 127.950 910.050 132.000 ;
        RECT 913.950 130.950 916.050 133.050 ;
        RECT 905.400 109.050 906.450 127.950 ;
        RECT 908.400 124.050 909.450 127.950 ;
        RECT 907.950 121.950 910.050 124.050 ;
        RECT 907.950 115.950 910.050 118.050 ;
        RECT 899.400 107.400 903.450 108.450 ;
        RECT 878.400 103.350 879.600 105.600 ;
        RECT 884.400 103.350 885.600 105.600 ;
        RECT 889.800 103.950 891.900 106.050 ;
        RECT 892.950 104.100 895.050 106.200 ;
        RECT 899.400 105.450 900.450 107.400 ;
        RECT 904.950 106.950 907.050 109.050 ;
        RECT 896.400 104.400 900.450 105.450 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 880.950 100.950 883.050 103.050 ;
        RECT 883.950 100.950 886.050 103.050 ;
        RECT 886.950 100.950 889.050 103.050 ;
        RECT 881.400 99.900 882.600 100.650 ;
        RECT 887.400 99.900 888.600 100.650 ;
        RECT 880.950 97.800 883.050 99.900 ;
        RECT 886.950 97.800 889.050 99.900 ;
        RECT 889.950 97.950 892.050 100.050 ;
        RECT 874.950 91.950 877.050 94.050 ;
        RECT 880.950 91.950 883.050 94.050 ;
        RECT 875.400 76.050 876.450 91.950 ;
        RECT 871.950 73.950 874.050 76.050 ;
        RECT 874.950 73.950 877.050 76.050 ;
        RECT 877.950 73.950 880.050 76.050 ;
        RECT 874.950 70.800 877.050 72.900 ;
        RECT 868.950 62.100 871.050 67.050 ;
        RECT 862.950 59.100 865.050 61.200 ;
        RECT 875.400 61.050 876.450 70.800 ;
        RECT 863.400 58.350 864.600 59.100 ;
        RECT 868.950 58.950 871.050 61.050 ;
        RECT 874.950 58.950 877.050 61.050 ;
        RECT 869.400 58.350 870.600 58.950 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 859.950 52.950 862.050 55.050 ;
        RECT 866.400 53.400 867.600 55.650 ;
        RECT 872.400 54.450 873.600 55.650 ;
        RECT 872.400 53.400 876.450 54.450 ;
        RECT 856.950 46.950 859.050 49.050 ;
        RECT 860.400 46.050 861.450 52.950 ;
        RECT 853.950 43.950 856.050 46.050 ;
        RECT 859.950 43.950 862.050 46.050 ;
        RECT 856.950 37.950 859.050 40.050 ;
        RECT 850.950 34.950 853.050 37.050 ;
        RECT 847.950 28.950 850.050 31.050 ;
        RECT 836.400 25.350 837.600 27.600 ;
        RECT 842.400 25.350 843.600 27.600 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 832.950 22.950 835.050 25.050 ;
        RECT 835.950 22.950 838.050 25.050 ;
        RECT 838.950 22.950 841.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 808.950 16.950 811.050 21.000 ;
        RECT 818.400 20.400 822.450 21.450 ;
        RECT 833.400 21.000 834.600 22.650 ;
        RECT 832.950 16.950 835.050 21.000 ;
        RECT 839.400 20.400 840.600 22.650 ;
        RECT 845.400 21.900 846.600 22.650 ;
        RECT 851.400 21.900 852.450 34.950 ;
        RECT 857.400 31.050 858.450 37.950 ;
        RECT 866.400 37.050 867.450 53.400 ;
        RECT 871.950 49.950 874.050 52.050 ;
        RECT 868.950 37.950 871.050 40.050 ;
        RECT 865.950 34.950 868.050 37.050 ;
        RECT 856.950 28.950 859.050 31.050 ;
        RECT 859.950 26.100 862.050 28.200 ;
        RECT 865.950 27.000 868.050 31.050 ;
        RECT 869.400 28.050 870.450 37.950 ;
        RECT 860.400 25.350 861.600 26.100 ;
        RECT 866.400 25.350 867.600 27.000 ;
        RECT 868.950 25.950 871.050 28.050 ;
        RECT 856.950 22.950 859.050 25.050 ;
        RECT 859.950 22.950 862.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 857.400 21.900 858.600 22.650 ;
        RECT 863.400 21.900 864.600 22.650 ;
        RECT 839.400 16.050 840.450 20.400 ;
        RECT 844.950 19.800 847.050 21.900 ;
        RECT 850.950 19.800 853.050 21.900 ;
        RECT 856.950 19.800 859.050 21.900 ;
        RECT 862.950 19.800 865.050 21.900 ;
        RECT 872.400 16.050 873.450 49.950 ;
        RECT 875.400 46.050 876.450 53.400 ;
        RECT 874.950 43.950 877.050 46.050 ;
        RECT 874.950 34.950 877.050 37.050 ;
        RECT 875.400 31.050 876.450 34.950 ;
        RECT 874.950 28.950 877.050 31.050 ;
        RECT 878.400 27.450 879.450 73.950 ;
        RECT 881.400 52.050 882.450 91.950 ;
        RECT 883.950 73.950 886.050 76.050 ;
        RECT 884.400 70.050 885.450 73.950 ;
        RECT 883.950 67.950 886.050 70.050 ;
        RECT 890.400 60.600 891.450 97.950 ;
        RECT 893.400 94.050 894.450 104.100 ;
        RECT 896.400 100.050 897.450 104.400 ;
        RECT 901.950 104.100 904.050 106.200 ;
        RECT 908.400 105.600 909.450 115.950 ;
        RECT 902.400 103.350 903.600 104.100 ;
        RECT 908.400 103.350 909.600 105.600 ;
        RECT 914.400 105.450 915.450 130.950 ;
        RECT 914.400 104.400 918.450 105.450 ;
        RECT 901.950 100.950 904.050 103.050 ;
        RECT 904.950 100.950 907.050 103.050 ;
        RECT 907.950 100.950 910.050 103.050 ;
        RECT 910.950 100.950 913.050 103.050 ;
        RECT 895.950 97.950 898.050 100.050 ;
        RECT 905.400 98.400 906.600 100.650 ;
        RECT 911.400 99.900 912.600 100.650 ;
        RECT 895.950 94.800 898.050 96.900 ;
        RECT 901.950 94.950 904.050 97.050 ;
        RECT 892.950 91.950 895.050 94.050 ;
        RECT 896.400 61.200 897.450 94.800 ;
        RECT 898.950 67.950 901.050 70.050 ;
        RECT 890.400 58.350 891.600 60.600 ;
        RECT 895.950 59.100 898.050 61.200 ;
        RECT 899.400 61.050 900.450 67.950 ;
        RECT 896.400 58.350 897.600 59.100 ;
        RECT 898.950 58.950 901.050 61.050 ;
        RECT 886.950 55.950 889.050 58.050 ;
        RECT 889.950 55.950 892.050 58.050 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 887.400 53.400 888.600 55.650 ;
        RECT 893.400 54.900 894.600 55.650 ;
        RECT 880.950 49.950 883.050 52.050 ;
        RECT 883.950 34.950 886.050 37.050 ;
        RECT 875.400 26.400 879.450 27.450 ;
        RECT 884.400 27.600 885.450 34.950 ;
        RECT 887.400 31.050 888.450 53.400 ;
        RECT 892.950 52.800 895.050 54.900 ;
        RECT 889.950 49.950 892.050 52.050 ;
        RECT 886.950 28.950 889.050 31.050 ;
        RECT 890.400 27.600 891.450 49.950 ;
        RECT 895.950 46.950 898.050 49.050 ;
        RECT 875.400 21.900 876.450 26.400 ;
        RECT 884.400 25.350 885.600 27.600 ;
        RECT 890.400 25.350 891.600 27.600 ;
        RECT 880.950 22.950 883.050 25.050 ;
        RECT 883.950 22.950 886.050 25.050 ;
        RECT 886.950 22.950 889.050 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 881.400 21.900 882.600 22.650 ;
        RECT 887.400 21.900 888.600 22.650 ;
        RECT 874.950 19.800 877.050 21.900 ;
        RECT 880.950 19.800 883.050 21.900 ;
        RECT 886.950 19.800 889.050 21.900 ;
        RECT 742.950 13.950 745.050 16.050 ;
        RECT 838.950 13.950 841.050 16.050 ;
        RECT 871.950 13.950 874.050 16.050 ;
        RECT 896.400 10.050 897.450 46.950 ;
        RECT 902.400 30.450 903.450 94.950 ;
        RECT 905.400 88.050 906.450 98.400 ;
        RECT 910.950 94.950 913.050 99.900 ;
        RECT 904.950 85.950 907.050 88.050 ;
        RECT 917.400 70.050 918.450 104.400 ;
        RECT 907.950 67.950 910.050 70.050 ;
        RECT 916.950 67.950 919.050 70.050 ;
        RECT 904.950 64.950 907.050 67.050 ;
        RECT 905.400 61.050 906.450 64.950 ;
        RECT 904.950 58.950 907.050 61.050 ;
        RECT 908.400 60.600 909.450 67.950 ;
        RECT 908.400 58.350 909.600 60.600 ;
        RECT 913.950 60.000 916.050 64.050 ;
        RECT 920.400 61.050 921.450 175.800 ;
        RECT 922.950 127.950 925.050 130.050 ;
        RECT 914.400 58.350 915.600 60.000 ;
        RECT 919.950 58.950 922.050 61.050 ;
        RECT 907.950 55.950 910.050 58.050 ;
        RECT 910.950 55.950 913.050 58.050 ;
        RECT 913.950 55.950 916.050 58.050 ;
        RECT 916.950 55.950 919.050 58.050 ;
        RECT 904.950 52.950 907.050 55.050 ;
        RECT 911.400 53.400 912.600 55.650 ;
        RECT 917.400 54.900 918.600 55.650 ;
        RECT 899.400 29.400 903.450 30.450 ;
        RECT 899.400 21.900 900.450 29.400 ;
        RECT 905.400 27.600 906.450 52.950 ;
        RECT 911.400 49.050 912.450 53.400 ;
        RECT 916.950 52.800 919.050 54.900 ;
        RECT 910.950 46.950 913.050 49.050 ;
        RECT 923.400 37.050 924.450 127.950 ;
        RECT 926.400 64.050 927.450 250.950 ;
        RECT 929.400 250.050 930.450 259.950 ;
        RECT 928.950 247.950 931.050 250.050 ;
        RECT 928.950 229.950 931.050 232.050 ;
        RECT 929.400 210.900 930.450 229.950 ;
        RECT 928.950 208.800 931.050 210.900 ;
        RECT 928.950 151.950 931.050 154.050 ;
        RECT 925.950 61.950 928.050 64.050 ;
        RECT 922.950 34.950 925.050 37.050 ;
        RECT 929.400 31.050 930.450 151.950 ;
        RECT 928.950 28.950 931.050 31.050 ;
        RECT 905.400 25.350 906.600 27.600 ;
        RECT 902.100 22.950 904.200 25.050 ;
        RECT 905.400 22.950 907.500 25.050 ;
        RECT 910.800 22.950 912.900 25.050 ;
        RECT 898.950 19.800 901.050 21.900 ;
        RECT 902.400 20.400 903.600 22.650 ;
        RECT 911.400 20.400 912.600 22.650 ;
        RECT 902.400 16.050 903.450 20.400 ;
        RECT 901.950 13.950 904.050 16.050 ;
        RECT 911.400 10.050 912.450 20.400 ;
        RECT 932.400 16.050 933.450 292.800 ;
        RECT 935.400 244.050 936.450 424.950 ;
        RECT 934.950 241.950 937.050 244.050 ;
        RECT 935.400 49.050 936.450 241.950 ;
        RECT 934.950 46.950 937.050 49.050 ;
        RECT 931.950 13.950 934.050 16.050 ;
        RECT 577.950 7.950 580.050 10.050 ;
        RECT 610.950 7.950 613.050 10.050 ;
        RECT 703.950 7.950 706.050 10.050 ;
        RECT 736.950 7.950 739.050 10.050 ;
        RECT 895.950 7.950 898.050 10.050 ;
        RECT 910.950 7.950 913.050 10.050 ;
        RECT 112.950 4.950 115.050 7.050 ;
        RECT 157.950 4.950 160.050 7.050 ;
        RECT 475.950 4.950 478.050 7.050 ;
        RECT 505.950 4.950 508.050 7.050 ;
      LAYER metal3 ;
        RECT 367.950 936.600 370.050 937.050 ;
        RECT 577.950 936.600 580.050 937.050 ;
        RECT 367.950 935.400 580.050 936.600 ;
        RECT 367.950 934.950 370.050 935.400 ;
        RECT 577.950 934.950 580.050 935.400 ;
        RECT 91.950 933.600 94.050 934.050 ;
        RECT 133.950 933.600 136.050 934.050 ;
        RECT 91.950 932.400 136.050 933.600 ;
        RECT 91.950 931.950 94.050 932.400 ;
        RECT 133.950 931.950 136.050 932.400 ;
        RECT 61.950 930.600 64.050 931.050 ;
        RECT 124.950 930.600 127.050 931.050 ;
        RECT 61.950 929.400 127.050 930.600 ;
        RECT 61.950 928.950 64.050 929.400 ;
        RECT 124.950 928.950 127.050 929.400 ;
        RECT 160.950 930.600 163.050 931.050 ;
        RECT 181.950 930.600 184.050 931.050 ;
        RECT 160.950 929.400 184.050 930.600 ;
        RECT 160.950 928.950 163.050 929.400 ;
        RECT 181.950 928.950 184.050 929.400 ;
        RECT 361.950 930.600 364.050 931.050 ;
        RECT 412.950 930.600 415.050 931.050 ;
        RECT 361.950 929.400 415.050 930.600 ;
        RECT 361.950 928.950 364.050 929.400 ;
        RECT 412.950 928.950 415.050 929.400 ;
        RECT 463.950 930.600 466.050 931.050 ;
        RECT 502.950 930.600 505.050 931.050 ;
        RECT 514.950 930.600 517.050 931.050 ;
        RECT 463.950 929.400 517.050 930.600 ;
        RECT 463.950 928.950 466.050 929.400 ;
        RECT 502.950 928.950 505.050 929.400 ;
        RECT 514.950 928.950 517.050 929.400 ;
        RECT 328.950 927.600 331.050 928.050 ;
        RECT 418.950 927.600 421.050 928.050 ;
        RECT 697.950 927.600 700.050 928.050 ;
        RECT 328.950 926.400 421.050 927.600 ;
        RECT 328.950 925.950 331.050 926.400 ;
        RECT 418.950 925.950 421.050 926.400 ;
        RECT 647.400 926.400 700.050 927.600 ;
        RECT 647.400 925.050 648.600 926.400 ;
        RECT 697.950 925.950 700.050 926.400 ;
        RECT 829.950 927.600 832.050 928.050 ;
        RECT 844.950 927.600 847.050 928.050 ;
        RECT 862.950 927.600 865.050 928.050 ;
        RECT 829.950 926.400 865.050 927.600 ;
        RECT 829.950 925.950 832.050 926.400 ;
        RECT 844.950 925.950 847.050 926.400 ;
        RECT 862.950 925.950 865.050 926.400 ;
        RECT 73.950 924.600 76.050 925.050 ;
        RECT 85.950 924.600 88.050 925.050 ;
        RECT 100.950 924.600 103.050 925.050 ;
        RECT 73.950 923.400 103.050 924.600 ;
        RECT 73.950 922.950 76.050 923.400 ;
        RECT 85.950 922.950 88.050 923.400 ;
        RECT 100.950 922.950 103.050 923.400 ;
        RECT 181.950 924.600 184.050 925.050 ;
        RECT 214.950 924.600 217.050 925.050 ;
        RECT 181.950 923.400 217.050 924.600 ;
        RECT 181.950 922.950 184.050 923.400 ;
        RECT 214.950 922.950 217.050 923.400 ;
        RECT 229.950 924.600 232.050 925.050 ;
        RECT 322.950 924.600 325.050 925.050 ;
        RECT 229.950 923.400 325.050 924.600 ;
        RECT 229.950 922.950 232.050 923.400 ;
        RECT 322.950 922.950 325.050 923.400 ;
        RECT 424.950 924.600 427.050 925.050 ;
        RECT 472.950 924.600 475.050 925.050 ;
        RECT 496.950 924.600 499.050 925.050 ;
        RECT 424.950 923.400 441.600 924.600 ;
        RECT 424.950 922.950 427.050 923.400 ;
        RECT 34.950 921.600 37.050 922.050 ;
        RECT 46.950 921.600 49.050 922.050 ;
        RECT 34.950 920.400 49.050 921.600 ;
        RECT 34.950 919.950 37.050 920.400 ;
        RECT 46.950 919.950 49.050 920.400 ;
        RECT 313.950 921.600 316.050 922.050 ;
        RECT 346.950 921.600 349.050 922.050 ;
        RECT 385.950 921.600 388.050 922.050 ;
        RECT 421.950 921.600 424.050 922.050 ;
        RECT 313.950 920.400 424.050 921.600 ;
        RECT 440.400 921.600 441.600 923.400 ;
        RECT 472.950 923.400 499.050 924.600 ;
        RECT 472.950 922.950 475.050 923.400 ;
        RECT 496.950 922.950 499.050 923.400 ;
        RECT 622.950 924.600 625.050 925.050 ;
        RECT 646.950 924.600 649.050 925.050 ;
        RECT 622.950 923.400 649.050 924.600 ;
        RECT 622.950 922.950 625.050 923.400 ;
        RECT 646.950 922.950 649.050 923.400 ;
        RECT 682.950 924.600 685.050 925.050 ;
        RECT 712.950 924.600 715.050 925.050 ;
        RECT 682.950 923.400 715.050 924.600 ;
        RECT 682.950 922.950 685.050 923.400 ;
        RECT 712.950 922.950 715.050 923.400 ;
        RECT 718.950 924.600 721.050 925.050 ;
        RECT 751.950 924.600 754.050 925.050 ;
        RECT 769.950 924.600 772.050 925.050 ;
        RECT 718.950 923.400 772.050 924.600 ;
        RECT 718.950 922.950 721.050 923.400 ;
        RECT 751.950 922.950 754.050 923.400 ;
        RECT 769.950 922.950 772.050 923.400 ;
        RECT 778.950 924.600 781.050 925.050 ;
        RECT 784.950 924.600 787.050 925.050 ;
        RECT 778.950 923.400 787.050 924.600 ;
        RECT 778.950 922.950 781.050 923.400 ;
        RECT 784.950 922.950 787.050 923.400 ;
        RECT 790.950 924.600 793.050 925.050 ;
        RECT 850.950 924.600 853.050 925.050 ;
        RECT 790.950 923.400 853.050 924.600 ;
        RECT 790.950 922.950 793.050 923.400 ;
        RECT 850.950 922.950 853.050 923.400 ;
        RECT 868.950 924.600 871.050 925.050 ;
        RECT 928.950 924.600 931.050 925.050 ;
        RECT 868.950 923.400 931.050 924.600 ;
        RECT 868.950 922.950 871.050 923.400 ;
        RECT 928.950 922.950 931.050 923.400 ;
        RECT 565.950 921.600 568.050 922.050 ;
        RECT 571.950 921.600 574.050 922.050 ;
        RECT 440.400 920.400 450.600 921.600 ;
        RECT 313.950 919.950 316.050 920.400 ;
        RECT 346.950 919.950 349.050 920.400 ;
        RECT 385.950 919.950 388.050 920.400 ;
        RECT 421.950 919.950 424.050 920.400 ;
        RECT 16.950 917.100 19.050 919.200 ;
        RECT 22.950 918.600 25.050 919.200 ;
        RECT 34.950 918.600 37.050 919.200 ;
        RECT 22.950 917.400 37.050 918.600 ;
        RECT 22.950 917.100 25.050 917.400 ;
        RECT 34.950 917.100 37.050 917.400 ;
        RECT 40.950 917.100 43.050 919.200 ;
        RECT 67.950 917.100 70.050 919.200 ;
        RECT 97.950 918.750 100.050 919.200 ;
        RECT 109.950 918.750 112.050 919.200 ;
        RECT 97.950 917.550 112.050 918.750 ;
        RECT 97.950 917.100 100.050 917.550 ;
        RECT 109.950 917.100 112.050 917.550 ;
        RECT 133.950 917.100 136.050 919.200 ;
        RECT 139.950 918.600 142.050 919.200 ;
        RECT 154.950 918.750 157.050 919.200 ;
        RECT 169.950 918.750 172.050 919.200 ;
        RECT 154.950 918.600 172.050 918.750 ;
        RECT 139.950 917.550 172.050 918.600 ;
        RECT 139.950 917.400 157.050 917.550 ;
        RECT 139.950 917.100 142.050 917.400 ;
        RECT 154.950 917.100 157.050 917.400 ;
        RECT 169.950 917.100 172.050 917.550 ;
        RECT 175.950 917.100 178.050 919.200 ;
        RECT 190.950 918.600 193.050 919.050 ;
        RECT 229.950 918.600 232.050 919.200 ;
        RECT 190.950 917.400 232.050 918.600 ;
        RECT 17.400 912.600 18.600 917.100 ;
        RECT 41.400 912.600 42.600 917.100 ;
        RECT 68.400 915.600 69.600 917.100 ;
        RECT 68.400 914.400 72.600 915.600 ;
        RECT 49.950 912.600 52.050 913.050 ;
        RECT 17.400 911.400 52.050 912.600 ;
        RECT 71.400 912.600 72.600 914.400 ;
        RECT 76.950 912.600 79.050 913.050 ;
        RECT 134.400 912.600 135.600 917.100 ;
        RECT 157.950 912.600 160.050 912.900 ;
        RECT 71.400 911.400 79.050 912.600 ;
        RECT 49.950 910.950 52.050 911.400 ;
        RECT 76.950 910.950 79.050 911.400 ;
        RECT 122.400 911.400 160.050 912.600 ;
        RECT 19.950 909.600 22.050 910.050 ;
        RECT 43.950 909.600 46.050 910.050 ;
        RECT 19.950 908.400 46.050 909.600 ;
        RECT 19.950 907.950 22.050 908.400 ;
        RECT 43.950 907.950 46.050 908.400 ;
        RECT 112.950 909.600 115.050 910.050 ;
        RECT 115.950 909.600 118.050 910.050 ;
        RECT 122.400 909.600 123.600 911.400 ;
        RECT 157.950 910.800 160.050 911.400 ;
        RECT 163.950 912.450 166.050 912.900 ;
        RECT 172.950 912.600 175.050 912.900 ;
        RECT 176.400 912.600 177.600 917.100 ;
        RECT 190.950 916.950 193.050 917.400 ;
        RECT 229.950 917.100 232.050 917.400 ;
        RECT 238.950 918.750 241.050 919.200 ;
        RECT 247.950 918.750 250.050 919.200 ;
        RECT 238.950 917.550 250.050 918.750 ;
        RECT 238.950 917.100 241.050 917.550 ;
        RECT 247.950 917.100 250.050 917.550 ;
        RECT 262.950 918.750 265.050 919.200 ;
        RECT 268.950 918.750 271.050 919.200 ;
        RECT 262.950 917.550 271.050 918.750 ;
        RECT 262.950 917.100 265.050 917.550 ;
        RECT 268.950 917.100 271.050 917.550 ;
        RECT 274.950 917.100 277.050 919.200 ;
        RECT 292.950 918.600 295.050 919.200 ;
        RECT 298.950 918.600 301.050 919.050 ;
        RECT 292.950 917.400 301.050 918.600 ;
        RECT 292.950 917.100 295.050 917.400 ;
        RECT 172.950 912.450 177.600 912.600 ;
        RECT 163.950 911.400 177.600 912.450 ;
        RECT 184.950 912.450 187.050 912.900 ;
        RECT 187.950 912.450 190.050 913.050 ;
        RECT 190.950 912.450 193.050 912.900 ;
        RECT 163.950 911.250 175.050 911.400 ;
        RECT 163.950 910.800 166.050 911.250 ;
        RECT 172.950 910.800 175.050 911.250 ;
        RECT 184.950 911.250 193.050 912.450 ;
        RECT 184.950 910.800 187.050 911.250 ;
        RECT 187.950 910.950 190.050 911.250 ;
        RECT 190.950 910.800 193.050 911.250 ;
        RECT 211.950 912.450 214.050 912.900 ;
        RECT 238.950 912.450 241.050 912.900 ;
        RECT 211.950 911.250 241.050 912.450 ;
        RECT 211.950 910.800 214.050 911.250 ;
        RECT 238.950 910.800 241.050 911.250 ;
        RECT 250.950 912.600 253.050 912.900 ;
        RECT 262.950 912.600 265.050 913.050 ;
        RECT 250.950 911.400 265.050 912.600 ;
        RECT 275.400 912.600 276.600 917.100 ;
        RECT 298.950 916.950 301.050 917.400 ;
        RECT 334.950 918.750 337.050 919.200 ;
        RECT 340.950 918.750 343.050 919.200 ;
        RECT 334.950 917.550 343.050 918.750 ;
        RECT 334.950 917.100 337.050 917.550 ;
        RECT 340.950 917.100 343.050 917.550 ;
        RECT 352.950 918.600 355.050 919.200 ;
        RECT 367.950 918.600 370.050 919.200 ;
        RECT 352.950 917.400 370.050 918.600 ;
        RECT 352.950 917.100 355.050 917.400 ;
        RECT 367.950 917.100 370.050 917.400 ;
        RECT 373.950 918.750 376.050 919.200 ;
        RECT 379.950 918.750 382.050 919.200 ;
        RECT 373.950 917.550 382.050 918.750 ;
        RECT 373.950 917.100 376.050 917.550 ;
        RECT 379.950 917.100 382.050 917.550 ;
        RECT 424.950 918.750 427.050 919.200 ;
        RECT 430.950 918.750 433.050 919.200 ;
        RECT 424.950 917.550 433.050 918.750 ;
        RECT 424.950 917.100 427.050 917.550 ;
        RECT 430.950 917.100 433.050 917.550 ;
        RECT 436.950 918.750 439.050 919.200 ;
        RECT 445.950 918.750 448.050 919.200 ;
        RECT 436.950 917.550 448.050 918.750 ;
        RECT 436.950 917.100 439.050 917.550 ;
        RECT 445.950 917.100 448.050 917.550 ;
        RECT 295.800 912.600 297.900 913.050 ;
        RECT 275.400 911.400 297.900 912.600 ;
        RECT 250.950 910.800 253.050 911.400 ;
        RECT 262.950 910.950 265.050 911.400 ;
        RECT 295.800 910.950 297.900 911.400 ;
        RECT 298.950 912.450 301.050 912.900 ;
        RECT 310.950 912.450 313.050 912.900 ;
        RECT 298.950 911.250 313.050 912.450 ;
        RECT 298.950 910.800 301.050 911.250 ;
        RECT 310.950 910.800 313.050 911.250 ;
        RECT 340.950 912.600 343.050 913.050 ;
        RECT 370.950 912.600 373.050 912.900 ;
        RECT 340.950 911.400 373.050 912.600 ;
        RECT 340.950 910.950 343.050 911.400 ;
        RECT 370.950 910.800 373.050 911.400 ;
        RECT 379.950 912.600 382.050 913.050 ;
        RECT 388.950 912.600 391.050 912.900 ;
        RECT 379.950 911.400 391.050 912.600 ;
        RECT 379.950 910.950 382.050 911.400 ;
        RECT 388.950 910.800 391.050 911.400 ;
        RECT 400.950 912.600 403.050 913.050 ;
        RECT 409.950 912.600 412.050 912.900 ;
        RECT 400.950 911.400 412.050 912.600 ;
        RECT 400.950 910.950 403.050 911.400 ;
        RECT 409.950 910.800 412.050 911.400 ;
        RECT 421.950 912.600 424.050 913.050 ;
        RECT 433.950 912.600 436.050 912.900 ;
        RECT 421.950 911.400 436.050 912.600 ;
        RECT 449.400 912.600 450.600 920.400 ;
        RECT 565.950 920.400 574.050 921.600 ;
        RECT 565.950 919.950 568.050 920.400 ;
        RECT 571.950 919.950 574.050 920.400 ;
        RECT 457.950 917.100 460.050 919.200 ;
        RECT 478.950 918.750 481.050 919.200 ;
        RECT 484.950 918.750 487.050 919.200 ;
        RECT 478.950 917.550 487.050 918.750 ;
        RECT 478.950 917.100 481.050 917.550 ;
        RECT 484.950 917.100 487.050 917.550 ;
        RECT 496.950 918.750 499.050 919.200 ;
        RECT 508.950 918.750 511.050 919.200 ;
        RECT 496.950 917.550 511.050 918.750 ;
        RECT 496.950 917.100 499.050 917.550 ;
        RECT 508.950 917.100 511.050 917.550 ;
        RECT 520.950 918.600 523.050 919.200 ;
        RECT 541.950 918.600 544.050 919.200 ;
        RECT 556.950 918.600 559.050 919.200 ;
        RECT 520.950 917.400 544.050 918.600 ;
        RECT 520.950 917.100 523.050 917.400 ;
        RECT 541.950 917.100 544.050 917.400 ;
        RECT 545.400 917.400 559.050 918.600 ;
        RECT 458.400 915.600 459.600 917.100 ;
        RECT 545.400 915.600 546.600 917.400 ;
        RECT 556.950 917.100 559.050 917.400 ;
        RECT 583.950 917.100 586.050 919.200 ;
        RECT 589.950 918.600 592.050 919.050 ;
        RECT 601.950 918.600 604.050 919.200 ;
        RECT 589.950 917.400 604.050 918.600 ;
        RECT 458.400 914.400 483.600 915.600 ;
        RECT 454.950 912.600 457.050 912.900 ;
        RECT 449.400 911.400 457.050 912.600 ;
        RECT 482.400 912.600 483.600 914.400 ;
        RECT 524.400 914.400 546.600 915.600 ;
        RECT 584.400 915.600 585.600 917.100 ;
        RECT 589.950 916.950 592.050 917.400 ;
        RECT 601.950 917.100 604.050 917.400 ;
        RECT 631.950 918.600 634.050 919.050 ;
        RECT 637.950 918.600 640.050 919.200 ;
        RECT 631.950 917.400 640.050 918.600 ;
        RECT 631.950 916.950 634.050 917.400 ;
        RECT 637.950 917.100 640.050 917.400 ;
        RECT 676.950 918.750 679.050 919.200 ;
        RECT 688.950 918.750 691.050 919.200 ;
        RECT 676.950 917.550 691.050 918.750 ;
        RECT 676.950 917.100 679.050 917.550 ;
        RECT 688.950 917.100 691.050 917.550 ;
        RECT 703.950 917.100 706.050 919.200 ;
        RECT 727.950 918.750 730.050 919.200 ;
        RECT 736.950 918.750 739.050 919.200 ;
        RECT 727.950 917.550 739.050 918.750 ;
        RECT 727.950 917.100 730.050 917.550 ;
        RECT 736.950 917.100 739.050 917.550 ;
        RECT 748.950 918.600 751.050 919.200 ;
        RECT 763.950 918.600 766.050 919.200 ;
        RECT 787.950 918.600 790.050 919.200 ;
        RECT 748.950 917.400 790.050 918.600 ;
        RECT 748.950 917.100 751.050 917.400 ;
        RECT 763.950 917.100 766.050 917.400 ;
        RECT 787.950 917.100 790.050 917.400 ;
        RECT 799.950 918.600 802.050 919.050 ;
        RECT 808.950 918.600 811.050 919.200 ;
        RECT 799.950 917.400 811.050 918.600 ;
        RECT 704.400 915.600 705.600 917.100 ;
        RECT 799.950 916.950 802.050 917.400 ;
        RECT 808.950 917.100 811.050 917.400 ;
        RECT 817.950 918.750 820.050 919.200 ;
        RECT 823.950 918.750 826.050 919.200 ;
        RECT 817.950 917.550 826.050 918.750 ;
        RECT 850.950 918.600 853.050 919.200 ;
        RECT 817.950 917.100 820.050 917.550 ;
        RECT 823.950 917.100 826.050 917.550 ;
        RECT 827.400 917.400 853.050 918.600 ;
        RECT 584.400 915.000 588.600 915.600 ;
        RECT 584.400 914.400 589.050 915.000 ;
        RECT 524.400 912.900 525.600 914.400 ;
        RECT 517.950 912.600 520.050 912.900 ;
        RECT 482.400 911.400 520.050 912.600 ;
        RECT 421.950 910.950 424.050 911.400 ;
        RECT 433.950 910.800 436.050 911.400 ;
        RECT 454.950 910.800 457.050 911.400 ;
        RECT 517.950 910.800 520.050 911.400 ;
        RECT 523.950 910.800 526.050 912.900 ;
        RECT 574.950 910.800 577.050 912.900 ;
        RECT 586.950 910.950 589.050 914.400 ;
        RECT 686.400 914.400 705.600 915.600 ;
        RECT 604.950 912.600 607.050 912.900 ;
        RECT 619.950 912.600 622.050 912.900 ;
        RECT 604.950 911.400 622.050 912.600 ;
        RECT 604.950 910.800 607.050 911.400 ;
        RECT 619.950 910.800 622.050 911.400 ;
        RECT 625.950 912.450 628.050 912.900 ;
        RECT 631.950 912.450 634.050 912.900 ;
        RECT 625.950 911.250 634.050 912.450 ;
        RECT 625.950 910.800 628.050 911.250 ;
        RECT 631.950 910.800 634.050 911.250 ;
        RECT 646.950 912.600 649.050 913.050 ;
        RECT 655.950 912.600 658.050 912.900 ;
        RECT 646.950 911.400 658.050 912.600 ;
        RECT 646.950 910.950 649.050 911.400 ;
        RECT 655.950 910.800 658.050 911.400 ;
        RECT 679.950 912.600 682.050 912.900 ;
        RECT 686.400 912.600 687.600 914.400 ;
        RECT 679.950 911.400 687.600 912.600 ;
        RECT 688.950 912.600 691.050 913.050 ;
        RECT 700.950 912.600 703.050 912.900 ;
        RECT 688.950 911.400 703.050 912.600 ;
        RECT 679.950 910.800 682.050 911.400 ;
        RECT 688.950 910.950 691.050 911.400 ;
        RECT 700.950 910.800 703.050 911.400 ;
        RECT 721.950 912.600 724.050 912.900 ;
        RECT 742.950 912.600 745.050 912.900 ;
        RECT 721.950 911.400 745.050 912.600 ;
        RECT 721.950 910.800 724.050 911.400 ;
        RECT 742.950 910.800 745.050 911.400 ;
        RECT 766.950 912.600 769.050 912.900 ;
        RECT 778.950 912.600 781.050 913.050 ;
        RECT 827.400 912.900 828.600 917.400 ;
        RECT 850.950 917.100 853.050 917.400 ;
        RECT 874.950 918.600 877.050 919.200 ;
        RECT 883.950 918.600 886.050 919.050 ;
        RECT 892.950 918.600 895.050 919.200 ;
        RECT 874.950 917.400 895.050 918.600 ;
        RECT 874.950 917.100 877.050 917.400 ;
        RECT 883.950 916.950 886.050 917.400 ;
        RECT 892.950 917.100 895.050 917.400 ;
        RECT 898.950 918.600 901.050 919.200 ;
        RECT 907.950 918.600 910.050 919.050 ;
        RECT 916.950 918.600 919.050 919.200 ;
        RECT 898.950 917.400 919.050 918.600 ;
        RECT 898.950 917.100 901.050 917.400 ;
        RECT 907.950 916.950 910.050 917.400 ;
        RECT 916.950 917.100 919.050 917.400 ;
        RECT 766.950 911.400 781.050 912.600 ;
        RECT 766.950 910.800 769.050 911.400 ;
        RECT 778.950 910.950 781.050 911.400 ;
        RECT 790.950 912.450 793.050 912.900 ;
        RECT 799.950 912.450 802.050 912.900 ;
        RECT 790.950 911.250 802.050 912.450 ;
        RECT 790.950 910.800 793.050 911.250 ;
        RECT 799.950 910.800 802.050 911.250 ;
        RECT 826.950 910.800 829.050 912.900 ;
        RECT 832.950 912.450 835.050 912.900 ;
        RECT 841.950 912.450 844.050 912.900 ;
        RECT 832.950 911.250 844.050 912.450 ;
        RECT 832.950 910.800 835.050 911.250 ;
        RECT 841.950 910.800 844.050 911.250 ;
        RECT 847.950 912.600 850.050 912.900 ;
        RECT 871.950 912.600 874.050 912.900 ;
        RECT 847.950 911.400 874.050 912.600 ;
        RECT 847.950 910.800 850.050 911.400 ;
        RECT 871.950 910.800 874.050 911.400 ;
        RECT 877.950 912.600 880.050 912.900 ;
        RECT 889.950 912.600 892.050 912.900 ;
        RECT 904.950 912.600 907.050 913.050 ;
        RECT 877.950 911.400 907.050 912.600 ;
        RECT 877.950 910.800 880.050 911.400 ;
        RECT 889.950 910.800 892.050 911.400 ;
        RECT 904.950 910.950 907.050 911.400 ;
        RECT 913.950 912.450 916.050 912.900 ;
        RECT 928.950 912.450 931.050 912.900 ;
        RECT 913.950 911.250 931.050 912.450 ;
        RECT 913.950 910.800 916.050 911.250 ;
        RECT 928.950 910.800 931.050 911.250 ;
        RECT 112.950 908.400 123.600 909.600 ;
        RECT 169.950 909.600 172.050 910.050 ;
        RECT 178.950 909.600 181.050 910.050 ;
        RECT 169.950 908.400 181.050 909.600 ;
        RECT 112.950 907.950 115.050 908.400 ;
        RECT 115.950 907.950 118.050 908.400 ;
        RECT 169.950 907.950 172.050 908.400 ;
        RECT 178.950 907.950 181.050 908.400 ;
        RECT 232.950 909.600 235.050 910.050 ;
        RECT 241.950 909.600 244.050 910.050 ;
        RECT 232.950 908.400 244.050 909.600 ;
        RECT 232.950 907.950 235.050 908.400 ;
        RECT 241.950 907.950 244.050 908.400 ;
        RECT 439.950 909.600 442.050 910.050 ;
        RECT 469.950 909.600 472.050 910.050 ;
        RECT 439.950 908.400 472.050 909.600 ;
        RECT 439.950 907.950 442.050 908.400 ;
        RECT 469.950 907.950 472.050 908.400 ;
        RECT 478.950 909.600 481.050 910.050 ;
        RECT 523.950 909.600 526.050 910.050 ;
        RECT 478.950 908.400 526.050 909.600 ;
        RECT 575.400 909.600 576.600 910.800 ;
        RECT 583.950 909.600 586.050 910.050 ;
        RECT 575.400 908.400 586.050 909.600 ;
        RECT 478.950 907.950 481.050 908.400 ;
        RECT 523.950 907.950 526.050 908.400 ;
        RECT 583.950 907.950 586.050 908.400 ;
        RECT 49.950 906.600 52.050 907.050 ;
        RECT 70.950 906.600 73.050 907.050 ;
        RECT 49.950 905.400 73.050 906.600 ;
        RECT 49.950 904.950 52.050 905.400 ;
        RECT 70.950 904.950 73.050 905.400 ;
        RECT 289.950 906.600 292.050 907.050 ;
        RECT 319.950 906.600 322.050 907.050 ;
        RECT 289.950 905.400 322.050 906.600 ;
        RECT 289.950 904.950 292.050 905.400 ;
        RECT 319.950 904.950 322.050 905.400 ;
        RECT 355.950 906.600 358.050 907.050 ;
        RECT 361.950 906.600 364.050 907.050 ;
        RECT 355.950 905.400 364.050 906.600 ;
        RECT 355.950 904.950 358.050 905.400 ;
        RECT 361.950 904.950 364.050 905.400 ;
        RECT 394.950 906.600 397.050 907.050 ;
        RECT 415.950 906.600 418.050 907.050 ;
        RECT 424.950 906.600 427.050 907.050 ;
        RECT 430.950 906.600 433.050 907.050 ;
        RECT 394.950 905.400 433.050 906.600 ;
        RECT 394.950 904.950 397.050 905.400 ;
        RECT 415.950 904.950 418.050 905.400 ;
        RECT 424.950 904.950 427.050 905.400 ;
        RECT 430.950 904.950 433.050 905.400 ;
        RECT 436.950 906.600 439.050 907.050 ;
        RECT 442.950 906.600 445.050 907.050 ;
        RECT 436.950 905.400 445.050 906.600 ;
        RECT 436.950 904.950 439.050 905.400 ;
        RECT 442.950 904.950 445.050 905.400 ;
        RECT 595.950 906.600 598.050 907.050 ;
        RECT 646.950 906.600 649.050 907.050 ;
        RECT 595.950 905.400 649.050 906.600 ;
        RECT 595.950 904.950 598.050 905.400 ;
        RECT 646.950 904.950 649.050 905.400 ;
        RECT 694.950 906.600 697.050 907.050 ;
        RECT 706.950 906.600 709.050 907.050 ;
        RECT 712.950 906.600 715.050 907.050 ;
        RECT 694.950 905.400 715.050 906.600 ;
        RECT 694.950 904.950 697.050 905.400 ;
        RECT 706.950 904.950 709.050 905.400 ;
        RECT 712.950 904.950 715.050 905.400 ;
        RECT 817.950 906.600 820.050 907.050 ;
        RECT 835.950 906.600 838.050 907.050 ;
        RECT 817.950 905.400 838.050 906.600 ;
        RECT 817.950 904.950 820.050 905.400 ;
        RECT 835.950 904.950 838.050 905.400 ;
        RECT 124.950 903.600 127.050 904.050 ;
        RECT 157.950 903.600 160.050 904.050 ;
        RECT 124.950 902.400 160.050 903.600 ;
        RECT 124.950 901.950 127.050 902.400 ;
        RECT 157.950 901.950 160.050 902.400 ;
        RECT 193.950 903.600 196.050 904.050 ;
        RECT 259.950 903.600 262.050 904.050 ;
        RECT 283.950 903.600 286.050 904.050 ;
        RECT 349.950 903.600 352.050 904.050 ;
        RECT 193.950 902.400 352.050 903.600 ;
        RECT 193.950 901.950 196.050 902.400 ;
        RECT 259.950 901.950 262.050 902.400 ;
        RECT 283.950 901.950 286.050 902.400 ;
        RECT 349.950 901.950 352.050 902.400 ;
        RECT 463.950 903.600 466.050 904.050 ;
        RECT 475.950 903.600 478.050 904.050 ;
        RECT 463.950 902.400 478.050 903.600 ;
        RECT 463.950 901.950 466.050 902.400 ;
        RECT 475.950 901.950 478.050 902.400 ;
        RECT 508.950 903.600 511.050 904.050 ;
        RECT 538.950 903.600 541.050 904.050 ;
        RECT 673.950 903.600 676.050 904.050 ;
        RECT 508.950 902.400 676.050 903.600 ;
        RECT 508.950 901.950 511.050 902.400 ;
        RECT 538.950 901.950 541.050 902.400 ;
        RECT 673.950 901.950 676.050 902.400 ;
        RECT 883.950 903.600 886.050 904.050 ;
        RECT 931.950 903.600 934.050 904.050 ;
        RECT 883.950 902.400 934.050 903.600 ;
        RECT 883.950 901.950 886.050 902.400 ;
        RECT 931.950 901.950 934.050 902.400 ;
        RECT 46.950 900.600 49.050 901.050 ;
        RECT 97.950 900.600 100.050 901.050 ;
        RECT 115.950 900.600 118.050 901.050 ;
        RECT 46.950 899.400 57.600 900.600 ;
        RECT 46.950 898.950 49.050 899.400 ;
        RECT 56.400 897.600 57.600 899.400 ;
        RECT 97.950 899.400 118.050 900.600 ;
        RECT 97.950 898.950 100.050 899.400 ;
        RECT 115.950 898.950 118.050 899.400 ;
        RECT 238.950 900.600 241.050 901.050 ;
        RECT 289.950 900.600 292.050 901.050 ;
        RECT 238.950 899.400 292.050 900.600 ;
        RECT 238.950 898.950 241.050 899.400 ;
        RECT 289.950 898.950 292.050 899.400 ;
        RECT 586.950 900.600 589.050 901.050 ;
        RECT 610.950 900.600 613.050 901.050 ;
        RECT 586.950 899.400 613.050 900.600 ;
        RECT 586.950 898.950 589.050 899.400 ;
        RECT 610.950 898.950 613.050 899.400 ;
        RECT 727.950 900.600 730.050 901.050 ;
        RECT 802.950 900.600 805.050 901.050 ;
        RECT 808.950 900.600 811.050 901.050 ;
        RECT 727.950 899.400 811.050 900.600 ;
        RECT 727.950 898.950 730.050 899.400 ;
        RECT 802.950 898.950 805.050 899.400 ;
        RECT 808.950 898.950 811.050 899.400 ;
        RECT 862.950 900.600 865.050 901.050 ;
        RECT 892.950 900.600 895.050 901.050 ;
        RECT 862.950 899.400 895.050 900.600 ;
        RECT 862.950 898.950 865.050 899.400 ;
        RECT 892.950 898.950 895.050 899.400 ;
        RECT 106.950 897.600 109.050 898.050 ;
        RECT 56.400 896.400 109.050 897.600 ;
        RECT 106.950 895.950 109.050 896.400 ;
        RECT 121.950 897.600 124.050 898.050 ;
        RECT 130.950 897.600 133.050 898.050 ;
        RECT 331.950 897.600 334.050 898.050 ;
        RECT 121.950 896.400 133.050 897.600 ;
        RECT 121.950 895.950 124.050 896.400 ;
        RECT 130.950 895.950 133.050 896.400 ;
        RECT 293.400 896.400 334.050 897.600 ;
        RECT 46.950 894.600 49.050 895.050 ;
        RECT 88.950 894.600 91.050 895.050 ;
        RECT 46.950 893.400 91.050 894.600 ;
        RECT 46.950 892.950 49.050 893.400 ;
        RECT 88.950 892.950 91.050 893.400 ;
        RECT 199.950 894.600 202.050 895.050 ;
        RECT 205.950 894.600 208.050 895.050 ;
        RECT 199.950 893.400 208.050 894.600 ;
        RECT 199.950 892.950 202.050 893.400 ;
        RECT 205.950 892.950 208.050 893.400 ;
        RECT 226.950 894.600 229.050 895.050 ;
        RECT 235.950 894.600 238.050 895.050 ;
        RECT 226.950 893.400 238.050 894.600 ;
        RECT 226.950 892.950 229.050 893.400 ;
        RECT 235.950 892.950 238.050 893.400 ;
        RECT 271.950 894.600 274.050 895.050 ;
        RECT 293.400 894.600 294.600 896.400 ;
        RECT 331.950 895.950 334.050 896.400 ;
        RECT 400.950 897.600 403.050 898.050 ;
        RECT 409.950 897.600 412.050 898.050 ;
        RECT 415.950 897.600 418.050 898.050 ;
        RECT 400.950 896.400 418.050 897.600 ;
        RECT 400.950 895.950 403.050 896.400 ;
        RECT 409.950 895.950 412.050 896.400 ;
        RECT 415.950 895.950 418.050 896.400 ;
        RECT 523.950 897.600 526.050 898.050 ;
        RECT 541.950 897.600 544.050 898.050 ;
        RECT 577.950 897.600 580.050 898.050 ;
        RECT 640.950 897.600 643.050 898.050 ;
        RECT 679.950 897.600 682.050 898.050 ;
        RECT 523.950 896.400 682.050 897.600 ;
        RECT 523.950 895.950 526.050 896.400 ;
        RECT 541.950 895.950 544.050 896.400 ;
        RECT 577.950 895.950 580.050 896.400 ;
        RECT 640.950 895.950 643.050 896.400 ;
        RECT 679.950 895.950 682.050 896.400 ;
        RECT 706.950 897.600 709.050 898.050 ;
        RECT 721.950 897.600 724.050 898.050 ;
        RECT 706.950 896.400 724.050 897.600 ;
        RECT 706.950 895.950 709.050 896.400 ;
        RECT 721.950 895.950 724.050 896.400 ;
        RECT 772.950 897.600 775.050 898.050 ;
        RECT 787.950 897.600 790.050 898.050 ;
        RECT 772.950 896.400 790.050 897.600 ;
        RECT 772.950 895.950 775.050 896.400 ;
        RECT 787.950 895.950 790.050 896.400 ;
        RECT 853.950 897.600 856.050 898.050 ;
        RECT 862.950 897.600 865.050 897.900 ;
        RECT 853.950 896.400 865.050 897.600 ;
        RECT 853.950 895.950 856.050 896.400 ;
        RECT 862.950 895.800 865.050 896.400 ;
        RECT 898.950 897.600 901.050 898.050 ;
        RECT 907.950 897.600 910.050 898.050 ;
        RECT 898.950 896.400 910.050 897.600 ;
        RECT 898.950 895.950 901.050 896.400 ;
        RECT 907.950 895.950 910.050 896.400 ;
        RECT 271.950 893.400 294.600 894.600 ;
        RECT 412.950 894.600 415.050 895.050 ;
        RECT 445.950 894.600 448.050 895.050 ;
        RECT 469.950 894.600 472.050 895.050 ;
        RECT 412.950 893.400 472.050 894.600 ;
        RECT 271.950 892.950 274.050 893.400 ;
        RECT 412.950 892.950 415.050 893.400 ;
        RECT 445.950 892.950 448.050 893.400 ;
        RECT 469.950 892.950 472.050 893.400 ;
        RECT 484.950 894.600 487.050 895.050 ;
        RECT 493.950 894.600 496.050 895.050 ;
        RECT 547.950 894.600 550.050 895.050 ;
        RECT 565.950 894.600 568.050 895.050 ;
        RECT 484.950 893.400 568.050 894.600 ;
        RECT 484.950 892.950 487.050 893.400 ;
        RECT 493.950 892.950 496.050 893.400 ;
        RECT 547.950 892.950 550.050 893.400 ;
        RECT 565.950 892.950 568.050 893.400 ;
        RECT 1.950 891.600 4.050 892.050 ;
        RECT 13.950 891.600 16.050 892.050 ;
        RECT 1.950 890.400 16.050 891.600 ;
        RECT 1.950 889.950 4.050 890.400 ;
        RECT 13.950 889.950 16.050 890.400 ;
        RECT 25.950 891.600 28.050 892.050 ;
        RECT 37.950 891.600 40.050 892.050 ;
        RECT 55.950 891.600 58.050 892.050 ;
        RECT 25.950 890.400 40.050 891.600 ;
        RECT 25.950 889.950 28.050 890.400 ;
        RECT 37.950 889.950 40.050 890.400 ;
        RECT 50.400 890.400 58.050 891.600 ;
        RECT 50.400 888.600 51.600 890.400 ;
        RECT 55.950 889.950 58.050 890.400 ;
        RECT 175.950 891.600 178.050 892.050 ;
        RECT 187.950 891.600 190.050 892.050 ;
        RECT 175.950 890.400 190.050 891.600 ;
        RECT 175.950 889.950 178.050 890.400 ;
        RECT 187.950 889.950 190.050 890.400 ;
        RECT 211.950 891.600 214.050 892.050 ;
        RECT 256.950 891.600 259.050 892.050 ;
        RECT 211.950 890.400 259.050 891.600 ;
        RECT 211.950 889.950 214.050 890.400 ;
        RECT 256.950 889.950 259.050 890.400 ;
        RECT 301.950 891.600 304.050 892.050 ;
        RECT 322.950 891.600 325.050 892.050 ;
        RECT 400.950 891.600 403.050 892.050 ;
        RECT 301.950 890.400 318.600 891.600 ;
        RECT 301.950 889.950 304.050 890.400 ;
        RECT 41.400 887.400 51.600 888.600 ;
        RECT 88.950 888.600 91.050 889.050 ;
        RECT 94.950 888.600 97.050 889.050 ;
        RECT 88.950 887.400 97.050 888.600 ;
        RECT 4.950 885.600 7.050 886.050 ;
        RECT 13.950 885.600 16.050 886.200 ;
        RECT 4.950 884.400 16.050 885.600 ;
        RECT 4.950 883.950 7.050 884.400 ;
        RECT 13.950 884.100 16.050 884.400 ;
        RECT 22.950 885.600 25.050 886.050 ;
        RECT 31.950 885.600 34.050 886.200 ;
        RECT 22.950 884.400 34.050 885.600 ;
        RECT 22.950 883.950 25.050 884.400 ;
        RECT 31.950 884.100 34.050 884.400 ;
        RECT 37.950 885.600 40.050 886.200 ;
        RECT 41.400 885.600 42.600 887.400 ;
        RECT 88.950 886.950 91.050 887.400 ;
        RECT 94.950 886.950 97.050 887.400 ;
        RECT 109.950 888.600 112.050 889.050 ;
        RECT 118.950 888.600 121.050 889.050 ;
        RECT 109.950 887.400 121.050 888.600 ;
        RECT 109.950 886.950 112.050 887.400 ;
        RECT 118.950 886.950 121.050 887.400 ;
        RECT 205.950 888.600 208.050 889.050 ;
        RECT 214.950 888.600 217.050 889.050 ;
        RECT 205.950 887.400 217.050 888.600 ;
        RECT 205.950 886.950 208.050 887.400 ;
        RECT 214.950 886.950 217.050 887.400 ;
        RECT 289.950 888.600 292.050 889.050 ;
        RECT 298.950 888.600 301.050 889.050 ;
        RECT 289.950 887.400 301.050 888.600 ;
        RECT 317.400 888.600 318.600 890.400 ;
        RECT 322.950 890.400 403.050 891.600 ;
        RECT 322.950 889.950 325.050 890.400 ;
        RECT 334.950 888.600 337.050 889.050 ;
        RECT 317.400 887.400 337.050 888.600 ;
        RECT 289.950 886.950 292.050 887.400 ;
        RECT 298.950 886.950 301.050 887.400 ;
        RECT 334.950 886.950 337.050 887.400 ;
        RECT 340.950 886.950 343.050 890.400 ;
        RECT 400.950 889.950 403.050 890.400 ;
        RECT 415.950 891.600 418.050 892.050 ;
        RECT 439.950 891.600 442.050 892.050 ;
        RECT 415.950 890.400 442.050 891.600 ;
        RECT 415.950 889.950 418.050 890.400 ;
        RECT 439.950 889.950 442.050 890.400 ;
        RECT 475.950 891.600 478.050 892.050 ;
        RECT 487.950 891.600 490.050 892.050 ;
        RECT 475.950 890.400 490.050 891.600 ;
        RECT 475.950 889.950 478.050 890.400 ;
        RECT 487.950 889.950 490.050 890.400 ;
        RECT 604.950 891.600 607.050 892.050 ;
        RECT 628.950 891.600 631.050 892.050 ;
        RECT 604.950 890.400 631.050 891.600 ;
        RECT 604.950 889.950 607.050 890.400 ;
        RECT 628.950 889.950 631.050 890.400 ;
        RECT 640.950 891.600 643.050 892.050 ;
        RECT 649.950 891.600 652.050 892.050 ;
        RECT 697.950 891.600 700.050 892.050 ;
        RECT 640.950 890.400 700.050 891.600 ;
        RECT 640.950 889.950 643.050 890.400 ;
        RECT 649.950 889.950 652.050 890.400 ;
        RECT 697.950 889.950 700.050 890.400 ;
        RECT 832.950 891.600 835.050 892.050 ;
        RECT 850.950 891.600 853.050 892.050 ;
        RECT 895.950 891.600 898.050 892.050 ;
        RECT 832.950 890.400 898.050 891.600 ;
        RECT 832.950 889.950 835.050 890.400 ;
        RECT 850.950 889.950 853.050 890.400 ;
        RECT 895.950 889.950 898.050 890.400 ;
        RECT 358.950 888.600 361.050 889.050 ;
        RECT 376.950 888.600 379.050 889.050 ;
        RECT 415.950 888.600 418.050 888.900 ;
        RECT 358.950 887.400 379.050 888.600 ;
        RECT 358.950 886.950 361.050 887.400 ;
        RECT 376.950 886.950 379.050 887.400 ;
        RECT 395.400 887.400 418.050 888.600 ;
        RECT 395.400 886.200 396.600 887.400 ;
        RECT 415.950 886.800 418.050 887.400 ;
        RECT 469.950 888.600 472.050 889.050 ;
        RECT 508.950 888.600 511.050 889.050 ;
        RECT 469.950 887.400 511.050 888.600 ;
        RECT 469.950 886.950 472.050 887.400 ;
        RECT 508.950 886.950 511.050 887.400 ;
        RECT 37.950 884.400 42.600 885.600 ;
        RECT 37.950 884.100 40.050 884.400 ;
        RECT 55.950 884.100 58.050 886.200 ;
        RECT 64.950 885.600 67.050 885.900 ;
        RECT 73.950 885.600 76.050 886.200 ;
        RECT 64.950 884.400 76.050 885.600 ;
        RECT 35.400 881.400 48.600 882.600 ;
        RECT 35.400 879.900 36.600 881.400 ;
        RECT 47.400 879.900 48.600 881.400 ;
        RECT 1.950 879.450 4.050 879.900 ;
        RECT 10.950 879.450 13.050 879.900 ;
        RECT 1.950 878.250 13.050 879.450 ;
        RECT 1.950 877.800 4.050 878.250 ;
        RECT 10.950 877.800 13.050 878.250 ;
        RECT 16.950 879.450 19.050 879.900 ;
        RECT 22.950 879.450 25.050 879.900 ;
        RECT 16.950 878.250 25.050 879.450 ;
        RECT 16.950 877.800 19.050 878.250 ;
        RECT 22.950 877.800 25.050 878.250 ;
        RECT 34.950 877.800 37.050 879.900 ;
        RECT 46.950 879.450 49.050 879.900 ;
        RECT 52.950 879.450 55.050 879.900 ;
        RECT 46.950 878.250 55.050 879.450 ;
        RECT 46.950 877.800 49.050 878.250 ;
        RECT 52.950 877.800 55.050 878.250 ;
        RECT 56.400 877.050 57.600 884.100 ;
        RECT 64.950 883.800 67.050 884.400 ;
        RECT 73.950 884.100 76.050 884.400 ;
        RECT 79.950 884.100 82.050 886.200 ;
        RECT 133.950 884.100 136.050 886.200 ;
        RECT 139.950 885.600 142.050 886.200 ;
        RECT 169.950 885.600 172.050 886.050 ;
        RECT 181.950 885.600 184.050 886.200 ;
        RECT 139.950 884.400 144.600 885.600 ;
        RECT 139.950 884.100 142.050 884.400 ;
        RECT 58.950 879.450 61.050 879.900 ;
        RECT 64.950 879.450 67.050 879.900 ;
        RECT 58.950 878.250 67.050 879.450 ;
        RECT 80.400 879.600 81.600 884.100 ;
        RECT 134.400 882.600 135.600 884.100 ;
        RECT 122.400 881.400 135.600 882.600 ;
        RECT 94.950 879.600 97.050 879.900 ;
        RECT 80.400 878.400 97.050 879.600 ;
        RECT 58.950 877.800 61.050 878.250 ;
        RECT 64.950 877.800 67.050 878.250 ;
        RECT 94.950 877.800 97.050 878.400 ;
        RECT 112.950 879.600 115.050 879.900 ;
        RECT 122.400 879.600 123.600 881.400 ;
        RECT 143.400 880.050 144.600 884.400 ;
        RECT 169.950 884.400 184.050 885.600 ;
        RECT 169.950 883.950 172.050 884.400 ;
        RECT 181.950 884.100 184.050 884.400 ;
        RECT 196.950 885.600 199.050 886.050 ;
        RECT 205.950 885.600 208.050 886.200 ;
        RECT 229.950 885.600 232.050 886.200 ;
        RECT 196.950 884.400 208.050 885.600 ;
        RECT 196.950 883.950 199.050 884.400 ;
        RECT 205.950 884.100 208.050 884.400 ;
        RECT 209.400 884.400 232.050 885.600 ;
        RECT 112.950 878.400 123.600 879.600 ;
        RECT 124.950 879.450 127.050 879.900 ;
        RECT 136.950 879.450 139.050 879.900 ;
        RECT 112.950 877.800 115.050 878.400 ;
        RECT 124.950 878.250 139.050 879.450 ;
        RECT 124.950 877.800 127.050 878.250 ;
        RECT 136.950 877.800 139.050 878.250 ;
        RECT 142.950 877.950 145.050 880.050 ;
        RECT 209.400 879.900 210.600 884.400 ;
        RECT 229.950 884.100 232.050 884.400 ;
        RECT 235.950 885.750 238.050 886.200 ;
        RECT 244.950 885.750 247.050 886.200 ;
        RECT 235.950 884.550 247.050 885.750 ;
        RECT 235.950 884.100 238.050 884.550 ;
        RECT 244.950 884.100 247.050 884.550 ;
        RECT 283.950 885.600 288.000 886.050 ;
        RECT 307.950 885.750 310.050 886.200 ;
        RECT 313.950 885.750 316.050 886.200 ;
        RECT 283.950 883.950 288.600 885.600 ;
        RECT 307.950 884.550 316.050 885.750 ;
        RECT 307.950 884.100 310.050 884.550 ;
        RECT 313.950 884.100 316.050 884.550 ;
        RECT 328.950 885.600 331.050 886.050 ;
        RECT 337.950 885.600 340.050 886.200 ;
        RECT 328.950 884.400 340.050 885.600 ;
        RECT 328.950 883.950 331.050 884.400 ;
        RECT 337.950 884.100 340.050 884.400 ;
        RECT 349.950 885.750 352.050 886.200 ;
        RECT 355.950 885.750 358.050 886.200 ;
        RECT 349.950 884.550 358.050 885.750 ;
        RECT 349.950 884.100 352.050 884.550 ;
        RECT 355.950 884.100 358.050 884.550 ;
        RECT 382.950 885.750 385.050 886.200 ;
        RECT 388.950 885.750 391.050 886.050 ;
        RECT 394.950 885.750 397.050 886.200 ;
        RECT 382.950 884.550 397.050 885.750 ;
        RECT 382.950 884.100 385.050 884.550 ;
        RECT 388.950 883.950 391.050 884.550 ;
        RECT 394.950 884.100 397.050 884.550 ;
        RECT 421.950 885.600 424.050 886.200 ;
        RECT 439.950 885.600 442.050 886.200 ;
        RECT 421.950 884.400 442.050 885.600 ;
        RECT 421.950 884.100 424.050 884.400 ;
        RECT 439.950 884.100 442.050 884.400 ;
        RECT 448.950 885.750 451.050 886.200 ;
        RECT 454.950 885.750 457.050 886.200 ;
        RECT 448.950 884.550 457.050 885.750 ;
        RECT 448.950 884.100 451.050 884.550 ;
        RECT 454.950 884.100 457.050 884.550 ;
        RECT 514.950 885.750 517.050 886.200 ;
        RECT 526.800 885.750 528.900 886.200 ;
        RECT 514.950 884.550 528.900 885.750 ;
        RECT 529.950 885.600 532.050 889.050 ;
        RECT 631.950 888.600 634.050 889.050 ;
        RECT 637.950 888.600 640.050 889.050 ;
        RECT 631.950 887.400 640.050 888.600 ;
        RECT 631.950 886.950 634.050 887.400 ;
        RECT 637.950 886.950 640.050 887.400 ;
        RECT 667.950 888.600 670.050 889.050 ;
        RECT 688.950 888.600 691.050 889.050 ;
        RECT 667.950 887.400 691.050 888.600 ;
        RECT 667.950 886.950 670.050 887.400 ;
        RECT 688.950 886.950 691.050 887.400 ;
        RECT 736.950 888.600 739.050 889.050 ;
        RECT 748.950 888.600 751.050 889.050 ;
        RECT 736.950 887.400 751.050 888.600 ;
        RECT 736.950 886.950 739.050 887.400 ;
        RECT 748.950 886.950 751.050 887.400 ;
        RECT 754.950 888.600 757.050 889.050 ;
        RECT 760.950 888.600 763.050 889.050 ;
        RECT 754.950 887.400 763.050 888.600 ;
        RECT 754.950 886.950 757.050 887.400 ;
        RECT 760.950 886.950 763.050 887.400 ;
        RECT 535.950 885.600 538.050 886.200 ;
        RECT 529.950 885.000 538.050 885.600 ;
        RECT 514.950 884.100 517.050 884.550 ;
        RECT 526.800 884.100 528.900 884.550 ;
        RECT 530.400 884.400 538.050 885.000 ;
        RECT 535.950 884.100 538.050 884.400 ;
        RECT 559.950 885.600 562.050 886.200 ;
        RECT 571.950 885.600 574.050 886.050 ;
        RECT 604.950 885.600 607.050 886.200 ;
        RECT 559.950 884.400 574.050 885.600 ;
        RECT 559.950 884.100 562.050 884.400 ;
        RECT 571.950 883.950 574.050 884.400 ;
        RECT 587.400 884.400 607.050 885.600 ;
        RECT 184.950 879.450 187.050 879.900 ;
        RECT 196.950 879.450 199.050 879.900 ;
        RECT 184.950 878.250 199.050 879.450 ;
        RECT 184.950 877.800 187.050 878.250 ;
        RECT 196.950 877.800 199.050 878.250 ;
        RECT 208.950 877.800 211.050 879.900 ;
        RECT 214.950 879.600 217.050 879.900 ;
        RECT 247.950 879.600 250.050 879.900 ;
        RECT 259.950 879.600 262.050 880.050 ;
        RECT 287.400 879.900 288.600 883.950 ;
        RECT 214.950 878.400 262.050 879.600 ;
        RECT 214.950 877.800 217.050 878.400 ;
        RECT 247.950 877.800 250.050 878.400 ;
        RECT 259.950 877.950 262.050 878.400 ;
        RECT 286.950 877.800 289.050 879.900 ;
        RECT 316.950 879.600 319.050 879.900 ;
        RECT 340.950 879.600 343.050 879.900 ;
        RECT 349.950 879.600 352.050 880.050 ;
        RECT 316.950 878.400 352.050 879.600 ;
        RECT 316.950 877.800 319.050 878.400 ;
        RECT 340.950 877.800 343.050 878.400 ;
        RECT 349.950 877.950 352.050 878.400 ;
        RECT 358.950 879.600 361.050 879.900 ;
        RECT 373.950 879.600 376.050 879.900 ;
        RECT 358.950 878.400 376.050 879.600 ;
        RECT 358.950 877.800 361.050 878.400 ;
        RECT 373.950 877.800 376.050 878.400 ;
        RECT 436.950 879.600 439.050 880.050 ;
        RECT 442.950 879.600 445.050 879.900 ;
        RECT 436.950 878.400 445.050 879.600 ;
        RECT 436.950 877.950 439.050 878.400 ;
        RECT 442.950 877.800 445.050 878.400 ;
        RECT 517.950 879.450 520.050 879.900 ;
        RECT 523.800 879.450 525.900 879.900 ;
        RECT 517.950 878.250 525.900 879.450 ;
        RECT 517.950 877.800 520.050 878.250 ;
        RECT 523.800 877.800 525.900 878.250 ;
        RECT 526.950 879.600 529.050 880.050 ;
        RECT 587.400 879.900 588.600 884.400 ;
        RECT 604.950 884.100 607.050 884.400 ;
        RECT 616.950 885.750 619.050 886.200 ;
        RECT 622.950 885.750 625.050 886.200 ;
        RECT 616.950 884.550 625.050 885.750 ;
        RECT 616.950 884.100 619.050 884.550 ;
        RECT 622.950 884.100 625.050 884.550 ;
        RECT 715.950 885.600 718.050 886.050 ;
        RECT 721.950 885.600 724.050 886.200 ;
        RECT 715.950 884.400 724.050 885.600 ;
        RECT 715.950 883.950 718.050 884.400 ;
        RECT 721.950 884.100 724.050 884.400 ;
        RECT 766.950 885.600 769.050 886.200 ;
        RECT 772.950 885.600 775.050 889.050 ;
        RECT 778.950 888.600 781.050 889.050 ;
        RECT 784.800 888.600 786.900 889.050 ;
        RECT 778.950 887.400 786.900 888.600 ;
        RECT 778.950 886.950 781.050 887.400 ;
        RECT 784.800 886.950 786.900 887.400 ;
        RECT 787.950 888.600 790.050 889.050 ;
        RECT 811.950 888.600 814.050 889.050 ;
        RECT 787.950 887.400 814.050 888.600 ;
        RECT 787.950 886.950 790.050 887.400 ;
        RECT 811.950 886.950 814.050 887.400 ;
        RECT 766.950 885.000 775.050 885.600 ;
        RECT 814.950 885.600 817.050 886.200 ;
        RECT 820.950 885.600 823.050 886.050 ;
        RECT 766.950 884.400 774.600 885.000 ;
        RECT 814.950 884.400 823.050 885.600 ;
        RECT 766.950 884.100 769.050 884.400 ;
        RECT 814.950 884.100 817.050 884.400 ;
        RECT 820.950 883.950 823.050 884.400 ;
        RECT 826.950 885.600 829.050 886.200 ;
        RECT 856.950 885.600 859.050 886.200 ;
        RECT 865.950 885.600 868.050 886.050 ;
        RECT 871.950 885.600 874.050 886.200 ;
        RECT 826.950 884.400 855.600 885.600 ;
        RECT 826.950 884.100 829.050 884.400 ;
        RECT 854.400 882.600 855.600 884.400 ;
        RECT 856.950 884.400 868.050 885.600 ;
        RECT 856.950 884.100 859.050 884.400 ;
        RECT 865.950 883.950 868.050 884.400 ;
        RECT 869.400 884.400 874.050 885.600 ;
        RECT 755.400 881.400 813.600 882.600 ;
        RECT 854.400 882.000 861.600 882.600 ;
        RECT 854.400 881.400 862.050 882.000 ;
        RECT 755.400 880.050 756.600 881.400 ;
        RECT 538.950 879.600 541.050 879.900 ;
        RECT 526.950 878.400 541.050 879.600 ;
        RECT 526.950 877.950 529.050 878.400 ;
        RECT 538.950 877.800 541.050 878.400 ;
        RECT 586.950 877.800 589.050 879.900 ;
        RECT 625.950 879.450 628.050 879.900 ;
        RECT 637.950 879.450 640.050 879.900 ;
        RECT 625.950 878.250 640.050 879.450 ;
        RECT 625.950 877.800 628.050 878.250 ;
        RECT 637.950 877.800 640.050 878.250 ;
        RECT 730.950 879.450 733.050 879.900 ;
        RECT 736.950 879.450 739.050 879.900 ;
        RECT 730.950 878.250 739.050 879.450 ;
        RECT 730.950 877.800 733.050 878.250 ;
        RECT 736.950 877.800 739.050 878.250 ;
        RECT 745.950 879.600 748.050 879.900 ;
        RECT 754.950 879.600 757.050 880.050 ;
        RECT 745.950 878.400 757.050 879.600 ;
        RECT 745.950 877.800 748.050 878.400 ;
        RECT 754.950 877.950 757.050 878.400 ;
        RECT 769.950 879.450 772.050 879.900 ;
        RECT 775.950 879.450 778.050 880.050 ;
        RECT 812.400 879.900 813.600 881.400 ;
        RECT 769.950 878.250 778.050 879.450 ;
        RECT 769.950 877.800 772.050 878.250 ;
        RECT 775.950 877.950 778.050 878.250 ;
        RECT 799.950 879.450 802.050 879.900 ;
        RECT 805.950 879.450 808.050 879.900 ;
        RECT 799.950 878.250 808.050 879.450 ;
        RECT 799.950 877.800 802.050 878.250 ;
        RECT 805.950 877.800 808.050 878.250 ;
        RECT 811.950 877.800 814.050 879.900 ;
        RECT 820.950 879.450 823.050 879.900 ;
        RECT 829.950 879.600 832.050 879.900 ;
        RECT 847.950 879.600 850.050 879.900 ;
        RECT 829.950 879.450 850.050 879.600 ;
        RECT 820.950 878.400 850.050 879.450 ;
        RECT 820.950 878.250 832.050 878.400 ;
        RECT 820.950 877.800 823.050 878.250 ;
        RECT 829.950 877.800 832.050 878.250 ;
        RECT 847.950 877.800 850.050 878.400 ;
        RECT 859.950 877.950 862.050 881.400 ;
        RECT 869.400 880.050 870.600 884.400 ;
        RECT 871.950 884.100 874.050 884.400 ;
        RECT 877.950 885.600 880.050 886.200 ;
        RECT 886.800 885.600 888.900 886.050 ;
        RECT 877.950 884.400 888.900 885.600 ;
        RECT 889.950 885.600 892.050 889.050 ;
        RECT 907.950 888.600 910.050 889.050 ;
        RECT 922.950 888.600 925.050 889.050 ;
        RECT 907.950 887.400 925.050 888.600 ;
        RECT 907.950 886.950 910.050 887.400 ;
        RECT 922.950 886.950 925.050 887.400 ;
        RECT 898.950 885.600 901.050 886.200 ;
        RECT 889.950 885.000 901.050 885.600 ;
        RECT 890.400 884.400 901.050 885.000 ;
        RECT 877.950 884.100 880.050 884.400 ;
        RECT 886.800 883.950 888.900 884.400 ;
        RECT 898.950 884.100 901.050 884.400 ;
        RECT 916.950 884.100 919.050 886.200 ;
        RECT 868.950 877.950 871.050 880.050 ;
        RECT 886.950 879.450 889.050 879.900 ;
        RECT 901.950 879.600 904.050 879.900 ;
        RECT 917.400 879.600 918.600 884.100 ;
        RECT 901.950 879.450 918.600 879.600 ;
        RECT 886.950 878.400 918.600 879.450 ;
        RECT 886.950 878.250 904.050 878.400 ;
        RECT 886.950 877.800 889.050 878.250 ;
        RECT 901.950 877.800 904.050 878.250 ;
        RECT 55.950 874.950 58.050 877.050 ;
        RECT 262.950 876.600 265.050 877.050 ;
        RECT 367.950 876.600 370.050 877.050 ;
        RECT 379.950 876.600 382.050 877.050 ;
        RECT 418.950 876.600 421.050 877.050 ;
        RECT 262.950 875.400 421.050 876.600 ;
        RECT 262.950 874.950 265.050 875.400 ;
        RECT 367.950 874.950 370.050 875.400 ;
        RECT 379.950 874.950 382.050 875.400 ;
        RECT 418.950 874.950 421.050 875.400 ;
        RECT 424.950 876.600 427.050 877.050 ;
        RECT 454.950 876.600 457.050 877.050 ;
        RECT 466.950 876.600 469.050 877.050 ;
        RECT 424.950 875.400 469.050 876.600 ;
        RECT 424.950 874.950 427.050 875.400 ;
        RECT 454.950 874.950 457.050 875.400 ;
        RECT 466.950 874.950 469.050 875.400 ;
        RECT 565.950 876.600 568.050 877.050 ;
        RECT 580.950 876.600 583.050 877.050 ;
        RECT 595.950 876.600 598.050 877.050 ;
        RECT 565.950 875.400 598.050 876.600 ;
        RECT 565.950 874.950 568.050 875.400 ;
        RECT 580.950 874.950 583.050 875.400 ;
        RECT 595.950 874.950 598.050 875.400 ;
        RECT 697.950 876.600 700.050 877.050 ;
        RECT 724.950 876.600 727.050 877.050 ;
        RECT 697.950 875.400 727.050 876.600 ;
        RECT 697.950 874.950 700.050 875.400 ;
        RECT 724.950 874.950 727.050 875.400 ;
        RECT 40.950 873.600 43.050 874.050 ;
        RECT 58.950 873.600 61.050 874.050 ;
        RECT 40.950 872.400 61.050 873.600 ;
        RECT 40.950 871.950 43.050 872.400 ;
        RECT 58.950 871.950 61.050 872.400 ;
        RECT 106.950 873.600 109.050 874.050 ;
        RECT 130.950 873.600 133.050 874.050 ;
        RECT 106.950 872.400 133.050 873.600 ;
        RECT 106.950 871.950 109.050 872.400 ;
        RECT 130.950 871.950 133.050 872.400 ;
        RECT 232.950 873.600 235.050 874.050 ;
        RECT 256.950 873.600 259.050 874.050 ;
        RECT 349.950 873.600 352.050 874.050 ;
        RECT 232.950 872.400 352.050 873.600 ;
        RECT 232.950 871.950 235.050 872.400 ;
        RECT 256.950 871.950 259.050 872.400 ;
        RECT 349.950 871.950 352.050 872.400 ;
        RECT 430.950 873.600 433.050 874.050 ;
        RECT 448.950 873.600 451.050 874.050 ;
        RECT 430.950 872.400 451.050 873.600 ;
        RECT 430.950 871.950 433.050 872.400 ;
        RECT 448.950 871.950 451.050 872.400 ;
        RECT 544.950 873.600 547.050 874.050 ;
        RECT 553.950 873.600 556.050 874.050 ;
        RECT 586.950 873.600 589.050 874.050 ;
        RECT 544.950 872.400 552.600 873.600 ;
        RECT 544.950 871.950 547.050 872.400 ;
        RECT 298.950 870.600 301.050 871.050 ;
        RECT 307.950 870.600 310.050 871.050 ;
        RECT 334.950 870.600 337.050 871.050 ;
        RECT 469.950 870.600 472.050 871.050 ;
        RECT 298.950 869.400 472.050 870.600 ;
        RECT 551.400 870.600 552.600 872.400 ;
        RECT 553.950 872.400 589.050 873.600 ;
        RECT 553.950 871.950 556.050 872.400 ;
        RECT 586.950 871.950 589.050 872.400 ;
        RECT 631.950 873.600 634.050 874.050 ;
        RECT 664.950 873.600 667.050 874.050 ;
        RECT 631.950 872.400 667.050 873.600 ;
        RECT 631.950 871.950 634.050 872.400 ;
        RECT 664.950 871.950 667.050 872.400 ;
        RECT 889.950 873.600 892.050 874.050 ;
        RECT 913.950 873.600 916.050 874.050 ;
        RECT 889.950 872.400 916.050 873.600 ;
        RECT 889.950 871.950 892.050 872.400 ;
        RECT 913.950 871.950 916.050 872.400 ;
        RECT 643.950 870.600 646.050 871.050 ;
        RECT 551.400 869.400 646.050 870.600 ;
        RECT 298.950 868.950 301.050 869.400 ;
        RECT 307.950 868.950 310.050 869.400 ;
        RECT 334.950 868.950 337.050 869.400 ;
        RECT 469.950 868.950 472.050 869.400 ;
        RECT 643.950 868.950 646.050 869.400 ;
        RECT 865.950 870.600 868.050 871.050 ;
        RECT 877.950 870.600 880.050 871.050 ;
        RECT 865.950 869.400 880.050 870.600 ;
        RECT 865.950 868.950 868.050 869.400 ;
        RECT 877.950 868.950 880.050 869.400 ;
        RECT 907.950 870.600 910.050 871.050 ;
        RECT 919.950 870.600 922.050 871.050 ;
        RECT 907.950 869.400 922.050 870.600 ;
        RECT 907.950 868.950 910.050 869.400 ;
        RECT 919.950 868.950 922.050 869.400 ;
        RECT 193.950 867.600 196.050 868.050 ;
        RECT 277.950 867.600 280.050 868.050 ;
        RECT 193.950 866.400 280.050 867.600 ;
        RECT 193.950 865.950 196.050 866.400 ;
        RECT 277.950 865.950 280.050 866.400 ;
        RECT 337.950 867.600 340.050 868.050 ;
        RECT 475.950 867.600 478.050 868.050 ;
        RECT 337.950 866.400 478.050 867.600 ;
        RECT 337.950 865.950 340.050 866.400 ;
        RECT 475.950 865.950 478.050 866.400 ;
        RECT 547.950 867.600 550.050 868.050 ;
        RECT 583.950 867.600 586.050 868.050 ;
        RECT 547.950 866.400 586.050 867.600 ;
        RECT 547.950 865.950 550.050 866.400 ;
        RECT 583.950 865.950 586.050 866.400 ;
        RECT 646.950 867.600 649.050 868.050 ;
        RECT 709.950 867.600 712.050 868.050 ;
        RECT 787.950 867.600 790.050 868.050 ;
        RECT 646.950 866.400 790.050 867.600 ;
        RECT 646.950 865.950 649.050 866.400 ;
        RECT 709.950 865.950 712.050 866.400 ;
        RECT 787.950 865.950 790.050 866.400 ;
        RECT 835.950 867.600 838.050 868.050 ;
        RECT 853.950 867.600 856.050 868.050 ;
        RECT 868.950 867.600 871.050 868.050 ;
        RECT 835.950 866.400 871.050 867.600 ;
        RECT 835.950 865.950 838.050 866.400 ;
        RECT 853.950 865.950 856.050 866.400 ;
        RECT 868.950 865.950 871.050 866.400 ;
        RECT 172.950 864.600 175.050 865.050 ;
        RECT 190.950 864.600 193.050 865.050 ;
        RECT 511.950 864.600 514.050 865.050 ;
        RECT 172.950 863.400 514.050 864.600 ;
        RECT 172.950 862.950 175.050 863.400 ;
        RECT 190.950 862.950 193.050 863.400 ;
        RECT 511.950 862.950 514.050 863.400 ;
        RECT 532.950 864.600 535.050 865.050 ;
        RECT 565.950 864.600 568.050 865.050 ;
        RECT 532.950 863.400 568.050 864.600 ;
        RECT 532.950 862.950 535.050 863.400 ;
        RECT 565.950 862.950 568.050 863.400 ;
        RECT 589.950 864.600 592.050 865.050 ;
        RECT 647.400 864.600 648.600 865.950 ;
        RECT 589.950 863.400 648.600 864.600 ;
        RECT 808.950 864.600 811.050 865.050 ;
        RECT 880.950 864.600 883.050 865.050 ;
        RECT 928.950 864.600 931.050 865.050 ;
        RECT 808.950 863.400 931.050 864.600 ;
        RECT 589.950 862.950 592.050 863.400 ;
        RECT 808.950 862.950 811.050 863.400 ;
        RECT 880.950 862.950 883.050 863.400 ;
        RECT 928.950 862.950 931.050 863.400 ;
        RECT 82.950 861.600 85.050 862.050 ;
        RECT 112.950 861.600 115.050 862.050 ;
        RECT 121.950 861.600 124.050 862.050 ;
        RECT 82.950 860.400 124.050 861.600 ;
        RECT 82.950 859.950 85.050 860.400 ;
        RECT 112.950 859.950 115.050 860.400 ;
        RECT 121.950 859.950 124.050 860.400 ;
        RECT 196.950 861.600 199.050 862.050 ;
        RECT 436.950 861.600 439.050 862.050 ;
        RECT 196.950 860.400 439.050 861.600 ;
        RECT 196.950 859.950 199.050 860.400 ;
        RECT 436.950 859.950 439.050 860.400 ;
        RECT 475.950 861.600 478.050 862.050 ;
        RECT 586.950 861.600 589.050 862.050 ;
        RECT 724.950 861.600 727.050 862.050 ;
        RECT 784.950 861.600 787.050 862.050 ;
        RECT 475.950 860.400 549.600 861.600 ;
        RECT 475.950 859.950 478.050 860.400 ;
        RECT 73.950 858.600 76.050 859.050 ;
        RECT 103.950 858.600 106.050 859.050 ;
        RECT 73.950 857.400 106.050 858.600 ;
        RECT 73.950 856.950 76.050 857.400 ;
        RECT 103.950 856.950 106.050 857.400 ;
        RECT 133.950 858.600 136.050 859.050 ;
        RECT 175.950 858.600 178.050 859.050 ;
        RECT 133.950 857.400 178.050 858.600 ;
        RECT 133.950 856.950 136.050 857.400 ;
        RECT 175.950 856.950 178.050 857.400 ;
        RECT 226.950 858.600 229.050 859.050 ;
        RECT 241.950 858.600 244.050 859.050 ;
        RECT 262.950 858.600 265.050 859.050 ;
        RECT 226.950 857.400 265.050 858.600 ;
        RECT 226.950 856.950 229.050 857.400 ;
        RECT 241.950 856.950 244.050 857.400 ;
        RECT 262.950 856.950 265.050 857.400 ;
        RECT 376.950 858.600 379.050 859.050 ;
        RECT 472.950 858.600 475.050 859.050 ;
        RECT 544.950 858.600 547.050 859.050 ;
        RECT 376.950 857.400 547.050 858.600 ;
        RECT 548.400 858.600 549.600 860.400 ;
        RECT 586.950 860.400 787.050 861.600 ;
        RECT 586.950 859.950 589.050 860.400 ;
        RECT 724.950 859.950 727.050 860.400 ;
        RECT 784.950 859.950 787.050 860.400 ;
        RECT 841.950 861.600 844.050 862.050 ;
        RECT 871.950 861.600 874.050 862.050 ;
        RECT 841.950 860.400 874.050 861.600 ;
        RECT 841.950 859.950 844.050 860.400 ;
        RECT 871.950 859.950 874.050 860.400 ;
        RECT 565.950 858.600 568.050 859.050 ;
        RECT 548.400 857.400 568.050 858.600 ;
        RECT 376.950 856.950 379.050 857.400 ;
        RECT 472.950 856.950 475.050 857.400 ;
        RECT 544.950 856.950 547.050 857.400 ;
        RECT 565.950 856.950 568.050 857.400 ;
        RECT 571.950 858.600 574.050 859.050 ;
        RECT 601.950 858.600 604.050 859.050 ;
        RECT 571.950 857.400 604.050 858.600 ;
        RECT 571.950 856.950 574.050 857.400 ;
        RECT 601.950 856.950 604.050 857.400 ;
        RECT 643.950 858.600 646.050 859.050 ;
        RECT 709.950 858.600 712.050 859.050 ;
        RECT 790.950 858.600 793.050 859.050 ;
        RECT 802.950 858.600 805.050 859.050 ;
        RECT 643.950 857.400 805.050 858.600 ;
        RECT 643.950 856.950 646.050 857.400 ;
        RECT 709.950 856.950 712.050 857.400 ;
        RECT 790.950 856.950 793.050 857.400 ;
        RECT 802.950 856.950 805.050 857.400 ;
        RECT 154.950 855.600 157.050 856.050 ;
        RECT 247.950 855.600 250.050 856.050 ;
        RECT 154.950 854.400 250.050 855.600 ;
        RECT 154.950 853.950 157.050 854.400 ;
        RECT 247.950 853.950 250.050 854.400 ;
        RECT 334.950 855.600 337.050 856.050 ;
        RECT 377.400 855.600 378.600 856.950 ;
        RECT 334.950 854.400 378.600 855.600 ;
        RECT 427.950 855.600 430.050 856.050 ;
        RECT 454.950 855.600 457.050 856.050 ;
        RECT 589.950 855.600 592.050 856.050 ;
        RECT 427.950 854.400 592.050 855.600 ;
        RECT 334.950 853.950 337.050 854.400 ;
        RECT 427.950 853.950 430.050 854.400 ;
        RECT 454.950 853.950 457.050 854.400 ;
        RECT 589.950 853.950 592.050 854.400 ;
        RECT 832.950 855.600 835.050 856.050 ;
        RECT 886.950 855.600 889.050 856.050 ;
        RECT 832.950 854.400 889.050 855.600 ;
        RECT 832.950 853.950 835.050 854.400 ;
        RECT 886.950 853.950 889.050 854.400 ;
        RECT 292.950 852.600 295.050 853.050 ;
        RECT 313.950 852.600 316.050 853.050 ;
        RECT 292.950 851.400 316.050 852.600 ;
        RECT 292.950 850.950 295.050 851.400 ;
        RECT 313.950 850.950 316.050 851.400 ;
        RECT 610.950 852.600 613.050 853.050 ;
        RECT 817.950 852.600 820.050 853.050 ;
        RECT 610.950 851.400 820.050 852.600 ;
        RECT 610.950 850.950 613.050 851.400 ;
        RECT 817.950 850.950 820.050 851.400 ;
        RECT 4.950 849.600 7.050 850.050 ;
        RECT 58.950 849.600 61.050 850.050 ;
        RECT 4.950 848.400 61.050 849.600 ;
        RECT 4.950 847.950 7.050 848.400 ;
        RECT 58.950 847.950 61.050 848.400 ;
        RECT 223.950 849.600 226.050 850.050 ;
        RECT 232.950 849.600 235.050 850.050 ;
        RECT 223.950 848.400 235.050 849.600 ;
        RECT 223.950 847.950 226.050 848.400 ;
        RECT 232.950 847.950 235.050 848.400 ;
        RECT 262.950 849.600 265.050 850.050 ;
        RECT 274.950 849.600 277.050 850.050 ;
        RECT 262.950 848.400 277.050 849.600 ;
        RECT 262.950 847.950 265.050 848.400 ;
        RECT 274.950 847.950 277.050 848.400 ;
        RECT 421.950 849.600 424.050 850.050 ;
        RECT 532.950 849.600 535.050 850.050 ;
        RECT 421.950 848.400 535.050 849.600 ;
        RECT 421.950 847.950 424.050 848.400 ;
        RECT 532.950 847.950 535.050 848.400 ;
        RECT 547.950 849.600 550.050 850.050 ;
        RECT 562.800 849.600 564.900 849.900 ;
        RECT 547.950 848.400 564.900 849.600 ;
        RECT 547.950 847.950 550.050 848.400 ;
        RECT 562.800 847.800 564.900 848.400 ;
        RECT 565.950 849.600 568.050 850.050 ;
        RECT 589.950 849.600 592.050 850.050 ;
        RECT 565.950 848.400 592.050 849.600 ;
        RECT 565.950 847.950 568.050 848.400 ;
        RECT 589.950 847.950 592.050 848.400 ;
        RECT 601.950 849.600 604.050 850.050 ;
        RECT 616.950 849.600 619.050 850.050 ;
        RECT 637.950 849.600 640.050 850.050 ;
        RECT 601.950 848.400 640.050 849.600 ;
        RECT 601.950 847.950 604.050 848.400 ;
        RECT 616.950 847.950 619.050 848.400 ;
        RECT 637.950 847.950 640.050 848.400 ;
        RECT 715.950 849.600 718.050 850.050 ;
        RECT 739.950 849.600 742.050 850.050 ;
        RECT 811.950 849.600 814.050 850.050 ;
        RECT 715.950 848.400 814.050 849.600 ;
        RECT 715.950 847.950 718.050 848.400 ;
        RECT 739.950 847.950 742.050 848.400 ;
        RECT 811.950 847.950 814.050 848.400 ;
        RECT 826.950 849.600 829.050 850.050 ;
        RECT 913.950 849.600 916.050 850.050 ;
        RECT 826.950 848.400 916.050 849.600 ;
        RECT 826.950 847.950 829.050 848.400 ;
        RECT 913.950 847.950 916.050 848.400 ;
        RECT 55.950 846.600 58.050 847.050 ;
        RECT 79.950 846.600 82.050 847.050 ;
        RECT 115.950 846.600 118.050 847.050 ;
        RECT 55.950 845.400 118.050 846.600 ;
        RECT 55.950 844.950 58.050 845.400 ;
        RECT 79.950 844.950 82.050 845.400 ;
        RECT 115.950 844.950 118.050 845.400 ;
        RECT 142.950 846.600 145.050 847.050 ;
        RECT 148.950 846.600 151.050 847.050 ;
        RECT 142.950 845.400 151.050 846.600 ;
        RECT 142.950 844.950 145.050 845.400 ;
        RECT 148.950 844.950 151.050 845.400 ;
        RECT 202.950 846.600 205.050 847.050 ;
        RECT 310.950 846.600 313.050 847.050 ;
        RECT 202.950 845.400 313.050 846.600 ;
        RECT 202.950 844.950 205.050 845.400 ;
        RECT 310.950 844.950 313.050 845.400 ;
        RECT 349.950 846.600 352.050 847.050 ;
        RECT 382.950 846.600 385.050 847.050 ;
        RECT 349.950 845.400 385.050 846.600 ;
        RECT 349.950 844.950 352.050 845.400 ;
        RECT 382.950 844.950 385.050 845.400 ;
        RECT 445.950 846.600 448.050 847.050 ;
        RECT 475.950 846.600 478.050 847.050 ;
        RECT 445.950 845.400 478.050 846.600 ;
        RECT 445.950 844.950 448.050 845.400 ;
        RECT 475.950 844.950 478.050 845.400 ;
        RECT 571.950 846.600 574.050 847.050 ;
        RECT 580.950 846.600 583.050 847.050 ;
        RECT 571.950 845.400 583.050 846.600 ;
        RECT 571.950 844.950 574.050 845.400 ;
        RECT 580.950 844.950 583.050 845.400 ;
        RECT 703.950 846.600 706.050 847.050 ;
        RECT 721.950 846.600 724.050 847.050 ;
        RECT 703.950 845.400 724.050 846.600 ;
        RECT 703.950 844.950 706.050 845.400 ;
        RECT 721.950 844.950 724.050 845.400 ;
        RECT 874.950 846.600 877.050 847.050 ;
        RECT 892.950 846.600 895.050 847.050 ;
        RECT 895.950 846.600 898.050 847.050 ;
        RECT 904.950 846.600 907.050 847.050 ;
        RECT 874.950 845.400 907.050 846.600 ;
        RECT 874.950 844.950 877.050 845.400 ;
        RECT 892.950 844.950 895.050 845.400 ;
        RECT 895.950 844.950 898.050 845.400 ;
        RECT 904.950 844.950 907.050 845.400 ;
        RECT 274.950 843.600 277.050 844.050 ;
        RECT 283.950 843.600 286.050 844.050 ;
        RECT 346.950 843.600 349.050 844.050 ;
        RECT 146.400 842.400 189.600 843.600 ;
        RECT 16.950 838.950 19.050 841.050 ;
        RECT 22.950 838.950 25.050 841.050 ;
        RECT 40.950 840.750 43.050 841.200 ;
        RECT 46.950 840.750 49.050 841.200 ;
        RECT 40.950 839.550 49.050 840.750 ;
        RECT 40.950 839.100 43.050 839.550 ;
        RECT 46.950 839.100 49.050 839.550 ;
        RECT 73.950 838.950 76.050 841.050 ;
        RECT 94.950 840.750 97.050 841.200 ;
        RECT 100.950 840.750 103.050 841.200 ;
        RECT 94.950 839.550 103.050 840.750 ;
        RECT 94.950 839.100 97.050 839.550 ;
        RECT 100.950 839.100 103.050 839.550 ;
        RECT 106.950 839.100 109.050 841.200 ;
        RECT 1.950 834.450 4.050 834.900 ;
        RECT 13.950 834.450 16.050 834.900 ;
        RECT 1.950 833.250 16.050 834.450 ;
        RECT 1.950 832.800 4.050 833.250 ;
        RECT 13.950 832.800 16.050 833.250 ;
        RECT 17.400 832.050 18.600 838.950 ;
        RECT 23.400 835.050 24.600 838.950 ;
        RECT 74.400 835.050 75.600 838.950 ;
        RECT 107.400 837.600 108.600 839.100 ;
        RECT 118.950 838.950 121.050 841.050 ;
        RECT 124.950 840.600 127.050 841.200 ;
        RECT 130.950 840.600 133.050 841.050 ;
        RECT 124.950 839.400 133.050 840.600 ;
        RECT 124.950 839.100 127.050 839.400 ;
        RECT 130.950 838.950 133.050 839.400 ;
        RECT 136.950 839.100 139.050 841.200 ;
        RECT 142.950 840.600 145.050 841.200 ;
        RECT 146.400 840.600 147.600 842.400 ;
        RECT 142.950 839.400 147.600 840.600 ;
        RECT 148.950 840.750 151.050 841.200 ;
        RECT 157.950 840.750 160.050 841.200 ;
        RECT 148.950 839.550 160.050 840.750 ;
        RECT 142.950 839.100 145.050 839.400 ;
        RECT 148.950 839.100 151.050 839.550 ;
        RECT 157.950 839.100 160.050 839.550 ;
        RECT 188.400 840.600 189.600 842.400 ;
        RECT 274.950 842.400 349.050 843.600 ;
        RECT 274.950 841.950 277.050 842.400 ;
        RECT 283.950 841.950 286.050 842.400 ;
        RECT 346.950 841.950 349.050 842.400 ;
        RECT 394.950 843.600 397.050 844.050 ;
        RECT 403.950 843.600 406.050 844.050 ;
        RECT 394.950 842.400 406.050 843.600 ;
        RECT 394.950 841.950 397.050 842.400 ;
        RECT 403.950 841.950 406.050 842.400 ;
        RECT 562.950 843.600 565.050 844.050 ;
        RECT 574.950 843.600 577.050 844.050 ;
        RECT 562.950 842.400 577.050 843.600 ;
        RECT 562.950 841.950 565.050 842.400 ;
        RECT 574.950 841.950 577.050 842.400 ;
        RECT 631.950 843.600 634.050 844.050 ;
        RECT 640.950 843.600 643.050 844.050 ;
        RECT 631.950 842.400 643.050 843.600 ;
        RECT 631.950 841.950 634.050 842.400 ;
        RECT 640.950 841.950 643.050 842.400 ;
        RECT 760.950 843.600 763.050 844.050 ;
        RECT 778.950 843.600 781.050 844.050 ;
        RECT 760.950 842.400 781.050 843.600 ;
        RECT 760.950 841.950 763.050 842.400 ;
        RECT 778.950 841.950 781.050 842.400 ;
        RECT 886.950 843.600 889.050 844.050 ;
        RECT 931.950 843.600 934.050 844.050 ;
        RECT 886.950 842.400 934.050 843.600 ;
        RECT 886.950 841.950 889.050 842.400 ;
        RECT 931.950 841.950 934.050 842.400 ;
        RECT 208.950 840.750 211.050 841.200 ;
        RECT 220.950 840.750 223.050 841.200 ;
        RECT 188.400 839.400 201.600 840.600 ;
        RECT 107.400 837.000 111.600 837.600 ;
        RECT 107.400 836.400 112.050 837.000 ;
        RECT 22.950 832.950 25.050 835.050 ;
        RECT 28.950 834.450 31.050 834.900 ;
        RECT 37.950 834.450 40.050 834.900 ;
        RECT 28.950 833.250 40.050 834.450 ;
        RECT 28.950 832.800 31.050 833.250 ;
        RECT 37.950 832.800 40.050 833.250 ;
        RECT 73.950 832.950 76.050 835.050 ;
        RECT 109.950 832.950 112.050 836.400 ;
        RECT 119.400 835.050 120.600 838.950 ;
        RECT 118.950 832.950 121.050 835.050 ;
        RECT 127.950 834.600 130.050 835.050 ;
        RECT 137.400 834.600 138.600 839.100 ;
        RECT 143.400 834.600 144.600 839.100 ;
        RECT 175.950 837.600 178.050 838.050 ;
        RECT 196.950 837.600 199.050 838.050 ;
        RECT 175.950 836.400 199.050 837.600 ;
        RECT 175.950 835.950 178.050 836.400 ;
        RECT 196.950 835.950 199.050 836.400 ;
        RECT 127.950 833.400 138.600 834.600 ;
        RECT 140.400 833.400 144.600 834.600 ;
        RECT 200.400 834.600 201.600 839.400 ;
        RECT 208.950 839.550 223.050 840.750 ;
        RECT 208.950 839.100 211.050 839.550 ;
        RECT 220.950 839.100 223.050 839.550 ;
        RECT 247.950 839.100 250.050 841.200 ;
        RECT 253.950 840.600 256.050 841.200 ;
        RECT 271.950 840.600 274.050 841.200 ;
        RECT 253.950 839.400 274.050 840.600 ;
        RECT 253.950 839.100 256.050 839.400 ;
        RECT 271.950 839.100 274.050 839.400 ;
        RECT 248.400 837.600 249.600 839.100 ;
        RECT 277.950 837.600 280.050 841.050 ;
        RECT 286.950 840.750 289.050 841.200 ;
        RECT 313.950 840.750 316.050 841.200 ;
        RECT 286.950 839.550 316.050 840.750 ;
        RECT 286.950 839.100 289.050 839.550 ;
        RECT 313.950 839.100 316.050 839.550 ;
        RECT 352.950 840.750 355.050 841.200 ;
        RECT 361.950 840.750 364.050 841.200 ;
        RECT 352.950 839.550 364.050 840.750 ;
        RECT 388.950 840.600 391.050 841.200 ;
        RECT 352.950 839.100 355.050 839.550 ;
        RECT 361.950 839.100 364.050 839.550 ;
        RECT 377.400 839.400 391.050 840.600 ;
        RECT 248.400 836.400 252.600 837.600 ;
        RECT 205.950 834.600 208.050 834.900 ;
        RECT 200.400 833.400 208.050 834.600 ;
        RECT 127.950 832.950 130.050 833.400 ;
        RECT 140.400 832.050 141.600 833.400 ;
        RECT 205.950 832.800 208.050 833.400 ;
        RECT 220.950 834.600 223.050 835.050 ;
        RECT 229.950 834.600 232.050 834.900 ;
        RECT 220.950 833.400 232.050 834.600 ;
        RECT 251.400 834.600 252.600 836.400 ;
        RECT 269.400 837.000 280.050 837.600 ;
        RECT 340.950 837.600 343.050 838.050 ;
        RECT 269.400 836.400 279.600 837.000 ;
        RECT 340.950 836.400 354.600 837.600 ;
        RECT 269.400 834.900 270.600 836.400 ;
        RECT 340.950 835.950 343.050 836.400 ;
        RECT 251.400 833.400 264.600 834.600 ;
        RECT 220.950 832.950 223.050 833.400 ;
        RECT 229.950 832.800 232.050 833.400 ;
        RECT 16.950 829.950 19.050 832.050 ;
        RECT 49.950 831.600 52.050 832.050 ;
        RECT 82.800 831.600 84.900 832.050 ;
        RECT 49.950 830.400 84.900 831.600 ;
        RECT 49.950 829.950 52.050 830.400 ;
        RECT 82.800 829.950 84.900 830.400 ;
        RECT 106.950 831.600 109.050 832.050 ;
        RECT 112.950 831.600 115.050 832.050 ;
        RECT 106.950 830.400 115.050 831.600 ;
        RECT 106.950 829.950 109.050 830.400 ;
        RECT 112.950 829.950 115.050 830.400 ;
        RECT 136.950 830.400 141.600 832.050 ;
        RECT 154.950 831.600 157.050 832.050 ;
        RECT 175.950 831.600 178.050 832.050 ;
        RECT 154.950 830.400 178.050 831.600 ;
        RECT 136.950 829.950 141.000 830.400 ;
        RECT 154.950 829.950 157.050 830.400 ;
        RECT 175.950 829.950 178.050 830.400 ;
        RECT 235.950 831.600 238.050 832.050 ;
        RECT 259.950 831.600 262.050 832.050 ;
        RECT 235.950 830.400 262.050 831.600 ;
        RECT 263.400 831.600 264.600 833.400 ;
        RECT 268.950 832.800 271.050 834.900 ;
        RECT 304.950 834.450 307.050 834.900 ;
        RECT 331.950 834.450 334.050 834.900 ;
        RECT 304.950 833.250 334.050 834.450 ;
        RECT 353.400 834.600 354.600 836.400 ;
        RECT 355.950 834.600 358.050 834.900 ;
        RECT 353.400 833.400 358.050 834.600 ;
        RECT 304.950 832.800 307.050 833.250 ;
        RECT 331.950 832.800 334.050 833.250 ;
        RECT 355.950 832.800 358.050 833.400 ;
        RECT 361.950 834.600 364.050 835.050 ;
        RECT 377.400 834.900 378.600 839.400 ;
        RECT 388.950 839.100 391.050 839.400 ;
        RECT 406.950 840.750 409.050 841.200 ;
        RECT 415.950 840.750 418.050 841.200 ;
        RECT 406.950 839.550 418.050 840.750 ;
        RECT 406.950 839.100 409.050 839.550 ;
        RECT 415.950 839.100 418.050 839.550 ;
        RECT 466.950 840.750 469.050 841.200 ;
        RECT 475.950 840.750 478.050 841.200 ;
        RECT 466.950 839.550 478.050 840.750 ;
        RECT 466.950 839.100 469.050 839.550 ;
        RECT 475.950 839.100 478.050 839.550 ;
        RECT 490.950 840.750 493.050 841.200 ;
        RECT 496.950 840.750 499.050 841.200 ;
        RECT 490.950 839.550 499.050 840.750 ;
        RECT 490.950 839.100 493.050 839.550 ;
        RECT 496.950 839.100 499.050 839.550 ;
        RECT 502.950 840.600 505.050 841.200 ;
        RECT 523.950 840.600 526.050 841.200 ;
        RECT 538.950 840.600 541.050 841.200 ;
        RECT 502.950 839.400 526.050 840.600 ;
        RECT 502.950 839.100 505.050 839.400 ;
        RECT 523.950 839.100 526.050 839.400 ;
        RECT 527.400 839.400 541.050 840.600 ;
        RECT 491.400 837.600 492.600 839.100 ;
        RECT 434.400 836.400 492.600 837.600 ;
        RECT 434.400 834.900 435.600 836.400 ;
        RECT 370.950 834.600 373.050 834.900 ;
        RECT 361.950 833.400 373.050 834.600 ;
        RECT 361.950 832.950 364.050 833.400 ;
        RECT 370.950 832.800 373.050 833.400 ;
        RECT 376.950 832.800 379.050 834.900 ;
        RECT 391.950 834.450 394.050 834.900 ;
        RECT 409.950 834.450 412.050 834.900 ;
        RECT 391.950 833.250 412.050 834.450 ;
        RECT 391.950 832.800 394.050 833.250 ;
        RECT 409.950 832.800 412.050 833.250 ;
        RECT 433.950 832.800 436.050 834.900 ;
        RECT 439.950 834.450 442.050 834.900 ;
        RECT 445.950 834.450 448.050 834.900 ;
        RECT 439.950 833.250 448.050 834.450 ;
        RECT 439.950 832.800 442.050 833.250 ;
        RECT 445.950 832.800 448.050 833.250 ;
        RECT 457.950 834.600 460.050 834.900 ;
        RECT 466.800 834.600 468.900 835.050 ;
        RECT 457.950 833.400 468.900 834.600 ;
        RECT 457.950 832.800 460.050 833.400 ;
        RECT 466.800 832.950 468.900 833.400 ;
        RECT 469.950 834.600 472.050 835.050 ;
        RECT 478.950 834.600 481.050 834.900 ;
        RECT 469.950 833.400 481.050 834.600 ;
        RECT 469.950 832.950 472.050 833.400 ;
        RECT 478.950 832.800 481.050 833.400 ;
        RECT 493.950 834.600 496.050 835.050 ;
        RECT 527.400 834.900 528.600 839.400 ;
        RECT 538.950 839.100 541.050 839.400 ;
        RECT 544.950 838.950 547.050 841.050 ;
        RECT 553.950 839.100 556.050 841.200 ;
        RECT 559.950 839.100 562.050 841.200 ;
        RECT 583.950 840.600 586.050 841.050 ;
        RECT 578.400 839.400 586.050 840.600 ;
        RECT 545.400 835.050 546.600 838.950 ;
        RECT 554.400 835.050 555.600 839.100 ;
        RECT 499.950 834.600 502.050 834.900 ;
        RECT 493.950 833.400 502.050 834.600 ;
        RECT 493.950 832.950 496.050 833.400 ;
        RECT 499.950 832.800 502.050 833.400 ;
        RECT 526.950 832.800 529.050 834.900 ;
        RECT 544.950 832.950 547.050 835.050 ;
        RECT 550.950 833.400 555.600 835.050 ;
        RECT 560.400 835.050 561.600 839.100 ;
        RECT 560.400 833.400 565.050 835.050 ;
        RECT 578.400 834.900 579.600 839.400 ;
        RECT 583.950 838.950 586.050 839.400 ;
        RECT 589.950 840.750 592.050 841.200 ;
        RECT 595.950 840.750 598.050 841.200 ;
        RECT 589.950 839.550 598.050 840.750 ;
        RECT 589.950 839.100 592.050 839.550 ;
        RECT 595.950 839.100 598.050 839.550 ;
        RECT 607.950 838.950 610.050 841.050 ;
        RECT 622.950 840.750 625.050 841.200 ;
        RECT 628.950 840.750 631.050 841.200 ;
        RECT 622.950 839.550 631.050 840.750 ;
        RECT 622.950 839.100 625.050 839.550 ;
        RECT 628.950 839.100 631.050 839.550 ;
        RECT 637.950 839.100 640.050 841.200 ;
        RECT 661.950 840.600 664.050 841.200 ;
        RECT 676.950 840.600 679.050 841.200 ;
        RECT 661.950 839.400 679.050 840.600 ;
        RECT 661.950 839.100 664.050 839.400 ;
        RECT 676.950 839.100 679.050 839.400 ;
        RECT 682.950 840.750 685.050 841.200 ;
        RECT 694.950 840.750 697.050 841.200 ;
        RECT 682.950 839.550 697.050 840.750 ;
        RECT 682.950 839.100 685.050 839.550 ;
        RECT 694.950 839.100 697.050 839.550 ;
        RECT 721.950 840.600 724.050 841.200 ;
        RECT 730.950 840.600 733.050 841.050 ;
        RECT 721.950 839.400 733.050 840.600 ;
        RECT 721.950 839.100 724.050 839.400 ;
        RECT 550.950 832.950 555.000 833.400 ;
        RECT 561.000 832.950 565.050 833.400 ;
        RECT 577.950 832.800 580.050 834.900 ;
        RECT 608.400 834.600 609.600 838.950 ;
        RECT 638.400 837.600 639.600 839.100 ;
        RECT 730.950 838.950 733.050 839.400 ;
        RECT 745.950 840.750 748.050 841.200 ;
        RECT 754.950 840.750 757.050 841.200 ;
        RECT 745.950 839.550 757.050 840.750 ;
        RECT 745.950 839.100 748.050 839.550 ;
        RECT 754.950 839.100 757.050 839.550 ;
        RECT 766.950 840.600 769.050 841.050 ;
        RECT 775.950 840.600 778.050 841.200 ;
        RECT 796.950 840.600 799.050 841.200 ;
        RECT 766.950 839.400 778.050 840.600 ;
        RECT 766.950 838.950 769.050 839.400 ;
        RECT 775.950 839.100 778.050 839.400 ;
        RECT 794.400 839.400 799.050 840.600 ;
        RECT 769.950 837.600 772.050 838.050 ;
        RECT 794.400 837.600 795.600 839.400 ;
        RECT 796.950 839.100 799.050 839.400 ;
        RECT 841.950 840.600 844.050 841.200 ;
        RECT 865.950 840.600 868.050 841.200 ;
        RECT 841.950 839.400 868.050 840.600 ;
        RECT 841.950 839.100 844.050 839.400 ;
        RECT 865.950 839.100 868.050 839.400 ;
        RECT 871.950 839.100 874.050 841.200 ;
        RECT 638.400 836.400 657.600 837.600 ;
        RECT 656.400 834.900 657.600 836.400 ;
        RECT 769.950 836.400 795.600 837.600 ;
        RECT 769.950 835.950 772.050 836.400 ;
        RECT 872.400 835.050 873.600 839.100 ;
        RECT 619.950 834.600 622.050 834.900 ;
        RECT 608.400 833.400 622.050 834.600 ;
        RECT 619.950 832.800 622.050 833.400 ;
        RECT 655.800 832.800 657.900 834.900 ;
        RECT 658.950 834.600 661.050 835.050 ;
        RECT 679.950 834.600 682.050 834.900 ;
        RECT 658.950 833.400 682.050 834.600 ;
        RECT 658.950 832.950 661.050 833.400 ;
        RECT 679.950 832.800 682.050 833.400 ;
        RECT 697.950 834.600 700.050 834.900 ;
        RECT 715.950 834.600 718.050 834.900 ;
        RECT 697.950 833.400 718.050 834.600 ;
        RECT 697.950 832.800 700.050 833.400 ;
        RECT 715.950 832.800 718.050 833.400 ;
        RECT 730.950 834.450 733.050 834.900 ;
        RECT 736.950 834.450 739.050 834.900 ;
        RECT 730.950 833.250 739.050 834.450 ;
        RECT 730.950 832.800 733.050 833.250 ;
        RECT 736.950 832.800 739.050 833.250 ;
        RECT 757.950 834.450 760.050 834.900 ;
        RECT 766.950 834.450 769.050 834.900 ;
        RECT 757.950 833.250 769.050 834.450 ;
        RECT 757.950 832.800 760.050 833.250 ;
        RECT 766.950 832.800 769.050 833.250 ;
        RECT 799.950 834.450 802.050 834.900 ;
        RECT 808.950 834.450 811.050 834.900 ;
        RECT 799.950 833.250 811.050 834.450 ;
        RECT 799.950 832.800 802.050 833.250 ;
        RECT 808.950 832.800 811.050 833.250 ;
        RECT 823.950 834.450 826.050 834.900 ;
        RECT 832.950 834.450 835.050 834.900 ;
        RECT 823.950 833.250 835.050 834.450 ;
        RECT 823.950 832.800 826.050 833.250 ;
        RECT 832.950 832.800 835.050 833.250 ;
        RECT 856.950 834.450 859.050 834.900 ;
        RECT 862.950 834.450 865.050 834.900 ;
        RECT 856.950 833.250 865.050 834.450 ;
        RECT 872.400 833.400 877.050 835.050 ;
        RECT 856.950 832.800 859.050 833.250 ;
        RECT 862.950 832.800 865.050 833.250 ;
        RECT 873.000 832.950 877.050 833.400 ;
        RECT 889.950 834.450 892.050 834.900 ;
        RECT 898.950 834.450 901.050 834.900 ;
        RECT 889.950 833.250 901.050 834.450 ;
        RECT 889.950 832.800 892.050 833.250 ;
        RECT 898.950 832.800 901.050 833.250 ;
        RECT 292.950 831.600 295.050 832.050 ;
        RECT 263.400 830.400 295.050 831.600 ;
        RECT 235.950 829.950 238.050 830.400 ;
        RECT 259.950 829.950 262.050 830.400 ;
        RECT 292.950 829.950 295.050 830.400 ;
        RECT 403.950 831.600 406.050 832.050 ;
        RECT 418.950 831.600 421.050 832.050 ;
        RECT 403.950 830.400 421.050 831.600 ;
        RECT 403.950 829.950 406.050 830.400 ;
        RECT 418.950 829.950 421.050 830.400 ;
        RECT 448.950 831.600 451.050 832.050 ;
        RECT 454.950 831.600 457.050 832.050 ;
        RECT 448.950 830.400 457.050 831.600 ;
        RECT 448.950 829.950 451.050 830.400 ;
        RECT 454.950 829.950 457.050 830.400 ;
        RECT 547.950 831.600 550.050 832.050 ;
        RECT 556.950 831.600 559.050 832.050 ;
        RECT 547.950 830.400 559.050 831.600 ;
        RECT 547.950 829.950 550.050 830.400 ;
        RECT 556.950 829.950 559.050 830.400 ;
        RECT 19.950 828.600 22.050 829.050 ;
        RECT 25.950 828.600 28.050 829.050 ;
        RECT 19.950 827.400 28.050 828.600 ;
        RECT 19.950 826.950 22.050 827.400 ;
        RECT 25.950 826.950 28.050 827.400 ;
        RECT 61.950 828.600 64.050 829.050 ;
        RECT 79.950 828.600 82.050 829.050 ;
        RECT 61.950 827.400 82.050 828.600 ;
        RECT 61.950 826.950 64.050 827.400 ;
        RECT 79.950 826.950 82.050 827.400 ;
        RECT 97.950 828.600 100.050 829.050 ;
        RECT 130.800 828.600 132.900 829.050 ;
        RECT 97.950 827.400 132.900 828.600 ;
        RECT 97.950 826.950 100.050 827.400 ;
        RECT 130.800 826.950 132.900 827.400 ;
        RECT 133.950 828.600 136.050 829.050 ;
        RECT 145.950 828.600 148.050 829.050 ;
        RECT 133.950 827.400 148.050 828.600 ;
        RECT 133.950 826.950 136.050 827.400 ;
        RECT 145.950 826.950 148.050 827.400 ;
        RECT 151.950 828.600 154.050 829.050 ;
        RECT 187.950 828.600 190.050 829.050 ;
        RECT 151.950 827.400 190.050 828.600 ;
        RECT 151.950 826.950 154.050 827.400 ;
        RECT 187.950 826.950 190.050 827.400 ;
        RECT 232.950 828.600 235.050 829.050 ;
        RECT 262.950 828.600 265.050 829.050 ;
        RECT 472.950 828.600 475.050 829.050 ;
        RECT 484.950 828.600 487.050 829.050 ;
        RECT 232.950 828.000 294.450 828.600 ;
        RECT 232.950 827.400 295.050 828.000 ;
        RECT 232.950 826.950 235.050 827.400 ;
        RECT 262.950 826.950 265.050 827.400 ;
        RECT 55.950 825.600 58.050 826.050 ;
        RECT 98.400 825.600 99.600 826.950 ;
        RECT 292.950 826.050 295.050 827.400 ;
        RECT 472.950 827.400 487.050 828.600 ;
        RECT 472.950 826.950 475.050 827.400 ;
        RECT 484.950 826.950 487.050 827.400 ;
        RECT 568.950 828.600 571.050 829.050 ;
        RECT 583.950 828.600 586.050 829.050 ;
        RECT 568.950 827.400 586.050 828.600 ;
        RECT 568.950 826.950 571.050 827.400 ;
        RECT 583.950 826.950 586.050 827.400 ;
        RECT 628.950 828.600 631.050 829.050 ;
        RECT 658.950 828.600 661.050 829.050 ;
        RECT 628.950 827.400 661.050 828.600 ;
        RECT 628.950 826.950 631.050 827.400 ;
        RECT 658.950 826.950 661.050 827.400 ;
        RECT 670.950 828.600 673.050 829.050 ;
        RECT 697.950 828.600 700.050 829.050 ;
        RECT 670.950 827.400 700.050 828.600 ;
        RECT 670.950 826.950 673.050 827.400 ;
        RECT 697.950 826.950 700.050 827.400 ;
        RECT 703.950 828.600 706.050 829.050 ;
        RECT 727.950 828.600 730.050 829.050 ;
        RECT 703.950 827.400 730.050 828.600 ;
        RECT 703.950 826.950 706.050 827.400 ;
        RECT 727.950 826.950 730.050 827.400 ;
        RECT 787.950 828.600 790.050 829.050 ;
        RECT 811.950 828.600 814.050 829.050 ;
        RECT 787.950 827.400 814.050 828.600 ;
        RECT 787.950 826.950 790.050 827.400 ;
        RECT 811.950 826.950 814.050 827.400 ;
        RECT 838.950 828.600 841.050 829.050 ;
        RECT 853.950 828.600 856.050 829.050 ;
        RECT 838.950 827.400 856.050 828.600 ;
        RECT 838.950 826.950 841.050 827.400 ;
        RECT 853.950 826.950 856.050 827.400 ;
        RECT 883.950 828.600 886.050 829.050 ;
        RECT 928.950 828.600 931.050 829.050 ;
        RECT 883.950 827.400 931.050 828.600 ;
        RECT 883.950 826.950 886.050 827.400 ;
        RECT 928.950 826.950 931.050 827.400 ;
        RECT 55.950 824.400 99.600 825.600 ;
        RECT 130.950 825.600 133.050 825.900 ;
        RECT 250.950 825.600 253.050 826.050 ;
        RECT 130.950 824.400 253.050 825.600 ;
        RECT 55.950 823.950 58.050 824.400 ;
        RECT 130.950 823.800 133.050 824.400 ;
        RECT 250.950 823.950 253.050 824.400 ;
        RECT 274.950 825.600 277.050 826.050 ;
        RECT 286.950 825.600 289.050 826.050 ;
        RECT 274.950 824.400 289.050 825.600 ;
        RECT 274.950 823.950 277.050 824.400 ;
        RECT 286.950 823.950 289.050 824.400 ;
        RECT 292.800 825.000 295.050 826.050 ;
        RECT 295.950 825.600 298.050 826.050 ;
        RECT 337.950 825.600 340.050 826.050 ;
        RECT 292.800 823.950 294.900 825.000 ;
        RECT 295.950 824.400 340.050 825.600 ;
        RECT 295.950 823.950 298.050 824.400 ;
        RECT 337.950 823.950 340.050 824.400 ;
        RECT 382.950 825.600 385.050 826.050 ;
        RECT 406.950 825.600 409.050 826.050 ;
        RECT 382.950 824.400 409.050 825.600 ;
        RECT 382.950 823.950 385.050 824.400 ;
        RECT 406.950 823.950 409.050 824.400 ;
        RECT 562.950 825.600 565.050 826.050 ;
        RECT 598.950 825.600 601.050 826.050 ;
        RECT 562.950 824.400 601.050 825.600 ;
        RECT 562.950 823.950 565.050 824.400 ;
        RECT 598.950 823.950 601.050 824.400 ;
        RECT 688.950 825.600 691.050 826.050 ;
        RECT 745.950 825.600 748.050 826.050 ;
        RECT 778.950 825.600 781.050 826.050 ;
        RECT 688.950 824.400 781.050 825.600 ;
        RECT 688.950 823.950 691.050 824.400 ;
        RECT 745.950 823.950 748.050 824.400 ;
        RECT 778.950 823.950 781.050 824.400 ;
        RECT 784.950 825.600 787.050 826.050 ;
        RECT 814.950 825.600 817.050 826.050 ;
        RECT 784.950 824.400 817.050 825.600 ;
        RECT 784.950 823.950 787.050 824.400 ;
        RECT 814.950 823.950 817.050 824.400 ;
        RECT 832.950 825.600 835.050 826.050 ;
        RECT 868.950 825.600 871.050 826.050 ;
        RECT 832.950 824.400 871.050 825.600 ;
        RECT 832.950 823.950 835.050 824.400 ;
        RECT 868.950 823.950 871.050 824.400 ;
        RECT 46.950 822.600 49.050 823.050 ;
        RECT 58.950 822.600 61.050 823.050 ;
        RECT 46.950 821.400 61.050 822.600 ;
        RECT 46.950 820.950 49.050 821.400 ;
        RECT 58.950 820.950 61.050 821.400 ;
        RECT 124.950 822.600 127.050 823.050 ;
        RECT 169.950 822.600 172.050 823.050 ;
        RECT 124.950 821.400 172.050 822.600 ;
        RECT 124.950 820.950 127.050 821.400 ;
        RECT 169.950 820.950 172.050 821.400 ;
        RECT 238.950 822.600 241.050 823.050 ;
        RECT 298.950 822.600 301.050 823.050 ;
        RECT 238.950 821.400 301.050 822.600 ;
        RECT 238.950 820.950 241.050 821.400 ;
        RECT 298.950 820.950 301.050 821.400 ;
        RECT 376.950 822.600 379.050 823.050 ;
        RECT 412.950 822.600 415.050 823.050 ;
        RECT 376.950 821.400 415.050 822.600 ;
        RECT 376.950 820.950 379.050 821.400 ;
        RECT 412.950 820.950 415.050 821.400 ;
        RECT 439.950 822.600 442.050 823.050 ;
        RECT 472.950 822.600 475.050 823.050 ;
        RECT 439.950 821.400 475.050 822.600 ;
        RECT 439.950 820.950 442.050 821.400 ;
        RECT 472.950 820.950 475.050 821.400 ;
        RECT 694.950 822.600 697.050 823.050 ;
        RECT 700.950 822.600 703.050 823.050 ;
        RECT 694.950 821.400 703.050 822.600 ;
        RECT 694.950 820.950 697.050 821.400 ;
        RECT 700.950 820.950 703.050 821.400 ;
        RECT 805.950 822.600 808.050 823.050 ;
        RECT 817.950 822.600 820.050 823.050 ;
        RECT 826.950 822.600 829.050 823.050 ;
        RECT 805.950 821.400 829.050 822.600 ;
        RECT 805.950 820.950 808.050 821.400 ;
        RECT 817.950 820.950 820.050 821.400 ;
        RECT 826.950 820.950 829.050 821.400 ;
        RECT 880.950 822.600 883.050 823.050 ;
        RECT 919.950 822.600 922.050 823.050 ;
        RECT 880.950 821.400 922.050 822.600 ;
        RECT 880.950 820.950 883.050 821.400 ;
        RECT 919.950 820.950 922.050 821.400 ;
        RECT 7.950 819.600 10.050 820.050 ;
        RECT 70.950 819.600 73.050 820.050 ;
        RECT 166.950 819.600 169.050 820.050 ;
        RECT 7.950 818.400 169.050 819.600 ;
        RECT 7.950 817.950 10.050 818.400 ;
        RECT 70.950 817.950 73.050 818.400 ;
        RECT 166.950 817.950 169.050 818.400 ;
        RECT 268.950 819.600 271.050 820.050 ;
        RECT 280.950 819.600 283.050 820.050 ;
        RECT 268.950 818.400 283.050 819.600 ;
        RECT 268.950 817.950 271.050 818.400 ;
        RECT 280.950 817.950 283.050 818.400 ;
        RECT 286.950 819.600 289.050 820.050 ;
        RECT 295.950 819.600 298.050 820.050 ;
        RECT 286.950 818.400 298.050 819.600 ;
        RECT 286.950 817.950 289.050 818.400 ;
        RECT 295.950 817.950 298.050 818.400 ;
        RECT 424.950 819.600 427.050 820.050 ;
        RECT 487.800 819.600 489.900 820.050 ;
        RECT 424.950 818.400 489.900 819.600 ;
        RECT 424.950 817.950 427.050 818.400 ;
        RECT 487.800 817.950 489.900 818.400 ;
        RECT 490.950 819.600 493.050 820.050 ;
        RECT 523.950 819.600 526.050 820.050 ;
        RECT 550.800 819.600 552.900 820.050 ;
        RECT 490.950 818.400 552.900 819.600 ;
        RECT 490.950 817.950 493.050 818.400 ;
        RECT 523.950 817.950 526.050 818.400 ;
        RECT 550.800 817.950 552.900 818.400 ;
        RECT 628.950 819.600 631.050 820.050 ;
        RECT 640.950 819.600 643.050 820.050 ;
        RECT 691.950 819.600 694.050 820.050 ;
        RECT 628.950 818.400 694.050 819.600 ;
        RECT 628.950 817.950 631.050 818.400 ;
        RECT 640.950 817.950 643.050 818.400 ;
        RECT 691.950 817.950 694.050 818.400 ;
        RECT 766.950 819.600 769.050 820.050 ;
        RECT 856.950 819.600 859.050 820.050 ;
        RECT 766.950 818.400 859.050 819.600 ;
        RECT 766.950 817.950 769.050 818.400 ;
        RECT 856.950 817.950 859.050 818.400 ;
        RECT 106.950 816.600 109.050 817.050 ;
        RECT 139.950 816.600 142.050 817.050 ;
        RECT 205.950 816.600 208.050 817.050 ;
        RECT 106.950 815.400 142.050 816.600 ;
        RECT 106.950 814.950 109.050 815.400 ;
        RECT 139.950 814.950 142.050 815.400 ;
        RECT 194.400 815.400 208.050 816.600 ;
        RECT 194.400 814.050 195.600 815.400 ;
        RECT 205.950 814.950 208.050 815.400 ;
        RECT 277.950 816.600 280.050 817.050 ;
        RECT 283.950 816.600 286.050 817.050 ;
        RECT 277.950 815.400 286.050 816.600 ;
        RECT 277.950 814.950 280.050 815.400 ;
        RECT 283.950 814.950 286.050 815.400 ;
        RECT 304.950 816.600 307.050 817.050 ;
        RECT 373.950 816.600 376.050 817.050 ;
        RECT 304.950 815.400 376.050 816.600 ;
        RECT 304.950 814.950 307.050 815.400 ;
        RECT 373.950 814.950 376.050 815.400 ;
        RECT 445.950 816.600 448.050 817.050 ;
        RECT 508.950 816.600 511.050 817.050 ;
        RECT 445.950 815.400 511.050 816.600 ;
        RECT 445.950 814.950 448.050 815.400 ;
        RECT 508.950 814.950 511.050 815.400 ;
        RECT 571.950 816.600 574.050 817.050 ;
        RECT 625.950 816.600 628.050 817.050 ;
        RECT 571.950 815.400 628.050 816.600 ;
        RECT 571.950 814.950 574.050 815.400 ;
        RECT 625.950 814.950 628.050 815.400 ;
        RECT 718.950 816.600 721.050 817.050 ;
        RECT 733.950 816.600 736.050 817.050 ;
        RECT 718.950 815.400 736.050 816.600 ;
        RECT 718.950 814.950 721.050 815.400 ;
        RECT 733.950 814.950 736.050 815.400 ;
        RECT 751.950 816.600 754.050 817.050 ;
        RECT 784.950 816.600 787.050 817.050 ;
        RECT 751.950 815.400 787.050 816.600 ;
        RECT 751.950 814.950 754.050 815.400 ;
        RECT 784.950 814.950 787.050 815.400 ;
        RECT 796.950 816.600 799.050 817.050 ;
        RECT 847.950 816.600 850.050 817.050 ;
        RECT 796.950 815.400 850.050 816.600 ;
        RECT 796.950 814.950 799.050 815.400 ;
        RECT 847.950 814.950 850.050 815.400 ;
        RECT 31.950 813.600 34.050 814.050 ;
        RECT 64.950 813.600 67.050 814.050 ;
        RECT 31.950 812.400 67.050 813.600 ;
        RECT 31.950 811.950 34.050 812.400 ;
        RECT 64.950 811.950 67.050 812.400 ;
        RECT 139.950 813.600 142.050 813.900 ;
        RECT 193.950 813.600 196.050 814.050 ;
        RECT 139.950 812.400 196.050 813.600 ;
        RECT 139.950 811.800 142.050 812.400 ;
        RECT 193.950 811.950 196.050 812.400 ;
        RECT 217.950 813.600 220.050 814.050 ;
        RECT 223.950 813.600 226.050 814.050 ;
        RECT 238.950 813.600 241.050 814.050 ;
        RECT 217.950 812.400 226.050 813.600 ;
        RECT 217.950 811.950 220.050 812.400 ;
        RECT 223.950 811.950 226.050 812.400 ;
        RECT 227.400 812.400 241.050 813.600 ;
        RECT 22.950 811.050 25.050 811.200 ;
        RECT 21.000 810.600 25.050 811.050 ;
        RECT 20.400 809.100 25.050 810.600 ;
        RECT 82.950 810.600 85.050 811.050 ;
        RECT 118.950 810.600 121.050 811.050 ;
        RECT 136.950 810.600 139.050 811.050 ;
        RECT 82.950 809.400 121.050 810.600 ;
        RECT 20.400 808.950 24.000 809.100 ;
        RECT 82.950 808.950 85.050 809.400 ;
        RECT 16.950 806.100 19.050 808.200 ;
        RECT 10.950 801.600 13.050 802.050 ;
        RECT 17.400 801.600 18.600 806.100 ;
        RECT 20.400 801.900 21.600 808.950 ;
        RECT 22.950 807.600 25.050 808.050 ;
        RECT 40.950 807.600 43.050 808.200 ;
        RECT 22.950 806.400 43.050 807.600 ;
        RECT 22.950 805.950 25.050 806.400 ;
        RECT 40.950 806.100 43.050 806.400 ;
        RECT 58.950 807.600 61.050 808.200 ;
        RECT 64.950 807.600 67.050 808.050 ;
        RECT 97.950 807.600 100.050 808.200 ;
        RECT 58.950 806.400 67.050 807.600 ;
        RECT 58.950 806.100 61.050 806.400 ;
        RECT 64.950 805.950 67.050 806.400 ;
        RECT 92.400 806.400 100.050 807.600 ;
        RECT 92.400 802.050 93.600 806.400 ;
        RECT 97.950 806.100 100.050 806.400 ;
        RECT 10.950 800.400 18.600 801.600 ;
        RECT 10.950 799.950 13.050 800.400 ;
        RECT 19.950 799.800 22.050 801.900 ;
        RECT 37.950 801.450 40.050 801.900 ;
        RECT 49.800 801.450 51.900 801.900 ;
        RECT 37.950 800.250 51.900 801.450 ;
        RECT 37.950 799.800 40.050 800.250 ;
        RECT 49.800 799.800 51.900 800.250 ;
        RECT 61.950 801.600 64.050 801.900 ;
        RECT 79.950 801.600 82.050 801.900 ;
        RECT 61.950 800.400 82.050 801.600 ;
        RECT 61.950 799.800 64.050 800.400 ;
        RECT 79.950 799.800 82.050 800.400 ;
        RECT 91.950 799.950 94.050 802.050 ;
        RECT 101.400 801.900 102.600 809.400 ;
        RECT 118.950 808.950 121.050 809.400 ;
        RECT 125.400 809.400 139.050 810.600 ;
        RECT 125.400 807.600 126.600 809.400 ;
        RECT 136.950 808.950 139.050 809.400 ;
        RECT 196.950 810.600 199.050 811.050 ;
        RECT 227.400 810.600 228.600 812.400 ;
        RECT 238.950 811.950 241.050 812.400 ;
        RECT 250.950 813.600 253.050 814.050 ;
        RECT 262.950 813.600 265.050 814.050 ;
        RECT 325.950 813.600 328.050 814.050 ;
        RECT 250.950 812.400 265.050 813.600 ;
        RECT 250.950 811.950 253.050 812.400 ;
        RECT 262.950 811.950 265.050 812.400 ;
        RECT 287.400 812.400 328.050 813.600 ;
        RECT 231.000 810.600 235.050 811.050 ;
        RECT 287.400 810.600 288.600 812.400 ;
        RECT 325.950 811.950 328.050 812.400 ;
        RECT 385.950 813.600 388.050 814.050 ;
        RECT 397.950 813.600 400.050 814.050 ;
        RECT 385.950 812.400 400.050 813.600 ;
        RECT 385.950 811.950 388.050 812.400 ;
        RECT 397.950 811.950 400.050 812.400 ;
        RECT 487.950 813.600 490.050 814.050 ;
        RECT 520.950 813.600 523.050 814.050 ;
        RECT 487.950 812.400 523.050 813.600 ;
        RECT 487.950 811.950 490.050 812.400 ;
        RECT 520.950 811.950 523.050 812.400 ;
        RECT 529.950 813.600 532.050 814.050 ;
        RECT 559.950 813.600 562.050 814.050 ;
        RECT 529.950 812.400 562.050 813.600 ;
        RECT 529.950 811.950 532.050 812.400 ;
        RECT 559.950 811.950 562.050 812.400 ;
        RECT 601.950 813.600 604.050 814.050 ;
        RECT 613.950 813.600 616.050 814.050 ;
        RECT 601.950 812.400 616.050 813.600 ;
        RECT 601.950 811.950 604.050 812.400 ;
        RECT 613.950 811.950 616.050 812.400 ;
        RECT 673.950 813.600 676.050 814.050 ;
        RECT 703.950 813.600 706.050 814.050 ;
        RECT 673.950 812.400 706.050 813.600 ;
        RECT 673.950 811.950 676.050 812.400 ;
        RECT 703.950 811.950 706.050 812.400 ;
        RECT 196.950 809.400 228.600 810.600 ;
        RECT 196.950 808.950 199.050 809.400 ;
        RECT 230.400 808.950 235.050 810.600 ;
        RECT 254.400 809.400 288.600 810.600 ;
        RECT 301.950 810.600 304.050 811.050 ;
        RECT 313.950 810.600 316.050 811.050 ;
        RECT 301.950 809.400 316.050 810.600 ;
        RECT 122.400 806.400 126.600 807.600 ;
        RECT 148.950 807.750 151.050 808.200 ;
        RECT 157.950 807.750 160.050 808.200 ;
        RECT 148.950 806.550 160.050 807.750 ;
        RECT 122.400 801.900 123.600 806.400 ;
        RECT 148.950 806.100 151.050 806.550 ;
        RECT 157.950 806.100 160.050 806.550 ;
        RECT 163.950 807.750 166.050 808.200 ;
        RECT 184.950 807.750 187.050 808.200 ;
        RECT 163.950 806.550 187.050 807.750 ;
        RECT 163.950 806.100 166.050 806.550 ;
        RECT 184.950 806.100 187.050 806.550 ;
        RECT 205.950 807.600 210.000 808.050 ;
        RECT 211.950 807.600 214.050 808.050 ;
        RECT 230.400 807.600 231.600 808.950 ;
        RECT 205.950 805.950 210.600 807.600 ;
        RECT 211.950 806.400 231.600 807.600 ;
        RECT 238.950 807.600 241.050 808.200 ;
        RECT 254.400 807.600 255.600 809.400 ;
        RECT 301.950 808.950 304.050 809.400 ;
        RECT 313.950 808.950 316.050 809.400 ;
        RECT 427.950 810.600 430.050 811.050 ;
        RECT 433.950 810.600 436.050 811.050 ;
        RECT 427.950 809.400 436.050 810.600 ;
        RECT 427.950 808.950 430.050 809.400 ;
        RECT 433.950 808.950 436.050 809.400 ;
        RECT 481.950 808.950 484.050 811.050 ;
        RECT 535.950 810.600 538.050 811.200 ;
        RECT 541.950 810.600 544.050 811.050 ;
        RECT 535.950 809.400 544.050 810.600 ;
        RECT 535.950 809.100 538.050 809.400 ;
        RECT 541.950 808.950 544.050 809.400 ;
        RECT 586.950 810.600 589.050 811.050 ;
        RECT 595.950 810.600 598.050 811.050 ;
        RECT 586.950 809.400 598.050 810.600 ;
        RECT 586.950 808.950 589.050 809.400 ;
        RECT 595.950 808.950 598.050 809.400 ;
        RECT 727.950 810.600 730.050 811.050 ;
        RECT 757.950 810.600 760.050 811.050 ;
        RECT 727.950 809.400 760.050 810.600 ;
        RECT 727.950 808.950 730.050 809.400 ;
        RECT 757.950 808.950 760.050 809.400 ;
        RECT 826.950 810.600 829.050 811.050 ;
        RECT 841.800 810.600 843.900 811.050 ;
        RECT 826.950 809.400 843.900 810.600 ;
        RECT 826.950 808.950 829.050 809.400 ;
        RECT 841.800 808.950 843.900 809.400 ;
        RECT 844.950 808.950 847.050 811.050 ;
        RECT 895.950 810.600 898.050 811.050 ;
        RECT 904.950 810.600 907.050 811.050 ;
        RECT 895.950 809.400 907.050 810.600 ;
        RECT 895.950 808.950 898.050 809.400 ;
        RECT 904.950 808.950 907.050 809.400 ;
        RECT 910.950 810.600 913.050 811.050 ;
        RECT 922.950 810.600 925.050 811.050 ;
        RECT 910.950 809.400 925.050 810.600 ;
        RECT 910.950 808.950 913.050 809.400 ;
        RECT 922.950 808.950 925.050 809.400 ;
        RECT 238.950 806.400 255.600 807.600 ;
        RECT 211.950 805.950 214.050 806.400 ;
        RECT 238.950 806.100 241.050 806.400 ;
        RECT 256.950 806.100 259.050 808.200 ;
        RECT 209.400 804.600 210.600 805.950 ;
        RECT 239.400 804.600 240.600 806.100 ;
        RECT 209.400 803.400 237.600 804.600 ;
        RECT 239.400 803.400 246.600 804.600 ;
        RECT 100.950 799.800 103.050 801.900 ;
        RECT 106.950 801.450 109.050 801.900 ;
        RECT 115.950 801.450 118.050 801.900 ;
        RECT 106.950 800.250 118.050 801.450 ;
        RECT 106.950 799.800 109.050 800.250 ;
        RECT 115.950 799.800 118.050 800.250 ;
        RECT 121.950 799.800 124.050 801.900 ;
        RECT 136.950 801.600 139.050 801.900 ;
        RECT 154.950 801.600 157.050 801.900 ;
        RECT 136.950 800.400 157.050 801.600 ;
        RECT 136.950 799.800 139.050 800.400 ;
        RECT 154.950 799.800 157.050 800.400 ;
        RECT 160.950 801.450 163.050 801.900 ;
        RECT 172.950 801.450 175.050 801.900 ;
        RECT 160.950 800.250 175.050 801.450 ;
        RECT 160.950 799.800 163.050 800.250 ;
        RECT 172.950 799.800 175.050 800.250 ;
        RECT 187.950 801.600 190.050 802.050 ;
        RECT 236.400 801.900 237.600 803.400 ;
        RECT 193.950 801.600 196.050 801.900 ;
        RECT 187.950 800.400 196.050 801.600 ;
        RECT 187.950 799.950 190.050 800.400 ;
        RECT 193.950 799.800 196.050 800.400 ;
        RECT 202.950 801.450 205.050 801.900 ;
        RECT 208.950 801.450 211.050 801.900 ;
        RECT 202.950 800.250 211.050 801.450 ;
        RECT 202.950 799.800 205.050 800.250 ;
        RECT 208.950 799.800 211.050 800.250 ;
        RECT 235.950 799.800 238.050 801.900 ;
        RECT 241.950 799.800 244.050 801.900 ;
        RECT 245.400 801.600 246.600 803.400 ;
        RECT 253.950 801.600 256.050 802.050 ;
        RECT 245.400 800.400 256.050 801.600 ;
        RECT 253.950 799.950 256.050 800.400 ;
        RECT 223.950 798.600 226.050 799.050 ;
        RECT 242.400 798.600 243.600 799.800 ;
        RECT 250.950 798.600 253.050 799.050 ;
        RECT 223.950 797.400 243.600 798.600 ;
        RECT 245.400 797.400 253.050 798.600 ;
        RECT 257.400 798.600 258.600 806.100 ;
        RECT 277.950 805.950 280.050 808.050 ;
        RECT 289.950 807.750 292.050 808.200 ;
        RECT 295.950 807.750 298.050 808.200 ;
        RECT 289.950 806.550 298.050 807.750 ;
        RECT 289.950 806.100 292.050 806.550 ;
        RECT 295.950 806.100 298.050 806.550 ;
        RECT 328.950 807.600 331.050 808.200 ;
        RECT 340.950 807.600 343.050 808.050 ;
        RECT 328.950 806.400 343.050 807.600 ;
        RECT 328.950 806.100 331.050 806.400 ;
        RECT 268.950 798.600 271.050 799.050 ;
        RECT 257.400 797.400 271.050 798.600 ;
        RECT 278.400 798.600 279.600 805.950 ;
        RECT 296.400 804.600 297.600 806.100 ;
        RECT 340.950 805.950 343.050 806.400 ;
        RECT 349.950 806.100 352.050 808.200 ;
        RECT 355.950 807.750 358.050 808.200 ;
        RECT 364.950 807.750 367.050 808.200 ;
        RECT 355.950 806.550 367.050 807.750 ;
        RECT 397.950 807.600 400.050 808.200 ;
        RECT 355.950 806.100 358.050 806.550 ;
        RECT 364.950 806.100 367.050 806.550 ;
        RECT 371.400 806.400 400.050 807.600 ;
        RECT 296.400 803.400 333.600 804.600 ;
        RECT 332.400 801.900 333.600 803.400 ;
        RECT 286.950 801.600 289.050 801.900 ;
        RECT 325.950 801.600 328.050 801.900 ;
        RECT 286.950 800.400 328.050 801.600 ;
        RECT 286.950 799.800 289.050 800.400 ;
        RECT 325.950 799.800 328.050 800.400 ;
        RECT 331.950 799.800 334.050 801.900 ;
        RECT 340.950 801.450 343.050 801.900 ;
        RECT 346.950 801.450 349.050 801.900 ;
        RECT 340.950 800.250 349.050 801.450 ;
        RECT 350.400 801.600 351.600 806.100 ;
        RECT 361.950 801.600 364.050 802.050 ;
        RECT 371.400 801.900 372.600 806.400 ;
        RECT 397.950 806.100 400.050 806.400 ;
        RECT 406.950 807.600 409.050 808.050 ;
        RECT 415.950 807.750 418.050 808.200 ;
        RECT 424.950 807.750 427.050 808.200 ;
        RECT 415.950 807.600 427.050 807.750 ;
        RECT 406.950 806.550 427.050 807.600 ;
        RECT 406.950 806.400 418.050 806.550 ;
        RECT 406.950 805.950 409.050 806.400 ;
        RECT 415.950 806.100 418.050 806.400 ;
        RECT 424.950 806.100 427.050 806.550 ;
        RECT 463.950 807.600 466.050 808.200 ;
        RECT 475.950 807.600 478.050 808.050 ;
        RECT 463.950 806.400 478.050 807.600 ;
        RECT 463.950 806.100 466.050 806.400 ;
        RECT 475.950 805.950 478.050 806.400 ;
        RECT 350.400 800.400 364.050 801.600 ;
        RECT 340.950 799.800 343.050 800.250 ;
        RECT 346.950 799.800 349.050 800.250 ;
        RECT 361.950 799.950 364.050 800.400 ;
        RECT 370.950 799.800 373.050 801.900 ;
        RECT 388.950 801.450 391.050 801.900 ;
        RECT 394.950 801.450 397.050 801.900 ;
        RECT 388.950 800.250 397.050 801.450 ;
        RECT 388.950 799.800 391.050 800.250 ;
        RECT 394.950 799.800 397.050 800.250 ;
        RECT 406.950 801.600 409.050 802.050 ;
        RECT 415.950 801.600 418.050 802.050 ;
        RECT 406.950 800.400 418.050 801.600 ;
        RECT 406.950 799.950 409.050 800.400 ;
        RECT 415.950 799.950 418.050 800.400 ;
        RECT 427.950 801.600 430.050 801.900 ;
        RECT 442.950 801.600 445.050 801.900 ;
        RECT 427.950 800.400 445.050 801.600 ;
        RECT 482.400 801.600 483.600 808.950 ;
        RECT 490.950 807.750 493.050 808.200 ;
        RECT 499.950 807.750 502.050 808.200 ;
        RECT 490.950 807.600 502.050 807.750 ;
        RECT 535.950 807.600 538.050 808.050 ;
        RECT 490.950 806.550 538.050 807.600 ;
        RECT 490.950 806.100 493.050 806.550 ;
        RECT 499.950 806.400 538.050 806.550 ;
        RECT 499.950 806.100 502.050 806.400 ;
        RECT 535.950 805.950 538.050 806.400 ;
        RECT 550.950 807.750 553.050 808.200 ;
        RECT 577.950 807.750 580.050 808.200 ;
        RECT 550.950 807.600 580.050 807.750 ;
        RECT 583.950 807.600 586.050 808.050 ;
        RECT 550.950 806.550 586.050 807.600 ;
        RECT 550.950 806.100 553.050 806.550 ;
        RECT 577.950 806.400 586.050 806.550 ;
        RECT 577.950 806.100 580.050 806.400 ;
        RECT 583.950 805.950 586.050 806.400 ;
        RECT 610.950 807.600 613.050 807.900 ;
        RECT 619.950 807.600 622.050 808.200 ;
        RECT 640.950 807.600 643.050 808.200 ;
        RECT 610.950 806.400 643.050 807.600 ;
        RECT 610.950 805.800 613.050 806.400 ;
        RECT 619.950 806.100 622.050 806.400 ;
        RECT 640.950 806.100 643.050 806.400 ;
        RECT 646.950 807.600 649.050 808.200 ;
        RECT 679.950 807.600 682.050 808.200 ;
        RECT 691.950 807.600 694.050 808.050 ;
        RECT 706.950 807.600 709.050 808.050 ;
        RECT 646.950 806.400 687.600 807.600 ;
        RECT 646.950 806.100 649.050 806.400 ;
        RECT 679.950 806.100 682.050 806.400 ;
        RECT 686.400 802.050 687.600 806.400 ;
        RECT 691.950 806.400 709.050 807.600 ;
        RECT 691.950 805.950 694.050 806.400 ;
        RECT 706.950 805.950 709.050 806.400 ;
        RECT 748.950 807.600 751.050 808.050 ;
        RECT 778.950 807.600 781.050 808.200 ;
        RECT 748.950 806.400 781.050 807.600 ;
        RECT 748.950 805.950 751.050 806.400 ;
        RECT 778.950 806.100 781.050 806.400 ;
        RECT 793.950 807.600 796.050 808.050 ;
        RECT 799.950 807.600 802.050 808.200 ;
        RECT 793.950 806.400 802.050 807.600 ;
        RECT 793.950 805.950 796.050 806.400 ;
        RECT 799.950 806.100 802.050 806.400 ;
        RECT 811.950 807.750 814.050 808.200 ;
        RECT 820.950 807.750 823.050 808.200 ;
        RECT 811.950 806.550 823.050 807.750 ;
        RECT 811.950 806.100 814.050 806.550 ;
        RECT 814.950 804.600 817.050 805.050 ;
        RECT 803.400 803.400 817.050 804.600 ;
        RECT 487.950 801.600 490.050 801.900 ;
        RECT 538.950 801.600 541.050 801.900 ;
        RECT 482.400 800.400 490.050 801.600 ;
        RECT 427.950 799.800 430.050 800.400 ;
        RECT 442.950 799.800 445.050 800.400 ;
        RECT 487.950 799.800 490.050 800.400 ;
        RECT 530.400 800.400 541.050 801.600 ;
        RECT 283.950 798.600 286.050 799.050 ;
        RECT 278.400 797.400 286.050 798.600 ;
        RECT 223.950 796.950 226.050 797.400 ;
        RECT 94.950 795.600 97.050 796.050 ;
        RECT 103.950 795.600 106.050 796.050 ;
        RECT 94.950 794.400 106.050 795.600 ;
        RECT 94.950 793.950 97.050 794.400 ;
        RECT 103.950 793.950 106.050 794.400 ;
        RECT 181.950 795.600 184.050 796.050 ;
        RECT 214.950 795.600 217.050 796.050 ;
        RECT 181.950 794.400 217.050 795.600 ;
        RECT 181.950 793.950 184.050 794.400 ;
        RECT 214.950 793.950 217.050 794.400 ;
        RECT 229.950 795.600 232.050 796.050 ;
        RECT 245.400 795.600 246.600 797.400 ;
        RECT 250.950 796.950 253.050 797.400 ;
        RECT 268.950 796.950 271.050 797.400 ;
        RECT 283.950 796.950 286.050 797.400 ;
        RECT 376.950 798.600 379.050 799.050 ;
        RECT 385.950 798.600 388.050 799.050 ;
        RECT 376.950 797.400 388.050 798.600 ;
        RECT 376.950 796.950 379.050 797.400 ;
        RECT 385.950 796.950 388.050 797.400 ;
        RECT 466.950 798.600 469.050 799.050 ;
        RECT 472.950 798.600 475.050 799.050 ;
        RECT 466.950 797.400 475.050 798.600 ;
        RECT 466.950 796.950 469.050 797.400 ;
        RECT 472.950 796.950 475.050 797.400 ;
        RECT 481.950 798.600 484.050 799.050 ;
        RECT 514.950 798.600 517.050 799.050 ;
        RECT 481.950 797.400 517.050 798.600 ;
        RECT 481.950 796.950 484.050 797.400 ;
        RECT 514.950 796.950 517.050 797.400 ;
        RECT 229.950 794.400 246.600 795.600 ;
        RECT 298.950 795.600 301.050 796.050 ;
        RECT 328.950 795.600 331.050 796.050 ;
        RECT 298.950 794.400 331.050 795.600 ;
        RECT 386.400 795.600 387.600 796.950 ;
        RECT 400.950 795.600 403.050 796.050 ;
        RECT 386.400 794.400 403.050 795.600 ;
        RECT 229.950 793.950 232.050 794.400 ;
        RECT 298.950 793.950 301.050 794.400 ;
        RECT 328.950 793.950 331.050 794.400 ;
        RECT 400.950 793.950 403.050 794.400 ;
        RECT 418.950 795.600 421.050 796.050 ;
        RECT 439.800 795.600 441.900 796.050 ;
        RECT 418.950 794.400 441.900 795.600 ;
        RECT 418.950 793.950 421.050 794.400 ;
        RECT 439.800 793.950 441.900 794.400 ;
        RECT 442.950 795.600 445.050 796.050 ;
        RECT 460.950 795.600 463.050 796.050 ;
        RECT 442.950 794.400 463.050 795.600 ;
        RECT 442.950 793.950 445.050 794.400 ;
        RECT 460.950 793.950 463.050 794.400 ;
        RECT 475.950 795.600 478.050 796.050 ;
        RECT 482.400 795.600 483.600 796.950 ;
        RECT 530.400 795.600 531.600 800.400 ;
        RECT 538.950 799.800 541.050 800.400 ;
        RECT 574.950 801.600 577.050 801.900 ;
        RECT 586.950 801.600 589.050 802.050 ;
        RECT 574.950 800.400 589.050 801.600 ;
        RECT 574.950 799.800 577.050 800.400 ;
        RECT 586.950 799.950 589.050 800.400 ;
        RECT 592.950 801.450 595.050 801.900 ;
        RECT 610.950 801.450 613.050 801.900 ;
        RECT 592.950 800.250 613.050 801.450 ;
        RECT 592.950 799.800 595.050 800.250 ;
        RECT 610.950 799.800 613.050 800.250 ;
        RECT 622.950 801.450 625.050 801.900 ;
        RECT 628.950 801.600 631.050 802.050 ;
        RECT 649.950 801.600 652.050 801.900 ;
        RECT 628.950 801.450 652.050 801.600 ;
        RECT 622.950 800.400 652.050 801.450 ;
        RECT 622.950 800.250 631.050 800.400 ;
        RECT 622.950 799.800 625.050 800.250 ;
        RECT 628.950 799.950 631.050 800.250 ;
        RECT 649.950 799.800 652.050 800.400 ;
        RECT 685.950 799.950 688.050 802.050 ;
        RECT 691.950 801.450 694.050 801.900 ;
        RECT 697.950 801.450 700.050 801.900 ;
        RECT 691.950 800.250 700.050 801.450 ;
        RECT 691.950 799.800 694.050 800.250 ;
        RECT 697.950 799.800 700.050 800.250 ;
        RECT 712.950 801.450 715.050 801.900 ;
        RECT 727.950 801.600 730.050 801.900 ;
        RECT 736.950 801.600 739.050 802.050 ;
        RECT 803.400 801.900 804.600 803.400 ;
        RECT 814.950 802.950 817.050 803.400 ;
        RECT 727.950 801.450 739.050 801.600 ;
        RECT 712.950 800.400 739.050 801.450 ;
        RECT 712.950 800.250 730.050 800.400 ;
        RECT 712.950 799.800 715.050 800.250 ;
        RECT 727.950 799.800 730.050 800.250 ;
        RECT 736.950 799.950 739.050 800.400 ;
        RECT 802.950 799.800 805.050 801.900 ;
        RECT 808.950 801.600 811.050 801.900 ;
        RECT 818.400 801.600 819.600 806.550 ;
        RECT 820.950 806.100 823.050 806.550 ;
        RECT 808.950 800.400 819.600 801.600 ;
        RECT 829.950 801.600 832.050 802.050 ;
        RECT 845.400 801.900 846.600 808.950 ;
        RECT 850.950 805.950 853.050 808.050 ;
        RECT 856.950 807.600 859.050 808.050 ;
        RECT 862.950 807.600 865.050 808.200 ;
        RECT 856.950 806.400 865.050 807.600 ;
        RECT 856.950 805.950 859.050 806.400 ;
        RECT 862.950 806.100 865.050 806.400 ;
        RECT 868.950 807.750 871.050 808.200 ;
        RECT 877.950 807.750 880.050 808.050 ;
        RECT 868.950 807.600 880.050 807.750 ;
        RECT 889.950 807.600 892.050 808.200 ;
        RECT 868.950 806.550 892.050 807.600 ;
        RECT 868.950 806.100 871.050 806.550 ;
        RECT 877.950 806.400 892.050 806.550 ;
        RECT 877.950 805.950 880.050 806.400 ;
        RECT 889.950 806.100 892.050 806.400 ;
        RECT 898.950 805.950 901.050 808.050 ;
        RECT 851.400 802.050 852.600 805.950 ;
        RECT 899.400 802.050 900.600 805.950 ;
        RECT 844.950 801.600 847.050 801.900 ;
        RECT 829.950 800.400 847.050 801.600 ;
        RECT 808.950 799.800 811.050 800.400 ;
        RECT 829.950 799.950 832.050 800.400 ;
        RECT 844.950 799.800 847.050 800.400 ;
        RECT 850.950 799.950 853.050 802.050 ;
        RECT 865.950 801.600 868.050 801.900 ;
        RECT 877.950 801.600 880.050 802.050 ;
        RECT 865.950 800.400 880.050 801.600 ;
        RECT 865.950 799.800 868.050 800.400 ;
        RECT 877.950 799.950 880.050 800.400 ;
        RECT 898.800 799.950 900.900 802.050 ;
        RECT 901.950 801.450 904.050 801.900 ;
        RECT 913.950 801.450 916.050 801.900 ;
        RECT 901.950 800.250 916.050 801.450 ;
        RECT 901.950 799.800 904.050 800.250 ;
        RECT 913.950 799.800 916.050 800.250 ;
        RECT 634.950 798.600 637.050 799.050 ;
        RECT 643.950 798.600 646.050 799.050 ;
        RECT 634.950 797.400 646.050 798.600 ;
        RECT 634.950 796.950 637.050 797.400 ;
        RECT 643.950 796.950 646.050 797.400 ;
        RECT 661.950 798.600 664.050 799.050 ;
        RECT 676.950 798.600 679.050 799.050 ;
        RECT 661.950 797.400 679.050 798.600 ;
        RECT 661.950 796.950 664.050 797.400 ;
        RECT 676.950 796.950 679.050 797.400 ;
        RECT 745.950 798.600 748.050 799.050 ;
        RECT 775.950 798.600 778.050 799.050 ;
        RECT 793.950 798.600 796.050 799.050 ;
        RECT 745.950 797.400 796.050 798.600 ;
        RECT 745.950 796.950 748.050 797.400 ;
        RECT 775.950 796.950 778.050 797.400 ;
        RECT 793.950 796.950 796.050 797.400 ;
        RECT 856.950 798.600 859.050 799.050 ;
        RECT 880.950 798.600 883.050 799.050 ;
        RECT 856.950 797.400 883.050 798.600 ;
        RECT 856.950 796.950 859.050 797.400 ;
        RECT 880.950 796.950 883.050 797.400 ;
        RECT 475.950 794.400 483.600 795.600 ;
        RECT 527.400 794.400 531.600 795.600 ;
        RECT 697.950 795.600 700.050 796.050 ;
        RECT 703.950 795.600 706.050 796.050 ;
        RECT 697.950 794.400 706.050 795.600 ;
        RECT 475.950 793.950 478.050 794.400 ;
        RECT 7.950 792.600 10.050 793.050 ;
        RECT 28.950 792.600 31.050 793.050 ;
        RECT 7.950 791.400 31.050 792.600 ;
        RECT 7.950 790.950 10.050 791.400 ;
        RECT 28.950 790.950 31.050 791.400 ;
        RECT 73.950 792.600 76.050 793.050 ;
        RECT 106.950 792.600 109.050 793.050 ;
        RECT 73.950 791.400 109.050 792.600 ;
        RECT 73.950 790.950 76.050 791.400 ;
        RECT 106.950 790.950 109.050 791.400 ;
        RECT 280.950 792.600 283.050 793.050 ;
        RECT 310.800 792.600 312.900 793.050 ;
        RECT 280.950 791.400 312.900 792.600 ;
        RECT 280.950 790.950 283.050 791.400 ;
        RECT 310.800 790.950 312.900 791.400 ;
        RECT 313.950 792.600 316.050 793.050 ;
        RECT 367.950 792.600 370.050 793.050 ;
        RECT 313.950 791.400 370.050 792.600 ;
        RECT 313.950 790.950 316.050 791.400 ;
        RECT 367.950 790.950 370.050 791.400 ;
        RECT 430.950 792.600 433.050 793.050 ;
        RECT 436.950 792.600 439.050 793.050 ;
        RECT 448.950 792.600 451.050 793.050 ;
        RECT 430.950 791.400 451.050 792.600 ;
        RECT 430.950 790.950 433.050 791.400 ;
        RECT 436.950 790.950 439.050 791.400 ;
        RECT 448.950 790.950 451.050 791.400 ;
        RECT 478.950 792.600 481.050 793.050 ;
        RECT 520.950 792.600 523.050 793.050 ;
        RECT 478.950 791.400 523.050 792.600 ;
        RECT 478.950 790.950 481.050 791.400 ;
        RECT 520.950 790.950 523.050 791.400 ;
        RECT 193.950 789.600 196.050 790.050 ;
        RECT 292.950 789.600 295.050 790.050 ;
        RECT 304.950 789.600 307.050 790.050 ;
        RECT 193.950 788.400 225.600 789.600 ;
        RECT 193.950 787.950 196.050 788.400 ;
        RECT 112.950 786.600 115.050 787.050 ;
        RECT 145.950 786.600 148.050 787.050 ;
        RECT 112.950 785.400 148.050 786.600 ;
        RECT 112.950 784.950 115.050 785.400 ;
        RECT 145.950 784.950 148.050 785.400 ;
        RECT 205.950 786.600 208.050 787.050 ;
        RECT 217.950 786.600 220.050 787.050 ;
        RECT 205.950 785.400 220.050 786.600 ;
        RECT 224.400 786.600 225.600 788.400 ;
        RECT 292.950 788.400 307.050 789.600 ;
        RECT 292.950 787.950 295.050 788.400 ;
        RECT 304.950 787.950 307.050 788.400 ;
        RECT 316.950 789.600 319.050 790.050 ;
        RECT 352.950 789.600 355.050 790.050 ;
        RECT 316.950 788.400 355.050 789.600 ;
        RECT 316.950 787.950 319.050 788.400 ;
        RECT 352.950 787.950 355.050 788.400 ;
        RECT 370.950 789.600 373.050 790.050 ;
        RECT 472.950 789.600 475.050 790.050 ;
        RECT 370.950 788.400 475.050 789.600 ;
        RECT 370.950 787.950 373.050 788.400 ;
        RECT 472.950 787.950 475.050 788.400 ;
        RECT 508.950 789.600 511.050 790.050 ;
        RECT 517.950 789.600 520.050 790.050 ;
        RECT 508.950 788.400 520.050 789.600 ;
        RECT 527.400 789.600 528.600 794.400 ;
        RECT 697.950 793.950 700.050 794.400 ;
        RECT 703.950 793.950 706.050 794.400 ;
        RECT 736.950 795.600 739.050 796.050 ;
        RECT 754.950 795.600 757.050 796.050 ;
        RECT 736.950 794.400 757.050 795.600 ;
        RECT 736.950 793.950 739.050 794.400 ;
        RECT 754.950 793.950 757.050 794.400 ;
        RECT 841.950 795.600 844.050 796.050 ;
        RECT 904.950 795.600 907.050 796.050 ;
        RECT 841.950 794.400 907.050 795.600 ;
        RECT 841.950 793.950 844.050 794.400 ;
        RECT 904.950 793.950 907.050 794.400 ;
        RECT 595.950 792.600 598.050 793.050 ;
        RECT 616.950 792.600 619.050 793.050 ;
        RECT 595.950 791.400 619.050 792.600 ;
        RECT 595.950 790.950 598.050 791.400 ;
        RECT 616.950 790.950 619.050 791.400 ;
        RECT 691.950 792.600 694.050 793.050 ;
        RECT 715.950 792.600 718.050 793.050 ;
        RECT 691.950 791.400 718.050 792.600 ;
        RECT 691.950 790.950 694.050 791.400 ;
        RECT 715.950 790.950 718.050 791.400 ;
        RECT 733.950 792.600 736.050 793.050 ;
        RECT 763.950 792.600 766.050 793.050 ;
        RECT 769.950 792.600 772.050 793.050 ;
        RECT 733.950 791.400 772.050 792.600 ;
        RECT 733.950 790.950 736.050 791.400 ;
        RECT 763.950 790.950 766.050 791.400 ;
        RECT 769.950 790.950 772.050 791.400 ;
        RECT 781.950 792.600 784.050 793.050 ;
        RECT 823.800 792.600 825.900 793.050 ;
        RECT 781.950 791.400 825.900 792.600 ;
        RECT 781.950 790.950 784.050 791.400 ;
        RECT 823.800 790.950 825.900 791.400 ;
        RECT 826.950 792.600 831.000 793.050 ;
        RECT 850.950 792.600 853.050 793.050 ;
        RECT 892.950 792.600 895.050 793.050 ;
        RECT 826.950 790.950 831.600 792.600 ;
        RECT 850.950 791.400 895.050 792.600 ;
        RECT 850.950 790.950 853.050 791.400 ;
        RECT 892.950 790.950 895.050 791.400 ;
        RECT 553.950 789.600 556.050 790.050 ;
        RECT 574.950 789.600 577.050 790.050 ;
        RECT 527.400 789.000 531.600 789.600 ;
        RECT 527.400 788.400 532.050 789.000 ;
        RECT 508.950 787.950 511.050 788.400 ;
        RECT 517.950 787.950 520.050 788.400 ;
        RECT 259.950 786.600 262.050 787.050 ;
        RECT 224.400 785.400 262.050 786.600 ;
        RECT 205.950 784.950 208.050 785.400 ;
        RECT 217.950 784.950 220.050 785.400 ;
        RECT 259.950 784.950 262.050 785.400 ;
        RECT 265.950 786.600 268.050 787.050 ;
        RECT 313.950 786.600 316.050 787.050 ;
        RECT 265.950 785.400 316.050 786.600 ;
        RECT 265.950 784.950 268.050 785.400 ;
        RECT 313.950 784.950 316.050 785.400 ;
        RECT 367.950 786.600 370.050 787.050 ;
        RECT 385.950 786.600 388.050 787.050 ;
        RECT 367.950 785.400 388.050 786.600 ;
        RECT 367.950 784.950 370.050 785.400 ;
        RECT 385.950 784.950 388.050 785.400 ;
        RECT 415.950 786.600 418.050 787.050 ;
        RECT 430.950 786.600 433.050 787.050 ;
        RECT 415.950 785.400 433.050 786.600 ;
        RECT 415.950 784.950 418.050 785.400 ;
        RECT 430.950 784.950 433.050 785.400 ;
        RECT 439.950 786.600 442.050 787.050 ;
        RECT 466.950 786.600 469.050 787.050 ;
        RECT 496.950 786.600 499.050 787.050 ;
        RECT 439.950 785.400 499.050 786.600 ;
        RECT 439.950 784.950 442.050 785.400 ;
        RECT 466.950 784.950 469.050 785.400 ;
        RECT 496.950 784.950 499.050 785.400 ;
        RECT 514.950 786.600 517.050 787.050 ;
        RECT 520.950 786.600 523.050 786.900 ;
        RECT 514.950 785.400 523.050 786.600 ;
        RECT 514.950 784.950 517.050 785.400 ;
        RECT 73.950 783.600 76.050 784.050 ;
        RECT 130.950 783.600 133.050 784.050 ;
        RECT 73.950 782.400 133.050 783.600 ;
        RECT 146.400 783.600 147.600 784.950 ;
        RECT 520.950 784.800 523.050 785.400 ;
        RECT 529.950 784.950 532.050 788.400 ;
        RECT 553.950 788.400 577.050 789.600 ;
        RECT 553.950 787.950 556.050 788.400 ;
        RECT 574.950 787.950 577.050 788.400 ;
        RECT 619.950 789.600 622.050 790.050 ;
        RECT 649.950 789.600 652.050 790.050 ;
        RECT 619.950 788.400 652.050 789.600 ;
        RECT 830.400 789.600 831.600 790.950 ;
        RECT 865.950 789.600 868.050 790.050 ;
        RECT 830.400 788.400 868.050 789.600 ;
        RECT 619.950 787.950 622.050 788.400 ;
        RECT 649.950 787.950 652.050 788.400 ;
        RECT 865.950 787.950 868.050 788.400 ;
        RECT 583.950 786.600 586.050 787.050 ;
        RECT 661.950 786.600 664.050 787.050 ;
        RECT 583.950 785.400 664.050 786.600 ;
        RECT 583.950 784.950 586.050 785.400 ;
        RECT 661.950 784.950 664.050 785.400 ;
        RECT 709.950 786.600 712.050 787.050 ;
        RECT 739.950 786.600 742.050 787.050 ;
        RECT 709.950 785.400 742.050 786.600 ;
        RECT 709.950 784.950 712.050 785.400 ;
        RECT 739.950 784.950 742.050 785.400 ;
        RECT 772.950 786.600 775.050 787.050 ;
        RECT 808.950 786.600 811.050 787.050 ;
        RECT 772.950 785.400 811.050 786.600 ;
        RECT 772.950 784.950 775.050 785.400 ;
        RECT 808.950 784.950 811.050 785.400 ;
        RECT 817.950 786.600 820.050 787.050 ;
        RECT 871.950 786.600 874.050 787.050 ;
        RECT 886.950 786.600 889.050 787.050 ;
        RECT 817.950 785.400 889.050 786.600 ;
        RECT 817.950 784.950 820.050 785.400 ;
        RECT 871.950 784.950 874.050 785.400 ;
        RECT 886.950 784.950 889.050 785.400 ;
        RECT 250.800 783.600 252.900 784.050 ;
        RECT 146.400 782.400 252.900 783.600 ;
        RECT 73.950 781.950 76.050 782.400 ;
        RECT 130.950 781.950 133.050 782.400 ;
        RECT 250.800 781.950 252.900 782.400 ;
        RECT 253.950 783.600 256.050 784.050 ;
        RECT 292.950 783.600 295.050 784.050 ;
        RECT 364.950 783.600 367.050 784.050 ;
        RECT 253.950 782.400 367.050 783.600 ;
        RECT 253.950 781.950 256.050 782.400 ;
        RECT 292.950 781.950 295.050 782.400 ;
        RECT 364.950 781.950 367.050 782.400 ;
        RECT 373.950 783.600 376.050 784.050 ;
        RECT 418.950 783.600 421.050 784.050 ;
        RECT 373.950 782.400 421.050 783.600 ;
        RECT 373.950 781.950 376.050 782.400 ;
        RECT 418.950 781.950 421.050 782.400 ;
        RECT 424.950 783.600 427.050 784.050 ;
        RECT 499.950 783.600 502.050 784.050 ;
        RECT 559.950 783.600 562.050 784.050 ;
        RECT 424.950 782.400 562.050 783.600 ;
        RECT 424.950 781.950 427.050 782.400 ;
        RECT 499.950 781.950 502.050 782.400 ;
        RECT 559.950 781.950 562.050 782.400 ;
        RECT 568.950 783.600 571.050 784.050 ;
        RECT 619.950 783.600 622.050 784.050 ;
        RECT 568.950 782.400 622.050 783.600 ;
        RECT 568.950 781.950 571.050 782.400 ;
        RECT 619.950 781.950 622.050 782.400 ;
        RECT 676.950 783.600 679.050 784.050 ;
        RECT 706.950 783.600 709.050 784.050 ;
        RECT 676.950 782.400 709.050 783.600 ;
        RECT 676.950 781.950 679.050 782.400 ;
        RECT 706.950 781.950 709.050 782.400 ;
        RECT 148.950 780.600 151.050 781.050 ;
        RECT 160.950 780.600 163.050 781.050 ;
        RECT 148.950 779.400 163.050 780.600 ;
        RECT 148.950 778.950 151.050 779.400 ;
        RECT 160.950 778.950 163.050 779.400 ;
        RECT 169.950 780.600 172.050 781.050 ;
        RECT 229.950 780.600 232.050 781.050 ;
        RECT 169.950 779.400 232.050 780.600 ;
        RECT 169.950 778.950 172.050 779.400 ;
        RECT 229.950 778.950 232.050 779.400 ;
        RECT 307.950 780.600 310.050 781.050 ;
        RECT 325.800 780.600 327.900 781.050 ;
        RECT 307.950 779.400 327.900 780.600 ;
        RECT 307.950 778.950 310.050 779.400 ;
        RECT 325.800 778.950 327.900 779.400 ;
        RECT 328.950 780.600 331.050 781.050 ;
        RECT 370.950 780.600 373.050 781.050 ;
        RECT 328.950 779.400 373.050 780.600 ;
        RECT 328.950 778.950 331.050 779.400 ;
        RECT 370.950 778.950 373.050 779.400 ;
        RECT 376.950 780.600 379.050 781.050 ;
        RECT 397.950 780.600 400.050 781.050 ;
        RECT 376.950 779.400 400.050 780.600 ;
        RECT 376.950 778.950 379.050 779.400 ;
        RECT 397.950 778.950 400.050 779.400 ;
        RECT 523.950 780.600 526.050 781.050 ;
        RECT 556.950 780.600 559.050 781.050 ;
        RECT 523.950 779.400 559.050 780.600 ;
        RECT 523.950 778.950 526.050 779.400 ;
        RECT 556.950 778.950 559.050 779.400 ;
        RECT 589.950 780.600 592.050 781.050 ;
        RECT 664.950 780.600 667.050 781.050 ;
        RECT 589.950 779.400 667.050 780.600 ;
        RECT 589.950 778.950 592.050 779.400 ;
        RECT 664.950 778.950 667.050 779.400 ;
        RECT 757.950 780.600 760.050 781.050 ;
        RECT 817.950 780.600 820.050 781.050 ;
        RECT 757.950 779.400 820.050 780.600 ;
        RECT 757.950 778.950 760.050 779.400 ;
        RECT 817.950 778.950 820.050 779.400 ;
        RECT 838.950 780.600 841.050 781.050 ;
        RECT 859.950 780.600 862.050 781.050 ;
        RECT 838.950 779.400 862.050 780.600 ;
        RECT 838.950 778.950 841.050 779.400 ;
        RECT 859.950 778.950 862.050 779.400 ;
        RECT 13.950 777.600 16.050 778.050 ;
        RECT 25.950 777.600 28.050 778.050 ;
        RECT 91.950 777.600 94.050 778.050 ;
        RECT 316.950 777.600 319.050 778.050 ;
        RECT 13.950 776.400 94.050 777.600 ;
        RECT 13.950 775.950 16.050 776.400 ;
        RECT 25.950 775.950 28.050 776.400 ;
        RECT 91.950 775.950 94.050 776.400 ;
        RECT 311.400 776.400 319.050 777.600 ;
        RECT 79.950 774.600 82.050 775.050 ;
        RECT 85.950 774.600 88.050 775.050 ;
        RECT 79.950 773.400 88.050 774.600 ;
        RECT 79.950 772.950 82.050 773.400 ;
        RECT 85.950 772.950 88.050 773.400 ;
        RECT 154.950 774.600 157.050 775.050 ;
        RECT 193.950 774.600 196.050 775.050 ;
        RECT 154.950 773.400 196.050 774.600 ;
        RECT 154.950 772.950 157.050 773.400 ;
        RECT 193.950 772.950 196.050 773.400 ;
        RECT 214.950 774.600 217.050 775.050 ;
        RECT 226.950 774.600 229.050 775.050 ;
        RECT 214.950 773.400 229.050 774.600 ;
        RECT 214.950 772.950 217.050 773.400 ;
        RECT 226.950 772.950 229.050 773.400 ;
        RECT 298.950 774.600 301.050 775.050 ;
        RECT 311.400 774.600 312.600 776.400 ;
        RECT 316.950 775.950 319.050 776.400 ;
        RECT 379.950 777.600 382.050 778.050 ;
        RECT 430.950 777.600 433.050 778.050 ;
        RECT 475.950 777.600 478.050 778.050 ;
        RECT 379.950 776.400 433.050 777.600 ;
        RECT 379.950 775.950 382.050 776.400 ;
        RECT 430.950 775.950 433.050 776.400 ;
        RECT 461.400 776.400 478.050 777.600 ;
        RECT 298.950 773.400 312.600 774.600 ;
        RECT 322.950 774.600 325.050 775.050 ;
        RECT 373.950 774.600 376.050 775.050 ;
        RECT 322.950 773.400 376.050 774.600 ;
        RECT 298.950 772.950 301.050 773.400 ;
        RECT 322.950 772.950 325.050 773.400 ;
        RECT 373.950 772.950 376.050 773.400 ;
        RECT 385.950 774.600 388.050 775.050 ;
        RECT 461.400 774.600 462.600 776.400 ;
        RECT 475.950 775.950 478.050 776.400 ;
        RECT 526.950 777.600 529.050 778.050 ;
        RECT 532.950 777.600 535.050 778.050 ;
        RECT 526.950 776.400 535.050 777.600 ;
        RECT 526.950 775.950 529.050 776.400 ;
        RECT 532.950 775.950 535.050 776.400 ;
        RECT 625.950 777.600 628.050 778.050 ;
        RECT 631.950 777.600 634.050 778.050 ;
        RECT 625.950 776.400 634.050 777.600 ;
        RECT 625.950 775.950 628.050 776.400 ;
        RECT 631.950 775.950 634.050 776.400 ;
        RECT 694.950 777.600 697.050 778.050 ;
        RECT 712.950 777.600 715.050 778.050 ;
        RECT 694.950 776.400 715.050 777.600 ;
        RECT 694.950 775.950 697.050 776.400 ;
        RECT 712.950 775.950 715.050 776.400 ;
        RECT 718.950 777.600 721.050 778.050 ;
        RECT 748.950 777.600 751.050 778.050 ;
        RECT 718.950 776.400 751.050 777.600 ;
        RECT 718.950 775.950 721.050 776.400 ;
        RECT 748.950 775.950 751.050 776.400 ;
        RECT 796.950 777.600 799.050 778.050 ;
        RECT 826.950 777.600 829.050 778.050 ;
        RECT 796.950 776.400 829.050 777.600 ;
        RECT 796.950 775.950 799.050 776.400 ;
        RECT 826.950 775.950 829.050 776.400 ;
        RECT 874.950 777.600 877.050 778.050 ;
        RECT 916.950 777.600 919.050 778.050 ;
        RECT 874.950 776.400 919.050 777.600 ;
        RECT 874.950 775.950 877.050 776.400 ;
        RECT 916.950 775.950 919.050 776.400 ;
        RECT 385.950 773.400 462.600 774.600 ;
        RECT 517.950 774.600 520.050 775.050 ;
        RECT 529.950 774.600 532.050 775.050 ;
        RECT 517.950 773.400 532.050 774.600 ;
        RECT 385.950 772.950 388.050 773.400 ;
        RECT 517.950 772.950 520.050 773.400 ;
        RECT 529.950 772.950 532.050 773.400 ;
        RECT 658.950 774.600 661.050 775.050 ;
        RECT 676.950 774.600 679.050 775.050 ;
        RECT 658.950 773.400 679.050 774.600 ;
        RECT 658.950 772.950 661.050 773.400 ;
        RECT 676.950 772.950 679.050 773.400 ;
        RECT 742.950 774.600 745.050 775.050 ;
        RECT 766.950 774.600 769.050 775.050 ;
        RECT 742.950 773.400 769.050 774.600 ;
        RECT 742.950 772.950 745.050 773.400 ;
        RECT 766.950 772.950 769.050 773.400 ;
        RECT 790.950 774.600 793.050 775.050 ;
        RECT 835.950 774.600 838.050 775.050 ;
        RECT 790.950 773.400 838.050 774.600 ;
        RECT 790.950 772.950 793.050 773.400 ;
        RECT 835.950 772.950 838.050 773.400 ;
        RECT 889.950 774.600 892.050 775.050 ;
        RECT 898.950 774.600 901.050 775.050 ;
        RECT 913.950 774.600 916.050 775.050 ;
        RECT 889.950 773.400 916.050 774.600 ;
        RECT 889.950 772.950 892.050 773.400 ;
        RECT 898.950 772.950 901.050 773.400 ;
        RECT 913.950 772.950 916.050 773.400 ;
        RECT 181.950 771.600 184.050 772.050 ;
        RECT 158.400 770.400 184.050 771.600 ;
        RECT 79.950 768.600 82.050 769.050 ;
        RECT 97.950 768.600 100.050 769.050 ;
        RECT 79.950 767.400 100.050 768.600 ;
        RECT 79.950 766.950 82.050 767.400 ;
        RECT 97.950 766.950 100.050 767.400 ;
        RECT 124.950 768.600 127.050 769.050 ;
        RECT 142.950 768.600 145.050 769.050 ;
        RECT 124.950 767.400 145.050 768.600 ;
        RECT 124.950 766.950 127.050 767.400 ;
        RECT 142.950 766.950 145.050 767.400 ;
        RECT 151.950 768.600 154.050 769.050 ;
        RECT 158.400 768.600 159.600 770.400 ;
        RECT 181.950 769.950 184.050 770.400 ;
        RECT 217.950 771.600 220.050 772.050 ;
        RECT 253.950 771.600 256.050 772.050 ;
        RECT 217.950 770.400 256.050 771.600 ;
        RECT 217.950 769.950 220.050 770.400 ;
        RECT 253.950 769.950 256.050 770.400 ;
        RECT 448.950 771.600 451.050 772.050 ;
        RECT 469.950 771.600 472.050 772.050 ;
        RECT 448.950 770.400 472.050 771.600 ;
        RECT 448.950 769.950 451.050 770.400 ;
        RECT 469.950 769.950 472.050 770.400 ;
        RECT 478.950 771.600 481.050 772.050 ;
        RECT 508.950 771.600 511.050 772.050 ;
        RECT 478.950 770.400 511.050 771.600 ;
        RECT 478.950 769.950 481.050 770.400 ;
        RECT 508.950 769.950 511.050 770.400 ;
        RECT 559.950 771.600 562.050 772.050 ;
        RECT 628.950 771.600 631.050 772.050 ;
        RECT 559.950 770.400 631.050 771.600 ;
        RECT 559.950 769.950 562.050 770.400 ;
        RECT 628.950 769.950 631.050 770.400 ;
        RECT 643.950 771.600 646.050 772.050 ;
        RECT 724.950 771.600 727.050 772.050 ;
        RECT 772.800 771.600 774.900 772.050 ;
        RECT 643.950 770.400 681.600 771.600 ;
        RECT 643.950 769.950 646.050 770.400 ;
        RECT 680.400 769.050 681.600 770.400 ;
        RECT 724.950 770.400 774.900 771.600 ;
        RECT 724.950 769.950 727.050 770.400 ;
        RECT 772.800 769.950 774.900 770.400 ;
        RECT 775.950 771.600 778.050 772.050 ;
        RECT 811.950 771.600 814.050 772.050 ;
        RECT 775.950 770.400 814.050 771.600 ;
        RECT 775.950 769.950 778.050 770.400 ;
        RECT 811.950 769.950 814.050 770.400 ;
        RECT 151.950 767.400 159.600 768.600 ;
        RECT 184.950 768.600 187.050 769.050 ;
        RECT 262.950 768.600 265.050 769.050 ;
        RECT 313.950 768.600 316.050 769.050 ;
        RECT 184.950 767.400 213.600 768.600 ;
        RECT 151.950 766.950 154.050 767.400 ;
        RECT 184.950 766.950 187.050 767.400 ;
        RECT 109.800 763.950 111.900 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 212.400 765.600 213.600 767.400 ;
        RECT 239.400 767.400 316.050 768.600 ;
        RECT 212.400 764.400 216.600 765.600 ;
        RECT 10.950 760.950 13.050 763.050 ;
        RECT 19.950 762.600 22.050 763.200 ;
        RECT 34.950 762.600 37.050 763.200 ;
        RECT 19.950 761.400 37.050 762.600 ;
        RECT 19.950 761.100 22.050 761.400 ;
        RECT 34.950 761.100 37.050 761.400 ;
        RECT 40.950 761.100 43.050 763.200 ;
        RECT 46.950 762.750 49.050 763.200 ;
        RECT 52.950 762.750 55.050 763.200 ;
        RECT 46.950 761.550 55.050 762.750 ;
        RECT 46.950 761.100 49.050 761.550 ;
        RECT 52.950 761.100 55.050 761.550 ;
        RECT 91.950 761.100 94.050 763.200 ;
        RECT 100.950 762.600 103.050 763.050 ;
        RECT 106.950 762.600 109.050 763.200 ;
        RECT 100.950 761.400 109.050 762.600 ;
        RECT 11.400 756.600 12.600 760.950 ;
        RECT 41.400 759.600 42.600 761.100 ;
        RECT 29.400 759.000 42.600 759.600 ;
        RECT 28.950 758.400 42.600 759.000 ;
        RECT 22.950 756.600 25.050 757.050 ;
        RECT 11.400 755.400 25.050 756.600 ;
        RECT 22.950 754.950 25.050 755.400 ;
        RECT 28.950 754.950 31.050 758.400 ;
        RECT 92.400 757.050 93.600 761.100 ;
        RECT 100.950 760.950 103.050 761.400 ;
        RECT 106.950 761.100 109.050 761.400 ;
        RECT 67.950 756.600 70.050 756.900 ;
        RECT 82.950 756.600 85.050 756.900 ;
        RECT 67.950 755.400 85.050 756.600 ;
        RECT 92.400 755.400 97.050 757.050 ;
        RECT 67.950 754.800 70.050 755.400 ;
        RECT 82.950 754.800 85.050 755.400 ;
        RECT 93.000 754.950 97.050 755.400 ;
        RECT 110.250 754.050 111.450 763.950 ;
        RECT 113.400 756.900 114.600 763.950 ;
        RECT 130.950 761.100 133.050 763.200 ;
        RECT 136.950 761.100 139.050 763.200 ;
        RECT 169.950 762.600 172.050 763.050 ;
        RECT 175.950 762.600 178.050 763.200 ;
        RECT 169.950 761.400 178.050 762.600 ;
        RECT 131.400 757.050 132.600 761.100 ;
        RECT 112.950 756.600 115.050 756.900 ;
        RECT 112.950 755.400 126.600 756.600 ;
        RECT 112.950 754.800 115.050 755.400 ;
        RECT 7.950 753.600 10.050 754.050 ;
        RECT 19.950 753.600 22.050 754.050 ;
        RECT 7.950 752.400 22.050 753.600 ;
        RECT 7.950 751.950 10.050 752.400 ;
        RECT 19.950 751.950 22.050 752.400 ;
        RECT 109.800 751.950 111.900 754.050 ;
        RECT 125.400 753.600 126.600 755.400 ;
        RECT 127.950 755.400 132.600 757.050 ;
        RECT 137.400 756.600 138.600 761.100 ;
        RECT 169.950 760.950 172.050 761.400 ;
        RECT 175.950 761.100 178.050 761.400 ;
        RECT 181.950 762.600 184.050 763.050 ;
        RECT 199.950 762.600 202.050 763.050 ;
        RECT 181.950 761.400 202.050 762.600 ;
        RECT 181.950 760.950 184.050 761.400 ;
        RECT 199.950 760.950 202.050 761.400 ;
        RECT 208.950 761.100 211.050 763.200 ;
        RECT 142.950 756.600 145.050 757.050 ;
        RECT 137.400 755.400 145.050 756.600 ;
        RECT 127.950 754.950 132.000 755.400 ;
        RECT 142.950 754.950 145.050 755.400 ;
        RECT 157.950 756.450 160.050 756.900 ;
        RECT 169.950 756.450 172.050 756.900 ;
        RECT 157.950 755.250 172.050 756.450 ;
        RECT 157.950 754.800 160.050 755.250 ;
        RECT 169.950 754.800 172.050 755.250 ;
        RECT 178.950 756.450 181.050 756.900 ;
        RECT 184.950 756.450 187.050 756.900 ;
        RECT 178.950 755.250 187.050 756.450 ;
        RECT 178.950 754.800 181.050 755.250 ;
        RECT 184.950 754.800 187.050 755.250 ;
        RECT 196.950 756.600 199.050 756.900 ;
        RECT 209.400 756.600 210.600 761.100 ;
        RECT 215.400 759.600 216.600 764.400 ;
        RECT 223.950 762.750 226.050 763.200 ;
        RECT 229.950 762.750 232.050 763.200 ;
        RECT 223.950 761.550 232.050 762.750 ;
        RECT 223.950 761.100 226.050 761.550 ;
        RECT 229.950 761.100 232.050 761.550 ;
        RECT 215.400 758.400 234.600 759.600 ;
        RECT 218.400 756.900 219.600 758.400 ;
        RECT 233.400 756.900 234.600 758.400 ;
        RECT 239.400 756.900 240.600 767.400 ;
        RECT 262.950 766.950 265.050 767.400 ;
        RECT 313.950 766.950 316.050 767.400 ;
        RECT 322.950 768.600 325.050 769.050 ;
        RECT 349.950 768.600 352.050 769.050 ;
        RECT 322.950 767.400 352.050 768.600 ;
        RECT 322.950 766.950 325.050 767.400 ;
        RECT 349.950 766.950 352.050 767.400 ;
        RECT 361.950 768.600 364.050 769.050 ;
        RECT 421.950 768.600 424.050 769.050 ;
        RECT 445.950 768.600 448.050 769.050 ;
        RECT 457.950 768.600 460.050 769.050 ;
        RECT 361.950 767.400 387.600 768.600 ;
        RECT 361.950 766.950 364.050 767.400 ;
        RECT 386.400 766.050 387.600 767.400 ;
        RECT 421.950 767.400 460.050 768.600 ;
        RECT 421.950 766.950 424.050 767.400 ;
        RECT 445.950 766.950 448.050 767.400 ;
        RECT 457.950 766.950 460.050 767.400 ;
        RECT 499.950 768.600 502.050 769.050 ;
        RECT 505.950 768.600 508.050 768.900 ;
        RECT 499.950 767.400 508.050 768.600 ;
        RECT 499.950 766.950 502.050 767.400 ;
        RECT 505.950 766.800 508.050 767.400 ;
        RECT 520.950 768.600 523.050 769.050 ;
        RECT 541.950 768.600 544.050 769.050 ;
        RECT 520.950 767.400 544.050 768.600 ;
        RECT 520.950 766.950 523.050 767.400 ;
        RECT 541.950 766.950 544.050 767.400 ;
        RECT 565.950 768.600 568.050 769.050 ;
        RECT 583.950 768.600 586.050 769.050 ;
        RECT 565.950 767.400 586.050 768.600 ;
        RECT 565.950 766.950 568.050 767.400 ;
        RECT 583.950 766.950 586.050 767.400 ;
        RECT 613.950 768.600 616.050 769.050 ;
        RECT 628.950 768.600 631.050 768.900 ;
        RECT 613.950 767.400 631.050 768.600 ;
        RECT 613.950 766.950 616.050 767.400 ;
        RECT 628.950 766.800 631.050 767.400 ;
        RECT 655.950 768.600 658.050 769.050 ;
        RECT 679.950 768.600 682.050 769.050 ;
        RECT 721.950 768.600 724.050 769.050 ;
        RECT 655.950 767.400 678.600 768.600 ;
        RECT 655.950 766.950 658.050 767.400 ;
        RECT 250.950 759.600 253.050 763.050 ;
        RECT 256.950 761.100 259.050 763.200 ;
        RECT 271.950 762.750 274.050 763.200 ;
        RECT 277.950 762.750 280.050 763.200 ;
        RECT 271.950 761.550 280.050 762.750 ;
        RECT 271.950 761.100 274.050 761.550 ;
        RECT 277.950 761.100 280.050 761.550 ;
        RECT 283.950 762.600 286.050 763.200 ;
        RECT 289.950 762.600 292.050 763.050 ;
        RECT 283.950 761.400 292.050 762.600 ;
        RECT 304.950 762.600 307.050 766.050 ;
        RECT 385.950 765.600 388.050 766.050 ;
        RECT 424.950 765.600 427.050 766.050 ;
        RECT 385.950 764.400 427.050 765.600 ;
        RECT 385.950 763.950 388.050 764.400 ;
        RECT 424.950 763.950 427.050 764.400 ;
        RECT 508.950 765.600 511.050 766.050 ;
        RECT 544.950 765.600 547.050 766.050 ;
        RECT 568.950 765.600 571.050 766.050 ;
        RECT 595.950 765.600 598.050 766.050 ;
        RECT 508.950 764.400 571.050 765.600 ;
        RECT 508.950 763.950 511.050 764.400 ;
        RECT 544.950 763.950 547.050 764.400 ;
        RECT 568.950 763.950 571.050 764.400 ;
        RECT 572.400 764.400 598.050 765.600 ;
        RECT 310.950 762.600 313.050 762.900 ;
        RECT 304.950 762.000 313.050 762.600 ;
        RECT 305.400 761.400 313.050 762.000 ;
        RECT 283.950 761.100 286.050 761.400 ;
        RECT 250.950 759.000 255.600 759.600 ;
        RECT 251.400 758.400 255.600 759.000 ;
        RECT 254.400 756.900 255.600 758.400 ;
        RECT 196.950 755.400 210.600 756.600 ;
        RECT 196.950 754.800 199.050 755.400 ;
        RECT 217.950 754.800 220.050 756.900 ;
        RECT 232.950 754.800 235.050 756.900 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 253.950 754.800 256.050 756.900 ;
        RECT 257.400 756.600 258.600 761.100 ;
        RECT 289.950 760.950 292.050 761.400 ;
        RECT 310.950 760.800 313.050 761.400 ;
        RECT 328.950 762.750 331.050 763.200 ;
        RECT 334.950 762.750 337.050 763.200 ;
        RECT 328.950 761.550 337.050 762.750 ;
        RECT 328.950 761.100 331.050 761.550 ;
        RECT 334.950 761.100 337.050 761.550 ;
        RECT 355.950 762.600 358.050 763.200 ;
        RECT 358.950 762.600 361.050 763.050 ;
        RECT 367.950 762.600 370.050 763.200 ;
        RECT 355.950 761.400 370.050 762.600 ;
        RECT 355.950 761.100 358.050 761.400 ;
        RECT 358.950 760.950 361.050 761.400 ;
        RECT 367.950 761.100 370.050 761.400 ;
        RECT 388.950 762.600 393.000 763.050 ;
        RECT 433.950 762.750 436.050 763.200 ;
        RECT 439.950 762.750 442.050 763.200 ;
        RECT 388.950 760.950 393.600 762.600 ;
        RECT 433.950 761.550 442.050 762.750 ;
        RECT 433.950 761.100 436.050 761.550 ;
        RECT 439.950 761.100 442.050 761.550 ;
        RECT 448.950 762.600 451.050 763.050 ;
        RECT 454.950 762.600 457.050 763.050 ;
        RECT 448.950 761.400 457.050 762.600 ;
        RECT 448.950 760.950 451.050 761.400 ;
        RECT 454.950 760.950 457.050 761.400 ;
        RECT 478.950 761.100 481.050 763.200 ;
        RECT 484.950 762.750 487.050 763.200 ;
        RECT 493.950 762.750 496.050 762.900 ;
        RECT 484.950 761.550 496.050 762.750 ;
        RECT 484.950 761.100 487.050 761.550 ;
        RECT 274.950 756.600 277.050 756.900 ;
        RECT 257.400 755.400 277.050 756.600 ;
        RECT 274.950 754.800 277.050 755.400 ;
        RECT 292.950 756.450 295.050 756.900 ;
        RECT 304.950 756.450 307.050 756.900 ;
        RECT 292.950 755.250 307.050 756.450 ;
        RECT 292.950 754.800 295.050 755.250 ;
        RECT 304.950 754.800 307.050 755.250 ;
        RECT 313.950 756.600 316.050 757.050 ;
        RECT 325.950 756.600 328.050 756.900 ;
        RECT 313.950 755.400 328.050 756.600 ;
        RECT 313.950 754.950 316.050 755.400 ;
        RECT 325.950 754.800 328.050 755.400 ;
        RECT 331.950 756.600 334.050 757.050 ;
        RECT 337.950 756.600 340.050 760.050 ;
        RECT 347.400 758.400 387.600 759.600 ;
        RECT 347.400 756.900 348.600 758.400 ;
        RECT 331.950 756.000 340.050 756.600 ;
        RECT 331.950 755.400 339.600 756.000 ;
        RECT 331.950 754.950 334.050 755.400 ;
        RECT 346.950 754.800 349.050 756.900 ;
        RECT 376.950 756.450 379.050 756.900 ;
        RECT 382.950 756.450 385.050 757.050 ;
        RECT 386.400 756.900 387.600 758.400 ;
        RECT 385.950 756.450 388.050 756.900 ;
        RECT 376.950 755.250 388.050 756.450 ;
        RECT 392.400 756.600 393.600 760.950 ;
        RECT 394.950 756.600 397.050 756.900 ;
        RECT 392.400 755.400 397.050 756.600 ;
        RECT 376.950 754.800 379.050 755.250 ;
        RECT 382.950 754.950 385.050 755.250 ;
        RECT 385.950 754.800 388.050 755.250 ;
        RECT 394.950 754.800 397.050 755.400 ;
        RECT 400.950 756.600 403.050 756.900 ;
        RECT 418.950 756.600 421.050 756.900 ;
        RECT 400.950 755.400 421.050 756.600 ;
        RECT 400.950 754.800 403.050 755.400 ;
        RECT 418.950 754.800 421.050 755.400 ;
        RECT 424.950 756.450 427.050 756.900 ;
        RECT 433.950 756.450 436.050 756.900 ;
        RECT 424.950 755.250 436.050 756.450 ;
        RECT 424.950 754.800 427.050 755.250 ;
        RECT 433.950 754.800 436.050 755.250 ;
        RECT 479.400 754.050 480.600 761.100 ;
        RECT 493.950 760.800 496.050 761.550 ;
        RECT 523.950 761.100 526.050 763.200 ;
        RECT 550.950 762.600 553.050 763.050 ;
        RECT 572.400 762.600 573.600 764.400 ;
        RECT 595.950 763.950 598.050 764.400 ;
        RECT 640.950 765.600 643.050 766.050 ;
        RECT 646.950 765.600 649.050 766.050 ;
        RECT 640.950 764.400 649.050 765.600 ;
        RECT 677.400 765.600 678.600 767.400 ;
        RECT 679.950 767.400 724.050 768.600 ;
        RECT 679.950 766.950 682.050 767.400 ;
        RECT 721.950 766.950 724.050 767.400 ;
        RECT 781.950 768.600 784.050 769.050 ;
        RECT 829.950 768.600 832.050 769.050 ;
        RECT 781.950 767.400 832.050 768.600 ;
        RECT 781.950 766.950 784.050 767.400 ;
        RECT 829.950 766.950 832.050 767.400 ;
        RECT 847.950 768.600 850.050 769.050 ;
        RECT 901.950 768.600 904.050 769.050 ;
        RECT 847.950 767.400 904.050 768.600 ;
        RECT 847.950 766.950 850.050 767.400 ;
        RECT 901.950 766.950 904.050 767.400 ;
        RECT 685.950 765.600 688.050 766.050 ;
        RECT 677.400 764.400 688.050 765.600 ;
        RECT 640.950 763.950 643.050 764.400 ;
        RECT 646.950 763.950 649.050 764.400 ;
        RECT 685.950 763.950 688.050 764.400 ;
        RECT 727.950 765.600 730.050 766.050 ;
        RECT 745.950 765.600 748.050 766.050 ;
        RECT 727.950 764.400 748.050 765.600 ;
        RECT 727.950 763.950 730.050 764.400 ;
        RECT 745.950 763.950 748.050 764.400 ;
        RECT 754.950 765.600 757.050 766.050 ;
        RECT 766.950 765.600 769.050 766.050 ;
        RECT 754.950 764.400 769.050 765.600 ;
        RECT 754.950 763.950 757.050 764.400 ;
        RECT 766.950 763.950 769.050 764.400 ;
        RECT 844.950 765.600 849.000 766.050 ;
        RECT 922.950 765.600 925.050 766.050 ;
        RECT 934.950 765.600 937.050 766.050 ;
        RECT 844.950 763.950 849.600 765.600 ;
        RECT 922.950 764.400 937.050 765.600 ;
        RECT 922.950 763.950 925.050 764.400 ;
        RECT 934.950 763.950 937.050 764.400 ;
        RECT 550.950 761.400 573.600 762.600 ;
        RECT 493.950 756.600 496.050 757.050 ;
        RECT 505.950 756.600 508.050 757.050 ;
        RECT 493.950 755.400 508.050 756.600 ;
        RECT 524.400 756.600 525.600 761.100 ;
        RECT 550.950 760.950 553.050 761.400 ;
        RECT 589.950 760.950 592.050 763.050 ;
        RECT 631.950 761.100 634.050 763.200 ;
        RECT 646.950 762.750 649.050 762.900 ;
        RECT 655.950 762.750 658.050 763.200 ;
        RECT 646.950 761.550 658.050 762.750 ;
        RECT 541.950 756.600 544.050 756.900 ;
        RECT 524.400 755.400 544.050 756.600 ;
        RECT 493.950 754.950 496.050 755.400 ;
        RECT 505.950 754.950 508.050 755.400 ;
        RECT 541.950 754.800 544.050 755.400 ;
        RECT 577.950 756.600 580.050 757.050 ;
        RECT 590.400 756.600 591.600 760.950 ;
        RECT 625.950 759.600 628.050 759.900 ;
        RECT 632.400 759.600 633.600 761.100 ;
        RECT 646.950 760.800 649.050 761.550 ;
        RECT 655.950 761.100 658.050 761.550 ;
        RECT 709.950 762.600 712.050 763.200 ;
        RECT 709.950 761.400 714.600 762.600 ;
        RECT 709.950 761.100 712.050 761.400 ;
        RECT 667.950 759.600 670.050 760.050 ;
        RECT 625.950 758.400 670.050 759.600 ;
        RECT 625.950 757.800 628.050 758.400 ;
        RECT 667.950 757.950 670.050 758.400 ;
        RECT 713.400 757.050 714.600 761.400 ;
        RECT 727.950 761.100 730.050 763.200 ;
        RECT 733.950 762.750 736.050 763.200 ;
        RECT 739.950 762.750 742.050 763.200 ;
        RECT 733.950 761.550 742.050 762.750 ;
        RECT 733.950 761.100 736.050 761.550 ;
        RECT 739.950 761.100 742.050 761.550 ;
        RECT 802.950 762.600 805.050 763.200 ;
        RECT 802.950 761.400 807.600 762.600 ;
        RECT 802.950 761.100 805.050 761.400 ;
        RECT 577.950 755.400 591.600 756.600 ;
        RECT 595.950 756.600 598.050 757.050 ;
        RECT 616.950 756.600 619.050 756.900 ;
        RECT 595.950 755.400 619.050 756.600 ;
        RECT 577.950 754.950 580.050 755.400 ;
        RECT 595.950 754.950 598.050 755.400 ;
        RECT 616.950 754.800 619.050 755.400 ;
        RECT 682.950 756.600 685.050 756.900 ;
        RECT 691.950 756.600 694.050 757.050 ;
        RECT 682.950 755.400 694.050 756.600 ;
        RECT 682.950 754.800 685.050 755.400 ;
        RECT 691.950 754.950 694.050 755.400 ;
        RECT 712.950 754.950 715.050 757.050 ;
        RECT 728.400 754.050 729.600 761.100 ;
        RECT 790.950 759.600 793.050 760.050 ;
        RECT 779.400 758.400 801.600 759.600 ;
        RECT 739.950 756.600 742.050 757.050 ;
        RECT 754.950 756.600 757.050 756.900 ;
        RECT 739.950 755.400 757.050 756.600 ;
        RECT 739.950 754.950 742.050 755.400 ;
        RECT 754.950 754.800 757.050 755.400 ;
        RECT 760.950 756.600 763.050 757.050 ;
        RECT 779.400 756.900 780.600 758.400 ;
        RECT 790.950 757.950 793.050 758.400 ;
        RECT 800.400 756.900 801.600 758.400 ;
        RECT 772.950 756.600 775.050 756.900 ;
        RECT 760.950 755.400 775.050 756.600 ;
        RECT 760.950 754.950 763.050 755.400 ;
        RECT 772.950 754.800 775.050 755.400 ;
        RECT 778.950 754.800 781.050 756.900 ;
        RECT 799.950 754.800 802.050 756.900 ;
        RECT 806.400 756.600 807.600 761.400 ;
        RECT 808.950 761.100 811.050 763.200 ;
        RECT 814.950 762.600 817.050 763.050 ;
        RECT 829.950 762.600 832.050 763.200 ;
        RECT 814.950 761.400 832.050 762.600 ;
        RECT 809.400 759.600 810.600 761.100 ;
        RECT 814.950 760.950 817.050 761.400 ;
        RECT 829.950 761.100 832.050 761.400 ;
        RECT 841.950 760.950 844.050 763.050 ;
        RECT 848.400 762.600 849.600 763.950 ;
        RECT 859.950 762.750 862.050 763.200 ;
        RECT 868.950 762.750 871.050 763.200 ;
        RECT 848.400 761.400 855.600 762.600 ;
        RECT 842.400 759.600 843.600 760.950 ;
        RECT 809.400 758.400 816.600 759.600 ;
        RECT 842.400 758.400 849.600 759.600 ;
        RECT 811.950 756.600 814.050 757.050 ;
        RECT 806.400 755.400 814.050 756.600 ;
        RECT 815.400 756.600 816.600 758.400 ;
        RECT 826.950 756.600 829.050 756.900 ;
        RECT 844.950 756.600 847.050 756.900 ;
        RECT 815.400 755.400 847.050 756.600 ;
        RECT 848.400 756.600 849.600 758.400 ;
        RECT 854.400 756.600 855.600 761.400 ;
        RECT 859.950 761.550 871.050 762.750 ;
        RECT 859.950 761.100 862.050 761.550 ;
        RECT 868.950 761.100 871.050 761.550 ;
        RECT 895.950 762.600 898.050 763.200 ;
        RECT 904.950 762.600 907.050 763.050 ;
        RECT 895.950 761.400 907.050 762.600 ;
        RECT 895.950 761.100 898.050 761.400 ;
        RECT 904.950 760.950 907.050 761.400 ;
        RECT 919.950 762.750 922.050 763.200 ;
        RECT 925.950 762.750 928.050 763.200 ;
        RECT 919.950 761.550 928.050 762.750 ;
        RECT 919.950 761.100 922.050 761.550 ;
        RECT 925.950 761.100 928.050 761.550 ;
        RECT 865.950 756.600 868.050 756.900 ;
        RECT 848.400 755.400 852.600 756.600 ;
        RECT 854.400 755.400 868.050 756.600 ;
        RECT 811.950 754.950 814.050 755.400 ;
        RECT 826.950 754.800 829.050 755.400 ;
        RECT 844.950 754.800 847.050 755.400 ;
        RECT 136.950 753.600 139.050 754.050 ;
        RECT 125.400 752.400 139.050 753.600 ;
        RECT 136.950 751.950 139.050 752.400 ;
        RECT 205.950 753.600 208.050 754.050 ;
        RECT 211.950 753.600 214.050 754.050 ;
        RECT 205.950 752.400 214.050 753.600 ;
        RECT 205.950 751.950 208.050 752.400 ;
        RECT 211.950 751.950 214.050 752.400 ;
        RECT 430.950 753.600 433.050 754.050 ;
        RECT 442.950 753.600 445.050 754.050 ;
        RECT 430.950 752.400 445.050 753.600 ;
        RECT 430.950 751.950 433.050 752.400 ;
        RECT 442.950 751.950 445.050 752.400 ;
        RECT 478.950 751.950 481.050 754.050 ;
        RECT 496.950 753.600 499.050 754.050 ;
        RECT 514.950 753.600 517.050 754.050 ;
        RECT 496.950 752.400 517.050 753.600 ;
        RECT 496.950 751.950 499.050 752.400 ;
        RECT 514.950 751.950 517.050 752.400 ;
        RECT 598.950 753.600 601.050 754.050 ;
        RECT 604.800 753.600 606.900 754.050 ;
        RECT 598.950 752.400 606.900 753.600 ;
        RECT 598.950 751.950 601.050 752.400 ;
        RECT 604.800 751.950 606.900 752.400 ;
        RECT 607.950 753.600 610.050 754.050 ;
        RECT 658.950 753.600 661.050 754.050 ;
        RECT 694.950 753.600 697.050 754.050 ;
        RECT 607.950 752.400 661.050 753.600 ;
        RECT 607.950 751.950 610.050 752.400 ;
        RECT 658.950 751.950 661.050 752.400 ;
        RECT 677.400 752.400 697.050 753.600 ;
        RECT 97.950 750.600 100.050 751.050 ;
        RECT 115.950 750.600 118.050 751.050 ;
        RECT 97.950 749.400 118.050 750.600 ;
        RECT 97.950 748.950 100.050 749.400 ;
        RECT 115.950 748.950 118.050 749.400 ;
        RECT 121.950 750.600 124.050 751.050 ;
        RECT 136.950 750.600 139.050 750.900 ;
        RECT 121.950 749.400 139.050 750.600 ;
        RECT 121.950 748.950 124.050 749.400 ;
        RECT 136.950 748.800 139.050 749.400 ;
        RECT 196.950 750.600 199.050 751.050 ;
        RECT 223.950 750.600 226.050 751.050 ;
        RECT 256.950 750.600 259.050 751.050 ;
        RECT 196.950 749.400 259.050 750.600 ;
        RECT 196.950 748.950 199.050 749.400 ;
        RECT 223.950 748.950 226.050 749.400 ;
        RECT 256.950 748.950 259.050 749.400 ;
        RECT 304.950 750.600 307.050 751.050 ;
        RECT 352.950 750.600 355.050 751.050 ;
        RECT 304.950 749.400 355.050 750.600 ;
        RECT 304.950 748.950 307.050 749.400 ;
        RECT 352.950 748.950 355.050 749.400 ;
        RECT 367.950 750.600 370.050 751.050 ;
        RECT 406.950 750.600 409.050 751.050 ;
        RECT 367.950 749.400 409.050 750.600 ;
        RECT 367.950 748.950 370.050 749.400 ;
        RECT 406.950 748.950 409.050 749.400 ;
        RECT 451.950 750.600 454.050 751.050 ;
        RECT 520.950 750.600 523.050 751.050 ;
        RECT 451.950 749.400 523.050 750.600 ;
        RECT 605.400 750.600 606.600 751.950 ;
        RECT 677.400 750.600 678.600 752.400 ;
        RECT 694.950 751.950 697.050 752.400 ;
        RECT 727.950 751.950 730.050 754.050 ;
        RECT 802.950 753.600 805.050 754.050 ;
        RECT 820.950 753.600 823.050 754.050 ;
        RECT 802.950 752.400 823.050 753.600 ;
        RECT 851.400 753.600 852.600 755.400 ;
        RECT 865.950 754.800 868.050 755.400 ;
        RECT 871.950 756.600 874.050 756.900 ;
        RECT 910.950 756.600 913.050 756.900 ;
        RECT 871.950 755.400 913.050 756.600 ;
        RECT 871.950 754.800 874.050 755.400 ;
        RECT 910.950 754.800 913.050 755.400 ;
        RECT 851.400 752.400 867.600 753.600 ;
        RECT 802.950 751.950 805.050 752.400 ;
        RECT 820.950 751.950 823.050 752.400 ;
        RECT 605.400 749.400 678.600 750.600 ;
        RECT 706.950 750.600 709.050 751.050 ;
        RECT 715.950 750.600 718.050 751.050 ;
        RECT 706.950 749.400 718.050 750.600 ;
        RECT 451.950 748.950 454.050 749.400 ;
        RECT 520.950 748.950 523.050 749.400 ;
        RECT 706.950 748.950 709.050 749.400 ;
        RECT 715.950 748.950 718.050 749.400 ;
        RECT 730.950 750.600 733.050 751.050 ;
        RECT 742.950 750.600 745.050 751.050 ;
        RECT 730.950 749.400 745.050 750.600 ;
        RECT 730.950 748.950 733.050 749.400 ;
        RECT 742.950 748.950 745.050 749.400 ;
        RECT 766.950 750.600 769.050 751.050 ;
        RECT 841.950 750.600 844.050 751.050 ;
        RECT 862.950 750.600 865.050 751.050 ;
        RECT 766.950 749.400 844.050 750.600 ;
        RECT 766.950 748.950 769.050 749.400 ;
        RECT 841.950 748.950 844.050 749.400 ;
        RECT 851.400 749.400 865.050 750.600 ;
        RECT 866.400 750.600 867.600 752.400 ;
        RECT 874.800 750.600 876.900 751.050 ;
        RECT 866.400 749.400 876.900 750.600 ;
        RECT 851.400 748.050 852.600 749.400 ;
        RECT 862.950 748.950 865.050 749.400 ;
        RECT 874.800 748.950 876.900 749.400 ;
        RECT 877.950 750.600 880.050 751.050 ;
        RECT 889.950 750.600 892.050 751.050 ;
        RECT 877.950 749.400 892.050 750.600 ;
        RECT 877.950 748.950 880.050 749.400 ;
        RECT 889.950 748.950 892.050 749.400 ;
        RECT 904.950 750.600 907.050 751.050 ;
        RECT 916.950 750.600 919.050 751.050 ;
        RECT 904.950 749.400 919.050 750.600 ;
        RECT 904.950 748.950 907.050 749.400 ;
        RECT 916.950 748.950 919.050 749.400 ;
        RECT 25.950 747.600 28.050 748.050 ;
        RECT 37.950 747.600 40.050 748.050 ;
        RECT 25.950 746.400 40.050 747.600 ;
        RECT 25.950 745.950 28.050 746.400 ;
        RECT 37.950 745.950 40.050 746.400 ;
        RECT 52.950 747.600 55.050 748.050 ;
        RECT 115.800 747.600 117.900 747.900 ;
        RECT 52.950 746.400 117.900 747.600 ;
        RECT 52.950 745.950 55.050 746.400 ;
        RECT 115.800 745.800 117.900 746.400 ;
        RECT 118.950 747.600 121.050 748.050 ;
        RECT 142.950 747.600 145.050 748.050 ;
        RECT 205.950 747.600 208.050 748.050 ;
        RECT 118.950 746.400 208.050 747.600 ;
        RECT 118.950 745.950 121.050 746.400 ;
        RECT 142.950 745.950 145.050 746.400 ;
        RECT 205.950 745.950 208.050 746.400 ;
        RECT 259.950 747.600 262.050 748.050 ;
        RECT 295.950 747.600 298.050 748.050 ;
        RECT 259.950 746.400 298.050 747.600 ;
        RECT 259.950 745.950 262.050 746.400 ;
        RECT 295.950 745.950 298.050 746.400 ;
        RECT 505.950 747.600 508.050 748.050 ;
        RECT 520.950 747.600 523.050 747.900 ;
        RECT 550.950 747.600 553.050 748.050 ;
        RECT 505.950 746.400 553.050 747.600 ;
        RECT 505.950 745.950 508.050 746.400 ;
        RECT 520.950 745.800 523.050 746.400 ;
        RECT 550.950 745.950 553.050 746.400 ;
        RECT 577.950 747.600 580.050 748.050 ;
        RECT 592.950 747.600 595.050 748.050 ;
        RECT 577.950 746.400 595.050 747.600 ;
        RECT 577.950 745.950 580.050 746.400 ;
        RECT 592.950 745.950 595.050 746.400 ;
        RECT 616.950 747.600 619.050 748.050 ;
        RECT 628.950 747.600 631.050 748.050 ;
        RECT 616.950 746.400 631.050 747.600 ;
        RECT 616.950 745.950 619.050 746.400 ;
        RECT 628.950 745.950 631.050 746.400 ;
        RECT 658.950 747.600 661.050 748.050 ;
        RECT 676.950 747.600 679.050 748.050 ;
        RECT 658.950 746.400 679.050 747.600 ;
        RECT 658.950 745.950 661.050 746.400 ;
        RECT 676.950 745.950 679.050 746.400 ;
        RECT 682.950 747.600 685.050 748.050 ;
        RECT 763.950 747.600 766.050 748.050 ;
        RECT 682.950 746.400 766.050 747.600 ;
        RECT 682.950 745.950 685.050 746.400 ;
        RECT 763.950 745.950 766.050 746.400 ;
        RECT 787.950 747.600 790.050 748.050 ;
        RECT 850.950 747.600 853.050 748.050 ;
        RECT 787.950 746.400 853.050 747.600 ;
        RECT 787.950 745.950 790.050 746.400 ;
        RECT 850.950 745.950 853.050 746.400 ;
        RECT 97.950 744.600 100.050 745.050 ;
        RECT 109.950 744.600 112.050 745.050 ;
        RECT 97.950 743.400 112.050 744.600 ;
        RECT 97.950 742.950 100.050 743.400 ;
        RECT 109.950 742.950 112.050 743.400 ;
        RECT 130.950 744.600 133.050 745.050 ;
        RECT 268.950 744.600 271.050 745.050 ;
        RECT 130.950 743.400 271.050 744.600 ;
        RECT 130.950 742.950 133.050 743.400 ;
        RECT 268.950 742.950 271.050 743.400 ;
        RECT 370.950 744.600 373.050 745.050 ;
        RECT 409.950 744.600 412.050 745.050 ;
        RECT 460.950 744.600 463.050 745.050 ;
        RECT 370.950 743.400 438.600 744.600 ;
        RECT 370.950 742.950 373.050 743.400 ;
        RECT 409.950 742.950 412.050 743.400 ;
        RECT 94.950 741.600 97.050 742.050 ;
        RECT 131.400 741.600 132.600 742.950 ;
        RECT 94.950 740.400 132.600 741.600 ;
        RECT 136.950 741.600 139.050 742.050 ;
        RECT 151.950 741.600 154.050 742.050 ;
        RECT 136.950 740.400 154.050 741.600 ;
        RECT 94.950 739.950 97.050 740.400 ;
        RECT 136.950 739.950 139.050 740.400 ;
        RECT 151.950 739.950 154.050 740.400 ;
        RECT 265.950 741.600 268.050 742.050 ;
        RECT 310.800 741.600 312.900 742.050 ;
        RECT 265.950 740.400 312.900 741.600 ;
        RECT 265.950 739.950 268.050 740.400 ;
        RECT 310.800 739.950 312.900 740.400 ;
        RECT 313.950 741.600 316.050 742.050 ;
        RECT 328.950 741.600 331.050 742.050 ;
        RECT 376.950 741.600 379.050 742.050 ;
        RECT 313.950 740.400 331.050 741.600 ;
        RECT 313.950 739.950 316.050 740.400 ;
        RECT 328.950 739.950 331.050 740.400 ;
        RECT 332.400 740.400 379.050 741.600 ;
        RECT 437.400 741.600 438.600 743.400 ;
        RECT 449.400 743.400 463.050 744.600 ;
        RECT 449.400 741.600 450.600 743.400 ;
        RECT 460.950 742.950 463.050 743.400 ;
        RECT 502.950 744.600 505.050 745.050 ;
        RECT 547.950 744.600 550.050 745.050 ;
        RECT 502.950 743.400 550.050 744.600 ;
        RECT 502.950 742.950 505.050 743.400 ;
        RECT 547.950 742.950 550.050 743.400 ;
        RECT 595.950 744.600 598.050 745.050 ;
        RECT 646.950 744.600 649.050 745.050 ;
        RECT 595.950 743.400 649.050 744.600 ;
        RECT 595.950 742.950 598.050 743.400 ;
        RECT 646.950 742.950 649.050 743.400 ;
        RECT 703.950 744.600 706.050 745.050 ;
        RECT 721.950 744.600 724.050 745.050 ;
        RECT 760.950 744.600 763.050 745.050 ;
        RECT 703.950 743.400 763.050 744.600 ;
        RECT 703.950 742.950 706.050 743.400 ;
        RECT 721.950 742.950 724.050 743.400 ;
        RECT 760.950 742.950 763.050 743.400 ;
        RECT 790.950 744.600 793.050 745.050 ;
        RECT 805.950 744.600 808.050 745.050 ;
        RECT 790.950 743.400 808.050 744.600 ;
        RECT 790.950 742.950 793.050 743.400 ;
        RECT 805.950 742.950 808.050 743.400 ;
        RECT 829.950 744.600 832.050 745.050 ;
        RECT 841.950 744.600 844.050 745.050 ;
        RECT 883.950 744.600 886.050 745.050 ;
        RECT 829.950 743.400 886.050 744.600 ;
        RECT 829.950 742.950 832.050 743.400 ;
        RECT 841.950 742.950 844.050 743.400 ;
        RECT 883.950 742.950 886.050 743.400 ;
        RECT 892.950 744.600 895.050 745.050 ;
        RECT 913.950 744.600 916.050 745.050 ;
        RECT 925.950 744.600 928.050 745.050 ;
        RECT 892.950 743.400 928.050 744.600 ;
        RECT 892.950 742.950 895.050 743.400 ;
        RECT 913.950 742.950 916.050 743.400 ;
        RECT 925.950 742.950 928.050 743.400 ;
        RECT 437.400 740.400 450.600 741.600 ;
        RECT 454.950 741.600 457.050 742.050 ;
        RECT 481.950 741.600 484.050 742.050 ;
        RECT 454.950 740.400 484.050 741.600 ;
        RECT 70.950 738.600 73.050 739.050 ;
        RECT 82.950 738.600 85.050 739.050 ;
        RECT 70.950 737.400 85.050 738.600 ;
        RECT 70.950 736.950 73.050 737.400 ;
        RECT 82.950 736.950 85.050 737.400 ;
        RECT 211.950 738.600 214.050 739.050 ;
        RECT 332.400 738.600 333.600 740.400 ;
        RECT 376.950 739.950 379.050 740.400 ;
        RECT 454.950 739.950 457.050 740.400 ;
        RECT 481.950 739.950 484.050 740.400 ;
        RECT 529.950 741.600 532.050 742.050 ;
        RECT 562.950 741.600 565.050 742.050 ;
        RECT 529.950 740.400 565.050 741.600 ;
        RECT 529.950 739.950 532.050 740.400 ;
        RECT 562.950 739.950 565.050 740.400 ;
        RECT 649.950 741.600 652.050 742.050 ;
        RECT 682.950 741.600 685.050 742.050 ;
        RECT 649.950 740.400 685.050 741.600 ;
        RECT 649.950 739.950 652.050 740.400 ;
        RECT 682.950 739.950 685.050 740.400 ;
        RECT 688.950 741.600 691.050 742.050 ;
        RECT 748.950 741.600 751.050 742.050 ;
        RECT 688.950 740.400 751.050 741.600 ;
        RECT 688.950 739.950 691.050 740.400 ;
        RECT 748.950 739.950 751.050 740.400 ;
        RECT 763.950 741.600 766.050 742.050 ;
        RECT 784.950 741.600 787.050 742.050 ;
        RECT 763.950 740.400 787.050 741.600 ;
        RECT 763.950 739.950 766.050 740.400 ;
        RECT 784.950 739.950 787.050 740.400 ;
        RECT 844.950 741.600 847.050 742.050 ;
        RECT 856.950 741.600 859.050 742.050 ;
        RECT 844.950 740.400 859.050 741.600 ;
        RECT 844.950 739.950 847.050 740.400 ;
        RECT 856.950 739.950 859.050 740.400 ;
        RECT 880.950 741.600 883.050 742.050 ;
        RECT 880.950 740.400 888.600 741.600 ;
        RECT 880.950 739.950 883.050 740.400 ;
        RECT 211.950 737.400 333.600 738.600 ;
        RECT 361.950 738.600 364.050 739.050 ;
        RECT 379.950 738.600 382.050 739.050 ;
        RECT 361.950 737.400 382.050 738.600 ;
        RECT 211.950 736.950 214.050 737.400 ;
        RECT 361.950 736.950 364.050 737.400 ;
        RECT 379.950 736.950 382.050 737.400 ;
        RECT 499.950 738.600 502.050 739.050 ;
        RECT 526.950 738.600 529.050 739.050 ;
        RECT 499.950 737.400 529.050 738.600 ;
        RECT 499.950 736.950 502.050 737.400 ;
        RECT 526.950 736.950 529.050 737.400 ;
        RECT 586.950 738.600 589.050 739.050 ;
        RECT 607.950 738.600 610.050 739.050 ;
        RECT 586.950 737.400 610.050 738.600 ;
        RECT 586.950 736.950 589.050 737.400 ;
        RECT 607.950 736.950 610.050 737.400 ;
        RECT 619.950 738.600 622.050 739.050 ;
        RECT 625.950 738.600 628.050 739.050 ;
        RECT 619.950 737.400 628.050 738.600 ;
        RECT 619.950 736.950 622.050 737.400 ;
        RECT 625.950 736.950 628.050 737.400 ;
        RECT 766.950 738.600 769.050 739.050 ;
        RECT 781.950 738.600 784.050 739.050 ;
        RECT 766.950 737.400 784.050 738.600 ;
        RECT 766.950 736.950 769.050 737.400 ;
        RECT 781.950 736.950 784.050 737.400 ;
        RECT 793.950 736.950 799.050 739.050 ;
        RECT 862.950 738.600 865.050 739.050 ;
        RECT 877.950 738.600 880.050 739.050 ;
        RECT 862.950 737.400 880.050 738.600 ;
        RECT 887.400 738.600 888.600 740.400 ;
        RECT 898.950 738.600 901.050 739.050 ;
        RECT 887.400 737.400 901.050 738.600 ;
        RECT 862.950 736.950 865.050 737.400 ;
        RECT 877.950 736.950 880.050 737.400 ;
        RECT 898.950 736.950 901.050 737.400 ;
        RECT 28.950 735.600 31.050 736.050 ;
        RECT 61.950 735.600 64.050 736.050 ;
        RECT 85.950 735.600 88.050 736.050 ;
        RECT 28.950 734.400 88.050 735.600 ;
        RECT 28.950 733.950 31.050 734.400 ;
        RECT 61.950 733.950 64.050 734.400 ;
        RECT 85.950 733.950 88.050 734.400 ;
        RECT 115.950 735.600 118.050 736.050 ;
        RECT 121.950 735.600 124.050 736.050 ;
        RECT 148.950 735.600 151.050 736.050 ;
        RECT 115.950 734.400 124.050 735.600 ;
        RECT 115.950 733.950 118.050 734.400 ;
        RECT 121.950 733.950 124.050 734.400 ;
        RECT 140.400 734.400 151.050 735.600 ;
        RECT 82.950 732.600 85.050 733.050 ;
        RECT 109.950 732.600 112.050 733.050 ;
        RECT 140.400 732.600 141.600 734.400 ;
        RECT 148.950 733.950 151.050 734.400 ;
        RECT 160.950 735.600 163.050 736.050 ;
        RECT 166.950 735.600 169.050 736.050 ;
        RECT 175.950 735.600 178.050 736.050 ;
        RECT 160.950 734.400 178.050 735.600 ;
        RECT 160.950 733.950 163.050 734.400 ;
        RECT 166.950 733.950 169.050 734.400 ;
        RECT 175.950 733.950 178.050 734.400 ;
        RECT 223.950 735.600 226.050 736.050 ;
        RECT 247.950 735.600 250.050 736.050 ;
        RECT 223.950 734.400 250.050 735.600 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 247.950 733.950 250.050 734.400 ;
        RECT 268.950 735.600 271.050 736.050 ;
        RECT 355.950 735.600 358.050 736.050 ;
        RECT 400.950 735.600 403.050 736.050 ;
        RECT 268.950 734.400 358.050 735.600 ;
        RECT 268.950 733.950 271.050 734.400 ;
        RECT 355.950 733.950 358.050 734.400 ;
        RECT 359.400 734.400 403.050 735.600 ;
        RECT 157.950 732.600 160.050 733.050 ;
        RECT 82.950 731.400 112.050 732.600 ;
        RECT 82.950 730.950 85.050 731.400 ;
        RECT 109.950 730.950 112.050 731.400 ;
        RECT 131.400 731.400 141.600 732.600 ;
        RECT 143.400 731.400 160.050 732.600 ;
        RECT 19.950 729.600 22.050 730.050 ;
        RECT 31.950 729.600 34.050 730.200 ;
        RECT 19.950 728.400 34.050 729.600 ;
        RECT 19.950 727.950 22.050 728.400 ;
        RECT 31.950 728.100 34.050 728.400 ;
        RECT 52.950 729.750 55.050 730.200 ;
        RECT 58.950 729.750 61.050 730.200 ;
        RECT 52.950 728.550 61.050 729.750 ;
        RECT 52.950 728.100 55.050 728.550 ;
        RECT 58.950 728.100 61.050 728.550 ;
        RECT 79.950 727.950 82.050 730.050 ;
        RECT 109.950 729.600 112.050 730.200 ;
        RECT 124.950 729.600 127.050 730.200 ;
        RECT 109.950 728.400 127.050 729.600 ;
        RECT 109.950 728.100 112.050 728.400 ;
        RECT 124.950 728.100 127.050 728.400 ;
        RECT 67.950 723.600 70.050 723.900 ;
        RECT 80.400 723.600 81.600 727.950 ;
        RECT 131.400 726.600 132.600 731.400 ;
        RECT 143.400 730.200 144.600 731.400 ;
        RECT 157.950 730.950 160.050 731.400 ;
        RECT 211.950 732.600 214.050 733.050 ;
        RECT 253.950 732.600 256.050 733.050 ;
        RECT 265.950 732.600 268.050 733.050 ;
        RECT 211.950 731.400 237.600 732.600 ;
        RECT 211.950 730.950 214.050 731.400 ;
        RECT 133.950 727.950 136.050 730.050 ;
        RECT 142.950 728.100 145.050 730.200 ;
        RECT 193.950 729.750 196.050 730.200 ;
        RECT 202.950 729.750 205.050 730.200 ;
        RECT 193.950 728.550 205.050 729.750 ;
        RECT 193.950 728.100 196.050 728.550 ;
        RECT 202.950 728.100 205.050 728.550 ;
        RECT 220.950 729.600 223.050 730.050 ;
        RECT 232.950 729.600 235.050 730.200 ;
        RECT 220.950 728.400 235.050 729.600 ;
        RECT 220.950 727.950 223.050 728.400 ;
        RECT 232.950 728.100 235.050 728.400 ;
        RECT 119.400 726.000 132.600 726.600 ;
        RECT 118.950 725.400 132.600 726.000 ;
        RECT 67.950 722.400 81.600 723.600 ;
        RECT 82.950 723.450 85.050 723.900 ;
        RECT 91.950 723.450 94.050 723.900 ;
        RECT 67.950 721.800 70.050 722.400 ;
        RECT 82.950 722.250 94.050 723.450 ;
        RECT 82.950 721.800 85.050 722.250 ;
        RECT 91.950 721.800 94.050 722.250 ;
        RECT 100.950 723.450 103.050 723.900 ;
        RECT 112.950 723.450 115.050 723.900 ;
        RECT 100.950 722.250 115.050 723.450 ;
        RECT 100.950 721.800 103.050 722.250 ;
        RECT 112.950 721.800 115.050 722.250 ;
        RECT 118.950 721.950 121.050 725.400 ;
        RECT 134.400 723.600 135.600 727.950 ;
        RECT 236.400 723.900 237.600 731.400 ;
        RECT 253.950 731.400 268.050 732.600 ;
        RECT 253.950 730.950 256.050 731.400 ;
        RECT 265.950 730.950 268.050 731.400 ;
        RECT 280.950 732.600 283.050 733.050 ;
        RECT 280.950 731.400 288.600 732.600 ;
        RECT 280.950 730.950 283.050 731.400 ;
        RECT 238.950 729.600 241.050 730.200 ;
        RECT 244.950 729.600 247.050 730.050 ;
        RECT 277.950 729.600 280.050 730.200 ;
        RECT 238.950 728.400 280.050 729.600 ;
        RECT 287.400 729.600 288.600 731.400 ;
        RECT 316.950 730.950 319.050 733.050 ;
        RECT 334.950 732.600 337.050 733.050 ;
        RECT 359.400 732.600 360.600 734.400 ;
        RECT 400.950 733.950 403.050 734.400 ;
        RECT 433.950 735.600 436.050 736.050 ;
        RECT 448.950 735.600 451.050 736.050 ;
        RECT 511.950 735.600 514.050 736.050 ;
        RECT 433.950 734.400 451.050 735.600 ;
        RECT 433.950 733.950 436.050 734.400 ;
        RECT 448.950 733.950 451.050 734.400 ;
        RECT 503.400 734.400 514.050 735.600 ;
        RECT 334.950 731.400 360.600 732.600 ;
        RECT 379.950 732.600 382.050 733.050 ;
        RECT 412.950 732.600 415.050 733.050 ;
        RECT 379.950 731.400 415.050 732.600 ;
        RECT 334.950 730.950 337.050 731.400 ;
        RECT 379.950 730.950 382.050 731.400 ;
        RECT 412.950 730.950 415.050 731.400 ;
        RECT 298.950 729.750 301.050 730.200 ;
        RECT 304.950 729.750 307.050 730.200 ;
        RECT 298.950 729.600 307.050 729.750 ;
        RECT 287.400 728.550 307.050 729.600 ;
        RECT 287.400 728.400 301.050 728.550 ;
        RECT 238.950 728.100 241.050 728.400 ;
        RECT 244.950 727.950 247.050 728.400 ;
        RECT 277.950 728.100 280.050 728.400 ;
        RECT 298.950 728.100 301.050 728.400 ;
        RECT 304.950 728.100 307.050 728.550 ;
        RECT 317.400 726.600 318.600 730.950 ;
        RECT 364.950 729.600 367.050 730.050 ;
        RECT 376.950 729.600 379.050 730.200 ;
        RECT 364.950 728.400 375.600 729.600 ;
        RECT 364.950 727.950 367.050 728.400 ;
        RECT 317.400 725.400 324.600 726.600 ;
        RECT 323.400 723.900 324.600 725.400 ;
        RECT 374.400 723.900 375.600 728.400 ;
        RECT 376.950 728.400 381.600 729.600 ;
        RECT 376.950 728.100 379.050 728.400 ;
        RECT 125.400 722.400 135.600 723.600 ;
        RECT 208.950 723.450 211.050 723.900 ;
        RECT 220.950 723.450 223.050 723.900 ;
        RECT 125.400 721.050 126.600 722.400 ;
        RECT 208.950 722.250 223.050 723.450 ;
        RECT 208.950 721.800 211.050 722.250 ;
        RECT 220.950 721.800 223.050 722.250 ;
        RECT 235.950 721.800 238.050 723.900 ;
        RECT 250.950 723.450 253.050 723.900 ;
        RECT 265.950 723.450 268.050 723.900 ;
        RECT 250.950 722.250 268.050 723.450 ;
        RECT 250.950 721.800 253.050 722.250 ;
        RECT 265.950 721.800 268.050 722.250 ;
        RECT 307.950 723.450 310.050 723.900 ;
        RECT 316.950 723.450 319.050 723.900 ;
        RECT 307.950 722.250 319.050 723.450 ;
        RECT 307.950 721.800 310.050 722.250 ;
        RECT 316.950 721.800 319.050 722.250 ;
        RECT 322.950 723.450 325.050 723.900 ;
        RECT 343.950 723.450 346.050 723.900 ;
        RECT 322.950 722.250 346.050 723.450 ;
        RECT 322.950 721.800 325.050 722.250 ;
        RECT 343.950 721.800 346.050 722.250 ;
        RECT 373.950 721.800 376.050 723.900 ;
        RECT 380.400 721.050 381.600 728.400 ;
        RECT 388.800 727.950 390.900 730.050 ;
        RECT 391.950 729.600 394.050 730.050 ;
        RECT 421.950 729.600 424.050 730.200 ;
        RECT 391.950 728.400 424.050 729.600 ;
        RECT 391.950 727.950 394.050 728.400 ;
        RECT 421.950 728.100 424.050 728.400 ;
        RECT 436.950 727.950 439.050 730.050 ;
        RECT 442.950 729.600 445.050 730.200 ;
        RECT 454.950 729.600 457.050 730.050 ;
        RECT 442.950 728.400 457.050 729.600 ;
        RECT 442.950 728.100 445.050 728.400 ;
        RECT 454.950 727.950 457.050 728.400 ;
        RECT 463.950 729.750 466.050 730.200 ;
        RECT 475.950 729.750 478.050 730.200 ;
        RECT 463.950 728.550 478.050 729.750 ;
        RECT 463.950 728.100 466.050 728.550 ;
        RECT 475.950 728.100 478.050 728.550 ;
        RECT 487.950 729.600 490.050 730.200 ;
        RECT 503.400 729.600 504.600 734.400 ;
        RECT 511.950 733.950 514.050 734.400 ;
        RECT 613.950 735.600 616.050 736.050 ;
        RECT 625.950 735.600 628.050 735.900 ;
        RECT 613.950 734.400 628.050 735.600 ;
        RECT 613.950 733.950 616.050 734.400 ;
        RECT 625.950 733.800 628.050 734.400 ;
        RECT 676.950 735.600 679.050 736.050 ;
        RECT 700.950 735.600 703.050 736.050 ;
        RECT 676.950 734.400 703.050 735.600 ;
        RECT 676.950 733.950 679.050 734.400 ;
        RECT 700.950 733.950 703.050 734.400 ;
        RECT 733.950 735.600 736.050 736.050 ;
        RECT 763.950 735.600 766.050 736.050 ;
        RECT 733.950 734.400 766.050 735.600 ;
        RECT 733.950 733.950 736.050 734.400 ;
        RECT 763.950 733.950 766.050 734.400 ;
        RECT 784.950 735.600 787.050 735.900 ;
        RECT 799.800 735.600 801.900 736.050 ;
        RECT 784.950 734.400 801.900 735.600 ;
        RECT 610.950 732.600 613.050 732.900 ;
        RECT 616.950 732.600 619.050 733.050 ;
        RECT 610.950 731.400 619.050 732.600 ;
        RECT 610.950 730.800 613.050 731.400 ;
        RECT 616.950 730.950 619.050 731.400 ;
        RECT 622.950 732.600 625.050 733.050 ;
        RECT 646.950 732.600 649.050 733.050 ;
        RECT 677.400 732.600 678.600 733.950 ;
        RECT 784.950 733.800 787.050 734.400 ;
        RECT 799.800 733.950 801.900 734.400 ;
        RECT 802.950 735.600 805.050 736.050 ;
        RECT 811.950 735.600 814.050 736.050 ;
        RECT 802.950 734.400 814.050 735.600 ;
        RECT 802.950 733.950 805.050 734.400 ;
        RECT 811.950 733.950 814.050 734.400 ;
        RECT 820.950 735.600 823.050 736.050 ;
        RECT 826.950 735.600 829.050 736.050 ;
        RECT 850.950 735.600 853.050 736.050 ;
        RECT 820.950 734.400 853.050 735.600 ;
        RECT 820.950 733.950 823.050 734.400 ;
        RECT 826.950 733.950 829.050 734.400 ;
        RECT 850.950 733.950 853.050 734.400 ;
        RECT 856.950 733.950 859.050 736.050 ;
        RECT 904.950 735.600 907.050 736.050 ;
        RECT 884.400 734.400 907.050 735.600 ;
        RECT 622.950 731.400 649.050 732.600 ;
        RECT 622.950 730.950 625.050 731.400 ;
        RECT 646.950 730.950 649.050 731.400 ;
        RECT 656.400 731.400 678.600 732.600 ;
        RECT 505.950 729.600 508.050 730.200 ;
        RECT 487.950 728.400 508.050 729.600 ;
        RECT 487.950 728.100 490.050 728.400 ;
        RECT 505.950 728.100 508.050 728.400 ;
        RECT 511.950 729.600 514.050 730.200 ;
        RECT 532.950 729.750 535.050 730.200 ;
        RECT 541.950 729.750 544.050 730.200 ;
        RECT 532.950 729.600 544.050 729.750 ;
        RECT 547.950 729.600 550.050 730.200 ;
        RECT 511.950 728.550 544.050 729.600 ;
        RECT 511.950 728.400 535.050 728.550 ;
        RECT 511.950 728.100 514.050 728.400 ;
        RECT 532.950 728.100 535.050 728.400 ;
        RECT 541.950 728.100 544.050 728.550 ;
        RECT 545.400 728.400 550.050 729.600 ;
        RECT 389.250 724.050 390.450 727.950 ;
        RECT 388.800 721.950 390.900 724.050 ;
        RECT 403.950 723.600 406.050 723.900 ;
        RECT 418.950 723.600 421.050 723.900 ;
        RECT 437.400 723.600 438.600 727.950 ;
        RECT 439.950 723.600 442.050 723.900 ;
        RECT 403.950 722.400 421.050 723.600 ;
        RECT 403.950 721.800 406.050 722.400 ;
        RECT 418.950 721.800 421.050 722.400 ;
        RECT 434.400 722.400 442.050 723.600 ;
        RECT 10.950 720.600 13.050 721.050 ;
        RECT 22.950 720.600 25.050 721.050 ;
        RECT 10.950 719.400 25.050 720.600 ;
        RECT 10.950 718.950 13.050 719.400 ;
        RECT 22.950 718.950 25.050 719.400 ;
        RECT 106.950 720.600 109.050 721.050 ;
        RECT 115.950 720.600 118.050 721.050 ;
        RECT 106.950 719.400 118.050 720.600 ;
        RECT 106.950 718.950 109.050 719.400 ;
        RECT 115.950 718.950 118.050 719.400 ;
        RECT 121.950 719.400 126.600 721.050 ;
        RECT 169.950 720.600 172.050 721.050 ;
        RECT 190.950 720.600 193.050 721.050 ;
        RECT 169.950 719.400 193.050 720.600 ;
        RECT 121.950 718.950 126.000 719.400 ;
        RECT 169.950 718.950 172.050 719.400 ;
        RECT 190.950 718.950 193.050 719.400 ;
        RECT 229.950 720.600 232.050 721.050 ;
        RECT 241.950 720.600 244.050 721.050 ;
        RECT 268.950 720.600 271.050 721.050 ;
        RECT 229.950 719.400 271.050 720.600 ;
        RECT 380.400 719.400 385.050 721.050 ;
        RECT 229.950 718.950 232.050 719.400 ;
        RECT 241.950 718.950 244.050 719.400 ;
        RECT 268.950 718.950 271.050 719.400 ;
        RECT 381.000 718.950 385.050 719.400 ;
        RECT 394.950 720.600 397.050 721.050 ;
        RECT 434.400 720.600 435.600 722.400 ;
        RECT 439.950 721.800 442.050 722.400 ;
        RECT 445.950 723.600 448.050 723.900 ;
        RECT 460.950 723.600 463.050 723.900 ;
        RECT 478.950 723.600 481.050 727.050 ;
        RECT 545.400 726.600 546.600 728.400 ;
        RECT 547.950 728.100 550.050 728.400 ;
        RECT 601.950 728.100 604.050 730.200 ;
        RECT 602.400 726.600 603.600 728.100 ;
        RECT 539.400 726.000 546.600 726.600 ;
        RECT 538.950 725.400 546.600 726.000 ;
        RECT 596.400 725.400 603.600 726.600 ;
        RECT 445.950 722.400 463.050 723.600 ;
        RECT 445.950 721.800 448.050 722.400 ;
        RECT 460.950 721.800 463.050 722.400 ;
        RECT 467.400 723.000 481.050 723.600 ;
        RECT 496.950 723.600 499.050 724.050 ;
        RECT 508.950 723.600 511.050 723.900 ;
        RECT 467.400 722.400 480.600 723.000 ;
        RECT 496.950 722.400 511.050 723.600 ;
        RECT 394.950 719.400 435.600 720.600 ;
        RECT 442.950 720.600 445.050 721.050 ;
        RECT 467.400 720.600 468.600 722.400 ;
        RECT 496.950 721.950 499.050 722.400 ;
        RECT 508.950 721.800 511.050 722.400 ;
        RECT 520.950 723.450 523.050 723.900 ;
        RECT 529.950 723.450 532.050 723.900 ;
        RECT 520.950 722.250 532.050 723.450 ;
        RECT 520.950 721.800 523.050 722.250 ;
        RECT 529.950 721.800 532.050 722.250 ;
        RECT 538.950 721.950 541.050 725.400 ;
        RECT 596.400 723.600 597.600 725.400 ;
        RECT 656.400 723.900 657.600 731.400 ;
        RECT 658.950 729.600 661.050 730.200 ;
        RECT 682.950 729.600 685.050 730.200 ;
        RECT 691.950 729.600 694.050 733.050 ;
        RECT 709.950 732.600 712.050 733.050 ;
        RECT 718.950 732.600 721.050 733.050 ;
        RECT 709.950 731.400 721.050 732.600 ;
        RECT 709.950 730.950 712.050 731.400 ;
        RECT 718.950 730.950 721.050 731.400 ;
        RECT 772.950 732.600 775.050 733.050 ;
        RECT 808.950 732.600 811.050 733.050 ;
        RECT 847.950 732.600 850.050 733.050 ;
        RECT 772.950 731.400 850.050 732.600 ;
        RECT 772.950 730.950 775.050 731.400 ;
        RECT 808.950 730.950 811.050 731.400 ;
        RECT 847.950 730.950 850.050 731.400 ;
        RECT 697.950 729.600 700.050 730.200 ;
        RECT 712.950 729.600 715.050 730.050 ;
        RECT 724.800 729.600 726.900 730.050 ;
        RECT 658.950 728.400 666.600 729.600 ;
        RECT 658.950 728.100 661.050 728.400 ;
        RECT 665.400 724.050 666.600 728.400 ;
        RECT 682.950 728.400 690.600 729.600 ;
        RECT 691.950 729.000 700.050 729.600 ;
        RECT 692.400 728.400 700.050 729.000 ;
        RECT 682.950 728.100 685.050 728.400 ;
        RECT 689.400 726.600 690.600 728.400 ;
        RECT 697.950 728.100 700.050 728.400 ;
        RECT 707.400 728.400 715.050 729.600 ;
        RECT 689.400 725.400 696.600 726.600 ;
        RECT 584.400 723.000 597.600 723.600 ;
        RECT 583.950 722.400 597.600 723.000 ;
        RECT 442.950 719.400 468.600 720.600 ;
        RECT 394.950 718.950 397.050 719.400 ;
        RECT 442.950 718.950 445.050 719.400 ;
        RECT 583.950 718.950 586.050 722.400 ;
        RECT 655.950 721.800 658.050 723.900 ;
        RECT 664.950 721.950 667.050 724.050 ;
        RECT 695.400 723.900 696.600 725.400 ;
        RECT 707.400 724.050 708.600 728.400 ;
        RECT 712.950 727.950 715.050 728.400 ;
        RECT 716.400 728.400 726.900 729.600 ;
        RECT 716.400 726.600 717.600 728.400 ;
        RECT 724.800 727.950 726.900 728.400 ;
        RECT 727.950 726.600 730.050 730.050 ;
        RECT 754.950 729.600 757.050 730.200 ;
        RECT 778.950 729.600 781.050 730.200 ;
        RECT 802.950 729.600 805.050 730.200 ;
        RECT 814.950 729.600 817.050 730.200 ;
        RECT 754.950 728.400 781.050 729.600 ;
        RECT 754.950 728.100 757.050 728.400 ;
        RECT 778.950 728.100 781.050 728.400 ;
        RECT 791.400 728.400 805.050 729.600 ;
        RECT 713.400 726.000 717.600 726.600 ;
        RECT 712.950 725.400 717.600 726.000 ;
        RECT 719.400 726.000 730.050 726.600 ;
        RECT 719.400 725.400 729.600 726.000 ;
        RECT 694.950 721.800 697.050 723.900 ;
        RECT 706.950 721.950 709.050 724.050 ;
        RECT 712.950 721.950 715.050 725.400 ;
        RECT 719.400 723.900 720.600 725.400 ;
        RECT 791.400 724.050 792.600 728.400 ;
        RECT 802.950 728.100 805.050 728.400 ;
        RECT 806.400 728.400 817.050 729.600 ;
        RECT 806.400 726.600 807.600 728.400 ;
        RECT 814.950 728.100 817.050 728.400 ;
        RECT 800.400 725.400 807.600 726.600 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 757.950 723.450 760.050 723.900 ;
        RECT 763.950 723.450 766.050 723.900 ;
        RECT 757.950 722.250 766.050 723.450 ;
        RECT 757.950 721.800 760.050 722.250 ;
        RECT 763.950 721.800 766.050 722.250 ;
        RECT 775.950 723.450 778.050 723.900 ;
        RECT 784.950 723.450 787.050 723.900 ;
        RECT 775.950 722.250 787.050 723.450 ;
        RECT 775.950 721.800 778.050 722.250 ;
        RECT 784.950 721.800 787.050 722.250 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 800.400 723.900 801.600 725.400 ;
        RECT 857.400 724.050 858.600 733.950 ;
        RECT 859.950 732.600 862.050 733.050 ;
        RECT 865.950 732.600 868.050 733.050 ;
        RECT 859.950 731.400 868.050 732.600 ;
        RECT 859.950 730.950 862.050 731.400 ;
        RECT 865.950 730.950 868.050 731.400 ;
        RECT 865.950 729.600 868.050 730.200 ;
        RECT 877.950 729.600 880.050 730.050 ;
        RECT 865.950 728.400 880.050 729.600 ;
        RECT 865.950 728.100 868.050 728.400 ;
        RECT 877.950 727.950 880.050 728.400 ;
        RECT 884.400 726.600 885.600 734.400 ;
        RECT 904.950 733.950 907.050 734.400 ;
        RECT 886.800 730.950 888.900 733.050 ;
        RECT 889.950 732.600 892.050 733.050 ;
        RECT 895.950 732.600 898.050 733.050 ;
        RECT 889.950 731.400 898.050 732.600 ;
        RECT 889.950 730.950 892.050 731.400 ;
        RECT 895.950 730.950 898.050 731.400 ;
        RECT 878.400 726.000 885.600 726.600 ;
        RECT 877.950 725.400 885.600 726.000 ;
        RECT 887.400 729.600 888.600 730.950 ;
        RECT 901.950 729.600 904.050 730.050 ;
        RECT 887.400 728.400 904.050 729.600 ;
        RECT 799.950 721.800 802.050 723.900 ;
        RECT 823.950 723.450 826.050 723.900 ;
        RECT 829.950 723.450 832.050 723.900 ;
        RECT 823.950 722.250 832.050 723.450 ;
        RECT 823.950 721.800 826.050 722.250 ;
        RECT 829.950 721.800 832.050 722.250 ;
        RECT 856.950 721.950 859.050 724.050 ;
        RECT 877.950 721.950 880.050 725.400 ;
        RECT 887.400 723.900 888.600 728.400 ;
        RECT 901.950 727.950 904.050 728.400 ;
        RECT 907.950 729.750 910.050 730.200 ;
        RECT 919.950 729.750 922.050 730.200 ;
        RECT 907.950 728.550 922.050 729.750 ;
        RECT 907.950 728.100 910.050 728.550 ;
        RECT 919.950 728.100 922.050 728.550 ;
        RECT 886.950 721.800 889.050 723.900 ;
        RECT 598.950 720.600 601.050 721.050 ;
        RECT 607.950 720.600 610.050 721.050 ;
        RECT 598.950 719.400 610.050 720.600 ;
        RECT 598.950 718.950 601.050 719.400 ;
        RECT 607.950 718.950 610.050 719.400 ;
        RECT 616.950 720.600 619.050 721.050 ;
        RECT 622.950 720.600 625.050 721.050 ;
        RECT 634.950 720.600 637.050 721.050 ;
        RECT 616.950 719.400 637.050 720.600 ;
        RECT 616.950 718.950 619.050 719.400 ;
        RECT 622.950 718.950 625.050 719.400 ;
        RECT 634.950 718.950 637.050 719.400 ;
        RECT 838.950 720.600 841.050 721.050 ;
        RECT 853.950 720.600 856.050 721.050 ;
        RECT 838.950 719.400 856.050 720.600 ;
        RECT 838.950 718.950 841.050 719.400 ;
        RECT 853.950 718.950 856.050 719.400 ;
        RECT 862.950 720.600 865.050 721.050 ;
        RECT 871.950 720.600 874.050 720.900 ;
        RECT 901.950 720.600 904.050 721.050 ;
        RECT 862.950 719.400 874.050 720.600 ;
        RECT 862.950 718.950 865.050 719.400 ;
        RECT 871.950 718.800 874.050 719.400 ;
        RECT 890.400 719.400 904.050 720.600 ;
        RECT 274.950 717.600 277.050 718.050 ;
        RECT 304.950 717.600 307.050 718.050 ;
        RECT 331.950 717.600 334.050 718.050 ;
        RECT 274.950 716.400 334.050 717.600 ;
        RECT 274.950 715.950 277.050 716.400 ;
        RECT 304.950 715.950 307.050 716.400 ;
        RECT 331.950 715.950 334.050 716.400 ;
        RECT 352.950 717.600 355.050 718.050 ;
        RECT 376.950 717.600 379.050 717.900 ;
        RECT 352.950 716.400 379.050 717.600 ;
        RECT 352.950 715.950 355.050 716.400 ;
        RECT 376.950 715.800 379.050 716.400 ;
        RECT 424.950 717.600 427.050 718.050 ;
        RECT 445.950 717.600 448.050 718.050 ;
        RECT 424.950 716.400 448.050 717.600 ;
        RECT 424.950 715.950 427.050 716.400 ;
        RECT 445.950 715.950 448.050 716.400 ;
        RECT 484.950 717.600 487.050 718.050 ;
        RECT 514.950 717.600 517.050 718.050 ;
        RECT 538.950 717.600 541.050 718.050 ;
        RECT 574.950 717.600 577.050 718.050 ;
        RECT 484.950 716.400 577.050 717.600 ;
        RECT 484.950 715.950 487.050 716.400 ;
        RECT 514.950 715.950 517.050 716.400 ;
        RECT 538.950 715.950 541.050 716.400 ;
        RECT 574.950 715.950 577.050 716.400 ;
        RECT 700.950 717.600 703.050 718.050 ;
        RECT 721.950 717.600 724.050 718.050 ;
        RECT 730.950 717.600 733.050 718.050 ;
        RECT 700.950 716.400 733.050 717.600 ;
        RECT 700.950 715.950 703.050 716.400 ;
        RECT 721.950 715.950 724.050 716.400 ;
        RECT 730.950 715.950 733.050 716.400 ;
        RECT 772.950 717.600 775.050 718.050 ;
        RECT 793.950 717.600 796.050 718.050 ;
        RECT 772.950 716.400 796.050 717.600 ;
        RECT 772.950 715.950 775.050 716.400 ;
        RECT 793.950 715.950 796.050 716.400 ;
        RECT 853.950 717.600 856.050 717.900 ;
        RECT 880.800 717.600 882.900 717.900 ;
        RECT 853.950 716.400 882.900 717.600 ;
        RECT 853.950 715.800 856.050 716.400 ;
        RECT 880.800 715.800 882.900 716.400 ;
        RECT 883.950 717.600 886.050 718.050 ;
        RECT 890.400 717.600 891.600 719.400 ;
        RECT 901.950 718.950 904.050 719.400 ;
        RECT 910.950 720.600 913.050 721.050 ;
        RECT 916.950 720.600 919.050 721.050 ;
        RECT 910.950 719.400 919.050 720.600 ;
        RECT 910.950 718.950 913.050 719.400 ;
        RECT 916.950 718.950 919.050 719.400 ;
        RECT 883.950 716.400 891.600 717.600 ;
        RECT 883.950 715.950 886.050 716.400 ;
        RECT 214.950 714.600 217.050 715.050 ;
        RECT 244.950 714.600 247.050 715.050 ;
        RECT 277.950 714.600 280.050 715.050 ;
        RECT 214.950 713.400 280.050 714.600 ;
        RECT 214.950 712.950 217.050 713.400 ;
        RECT 244.950 712.950 247.050 713.400 ;
        RECT 277.950 712.950 280.050 713.400 ;
        RECT 307.950 714.600 310.050 715.050 ;
        RECT 325.950 714.600 328.050 715.050 ;
        RECT 307.950 713.400 328.050 714.600 ;
        RECT 307.950 712.950 310.050 713.400 ;
        RECT 325.950 712.950 328.050 713.400 ;
        RECT 343.950 714.600 346.050 715.050 ;
        RECT 394.950 714.600 397.050 715.050 ;
        RECT 343.950 713.400 397.050 714.600 ;
        RECT 343.950 712.950 346.050 713.400 ;
        RECT 394.950 712.950 397.050 713.400 ;
        RECT 412.950 714.600 415.050 715.050 ;
        RECT 442.950 714.600 445.050 715.050 ;
        RECT 412.950 713.400 445.050 714.600 ;
        RECT 412.950 712.950 415.050 713.400 ;
        RECT 442.950 712.950 445.050 713.400 ;
        RECT 469.950 714.600 472.050 715.050 ;
        RECT 520.950 714.600 523.050 715.050 ;
        RECT 469.950 713.400 523.050 714.600 ;
        RECT 469.950 712.950 472.050 713.400 ;
        RECT 520.950 712.950 523.050 713.400 ;
        RECT 550.950 714.600 553.050 715.050 ;
        RECT 562.950 714.600 565.050 715.050 ;
        RECT 550.950 713.400 565.050 714.600 ;
        RECT 550.950 712.950 553.050 713.400 ;
        RECT 562.950 712.950 565.050 713.400 ;
        RECT 589.950 714.600 592.050 715.050 ;
        RECT 598.950 714.600 601.050 715.050 ;
        RECT 619.950 714.600 622.050 715.050 ;
        RECT 589.950 713.400 622.050 714.600 ;
        RECT 589.950 712.950 592.050 713.400 ;
        RECT 598.950 712.950 601.050 713.400 ;
        RECT 619.950 712.950 622.050 713.400 ;
        RECT 661.950 714.600 664.050 715.050 ;
        RECT 679.950 714.600 682.050 715.050 ;
        RECT 709.950 714.600 712.050 715.050 ;
        RECT 661.950 713.400 712.050 714.600 ;
        RECT 661.950 712.950 664.050 713.400 ;
        RECT 679.950 712.950 682.050 713.400 ;
        RECT 709.950 712.950 712.050 713.400 ;
        RECT 733.950 714.600 736.050 715.050 ;
        RECT 802.950 714.600 805.050 715.050 ;
        RECT 733.950 713.400 805.050 714.600 ;
        RECT 733.950 712.950 736.050 713.400 ;
        RECT 802.950 712.950 805.050 713.400 ;
        RECT 868.950 714.600 871.050 715.050 ;
        RECT 892.950 714.600 895.050 715.050 ;
        RECT 868.950 713.400 895.050 714.600 ;
        RECT 868.950 712.950 871.050 713.400 ;
        RECT 892.950 712.950 895.050 713.400 ;
        RECT 901.950 714.600 904.050 715.050 ;
        RECT 922.950 714.600 925.050 715.050 ;
        RECT 901.950 713.400 925.050 714.600 ;
        RECT 901.950 712.950 904.050 713.400 ;
        RECT 922.950 712.950 925.050 713.400 ;
        RECT 58.950 711.600 61.050 712.050 ;
        RECT 97.950 711.600 100.050 712.050 ;
        RECT 109.950 711.600 112.050 712.050 ;
        RECT 58.950 710.400 112.050 711.600 ;
        RECT 58.950 709.950 61.050 710.400 ;
        RECT 97.950 709.950 100.050 710.400 ;
        RECT 109.950 709.950 112.050 710.400 ;
        RECT 328.950 711.600 331.050 712.050 ;
        RECT 340.950 711.600 343.050 712.050 ;
        RECT 391.950 711.600 394.050 712.050 ;
        RECT 328.950 710.400 394.050 711.600 ;
        RECT 328.950 709.950 331.050 710.400 ;
        RECT 340.950 709.950 343.050 710.400 ;
        RECT 391.950 709.950 394.050 710.400 ;
        RECT 418.950 711.600 421.050 712.050 ;
        RECT 436.950 711.600 439.050 712.050 ;
        RECT 418.950 710.400 439.050 711.600 ;
        RECT 418.950 709.950 421.050 710.400 ;
        RECT 436.950 709.950 439.050 710.400 ;
        RECT 457.950 711.600 460.050 712.050 ;
        RECT 472.950 711.600 475.050 712.050 ;
        RECT 457.950 710.400 475.050 711.600 ;
        RECT 457.950 709.950 460.050 710.400 ;
        RECT 472.950 709.950 475.050 710.400 ;
        RECT 496.950 711.600 499.050 712.050 ;
        RECT 541.950 711.600 544.050 712.050 ;
        RECT 496.950 710.400 544.050 711.600 ;
        RECT 496.950 709.950 499.050 710.400 ;
        RECT 541.950 709.950 544.050 710.400 ;
        RECT 637.950 711.600 640.050 712.050 ;
        RECT 646.950 711.600 649.050 712.050 ;
        RECT 637.950 710.400 649.050 711.600 ;
        RECT 637.950 709.950 640.050 710.400 ;
        RECT 646.950 709.950 649.050 710.400 ;
        RECT 871.950 711.600 874.050 712.050 ;
        RECT 889.950 711.600 892.050 712.050 ;
        RECT 871.950 710.400 892.050 711.600 ;
        RECT 871.950 709.950 874.050 710.400 ;
        RECT 889.950 709.950 892.050 710.400 ;
        RECT 175.950 708.600 178.050 709.050 ;
        RECT 268.950 708.600 271.050 709.050 ;
        RECT 175.950 707.400 271.050 708.600 ;
        RECT 175.950 706.950 178.050 707.400 ;
        RECT 268.950 706.950 271.050 707.400 ;
        RECT 316.950 708.600 319.050 709.050 ;
        RECT 424.950 708.600 427.050 709.050 ;
        RECT 316.950 707.400 427.050 708.600 ;
        RECT 316.950 706.950 319.050 707.400 ;
        RECT 424.950 706.950 427.050 707.400 ;
        RECT 454.950 708.600 457.050 709.050 ;
        RECT 475.950 708.600 478.050 709.050 ;
        RECT 454.950 707.400 478.050 708.600 ;
        RECT 454.950 706.950 457.050 707.400 ;
        RECT 475.950 706.950 478.050 707.400 ;
        RECT 652.950 708.600 655.050 709.050 ;
        RECT 667.950 708.600 670.050 709.050 ;
        RECT 652.950 707.400 670.050 708.600 ;
        RECT 652.950 706.950 655.050 707.400 ;
        RECT 667.950 706.950 670.050 707.400 ;
        RECT 730.950 708.600 733.050 709.050 ;
        RECT 742.950 708.600 745.050 709.050 ;
        RECT 769.950 708.600 772.050 709.050 ;
        RECT 730.950 707.400 772.050 708.600 ;
        RECT 730.950 706.950 733.050 707.400 ;
        RECT 742.950 706.950 745.050 707.400 ;
        RECT 769.950 706.950 772.050 707.400 ;
        RECT 880.950 708.600 883.050 709.050 ;
        RECT 919.950 708.600 922.050 709.050 ;
        RECT 880.950 707.400 922.050 708.600 ;
        RECT 880.950 706.950 883.050 707.400 ;
        RECT 919.950 706.950 922.050 707.400 ;
        RECT 172.950 705.600 175.050 706.050 ;
        RECT 211.950 705.600 214.050 706.050 ;
        RECT 172.950 704.400 214.050 705.600 ;
        RECT 172.950 703.950 175.050 704.400 ;
        RECT 211.950 703.950 214.050 704.400 ;
        RECT 265.950 705.600 268.050 706.050 ;
        RECT 289.950 705.600 292.050 706.050 ;
        RECT 265.950 704.400 292.050 705.600 ;
        RECT 265.950 703.950 268.050 704.400 ;
        RECT 289.950 703.950 292.050 704.400 ;
        RECT 313.950 705.600 316.050 706.050 ;
        RECT 442.950 705.600 445.050 706.050 ;
        RECT 313.950 704.400 445.050 705.600 ;
        RECT 313.950 703.950 316.050 704.400 ;
        RECT 442.950 703.950 445.050 704.400 ;
        RECT 448.950 705.600 451.050 706.050 ;
        RECT 646.950 705.600 649.050 706.050 ;
        RECT 694.950 705.600 697.050 706.050 ;
        RECT 448.950 704.400 633.600 705.600 ;
        RECT 448.950 703.950 451.050 704.400 ;
        RECT 268.950 702.600 271.050 703.050 ;
        RECT 316.950 702.600 319.050 703.050 ;
        RECT 268.950 701.400 319.050 702.600 ;
        RECT 268.950 700.950 271.050 701.400 ;
        RECT 316.950 700.950 319.050 701.400 ;
        RECT 322.950 702.600 325.050 703.050 ;
        RECT 346.950 702.600 349.050 703.050 ;
        RECT 322.950 701.400 349.050 702.600 ;
        RECT 322.950 700.950 325.050 701.400 ;
        RECT 346.950 700.950 349.050 701.400 ;
        RECT 382.950 702.600 385.050 703.050 ;
        RECT 421.950 702.600 424.050 703.050 ;
        RECT 382.950 701.400 424.050 702.600 ;
        RECT 382.950 700.950 385.050 701.400 ;
        RECT 421.950 700.950 424.050 701.400 ;
        RECT 535.950 702.600 538.050 703.050 ;
        RECT 568.950 702.600 571.050 703.050 ;
        RECT 535.950 701.400 571.050 702.600 ;
        RECT 535.950 700.950 538.050 701.400 ;
        RECT 568.950 700.950 571.050 701.400 ;
        RECT 574.950 702.600 577.050 703.050 ;
        RECT 583.950 702.600 586.050 703.050 ;
        RECT 574.950 701.400 586.050 702.600 ;
        RECT 632.400 702.600 633.600 704.400 ;
        RECT 646.950 704.400 697.050 705.600 ;
        RECT 646.950 703.950 649.050 704.400 ;
        RECT 694.950 703.950 697.050 704.400 ;
        RECT 796.950 705.600 799.050 706.050 ;
        RECT 805.950 705.600 808.050 706.050 ;
        RECT 862.950 705.600 865.050 706.050 ;
        RECT 796.950 704.400 865.050 705.600 ;
        RECT 796.950 703.950 799.050 704.400 ;
        RECT 805.950 703.950 808.050 704.400 ;
        RECT 862.950 703.950 865.050 704.400 ;
        RECT 895.950 705.600 898.050 706.050 ;
        RECT 901.950 705.600 904.050 706.050 ;
        RECT 895.950 704.400 904.050 705.600 ;
        RECT 895.950 703.950 898.050 704.400 ;
        RECT 901.950 703.950 904.050 704.400 ;
        RECT 655.950 702.600 658.050 703.050 ;
        RECT 632.400 701.400 658.050 702.600 ;
        RECT 574.950 700.950 577.050 701.400 ;
        RECT 583.950 700.950 586.050 701.400 ;
        RECT 655.950 700.950 658.050 701.400 ;
        RECT 763.950 702.600 766.050 703.050 ;
        RECT 871.950 702.600 874.050 703.050 ;
        RECT 928.950 702.600 931.050 703.050 ;
        RECT 763.950 701.400 858.600 702.600 ;
        RECT 763.950 700.950 766.050 701.400 ;
        RECT 301.950 699.600 304.050 700.050 ;
        RECT 310.950 699.600 313.050 700.050 ;
        RECT 301.950 698.400 313.050 699.600 ;
        RECT 301.950 697.950 304.050 698.400 ;
        RECT 310.950 697.950 313.050 698.400 ;
        RECT 424.950 699.600 427.050 700.050 ;
        RECT 448.950 699.600 451.050 700.050 ;
        RECT 424.950 698.400 451.050 699.600 ;
        RECT 424.950 697.950 427.050 698.400 ;
        RECT 448.950 697.950 451.050 698.400 ;
        RECT 475.950 699.600 478.050 700.050 ;
        RECT 520.950 699.600 523.050 700.050 ;
        RECT 475.950 698.400 523.050 699.600 ;
        RECT 475.950 697.950 478.050 698.400 ;
        RECT 520.950 697.950 523.050 698.400 ;
        RECT 526.950 699.600 529.050 700.050 ;
        RECT 607.950 699.600 610.050 700.050 ;
        RECT 526.950 698.400 610.050 699.600 ;
        RECT 526.950 697.950 529.050 698.400 ;
        RECT 607.950 697.950 610.050 698.400 ;
        RECT 628.950 699.600 631.050 700.050 ;
        RECT 664.950 699.600 667.050 700.050 ;
        RECT 628.950 698.400 667.050 699.600 ;
        RECT 628.950 697.950 631.050 698.400 ;
        RECT 664.950 697.950 667.050 698.400 ;
        RECT 814.950 699.600 817.050 700.050 ;
        RECT 857.400 699.600 858.600 701.400 ;
        RECT 871.950 701.400 931.050 702.600 ;
        RECT 871.950 700.950 874.050 701.400 ;
        RECT 928.950 700.950 931.050 701.400 ;
        RECT 934.950 699.600 937.050 700.050 ;
        RECT 814.950 698.400 855.600 699.600 ;
        RECT 857.400 698.400 937.050 699.600 ;
        RECT 814.950 697.950 817.050 698.400 ;
        RECT 268.950 696.600 271.050 697.050 ;
        RECT 325.950 696.600 328.050 697.050 ;
        RECT 268.950 695.400 328.050 696.600 ;
        RECT 268.950 694.950 271.050 695.400 ;
        RECT 325.950 694.950 328.050 695.400 ;
        RECT 451.950 696.600 454.050 697.050 ;
        RECT 514.950 696.600 517.050 697.050 ;
        RECT 616.950 696.600 619.050 697.050 ;
        RECT 451.950 695.400 619.050 696.600 ;
        RECT 451.950 694.950 454.050 695.400 ;
        RECT 514.950 694.950 517.050 695.400 ;
        RECT 616.950 694.950 619.050 695.400 ;
        RECT 661.950 696.600 664.050 697.050 ;
        RECT 685.950 696.600 688.050 697.050 ;
        RECT 661.950 695.400 688.050 696.600 ;
        RECT 661.950 694.950 664.050 695.400 ;
        RECT 685.950 694.950 688.050 695.400 ;
        RECT 736.950 696.600 739.050 697.050 ;
        RECT 766.950 696.600 769.050 697.050 ;
        RECT 799.950 696.600 802.050 697.050 ;
        RECT 736.950 695.400 802.050 696.600 ;
        RECT 854.400 696.600 855.600 698.400 ;
        RECT 934.950 697.950 937.050 698.400 ;
        RECT 865.950 696.600 868.050 697.050 ;
        RECT 854.400 695.400 868.050 696.600 ;
        RECT 736.950 694.950 739.050 695.400 ;
        RECT 766.950 694.950 769.050 695.400 ;
        RECT 799.950 694.950 802.050 695.400 ;
        RECT 865.950 694.950 868.050 695.400 ;
        RECT 895.950 696.600 898.050 697.050 ;
        RECT 904.950 696.600 907.050 697.050 ;
        RECT 895.950 695.400 907.050 696.600 ;
        RECT 895.950 694.950 898.050 695.400 ;
        RECT 904.950 694.950 907.050 695.400 ;
        RECT 7.950 693.600 10.050 694.050 ;
        RECT 13.950 693.600 16.050 694.050 ;
        RECT 7.950 692.400 16.050 693.600 ;
        RECT 7.950 691.950 10.050 692.400 ;
        RECT 13.950 691.950 16.050 692.400 ;
        RECT 76.950 693.600 79.050 694.050 ;
        RECT 94.950 693.600 97.050 694.050 ;
        RECT 76.950 692.400 97.050 693.600 ;
        RECT 76.950 691.950 79.050 692.400 ;
        RECT 94.950 691.950 97.050 692.400 ;
        RECT 112.950 693.600 115.050 694.050 ;
        RECT 139.950 693.600 142.050 694.050 ;
        RECT 112.950 692.400 142.050 693.600 ;
        RECT 112.950 691.950 115.050 692.400 ;
        RECT 139.950 691.950 142.050 692.400 ;
        RECT 202.950 693.600 205.050 694.050 ;
        RECT 238.950 693.600 241.050 694.050 ;
        RECT 202.950 692.400 241.050 693.600 ;
        RECT 202.950 691.950 205.050 692.400 ;
        RECT 238.950 691.950 241.050 692.400 ;
        RECT 310.950 693.600 313.050 694.050 ;
        RECT 322.950 693.600 325.050 694.050 ;
        RECT 310.950 692.400 325.050 693.600 ;
        RECT 310.950 691.950 313.050 692.400 ;
        RECT 322.950 691.950 325.050 692.400 ;
        RECT 421.950 693.600 424.050 694.050 ;
        RECT 454.950 693.600 457.050 694.050 ;
        RECT 421.950 692.400 457.050 693.600 ;
        RECT 421.950 691.950 424.050 692.400 ;
        RECT 454.950 691.950 457.050 692.400 ;
        RECT 469.950 693.600 472.050 694.050 ;
        RECT 496.950 693.600 499.050 694.050 ;
        RECT 469.950 692.400 499.050 693.600 ;
        RECT 469.950 691.950 472.050 692.400 ;
        RECT 496.950 691.950 499.050 692.400 ;
        RECT 520.950 693.600 523.050 694.050 ;
        RECT 556.950 693.600 559.050 694.050 ;
        RECT 520.950 692.400 559.050 693.600 ;
        RECT 520.950 691.950 523.050 692.400 ;
        RECT 556.950 691.950 559.050 692.400 ;
        RECT 676.950 693.600 679.050 694.050 ;
        RECT 706.950 693.600 709.050 694.050 ;
        RECT 676.950 692.400 709.050 693.600 ;
        RECT 676.950 691.950 679.050 692.400 ;
        RECT 706.950 691.950 709.050 692.400 ;
        RECT 748.950 693.600 751.050 694.050 ;
        RECT 796.950 693.600 799.050 694.050 ;
        RECT 748.950 692.400 799.050 693.600 ;
        RECT 748.950 691.950 751.050 692.400 ;
        RECT 796.950 691.950 799.050 692.400 ;
        RECT 835.950 693.600 838.050 694.050 ;
        RECT 877.950 693.600 880.050 694.050 ;
        RECT 835.950 692.400 880.050 693.600 ;
        RECT 835.950 691.950 838.050 692.400 ;
        RECT 877.950 691.950 880.050 692.400 ;
        RECT 1.950 690.600 4.050 691.050 ;
        RECT 22.950 690.600 25.050 691.050 ;
        RECT 1.950 689.400 25.050 690.600 ;
        RECT 1.950 688.950 4.050 689.400 ;
        RECT 22.950 688.950 25.050 689.400 ;
        RECT 145.950 690.600 148.050 691.050 ;
        RECT 175.950 690.600 178.050 691.050 ;
        RECT 145.950 689.400 178.050 690.600 ;
        RECT 145.950 688.950 148.050 689.400 ;
        RECT 175.950 688.950 178.050 689.400 ;
        RECT 280.950 690.600 283.050 691.050 ;
        RECT 307.950 690.600 310.050 691.050 ;
        RECT 280.950 689.400 310.050 690.600 ;
        RECT 280.950 688.950 283.050 689.400 ;
        RECT 307.950 688.950 310.050 689.400 ;
        RECT 367.950 688.950 370.050 691.050 ;
        RECT 607.950 690.600 610.050 691.050 ;
        RECT 673.950 690.600 676.050 691.050 ;
        RECT 733.950 690.600 736.050 691.050 ;
        RECT 607.950 689.400 676.050 690.600 ;
        RECT 607.950 688.950 610.050 689.400 ;
        RECT 673.950 688.950 676.050 689.400 ;
        RECT 689.400 689.400 736.050 690.600 ;
        RECT 55.950 687.600 58.050 688.050 ;
        RECT 61.950 687.600 64.050 688.050 ;
        RECT 55.950 686.400 64.050 687.600 ;
        RECT 55.950 685.950 58.050 686.400 ;
        RECT 61.950 685.950 64.050 686.400 ;
        RECT 76.950 687.600 79.050 688.050 ;
        RECT 85.950 687.600 88.050 688.050 ;
        RECT 76.950 686.400 88.050 687.600 ;
        RECT 76.950 685.950 79.050 686.400 ;
        RECT 85.950 685.950 88.050 686.400 ;
        RECT 211.800 685.950 213.900 688.050 ;
        RECT 214.950 687.600 217.050 688.200 ;
        RECT 319.950 687.600 322.050 688.050 ;
        RECT 214.950 686.400 322.050 687.600 ;
        RECT 214.950 686.100 217.050 686.400 ;
        RECT 46.800 683.100 48.900 685.200 ;
        RECT 49.950 684.600 52.050 685.050 ;
        RECT 73.950 684.600 76.050 684.900 ;
        RECT 49.950 683.400 76.050 684.600 ;
        RECT 47.400 681.600 48.600 683.100 ;
        RECT 49.950 682.950 52.050 683.400 ;
        RECT 73.950 682.800 76.050 683.400 ;
        RECT 88.950 684.600 91.050 685.050 ;
        RECT 103.950 684.600 106.050 685.200 ;
        RECT 118.950 684.600 121.050 685.200 ;
        RECT 88.950 683.400 106.050 684.600 ;
        RECT 88.950 682.950 91.050 683.400 ;
        RECT 103.950 683.100 106.050 683.400 ;
        RECT 110.400 683.400 121.050 684.600 ;
        RECT 70.950 681.600 73.050 682.050 ;
        RECT 47.400 680.400 73.050 681.600 ;
        RECT 70.950 679.950 73.050 680.400 ;
        RECT 10.950 678.600 13.050 679.050 ;
        RECT 16.950 678.600 19.050 678.900 ;
        RECT 10.950 677.400 19.050 678.600 ;
        RECT 10.950 676.950 13.050 677.400 ;
        RECT 16.950 676.800 19.050 677.400 ;
        RECT 82.950 678.450 85.050 678.900 ;
        RECT 88.950 678.450 91.050 678.900 ;
        RECT 82.950 677.250 91.050 678.450 ;
        RECT 82.950 676.800 85.050 677.250 ;
        RECT 88.950 676.800 91.050 677.250 ;
        RECT 94.950 678.450 97.050 678.900 ;
        RECT 100.950 678.450 103.050 678.900 ;
        RECT 94.950 677.250 103.050 678.450 ;
        RECT 94.950 676.800 97.050 677.250 ;
        RECT 100.950 676.800 103.050 677.250 ;
        RECT 106.950 678.600 109.050 678.900 ;
        RECT 110.400 678.600 111.600 683.400 ;
        RECT 118.950 683.100 121.050 683.400 ;
        RECT 124.950 683.100 127.050 685.200 ;
        RECT 154.950 684.600 157.050 685.050 ;
        RECT 163.950 684.600 166.050 685.050 ;
        RECT 154.950 683.400 166.050 684.600 ;
        RECT 106.950 677.400 111.600 678.600 ;
        RECT 112.950 678.600 115.050 679.050 ;
        RECT 121.950 678.600 124.050 678.900 ;
        RECT 112.950 677.400 124.050 678.600 ;
        RECT 125.400 678.600 126.600 683.100 ;
        RECT 154.950 682.950 157.050 683.400 ;
        RECT 163.950 682.950 166.050 683.400 ;
        RECT 169.950 681.600 172.050 685.050 ;
        RECT 181.950 684.750 184.050 685.200 ;
        RECT 196.950 684.750 199.050 685.200 ;
        RECT 181.950 683.550 199.050 684.750 ;
        RECT 181.950 683.100 184.050 683.550 ;
        RECT 196.950 683.100 199.050 683.550 ;
        RECT 202.950 683.100 205.050 685.200 ;
        RECT 167.400 681.000 172.050 681.600 ;
        RECT 167.400 680.400 171.600 681.000 ;
        RECT 167.400 678.900 168.600 680.400 ;
        RECT 148.950 678.600 151.050 678.900 ;
        RECT 125.400 677.400 151.050 678.600 ;
        RECT 106.950 676.800 109.050 677.400 ;
        RECT 112.950 676.950 115.050 677.400 ;
        RECT 121.950 676.800 124.050 677.400 ;
        RECT 148.950 676.800 151.050 677.400 ;
        RECT 166.950 676.800 169.050 678.900 ;
        RECT 178.950 678.600 181.050 678.900 ;
        RECT 170.400 678.450 181.050 678.600 ;
        RECT 199.950 678.600 202.050 678.900 ;
        RECT 203.400 678.600 204.600 683.100 ;
        RECT 212.400 679.050 213.600 685.950 ;
        RECT 215.400 682.050 216.600 686.100 ;
        RECT 319.950 685.950 322.050 686.400 ;
        RECT 325.950 687.600 328.050 688.050 ;
        RECT 325.950 686.400 333.600 687.600 ;
        RECT 325.950 685.950 328.050 686.400 ;
        RECT 238.950 684.750 241.050 685.200 ;
        RECT 295.800 684.750 297.900 685.200 ;
        RECT 238.950 683.550 297.900 684.750 ;
        RECT 238.950 683.100 241.050 683.550 ;
        RECT 295.800 683.100 297.900 683.550 ;
        RECT 215.400 680.400 220.050 682.050 ;
        RECT 216.000 679.950 220.050 680.400 ;
        RECT 238.950 681.600 241.050 682.050 ;
        RECT 262.950 681.600 265.050 682.050 ;
        RECT 238.950 680.400 265.050 681.600 ;
        RECT 238.950 679.950 241.050 680.400 ;
        RECT 262.950 679.950 265.050 680.400 ;
        RECT 271.950 681.600 274.050 682.050 ;
        RECT 271.950 680.400 297.600 681.600 ;
        RECT 271.950 679.950 274.050 680.400 ;
        RECT 199.950 678.450 204.600 678.600 ;
        RECT 170.400 677.400 204.600 678.450 ;
        RECT 151.950 675.600 154.050 676.050 ;
        RECT 170.400 675.600 171.600 677.400 ;
        RECT 178.950 677.250 202.050 677.400 ;
        RECT 178.950 676.800 181.050 677.250 ;
        RECT 199.950 676.800 202.050 677.250 ;
        RECT 211.950 676.950 214.050 679.050 ;
        RECT 280.950 678.600 283.050 679.050 ;
        RECT 292.950 678.600 295.050 678.900 ;
        RECT 280.950 677.400 295.050 678.600 ;
        RECT 296.400 678.600 297.600 680.400 ;
        RECT 310.950 678.600 313.050 678.900 ;
        RECT 296.400 677.400 313.050 678.600 ;
        RECT 280.950 676.950 283.050 677.400 ;
        RECT 292.950 676.800 295.050 677.400 ;
        RECT 310.950 676.800 313.050 677.400 ;
        RECT 332.400 676.050 333.600 686.400 ;
        RECT 346.950 680.100 349.050 682.200 ;
        RECT 347.400 678.600 348.600 680.100 ;
        RECT 368.400 678.600 369.600 688.950 ;
        RECT 595.950 687.600 598.050 688.050 ;
        RECT 689.400 687.600 690.600 689.400 ;
        RECT 733.950 688.950 736.050 689.400 ;
        RECT 874.950 690.600 877.050 691.050 ;
        RECT 898.950 690.600 901.050 691.050 ;
        RECT 874.950 689.400 901.050 690.600 ;
        RECT 874.950 688.950 877.050 689.400 ;
        RECT 898.950 688.950 901.050 689.400 ;
        RECT 919.950 690.600 922.050 691.050 ;
        RECT 931.950 690.600 934.050 691.050 ;
        RECT 919.950 689.400 934.050 690.600 ;
        RECT 919.950 688.950 922.050 689.400 ;
        RECT 931.950 688.950 934.050 689.400 ;
        RECT 595.950 686.400 690.600 687.600 ;
        RECT 694.950 687.600 697.050 688.050 ;
        RECT 709.950 687.600 712.050 688.050 ;
        RECT 694.950 686.400 712.050 687.600 ;
        RECT 595.950 685.950 598.050 686.400 ;
        RECT 694.950 685.950 697.050 686.400 ;
        RECT 709.950 685.950 712.050 686.400 ;
        RECT 739.950 687.600 742.050 688.050 ;
        RECT 745.950 687.600 748.050 688.050 ;
        RECT 867.000 687.600 871.050 688.050 ;
        RECT 739.950 686.400 748.050 687.600 ;
        RECT 739.950 685.950 742.050 686.400 ;
        RECT 745.950 685.950 748.050 686.400 ;
        RECT 866.400 685.950 871.050 687.600 ;
        RECT 391.950 684.750 394.050 685.200 ;
        RECT 397.950 684.750 400.050 685.200 ;
        RECT 391.950 683.550 400.050 684.750 ;
        RECT 451.950 684.600 454.050 685.200 ;
        RECT 391.950 683.100 394.050 683.550 ;
        RECT 397.950 683.100 400.050 683.550 ;
        RECT 428.400 683.400 454.050 684.600 ;
        RECT 370.950 681.600 373.050 682.050 ;
        RECT 376.950 681.600 379.050 682.050 ;
        RECT 370.950 680.400 379.050 681.600 ;
        RECT 370.950 679.950 373.050 680.400 ;
        RECT 376.950 679.950 379.050 680.400 ;
        RECT 376.950 678.600 379.050 678.900 ;
        RECT 347.400 677.400 354.600 678.600 ;
        RECT 368.400 677.400 379.050 678.600 ;
        RECT 151.950 674.400 171.600 675.600 ;
        RECT 193.950 675.600 196.050 676.050 ;
        RECT 205.950 675.600 208.050 676.050 ;
        RECT 193.950 674.400 208.050 675.600 ;
        RECT 151.950 673.950 154.050 674.400 ;
        RECT 193.950 673.950 196.050 674.400 ;
        RECT 205.950 673.950 208.050 674.400 ;
        RECT 265.950 675.600 268.050 676.050 ;
        RECT 295.950 675.600 298.050 676.050 ;
        RECT 265.950 674.400 298.050 675.600 ;
        RECT 265.950 673.950 268.050 674.400 ;
        RECT 295.950 673.950 298.050 674.400 ;
        RECT 328.950 674.400 333.600 676.050 ;
        RECT 353.400 675.600 354.600 677.400 ;
        RECT 376.950 676.800 379.050 677.400 ;
        RECT 388.950 678.600 391.050 679.050 ;
        RECT 400.950 678.600 403.050 678.900 ;
        RECT 388.950 677.400 403.050 678.600 ;
        RECT 388.950 676.950 391.050 677.400 ;
        RECT 400.950 676.800 403.050 677.400 ;
        RECT 412.950 678.600 415.050 679.050 ;
        RECT 428.400 678.900 429.600 683.400 ;
        RECT 451.950 683.100 454.050 683.400 ;
        RECT 463.950 684.750 466.050 685.200 ;
        RECT 475.950 684.750 478.050 685.200 ;
        RECT 463.950 683.550 478.050 684.750 ;
        RECT 463.950 683.100 466.050 683.550 ;
        RECT 475.950 683.100 478.050 683.550 ;
        RECT 484.950 683.100 487.050 685.200 ;
        RECT 502.950 684.600 505.050 685.200 ;
        RECT 562.950 684.600 565.050 685.200 ;
        RECT 580.950 684.600 583.050 685.050 ;
        RECT 502.950 683.400 583.050 684.600 ;
        RECT 502.950 683.100 505.050 683.400 ;
        RECT 562.950 683.100 565.050 683.400 ;
        RECT 421.950 678.600 424.050 678.900 ;
        RECT 412.950 677.400 424.050 678.600 ;
        RECT 412.950 676.950 415.050 677.400 ;
        RECT 421.950 676.800 424.050 677.400 ;
        RECT 427.950 676.800 430.050 678.900 ;
        RECT 454.950 678.600 457.050 679.050 ;
        RECT 460.950 678.600 463.050 679.050 ;
        RECT 454.950 677.400 463.050 678.600 ;
        RECT 454.950 676.950 457.050 677.400 ;
        RECT 460.950 676.950 463.050 677.400 ;
        RECT 478.950 678.600 481.050 679.050 ;
        RECT 485.400 678.600 486.600 683.100 ;
        RECT 580.950 682.950 583.050 683.400 ;
        RECT 592.950 681.600 595.050 685.050 ;
        RECT 622.950 683.100 625.050 685.200 ;
        RECT 634.950 684.750 637.050 685.200 ;
        RECT 640.950 684.750 643.050 685.200 ;
        RECT 634.950 683.550 643.050 684.750 ;
        RECT 634.950 683.100 637.050 683.550 ;
        RECT 640.950 683.100 643.050 683.550 ;
        RECT 667.950 684.600 670.050 685.200 ;
        RECT 682.950 684.600 685.050 685.200 ;
        RECT 667.950 683.400 685.050 684.600 ;
        RECT 667.950 683.100 670.050 683.400 ;
        RECT 682.950 683.100 685.050 683.400 ;
        RECT 691.950 684.600 694.050 685.050 ;
        RECT 700.950 684.600 703.050 685.200 ;
        RECT 691.950 683.400 703.050 684.600 ;
        RECT 584.400 681.000 595.050 681.600 ;
        RECT 584.400 680.400 594.600 681.000 ;
        RECT 478.950 677.400 486.600 678.600 ;
        RECT 529.950 678.600 532.050 678.900 ;
        RECT 559.950 678.600 562.050 678.900 ;
        RECT 584.400 678.600 585.600 680.400 ;
        RECT 529.950 677.400 562.050 678.600 ;
        RECT 581.400 678.000 585.600 678.600 ;
        RECT 478.950 676.950 481.050 677.400 ;
        RECT 529.950 676.800 532.050 677.400 ;
        RECT 559.950 676.800 562.050 677.400 ;
        RECT 580.950 677.400 585.600 678.000 ;
        RECT 604.950 678.600 607.050 678.900 ;
        RECT 623.400 678.600 624.600 683.100 ;
        RECT 691.950 682.950 694.050 683.400 ;
        RECT 700.950 683.100 703.050 683.400 ;
        RECT 694.950 681.600 697.050 682.050 ;
        RECT 712.950 681.600 715.050 685.050 ;
        RECT 718.950 681.600 721.050 685.050 ;
        RECT 724.950 684.750 727.050 684.900 ;
        RECT 730.950 684.750 733.050 685.200 ;
        RECT 724.950 683.550 733.050 684.750 ;
        RECT 724.950 682.800 727.050 683.550 ;
        RECT 730.950 683.100 733.050 683.550 ;
        RECT 757.950 684.600 760.050 685.200 ;
        RECT 772.950 684.600 775.050 685.200 ;
        RECT 757.950 683.400 775.050 684.600 ;
        RECT 757.950 683.100 760.050 683.400 ;
        RECT 772.950 683.100 775.050 683.400 ;
        RECT 778.950 684.750 781.050 685.200 ;
        RECT 784.950 684.750 787.050 685.200 ;
        RECT 778.950 683.550 787.050 684.750 ;
        RECT 778.950 683.100 781.050 683.550 ;
        RECT 784.950 683.100 787.050 683.550 ;
        RECT 811.950 684.600 814.050 685.050 ;
        RECT 817.950 684.600 820.050 685.200 ;
        RECT 811.950 683.400 820.050 684.600 ;
        RECT 811.950 682.950 814.050 683.400 ;
        RECT 817.950 683.100 820.050 683.400 ;
        RECT 823.950 684.600 826.050 685.200 ;
        RECT 829.950 684.600 832.050 685.050 ;
        RECT 823.950 683.400 832.050 684.600 ;
        RECT 823.950 683.100 826.050 683.400 ;
        RECT 829.950 682.950 832.050 683.400 ;
        RECT 838.950 682.950 841.050 685.050 ;
        RECT 694.950 681.000 715.050 681.600 ;
        RECT 716.400 681.000 721.050 681.600 ;
        RECT 694.950 680.400 714.600 681.000 ;
        RECT 716.400 680.400 720.600 681.000 ;
        RECT 694.950 679.950 697.050 680.400 ;
        RECT 604.950 677.400 624.600 678.600 ;
        RECT 625.950 678.600 628.050 678.900 ;
        RECT 634.950 678.600 637.050 679.050 ;
        RECT 625.950 677.400 637.050 678.600 ;
        RECT 442.950 675.600 445.050 676.050 ;
        RECT 475.950 675.600 478.050 676.050 ;
        RECT 353.400 674.400 357.600 675.600 ;
        RECT 328.950 673.950 333.000 674.400 ;
        RECT 70.950 672.600 73.050 673.050 ;
        RECT 85.950 672.600 88.050 673.050 ;
        RECT 70.950 671.400 88.050 672.600 ;
        RECT 70.950 670.950 73.050 671.400 ;
        RECT 85.950 670.950 88.050 671.400 ;
        RECT 91.950 672.600 94.050 673.050 ;
        RECT 103.950 672.600 106.050 673.050 ;
        RECT 91.950 671.400 106.050 672.600 ;
        RECT 91.950 670.950 94.050 671.400 ;
        RECT 103.950 670.950 106.050 671.400 ;
        RECT 223.950 672.600 226.050 673.050 ;
        RECT 271.950 672.600 274.050 673.050 ;
        RECT 223.950 671.400 274.050 672.600 ;
        RECT 223.950 670.950 226.050 671.400 ;
        RECT 271.950 670.950 274.050 671.400 ;
        RECT 283.950 672.600 286.050 673.050 ;
        RECT 298.950 672.600 301.050 673.050 ;
        RECT 283.950 671.400 301.050 672.600 ;
        RECT 356.400 672.600 357.600 674.400 ;
        RECT 442.950 674.400 478.050 675.600 ;
        RECT 442.950 673.950 445.050 674.400 ;
        RECT 475.950 673.950 478.050 674.400 ;
        RECT 580.950 673.950 583.050 677.400 ;
        RECT 604.950 676.800 607.050 677.400 ;
        RECT 625.950 676.800 628.050 677.400 ;
        RECT 634.950 676.950 637.050 677.400 ;
        RECT 655.950 678.600 658.050 679.050 ;
        RECT 716.400 678.900 717.600 680.400 ;
        RECT 664.950 678.600 667.050 678.900 ;
        RECT 655.950 677.400 667.050 678.600 ;
        RECT 655.950 676.950 658.050 677.400 ;
        RECT 664.950 676.800 667.050 677.400 ;
        RECT 685.950 678.450 688.050 678.900 ;
        RECT 691.950 678.450 694.050 678.900 ;
        RECT 685.950 677.250 694.050 678.450 ;
        RECT 685.950 676.800 688.050 677.250 ;
        RECT 691.950 676.800 694.050 677.250 ;
        RECT 715.950 676.800 718.050 678.900 ;
        RECT 724.950 678.600 727.050 679.050 ;
        RECT 742.950 678.600 745.050 678.900 ;
        RECT 724.950 678.450 745.050 678.600 ;
        RECT 754.950 678.450 757.050 678.900 ;
        RECT 724.950 677.400 757.050 678.450 ;
        RECT 724.950 676.950 727.050 677.400 ;
        RECT 742.950 677.250 757.050 677.400 ;
        RECT 742.950 676.800 745.050 677.250 ;
        RECT 754.950 676.800 757.050 677.250 ;
        RECT 787.950 678.600 790.050 679.050 ;
        RECT 826.950 678.600 829.050 678.900 ;
        RECT 787.950 677.400 829.050 678.600 ;
        RECT 787.950 676.950 790.050 677.400 ;
        RECT 826.950 676.800 829.050 677.400 ;
        RECT 839.400 676.050 840.600 682.950 ;
        RECT 850.950 678.600 853.050 679.050 ;
        RECT 862.950 678.600 865.050 678.900 ;
        RECT 866.400 678.600 867.600 685.950 ;
        RECT 871.950 684.750 874.050 685.200 ;
        RECT 880.950 684.750 883.050 685.200 ;
        RECT 871.950 683.550 883.050 684.750 ;
        RECT 871.950 683.100 874.050 683.550 ;
        RECT 880.950 683.100 883.050 683.550 ;
        RECT 889.950 682.950 892.050 685.050 ;
        RECT 895.950 682.950 898.050 685.050 ;
        RECT 913.950 684.750 916.050 685.200 ;
        RECT 925.950 684.750 928.050 685.200 ;
        RECT 913.950 683.550 928.050 684.750 ;
        RECT 913.950 683.100 916.050 683.550 ;
        RECT 925.950 683.100 928.050 683.550 ;
        RECT 931.950 683.100 934.050 685.200 ;
        RECT 850.950 677.400 867.600 678.600 ;
        RECT 850.950 676.950 853.050 677.400 ;
        RECT 862.950 676.800 865.050 677.400 ;
        RECT 586.950 675.600 589.050 676.050 ;
        RECT 595.950 675.600 598.050 676.050 ;
        RECT 586.950 674.400 598.050 675.600 ;
        RECT 586.950 673.950 589.050 674.400 ;
        RECT 595.950 673.950 598.050 674.400 ;
        RECT 775.950 675.600 778.050 676.050 ;
        RECT 808.950 675.600 811.050 676.050 ;
        RECT 775.950 674.400 811.050 675.600 ;
        RECT 775.950 673.950 778.050 674.400 ;
        RECT 808.950 673.950 811.050 674.400 ;
        RECT 838.950 673.950 841.050 676.050 ;
        RECT 880.950 675.600 883.050 676.050 ;
        RECT 890.400 675.600 891.600 682.950 ;
        RECT 896.400 679.050 897.600 682.950 ;
        RECT 932.400 679.050 933.600 683.100 ;
        RECT 895.950 676.950 898.050 679.050 ;
        RECT 907.950 678.600 910.050 678.900 ;
        RECT 928.950 678.600 931.050 678.900 ;
        RECT 907.950 677.400 931.050 678.600 ;
        RECT 932.400 677.400 937.050 679.050 ;
        RECT 907.950 676.800 910.050 677.400 ;
        RECT 928.950 676.800 931.050 677.400 ;
        RECT 933.000 676.950 937.050 677.400 ;
        RECT 901.950 675.600 904.050 676.050 ;
        RECT 880.950 674.400 904.050 675.600 ;
        RECT 880.950 673.950 883.050 674.400 ;
        RECT 901.950 673.950 904.050 674.400 ;
        RECT 400.950 672.600 403.050 673.050 ;
        RECT 356.400 671.400 403.050 672.600 ;
        RECT 283.950 670.950 286.050 671.400 ;
        RECT 298.950 670.950 301.050 671.400 ;
        RECT 400.950 670.950 403.050 671.400 ;
        RECT 409.950 672.600 412.050 673.050 ;
        RECT 418.950 672.600 421.050 673.050 ;
        RECT 409.950 671.400 421.050 672.600 ;
        RECT 409.950 670.950 412.050 671.400 ;
        RECT 418.950 670.950 421.050 671.400 ;
        RECT 433.950 672.600 436.050 673.050 ;
        RECT 445.950 672.600 448.050 673.050 ;
        RECT 466.950 672.600 469.050 673.050 ;
        RECT 499.950 672.600 502.050 673.050 ;
        RECT 433.950 671.400 502.050 672.600 ;
        RECT 433.950 670.950 436.050 671.400 ;
        RECT 445.950 670.950 448.050 671.400 ;
        RECT 466.950 670.950 469.050 671.400 ;
        RECT 499.950 670.950 502.050 671.400 ;
        RECT 667.950 672.600 670.050 673.050 ;
        RECT 694.950 672.600 697.050 673.050 ;
        RECT 667.950 671.400 697.050 672.600 ;
        RECT 667.950 670.950 670.050 671.400 ;
        RECT 694.950 670.950 697.050 671.400 ;
        RECT 739.950 672.600 742.050 673.050 ;
        RECT 790.950 672.600 793.050 673.050 ;
        RECT 739.950 671.400 793.050 672.600 ;
        RECT 739.950 670.950 742.050 671.400 ;
        RECT 790.950 670.950 793.050 671.400 ;
        RECT 811.950 672.600 814.050 673.050 ;
        RECT 841.950 672.600 844.050 673.050 ;
        RECT 811.950 671.400 844.050 672.600 ;
        RECT 811.950 670.950 814.050 671.400 ;
        RECT 841.950 670.950 844.050 671.400 ;
        RECT 847.950 672.600 850.050 673.050 ;
        RECT 868.950 672.600 871.050 673.050 ;
        RECT 847.950 671.400 871.050 672.600 ;
        RECT 847.950 670.950 850.050 671.400 ;
        RECT 868.950 670.950 871.050 671.400 ;
        RECT 925.950 672.600 928.050 673.050 ;
        RECT 934.950 672.600 937.050 673.050 ;
        RECT 925.950 671.400 937.050 672.600 ;
        RECT 925.950 670.950 928.050 671.400 ;
        RECT 934.950 670.950 937.050 671.400 ;
        RECT 325.950 669.600 328.050 670.050 ;
        RECT 331.950 669.600 334.050 670.050 ;
        RECT 403.950 669.600 406.050 670.050 ;
        RECT 325.950 668.400 334.050 669.600 ;
        RECT 325.950 667.950 328.050 668.400 ;
        RECT 331.950 667.950 334.050 668.400 ;
        RECT 335.400 668.400 406.050 669.600 ;
        RECT 115.950 666.600 118.050 667.050 ;
        RECT 142.800 666.600 144.900 667.050 ;
        RECT 115.950 665.400 144.900 666.600 ;
        RECT 115.950 664.950 118.050 665.400 ;
        RECT 142.800 664.950 144.900 665.400 ;
        RECT 145.950 666.600 148.050 667.050 ;
        RECT 151.950 666.600 154.050 667.050 ;
        RECT 244.950 666.600 247.050 667.050 ;
        RECT 145.950 665.400 247.050 666.600 ;
        RECT 145.950 664.950 148.050 665.400 ;
        RECT 151.950 664.950 154.050 665.400 ;
        RECT 244.950 664.950 247.050 665.400 ;
        RECT 253.950 666.600 256.050 667.050 ;
        RECT 259.950 666.600 262.050 667.050 ;
        RECT 274.950 666.600 277.050 667.050 ;
        RECT 253.950 665.400 277.050 666.600 ;
        RECT 253.950 664.950 256.050 665.400 ;
        RECT 259.950 664.950 262.050 665.400 ;
        RECT 274.950 664.950 277.050 665.400 ;
        RECT 319.950 666.600 322.050 667.050 ;
        RECT 335.400 666.600 336.600 668.400 ;
        RECT 403.950 667.950 406.050 668.400 ;
        RECT 421.950 669.600 424.050 670.050 ;
        RECT 523.950 669.600 526.050 670.050 ;
        RECT 421.950 668.400 526.050 669.600 ;
        RECT 421.950 667.950 424.050 668.400 ;
        RECT 523.950 667.950 526.050 668.400 ;
        RECT 535.950 669.600 538.050 670.050 ;
        RECT 544.950 669.600 547.050 670.050 ;
        RECT 535.950 668.400 547.050 669.600 ;
        RECT 535.950 667.950 538.050 668.400 ;
        RECT 544.950 667.950 547.050 668.400 ;
        RECT 571.950 669.600 574.050 670.050 ;
        RECT 643.950 669.600 646.050 670.050 ;
        RECT 571.950 668.400 646.050 669.600 ;
        RECT 571.950 667.950 574.050 668.400 ;
        RECT 643.950 667.950 646.050 668.400 ;
        RECT 763.950 669.600 766.050 670.050 ;
        RECT 775.950 669.600 778.050 670.050 ;
        RECT 829.950 669.600 832.050 670.050 ;
        RECT 763.950 668.400 778.050 669.600 ;
        RECT 763.950 667.950 766.050 668.400 ;
        RECT 775.950 667.950 778.050 668.400 ;
        RECT 815.400 668.400 832.050 669.600 ;
        RECT 412.950 666.600 415.050 667.050 ;
        RECT 319.950 665.400 336.600 666.600 ;
        RECT 356.400 665.400 415.050 666.600 ;
        RECT 319.950 664.950 322.050 665.400 ;
        RECT 55.950 663.600 58.050 664.050 ;
        RECT 121.950 663.600 124.050 664.050 ;
        RECT 55.950 662.400 124.050 663.600 ;
        RECT 55.950 661.950 58.050 662.400 ;
        RECT 121.950 661.950 124.050 662.400 ;
        RECT 217.950 663.600 220.050 664.050 ;
        RECT 232.800 663.600 234.900 664.050 ;
        RECT 217.950 662.400 234.900 663.600 ;
        RECT 217.950 661.950 220.050 662.400 ;
        RECT 232.800 661.950 234.900 662.400 ;
        RECT 235.950 663.600 238.050 664.050 ;
        RECT 268.950 663.600 271.050 664.050 ;
        RECT 235.950 662.400 271.050 663.600 ;
        RECT 235.950 661.950 238.050 662.400 ;
        RECT 268.950 661.950 271.050 662.400 ;
        RECT 277.950 663.600 280.050 664.050 ;
        RECT 295.950 663.600 298.050 664.050 ;
        RECT 277.950 662.400 298.050 663.600 ;
        RECT 277.950 661.950 280.050 662.400 ;
        RECT 295.950 661.950 298.050 662.400 ;
        RECT 328.950 663.600 331.050 664.050 ;
        RECT 356.400 663.600 357.600 665.400 ;
        RECT 412.950 664.950 415.050 665.400 ;
        RECT 448.950 666.600 451.050 667.050 ;
        RECT 478.950 666.600 481.050 667.050 ;
        RECT 484.950 666.600 487.050 667.050 ;
        RECT 448.950 665.400 487.050 666.600 ;
        RECT 448.950 664.950 451.050 665.400 ;
        RECT 478.950 664.950 481.050 665.400 ;
        RECT 484.950 664.950 487.050 665.400 ;
        RECT 547.950 666.600 550.050 667.050 ;
        RECT 562.950 666.600 565.050 667.050 ;
        RECT 547.950 665.400 565.050 666.600 ;
        RECT 547.950 664.950 550.050 665.400 ;
        RECT 562.950 664.950 565.050 665.400 ;
        RECT 679.950 666.600 682.050 667.050 ;
        RECT 724.950 666.600 727.050 667.050 ;
        RECT 679.950 665.400 727.050 666.600 ;
        RECT 679.950 664.950 682.050 665.400 ;
        RECT 724.950 664.950 727.050 665.400 ;
        RECT 739.950 666.600 742.050 667.050 ;
        RECT 748.950 666.600 751.050 667.050 ;
        RECT 739.950 665.400 751.050 666.600 ;
        RECT 739.950 664.950 742.050 665.400 ;
        RECT 748.950 664.950 751.050 665.400 ;
        RECT 799.950 666.600 802.050 667.050 ;
        RECT 815.400 666.600 816.600 668.400 ;
        RECT 829.950 667.950 832.050 668.400 ;
        RECT 853.950 669.600 856.050 670.050 ;
        RECT 862.950 669.600 865.050 670.050 ;
        RECT 853.950 668.400 865.050 669.600 ;
        RECT 853.950 667.950 856.050 668.400 ;
        RECT 862.950 667.950 865.050 668.400 ;
        RECT 871.950 669.600 874.050 670.050 ;
        RECT 910.800 669.600 912.900 670.050 ;
        RECT 871.950 668.400 912.900 669.600 ;
        RECT 871.950 667.950 874.050 668.400 ;
        RECT 910.800 667.950 912.900 668.400 ;
        RECT 913.950 669.600 916.050 670.050 ;
        RECT 934.950 669.600 937.050 669.900 ;
        RECT 913.950 668.400 937.050 669.600 ;
        RECT 913.950 667.950 916.050 668.400 ;
        RECT 934.950 667.800 937.050 668.400 ;
        RECT 799.950 665.400 816.600 666.600 ;
        RECT 832.950 666.600 835.050 667.050 ;
        RECT 853.950 666.600 856.050 666.900 ;
        RECT 832.950 665.400 856.050 666.600 ;
        RECT 799.950 664.950 802.050 665.400 ;
        RECT 832.950 664.950 835.050 665.400 ;
        RECT 853.950 664.800 856.050 665.400 ;
        RECT 328.950 662.400 357.600 663.600 ;
        RECT 358.950 663.600 361.050 664.050 ;
        RECT 370.950 663.600 373.050 664.050 ;
        RECT 358.950 662.400 373.050 663.600 ;
        RECT 328.950 661.950 331.050 662.400 ;
        RECT 358.950 661.950 361.050 662.400 ;
        RECT 370.950 661.950 373.050 662.400 ;
        RECT 391.950 663.600 394.050 664.050 ;
        RECT 397.800 663.600 399.900 664.050 ;
        RECT 391.950 662.400 399.900 663.600 ;
        RECT 391.950 661.950 394.050 662.400 ;
        RECT 397.800 661.950 399.900 662.400 ;
        RECT 400.950 663.600 403.050 664.050 ;
        RECT 409.950 663.600 412.050 664.050 ;
        RECT 400.950 662.400 412.050 663.600 ;
        RECT 400.950 661.950 403.050 662.400 ;
        RECT 409.950 661.950 412.050 662.400 ;
        RECT 415.950 663.600 418.050 664.050 ;
        RECT 445.950 663.600 448.050 664.050 ;
        RECT 583.950 663.600 586.050 664.050 ;
        RECT 595.950 663.600 598.050 664.050 ;
        RECT 415.950 662.400 448.050 663.600 ;
        RECT 415.950 661.950 418.050 662.400 ;
        RECT 445.950 661.950 448.050 662.400 ;
        RECT 581.400 662.400 598.050 663.600 ;
        RECT 43.950 660.600 46.050 661.050 ;
        RECT 49.950 660.600 52.050 661.050 ;
        RECT 43.950 659.400 52.050 660.600 ;
        RECT 43.950 658.950 46.050 659.400 ;
        RECT 49.950 658.950 52.050 659.400 ;
        RECT 133.950 660.600 136.050 661.050 ;
        RECT 178.950 660.600 181.050 661.050 ;
        RECT 133.950 659.400 181.050 660.600 ;
        RECT 133.950 658.950 136.050 659.400 ;
        RECT 178.950 658.950 181.050 659.400 ;
        RECT 184.950 660.600 187.050 661.050 ;
        RECT 214.950 660.600 217.050 661.050 ;
        RECT 184.950 659.400 217.050 660.600 ;
        RECT 184.950 658.950 187.050 659.400 ;
        RECT 214.950 658.950 217.050 659.400 ;
        RECT 250.950 660.600 253.050 661.050 ;
        RECT 298.950 660.600 301.050 661.050 ;
        RECT 373.950 660.600 376.050 661.050 ;
        RECT 250.950 659.400 301.050 660.600 ;
        RECT 250.950 658.950 253.050 659.400 ;
        RECT 298.950 658.950 301.050 659.400 ;
        RECT 326.400 659.400 376.050 660.600 ;
        RECT 154.950 657.600 157.050 658.050 ;
        RECT 163.950 657.600 166.050 658.050 ;
        RECT 154.950 656.400 166.050 657.600 ;
        RECT 154.950 655.950 157.050 656.400 ;
        RECT 163.950 655.950 166.050 656.400 ;
        RECT 208.950 657.600 211.050 658.050 ;
        RECT 235.950 657.600 238.050 658.050 ;
        RECT 208.950 656.400 238.050 657.600 ;
        RECT 208.950 655.950 211.050 656.400 ;
        RECT 235.950 655.950 238.050 656.400 ;
        RECT 301.950 657.600 304.050 658.050 ;
        RECT 319.950 657.600 322.050 658.050 ;
        RECT 326.400 657.600 327.600 659.400 ;
        RECT 373.950 658.950 376.050 659.400 ;
        RECT 412.950 660.600 415.050 661.050 ;
        RECT 421.950 660.600 424.050 661.050 ;
        RECT 412.950 659.400 424.050 660.600 ;
        RECT 412.950 658.950 415.050 659.400 ;
        RECT 421.950 658.950 424.050 659.400 ;
        RECT 568.950 660.600 571.050 661.050 ;
        RECT 581.400 660.600 582.600 662.400 ;
        RECT 583.950 661.950 586.050 662.400 ;
        RECT 595.950 661.950 598.050 662.400 ;
        RECT 649.950 663.600 652.050 664.050 ;
        RECT 676.950 663.600 679.050 664.050 ;
        RECT 649.950 662.400 679.050 663.600 ;
        RECT 649.950 661.950 652.050 662.400 ;
        RECT 676.950 661.950 679.050 662.400 ;
        RECT 835.950 663.600 838.050 664.050 ;
        RECT 883.950 663.600 886.050 664.050 ;
        RECT 835.950 662.400 886.050 663.600 ;
        RECT 835.950 661.950 838.050 662.400 ;
        RECT 883.950 661.950 886.050 662.400 ;
        RECT 568.950 659.400 582.600 660.600 ;
        RECT 598.950 660.600 601.050 661.050 ;
        RECT 607.950 660.600 610.050 661.050 ;
        RECT 670.950 660.600 673.050 661.050 ;
        RECT 598.950 659.400 610.050 660.600 ;
        RECT 568.950 658.950 571.050 659.400 ;
        RECT 598.950 658.950 601.050 659.400 ;
        RECT 607.950 658.950 610.050 659.400 ;
        RECT 653.400 659.400 673.050 660.600 ;
        RECT 653.400 658.050 654.600 659.400 ;
        RECT 670.950 658.950 673.050 659.400 ;
        RECT 301.950 656.400 327.600 657.600 ;
        RECT 559.950 657.600 562.050 658.050 ;
        RECT 652.950 657.600 655.050 658.050 ;
        RECT 559.950 656.400 655.050 657.600 ;
        RECT 301.950 655.950 304.050 656.400 ;
        RECT 319.950 655.950 322.050 656.400 ;
        RECT 559.950 655.950 562.050 656.400 ;
        RECT 652.950 655.950 655.050 656.400 ;
        RECT 751.950 657.600 754.050 658.050 ;
        RECT 784.950 657.600 787.050 658.050 ;
        RECT 751.950 656.400 787.050 657.600 ;
        RECT 751.950 655.950 754.050 656.400 ;
        RECT 784.950 655.950 787.050 656.400 ;
        RECT 820.950 657.600 823.050 658.050 ;
        RECT 838.950 657.600 841.050 658.050 ;
        RECT 877.950 657.600 880.050 658.050 ;
        RECT 820.950 656.400 880.050 657.600 ;
        RECT 820.950 655.950 823.050 656.400 ;
        RECT 838.950 655.950 841.050 656.400 ;
        RECT 877.950 655.950 880.050 656.400 ;
        RECT 913.950 657.600 916.050 658.050 ;
        RECT 922.950 657.600 925.050 657.900 ;
        RECT 913.950 656.400 925.050 657.600 ;
        RECT 913.950 655.950 916.050 656.400 ;
        RECT 922.950 655.800 925.050 656.400 ;
        RECT 223.950 654.600 226.050 655.050 ;
        RECT 229.950 654.600 232.050 655.050 ;
        RECT 223.950 653.400 232.050 654.600 ;
        RECT 223.950 652.950 226.050 653.400 ;
        RECT 229.950 652.950 232.050 653.400 ;
        RECT 244.950 654.600 247.050 655.050 ;
        RECT 304.950 654.600 307.050 655.050 ;
        RECT 244.950 653.400 307.050 654.600 ;
        RECT 244.950 652.950 247.050 653.400 ;
        RECT 304.950 652.950 307.050 653.400 ;
        RECT 433.950 654.600 436.050 655.050 ;
        RECT 478.950 654.600 481.050 655.050 ;
        RECT 433.950 653.400 481.050 654.600 ;
        RECT 433.950 652.950 436.050 653.400 ;
        RECT 478.950 652.950 481.050 653.400 ;
        RECT 490.950 654.600 493.050 655.050 ;
        RECT 502.950 654.600 505.050 655.050 ;
        RECT 490.950 653.400 505.050 654.600 ;
        RECT 490.950 652.950 493.050 653.400 ;
        RECT 502.950 652.950 505.050 653.400 ;
        RECT 508.950 654.600 511.050 655.050 ;
        RECT 643.950 654.600 646.050 655.050 ;
        RECT 652.950 654.600 655.050 654.900 ;
        RECT 508.950 653.400 546.600 654.600 ;
        RECT 508.950 652.950 511.050 653.400 ;
        RECT 7.950 651.750 10.050 652.200 ;
        RECT 13.950 651.750 16.050 652.200 ;
        RECT 7.950 650.550 16.050 651.750 ;
        RECT 7.950 650.100 10.050 650.550 ;
        RECT 13.950 650.100 16.050 650.550 ;
        RECT 19.950 651.750 22.050 652.200 ;
        RECT 25.950 651.750 28.050 652.200 ;
        RECT 19.950 650.550 28.050 651.750 ;
        RECT 19.950 650.100 22.050 650.550 ;
        RECT 25.950 650.100 28.050 650.550 ;
        RECT 55.950 651.600 58.050 652.200 ;
        RECT 64.950 651.600 67.050 652.050 ;
        RECT 55.950 650.400 67.050 651.600 ;
        RECT 55.950 650.100 58.050 650.400 ;
        RECT 64.950 649.950 67.050 650.400 ;
        RECT 85.950 650.100 88.050 652.200 ;
        RECT 127.950 651.600 130.050 652.200 ;
        RECT 142.950 651.600 145.050 652.200 ;
        RECT 127.950 650.400 145.050 651.600 ;
        RECT 127.950 650.100 130.050 650.400 ;
        RECT 142.950 650.100 145.050 650.400 ;
        RECT 148.950 651.600 151.050 652.050 ;
        RECT 157.950 651.600 160.050 652.200 ;
        RECT 184.950 651.600 187.050 652.200 ;
        RECT 199.950 651.600 202.050 652.200 ;
        RECT 148.950 650.400 160.050 651.600 ;
        RECT 70.950 645.600 73.050 645.900 ;
        RECT 86.400 645.600 87.600 650.100 ;
        RECT 148.950 649.950 151.050 650.400 ;
        RECT 157.950 650.100 160.050 650.400 ;
        RECT 164.400 650.400 187.050 651.600 ;
        RECT 97.950 645.600 100.050 646.050 ;
        RECT 70.950 644.400 100.050 645.600 ;
        RECT 70.950 643.800 73.050 644.400 ;
        RECT 97.950 643.950 100.050 644.400 ;
        RECT 124.950 645.600 127.050 645.900 ;
        RECT 133.950 645.600 136.050 646.050 ;
        RECT 124.950 644.400 136.050 645.600 ;
        RECT 124.950 643.800 127.050 644.400 ;
        RECT 133.950 643.950 136.050 644.400 ;
        RECT 139.950 645.450 142.050 645.900 ;
        RECT 148.950 645.450 151.050 645.900 ;
        RECT 139.950 644.250 151.050 645.450 ;
        RECT 139.950 643.800 142.050 644.250 ;
        RECT 148.950 643.800 151.050 644.250 ;
        RECT 160.950 645.600 163.050 645.900 ;
        RECT 164.400 645.600 165.600 650.400 ;
        RECT 184.950 650.100 187.050 650.400 ;
        RECT 191.400 650.400 202.050 651.600 ;
        RECT 191.400 648.600 192.600 650.400 ;
        RECT 199.950 650.100 202.050 650.400 ;
        RECT 211.950 651.750 214.050 652.200 ;
        RECT 238.950 651.750 241.050 652.200 ;
        RECT 211.950 650.550 241.050 651.750 ;
        RECT 211.950 650.100 214.050 650.550 ;
        RECT 238.950 650.100 241.050 650.550 ;
        RECT 250.950 649.950 253.050 652.050 ;
        RECT 188.400 647.400 192.600 648.600 ;
        RECT 160.950 644.400 165.600 645.600 ;
        RECT 172.950 645.600 175.050 646.050 ;
        RECT 188.400 645.600 189.600 647.400 ;
        RECT 172.950 644.400 189.600 645.600 ;
        RECT 160.950 643.800 163.050 644.400 ;
        RECT 172.950 643.950 175.050 644.400 ;
        RECT 251.400 643.050 252.600 649.950 ;
        RECT 253.950 645.600 256.050 649.050 ;
        RECT 259.950 648.600 262.050 652.050 ;
        RECT 307.950 651.600 310.050 652.050 ;
        RECT 337.950 651.600 340.050 652.200 ;
        RECT 307.950 650.400 340.050 651.600 ;
        RECT 307.950 649.950 310.050 650.400 ;
        RECT 337.950 650.100 340.050 650.400 ;
        RECT 376.950 649.950 379.050 652.050 ;
        RECT 388.950 651.600 391.050 652.200 ;
        RECT 400.950 651.600 403.050 652.050 ;
        RECT 388.950 650.400 403.050 651.600 ;
        RECT 388.950 650.100 391.050 650.400 ;
        RECT 400.950 649.950 403.050 650.400 ;
        RECT 469.950 651.600 472.050 652.200 ;
        RECT 545.400 652.050 546.600 653.400 ;
        RECT 643.950 653.400 655.050 654.600 ;
        RECT 643.950 652.950 646.050 653.400 ;
        RECT 652.950 652.800 655.050 653.400 ;
        RECT 661.950 654.600 664.050 655.050 ;
        RECT 679.950 654.600 682.050 655.050 ;
        RECT 661.950 653.400 682.050 654.600 ;
        RECT 661.950 652.950 664.050 653.400 ;
        RECT 679.950 652.950 682.050 653.400 ;
        RECT 712.950 654.600 715.050 655.050 ;
        RECT 745.950 654.600 748.050 655.050 ;
        RECT 712.950 653.400 748.050 654.600 ;
        RECT 712.950 652.950 715.050 653.400 ;
        RECT 745.950 652.950 748.050 653.400 ;
        RECT 811.950 654.600 814.050 655.200 ;
        RECT 817.950 654.600 820.050 655.050 ;
        RECT 811.950 653.400 820.050 654.600 ;
        RECT 811.950 653.100 814.050 653.400 ;
        RECT 817.950 652.950 820.050 653.400 ;
        RECT 844.950 654.600 847.050 655.050 ;
        RECT 850.950 654.600 853.050 655.050 ;
        RECT 844.950 653.400 853.050 654.600 ;
        RECT 844.950 652.950 847.050 653.400 ;
        RECT 850.950 652.950 853.050 653.400 ;
        RECT 910.950 654.600 913.050 655.050 ;
        RECT 916.950 654.600 919.050 655.050 ;
        RECT 910.950 653.400 919.050 654.600 ;
        RECT 910.950 652.950 913.050 653.400 ;
        RECT 916.950 652.950 919.050 653.400 ;
        RECT 475.950 651.600 478.050 652.050 ;
        RECT 469.950 650.400 478.050 651.600 ;
        RECT 469.950 650.100 472.050 650.400 ;
        RECT 475.950 649.950 478.050 650.400 ;
        RECT 479.400 650.400 528.600 651.600 ;
        RECT 545.400 650.400 550.050 652.050 ;
        RECT 565.950 651.600 568.050 652.050 ;
        RECT 271.950 648.600 274.050 649.050 ;
        RECT 259.950 648.000 274.050 648.600 ;
        RECT 260.400 647.400 274.050 648.000 ;
        RECT 271.950 646.950 274.050 647.400 ;
        RECT 253.950 645.000 258.600 645.600 ;
        RECT 254.400 644.400 258.600 645.000 ;
        RECT 25.950 642.600 28.050 643.050 ;
        RECT 58.950 642.600 61.050 643.050 ;
        RECT 94.950 642.600 97.050 643.050 ;
        RECT 139.950 642.600 142.050 643.050 ;
        RECT 25.950 641.400 142.050 642.600 ;
        RECT 251.400 641.400 256.050 643.050 ;
        RECT 25.950 640.950 28.050 641.400 ;
        RECT 58.950 640.950 61.050 641.400 ;
        RECT 94.950 640.950 97.050 641.400 ;
        RECT 139.950 640.950 142.050 641.400 ;
        RECT 252.000 640.950 256.050 641.400 ;
        RECT 199.950 639.600 202.050 640.050 ;
        RECT 208.950 639.600 211.050 640.050 ;
        RECT 199.950 638.400 211.050 639.600 ;
        RECT 257.400 639.600 258.600 644.400 ;
        RECT 304.950 645.450 307.050 646.050 ;
        RECT 328.950 645.450 331.050 645.900 ;
        RECT 304.950 644.250 331.050 645.450 ;
        RECT 304.950 643.950 307.050 644.250 ;
        RECT 328.950 643.800 331.050 644.250 ;
        RECT 271.950 642.600 274.050 643.050 ;
        RECT 304.950 642.600 307.050 642.900 ;
        RECT 271.950 641.400 307.050 642.600 ;
        RECT 271.950 640.950 274.050 641.400 ;
        RECT 304.950 640.800 307.050 641.400 ;
        RECT 361.950 642.600 364.050 643.050 ;
        RECT 377.400 642.600 378.600 649.950 ;
        RECT 421.950 648.600 424.050 649.050 ;
        RECT 479.400 648.600 480.600 650.400 ;
        RECT 421.950 647.400 480.600 648.600 ;
        RECT 502.950 648.600 505.050 649.050 ;
        RECT 523.950 648.600 526.050 648.900 ;
        RECT 502.950 647.400 526.050 648.600 ;
        RECT 527.400 648.600 528.600 650.400 ;
        RECT 546.000 649.950 550.050 650.400 ;
        RECT 551.400 650.400 568.050 651.600 ;
        RECT 551.400 648.600 552.600 650.400 ;
        RECT 565.950 649.950 568.050 650.400 ;
        RECT 574.950 651.600 577.050 652.200 ;
        RECT 586.950 651.600 589.050 652.050 ;
        RECT 574.950 650.400 589.050 651.600 ;
        RECT 574.950 650.100 577.050 650.400 ;
        RECT 586.950 649.950 589.050 650.400 ;
        RECT 601.950 651.600 604.050 652.200 ;
        RECT 628.950 651.750 631.050 652.200 ;
        RECT 637.950 651.750 640.050 652.200 ;
        RECT 628.950 651.600 640.050 651.750 ;
        RECT 601.950 650.550 640.050 651.600 ;
        RECT 601.950 650.400 631.050 650.550 ;
        RECT 601.950 650.100 604.050 650.400 ;
        RECT 628.950 650.100 631.050 650.400 ;
        RECT 637.950 650.100 640.050 650.550 ;
        RECT 667.950 649.950 670.050 652.050 ;
        RECT 676.950 651.600 679.050 652.200 ;
        RECT 674.400 650.400 679.050 651.600 ;
        RECT 527.400 647.400 552.600 648.600 ;
        RECT 641.400 647.400 651.600 648.600 ;
        RECT 421.950 646.950 424.050 647.400 ;
        RECT 502.950 646.950 505.050 647.400 ;
        RECT 523.950 646.800 526.050 647.400 ;
        RECT 641.400 645.900 642.600 647.400 ;
        RECT 650.400 645.900 651.600 647.400 ;
        RECT 400.950 645.450 403.050 645.900 ;
        RECT 406.950 645.450 409.050 645.900 ;
        RECT 400.950 644.250 409.050 645.450 ;
        RECT 400.950 643.800 403.050 644.250 ;
        RECT 406.950 643.800 409.050 644.250 ;
        RECT 481.950 645.450 484.050 645.900 ;
        RECT 493.950 645.450 496.050 645.900 ;
        RECT 481.950 644.250 496.050 645.450 ;
        RECT 481.950 643.800 484.050 644.250 ;
        RECT 493.950 643.800 496.050 644.250 ;
        RECT 592.950 645.450 595.050 645.900 ;
        RECT 607.950 645.450 610.050 645.900 ;
        RECT 592.950 644.250 610.050 645.450 ;
        RECT 592.950 643.800 595.050 644.250 ;
        RECT 607.950 643.800 610.050 644.250 ;
        RECT 640.950 643.800 643.050 645.900 ;
        RECT 649.950 645.450 652.050 645.900 ;
        RECT 664.950 645.450 667.050 645.900 ;
        RECT 649.950 644.250 667.050 645.450 ;
        RECT 649.950 643.800 652.050 644.250 ;
        RECT 664.950 643.800 667.050 644.250 ;
        RECT 361.950 641.400 378.600 642.600 ;
        RECT 379.950 642.600 382.050 643.050 ;
        RECT 385.950 642.600 388.050 643.050 ;
        RECT 397.950 642.600 400.050 643.050 ;
        RECT 379.950 641.400 400.050 642.600 ;
        RECT 361.950 640.950 364.050 641.400 ;
        RECT 379.950 640.950 382.050 641.400 ;
        RECT 385.950 640.950 388.050 641.400 ;
        RECT 397.950 640.950 400.050 641.400 ;
        RECT 424.950 642.600 427.050 643.050 ;
        RECT 451.950 642.600 454.050 643.050 ;
        RECT 424.950 641.400 454.050 642.600 ;
        RECT 424.950 640.950 427.050 641.400 ;
        RECT 451.950 640.950 454.050 641.400 ;
        RECT 469.950 642.450 472.050 642.900 ;
        RECT 499.950 642.600 502.050 642.900 ;
        RECT 523.950 642.600 526.050 643.050 ;
        RECT 499.950 642.450 526.050 642.600 ;
        RECT 469.950 641.400 526.050 642.450 ;
        RECT 469.950 641.250 502.050 641.400 ;
        RECT 469.950 640.800 472.050 641.250 ;
        RECT 499.950 640.800 502.050 641.250 ;
        RECT 523.950 640.950 526.050 641.400 ;
        RECT 643.950 642.600 646.050 643.050 ;
        RECT 652.950 642.600 655.050 643.050 ;
        RECT 643.950 641.400 655.050 642.600 ;
        RECT 643.950 640.950 646.050 641.400 ;
        RECT 652.950 640.950 655.050 641.400 ;
        RECT 661.950 642.600 664.050 643.050 ;
        RECT 668.400 642.600 669.600 649.950 ;
        RECT 674.400 646.050 675.600 650.400 ;
        RECT 676.950 650.100 679.050 650.400 ;
        RECT 682.950 651.600 685.050 652.200 ;
        RECT 700.950 651.600 703.050 652.200 ;
        RECT 682.950 650.400 703.050 651.600 ;
        RECT 682.950 650.100 685.050 650.400 ;
        RECT 700.950 650.100 703.050 650.400 ;
        RECT 706.950 651.600 709.050 652.200 ;
        RECT 715.950 651.600 718.050 652.050 ;
        RECT 721.950 651.600 724.050 652.200 ;
        RECT 706.950 650.400 718.050 651.600 ;
        RECT 706.950 650.100 709.050 650.400 ;
        RECT 715.950 649.950 718.050 650.400 ;
        RECT 719.400 650.400 724.050 651.600 ;
        RECT 719.400 648.600 720.600 650.400 ;
        RECT 721.950 650.100 724.050 650.400 ;
        RECT 763.950 651.750 766.050 652.200 ;
        RECT 769.950 651.750 772.050 652.200 ;
        RECT 763.950 650.550 772.050 651.750 ;
        RECT 763.950 650.100 766.050 650.550 ;
        RECT 769.950 650.100 772.050 650.550 ;
        RECT 775.950 651.600 778.050 652.200 ;
        RECT 793.950 651.600 796.050 652.200 ;
        RECT 775.950 650.400 796.050 651.600 ;
        RECT 775.950 650.100 778.050 650.400 ;
        RECT 793.950 650.100 796.050 650.400 ;
        RECT 739.950 648.600 742.050 648.900 ;
        RECT 776.400 648.600 777.600 650.100 ;
        RECT 811.950 649.950 814.050 652.050 ;
        RECT 841.950 651.750 844.050 652.200 ;
        RECT 847.950 651.750 850.050 652.200 ;
        RECT 841.950 650.550 850.050 651.750 ;
        RECT 841.950 650.100 844.050 650.550 ;
        RECT 847.950 650.100 850.050 650.550 ;
        RECT 862.950 651.600 865.050 652.050 ;
        RECT 874.950 651.600 877.050 652.200 ;
        RECT 862.950 650.400 877.050 651.600 ;
        RECT 862.950 649.950 865.050 650.400 ;
        RECT 874.950 650.100 877.050 650.400 ;
        RECT 880.950 649.950 883.050 652.050 ;
        RECT 892.950 651.600 895.050 652.050 ;
        RECT 907.950 651.600 910.050 652.200 ;
        RECT 892.950 650.400 910.050 651.600 ;
        RECT 892.950 649.950 895.050 650.400 ;
        RECT 698.400 647.400 742.050 648.600 ;
        RECT 767.400 648.000 777.600 648.600 ;
        RECT 673.950 643.950 676.050 646.050 ;
        RECT 698.400 645.900 699.600 647.400 ;
        RECT 739.950 646.800 742.050 647.400 ;
        RECT 766.950 647.400 777.600 648.000 ;
        RECT 812.400 648.600 813.600 649.950 ;
        RECT 826.950 648.600 829.050 649.050 ;
        RECT 812.400 647.400 829.050 648.600 ;
        RECT 685.950 645.600 688.050 645.900 ;
        RECT 697.950 645.600 700.050 645.900 ;
        RECT 685.950 644.400 700.050 645.600 ;
        RECT 685.950 643.800 688.050 644.400 ;
        RECT 697.950 643.800 700.050 644.400 ;
        RECT 724.950 645.450 727.050 645.900 ;
        RECT 736.950 645.450 739.050 645.900 ;
        RECT 724.950 644.250 739.050 645.450 ;
        RECT 724.950 643.800 727.050 644.250 ;
        RECT 736.950 643.800 739.050 644.250 ;
        RECT 748.950 645.450 751.050 645.900 ;
        RECT 760.950 645.450 763.050 645.900 ;
        RECT 748.950 644.250 763.050 645.450 ;
        RECT 748.950 643.800 751.050 644.250 ;
        RECT 760.950 643.800 763.050 644.250 ;
        RECT 766.950 643.950 769.050 647.400 ;
        RECT 826.950 646.950 829.050 647.400 ;
        RECT 881.400 646.050 882.600 649.950 ;
        RECT 896.400 646.050 897.600 650.400 ;
        RECT 907.950 650.100 910.050 650.400 ;
        RECT 820.950 645.600 823.050 645.900 ;
        RECT 835.950 645.600 838.050 645.900 ;
        RECT 820.950 645.450 838.050 645.600 ;
        RECT 862.950 645.450 865.050 645.900 ;
        RECT 820.950 644.400 865.050 645.450 ;
        RECT 820.950 643.800 823.050 644.400 ;
        RECT 835.950 644.250 865.050 644.400 ;
        RECT 835.950 643.800 838.050 644.250 ;
        RECT 862.950 643.800 865.050 644.250 ;
        RECT 880.950 643.950 883.050 646.050 ;
        RECT 895.950 643.950 898.050 646.050 ;
        RECT 917.400 645.900 918.600 652.950 ;
        RECT 919.950 651.600 922.050 652.050 ;
        RECT 928.950 651.600 931.050 651.900 ;
        RECT 919.950 650.400 931.050 651.600 ;
        RECT 919.950 649.950 922.050 650.400 ;
        RECT 928.950 649.800 931.050 650.400 ;
        RECT 916.950 643.800 919.050 645.900 ;
        RECT 661.950 641.400 669.600 642.600 ;
        RECT 754.950 642.600 757.050 643.050 ;
        RECT 805.950 642.600 808.050 643.050 ;
        RECT 817.950 642.600 820.050 643.050 ;
        RECT 754.950 641.400 820.050 642.600 ;
        RECT 661.950 640.950 664.050 641.400 ;
        RECT 754.950 640.950 757.050 641.400 ;
        RECT 805.950 640.950 808.050 641.400 ;
        RECT 817.950 640.950 820.050 641.400 ;
        RECT 310.950 639.600 313.050 640.050 ;
        RECT 257.400 638.400 313.050 639.600 ;
        RECT 199.950 637.950 202.050 638.400 ;
        RECT 208.950 637.950 211.050 638.400 ;
        RECT 310.950 637.950 313.050 638.400 ;
        RECT 391.950 639.600 394.050 640.050 ;
        RECT 412.950 639.600 415.050 640.050 ;
        RECT 391.950 638.400 415.050 639.600 ;
        RECT 391.950 637.950 394.050 638.400 ;
        RECT 412.950 637.950 415.050 638.400 ;
        RECT 577.950 639.600 580.050 640.050 ;
        RECT 598.950 639.600 601.050 640.050 ;
        RECT 577.950 638.400 601.050 639.600 ;
        RECT 577.950 637.950 580.050 638.400 ;
        RECT 598.950 637.950 601.050 638.400 ;
        RECT 631.950 639.600 634.050 640.050 ;
        RECT 682.950 639.600 685.050 640.050 ;
        RECT 631.950 638.400 685.050 639.600 ;
        RECT 631.950 637.950 634.050 638.400 ;
        RECT 682.950 637.950 685.050 638.400 ;
        RECT 697.950 639.600 700.050 640.050 ;
        RECT 733.950 639.600 736.050 640.050 ;
        RECT 697.950 638.400 736.050 639.600 ;
        RECT 697.950 637.950 700.050 638.400 ;
        RECT 733.950 637.950 736.050 638.400 ;
        RECT 796.950 639.600 799.050 640.050 ;
        RECT 805.950 639.600 808.050 639.900 ;
        RECT 796.950 638.400 808.050 639.600 ;
        RECT 796.950 637.950 799.050 638.400 ;
        RECT 805.950 637.800 808.050 638.400 ;
        RECT 883.950 639.600 886.050 640.050 ;
        RECT 892.950 639.600 895.050 640.050 ;
        RECT 883.950 638.400 895.050 639.600 ;
        RECT 883.950 637.950 886.050 638.400 ;
        RECT 892.950 637.950 895.050 638.400 ;
        RECT 52.950 636.600 55.050 637.050 ;
        RECT 58.950 636.600 61.050 637.050 ;
        RECT 52.950 635.400 61.050 636.600 ;
        RECT 52.950 634.950 55.050 635.400 ;
        RECT 58.950 634.950 61.050 635.400 ;
        RECT 112.950 636.600 115.050 637.050 ;
        RECT 139.950 636.600 142.050 637.050 ;
        RECT 112.950 635.400 142.050 636.600 ;
        RECT 112.950 634.950 115.050 635.400 ;
        RECT 139.950 634.950 142.050 635.400 ;
        RECT 235.950 636.600 238.050 637.050 ;
        RECT 250.950 636.600 253.050 637.050 ;
        RECT 235.950 635.400 253.050 636.600 ;
        RECT 235.950 634.950 238.050 635.400 ;
        RECT 250.950 634.950 253.050 635.400 ;
        RECT 418.950 636.600 421.050 637.050 ;
        RECT 439.950 636.600 442.050 637.050 ;
        RECT 418.950 635.400 442.050 636.600 ;
        RECT 418.950 634.950 421.050 635.400 ;
        RECT 439.950 634.950 442.050 635.400 ;
        RECT 448.950 636.600 451.050 637.050 ;
        RECT 457.950 636.600 460.050 637.050 ;
        RECT 448.950 635.400 460.050 636.600 ;
        RECT 448.950 634.950 451.050 635.400 ;
        RECT 457.950 634.950 460.050 635.400 ;
        RECT 496.950 636.600 499.050 637.050 ;
        RECT 622.950 636.600 625.050 637.050 ;
        RECT 688.950 636.600 691.050 637.050 ;
        RECT 790.950 636.600 793.050 637.050 ;
        RECT 808.950 636.600 811.050 637.050 ;
        RECT 496.950 635.400 811.050 636.600 ;
        RECT 496.950 634.950 499.050 635.400 ;
        RECT 622.950 634.950 625.050 635.400 ;
        RECT 688.950 634.950 691.050 635.400 ;
        RECT 790.950 634.950 793.050 635.400 ;
        RECT 808.950 634.950 811.050 635.400 ;
        RECT 865.950 636.600 868.050 637.050 ;
        RECT 884.400 636.600 885.600 637.950 ;
        RECT 865.950 635.400 885.600 636.600 ;
        RECT 913.950 636.600 916.050 637.050 ;
        RECT 919.950 636.600 922.050 637.050 ;
        RECT 913.950 635.400 922.050 636.600 ;
        RECT 865.950 634.950 868.050 635.400 ;
        RECT 913.950 634.950 916.050 635.400 ;
        RECT 919.950 634.950 922.050 635.400 ;
        RECT 196.950 633.600 199.050 634.050 ;
        RECT 298.950 633.600 301.050 634.050 ;
        RECT 196.950 632.400 301.050 633.600 ;
        RECT 196.950 631.950 199.050 632.400 ;
        RECT 298.950 631.950 301.050 632.400 ;
        RECT 307.950 633.600 310.050 634.050 ;
        RECT 313.950 633.600 316.050 634.050 ;
        RECT 307.950 632.400 316.050 633.600 ;
        RECT 307.950 631.950 310.050 632.400 ;
        RECT 313.950 631.950 316.050 632.400 ;
        RECT 328.950 633.600 331.050 634.050 ;
        RECT 352.950 633.600 355.050 634.050 ;
        RECT 328.950 632.400 355.050 633.600 ;
        RECT 328.950 631.950 331.050 632.400 ;
        RECT 352.950 631.950 355.050 632.400 ;
        RECT 373.950 633.600 376.050 634.050 ;
        RECT 391.950 633.600 394.050 634.050 ;
        RECT 373.950 632.400 394.050 633.600 ;
        RECT 373.950 631.950 376.050 632.400 ;
        RECT 391.950 631.950 394.050 632.400 ;
        RECT 397.950 633.600 400.050 634.050 ;
        RECT 442.950 633.600 445.050 634.050 ;
        RECT 460.950 633.600 463.050 634.050 ;
        RECT 397.950 632.400 463.050 633.600 ;
        RECT 397.950 631.950 400.050 632.400 ;
        RECT 442.950 631.950 445.050 632.400 ;
        RECT 460.950 631.950 463.050 632.400 ;
        RECT 466.950 633.600 469.050 634.050 ;
        RECT 487.950 633.600 490.050 634.050 ;
        RECT 466.950 632.400 490.050 633.600 ;
        RECT 466.950 631.950 469.050 632.400 ;
        RECT 487.950 631.950 490.050 632.400 ;
        RECT 544.950 633.600 547.050 634.050 ;
        RECT 619.950 633.600 622.050 634.050 ;
        RECT 667.950 633.600 670.050 634.050 ;
        RECT 544.950 632.400 670.050 633.600 ;
        RECT 544.950 631.950 547.050 632.400 ;
        RECT 619.950 631.950 622.050 632.400 ;
        RECT 667.950 631.950 670.050 632.400 ;
        RECT 730.950 633.600 733.050 634.050 ;
        RECT 781.950 633.600 784.050 634.050 ;
        RECT 799.950 633.600 802.050 634.050 ;
        RECT 730.950 632.400 802.050 633.600 ;
        RECT 730.950 631.950 733.050 632.400 ;
        RECT 781.950 631.950 784.050 632.400 ;
        RECT 799.950 631.950 802.050 632.400 ;
        RECT 814.950 633.600 817.050 634.050 ;
        RECT 826.950 633.600 829.050 634.050 ;
        RECT 841.950 633.600 844.050 634.050 ;
        RECT 877.950 633.600 880.050 634.050 ;
        RECT 889.950 633.600 892.050 634.050 ;
        RECT 898.950 633.600 901.050 634.050 ;
        RECT 814.950 632.400 855.600 633.600 ;
        RECT 814.950 631.950 817.050 632.400 ;
        RECT 826.950 631.950 829.050 632.400 ;
        RECT 841.950 631.950 844.050 632.400 ;
        RECT 34.950 630.600 37.050 631.050 ;
        RECT 181.950 630.600 184.050 631.050 ;
        RECT 34.950 629.400 184.050 630.600 ;
        RECT 34.950 628.950 37.050 629.400 ;
        RECT 181.950 628.950 184.050 629.400 ;
        RECT 364.950 630.600 367.050 631.050 ;
        RECT 394.950 630.600 397.050 631.050 ;
        RECT 364.950 629.400 397.050 630.600 ;
        RECT 364.950 628.950 367.050 629.400 ;
        RECT 394.950 628.950 397.050 629.400 ;
        RECT 409.950 630.600 412.050 631.050 ;
        RECT 472.950 630.600 475.050 631.050 ;
        RECT 496.950 630.600 499.050 631.050 ;
        RECT 409.950 629.400 499.050 630.600 ;
        RECT 409.950 628.950 412.050 629.400 ;
        RECT 472.950 628.950 475.050 629.400 ;
        RECT 496.950 628.950 499.050 629.400 ;
        RECT 562.950 630.600 565.050 631.050 ;
        RECT 577.950 630.600 580.050 631.050 ;
        RECT 562.950 629.400 580.050 630.600 ;
        RECT 562.950 628.950 565.050 629.400 ;
        RECT 577.950 628.950 580.050 629.400 ;
        RECT 610.950 630.600 613.050 631.050 ;
        RECT 625.950 630.600 628.050 631.050 ;
        RECT 610.950 629.400 628.050 630.600 ;
        RECT 610.950 628.950 613.050 629.400 ;
        RECT 625.950 628.950 628.050 629.400 ;
        RECT 811.950 630.600 814.050 631.050 ;
        RECT 850.950 630.600 853.050 631.050 ;
        RECT 811.950 629.400 853.050 630.600 ;
        RECT 854.400 630.600 855.600 632.400 ;
        RECT 877.950 632.400 901.050 633.600 ;
        RECT 877.950 631.950 880.050 632.400 ;
        RECT 889.950 631.950 892.050 632.400 ;
        RECT 898.950 631.950 901.050 632.400 ;
        RECT 854.400 629.400 873.600 630.600 ;
        RECT 811.950 628.950 814.050 629.400 ;
        RECT 850.950 628.950 853.050 629.400 ;
        RECT 175.950 627.600 178.050 628.050 ;
        RECT 217.950 627.600 220.050 628.050 ;
        RECT 175.950 626.400 220.050 627.600 ;
        RECT 175.950 625.950 178.050 626.400 ;
        RECT 217.950 625.950 220.050 626.400 ;
        RECT 223.950 627.600 226.050 628.050 ;
        RECT 340.950 627.600 343.050 628.050 ;
        RECT 223.950 626.400 343.050 627.600 ;
        RECT 223.950 625.950 226.050 626.400 ;
        RECT 340.950 625.950 343.050 626.400 ;
        RECT 538.950 627.600 541.050 628.050 ;
        RECT 553.950 627.600 556.050 628.050 ;
        RECT 538.950 626.400 556.050 627.600 ;
        RECT 538.950 625.950 541.050 626.400 ;
        RECT 553.950 625.950 556.050 626.400 ;
        RECT 628.950 627.600 631.050 628.050 ;
        RECT 640.950 627.600 643.050 628.050 ;
        RECT 628.950 626.400 643.050 627.600 ;
        RECT 628.950 625.950 631.050 626.400 ;
        RECT 640.950 625.950 643.050 626.400 ;
        RECT 649.950 627.600 652.050 628.050 ;
        RECT 697.950 627.600 700.050 628.050 ;
        RECT 649.950 626.400 700.050 627.600 ;
        RECT 649.950 625.950 652.050 626.400 ;
        RECT 697.950 625.950 700.050 626.400 ;
        RECT 772.950 627.600 775.050 628.050 ;
        RECT 812.400 627.600 813.600 628.950 ;
        RECT 772.950 626.400 813.600 627.600 ;
        RECT 872.400 627.600 873.600 629.400 ;
        RECT 895.950 627.600 898.050 628.050 ;
        RECT 872.400 626.400 898.050 627.600 ;
        RECT 772.950 625.950 775.050 626.400 ;
        RECT 895.950 625.950 898.050 626.400 ;
        RECT 919.950 627.600 922.050 628.050 ;
        RECT 928.950 627.600 931.050 628.050 ;
        RECT 919.950 626.400 931.050 627.600 ;
        RECT 919.950 625.950 922.050 626.400 ;
        RECT 928.950 625.950 931.050 626.400 ;
        RECT 64.950 624.600 67.050 625.050 ;
        RECT 124.950 624.600 127.050 625.050 ;
        RECT 64.950 623.400 127.050 624.600 ;
        RECT 64.950 622.950 67.050 623.400 ;
        RECT 124.950 622.950 127.050 623.400 ;
        RECT 403.950 624.600 406.050 625.050 ;
        RECT 463.950 624.600 466.050 625.050 ;
        RECT 403.950 623.400 466.050 624.600 ;
        RECT 403.950 622.950 406.050 623.400 ;
        RECT 463.950 622.950 466.050 623.400 ;
        RECT 508.950 624.600 511.050 625.050 ;
        RECT 514.950 624.600 517.050 625.050 ;
        RECT 508.950 623.400 517.050 624.600 ;
        RECT 508.950 622.950 511.050 623.400 ;
        RECT 514.950 622.950 517.050 623.400 ;
        RECT 523.950 624.600 526.050 625.050 ;
        RECT 574.950 624.600 577.050 625.050 ;
        RECT 523.950 623.400 577.050 624.600 ;
        RECT 523.950 622.950 526.050 623.400 ;
        RECT 574.950 622.950 577.050 623.400 ;
        RECT 898.950 624.600 901.050 625.050 ;
        RECT 922.950 624.600 925.050 625.050 ;
        RECT 898.950 623.400 925.050 624.600 ;
        RECT 898.950 622.950 901.050 623.400 ;
        RECT 922.950 622.950 925.050 623.400 ;
        RECT 106.950 621.600 109.050 622.050 ;
        RECT 142.950 621.600 145.050 622.050 ;
        RECT 106.950 620.400 145.050 621.600 ;
        RECT 106.950 619.950 109.050 620.400 ;
        RECT 142.950 619.950 145.050 620.400 ;
        RECT 241.950 621.600 244.050 622.050 ;
        RECT 367.950 621.600 370.050 622.050 ;
        RECT 421.950 621.600 424.050 622.050 ;
        RECT 700.950 621.600 703.050 622.050 ;
        RECT 241.950 620.400 370.050 621.600 ;
        RECT 241.950 619.950 244.050 620.400 ;
        RECT 367.950 619.950 370.050 620.400 ;
        RECT 371.400 620.400 424.050 621.600 ;
        RECT 37.950 618.600 40.050 619.050 ;
        RECT 55.950 618.600 58.050 619.050 ;
        RECT 37.950 617.400 58.050 618.600 ;
        RECT 37.950 616.950 40.050 617.400 ;
        RECT 55.950 616.950 58.050 617.400 ;
        RECT 88.950 618.600 91.050 619.050 ;
        RECT 178.950 618.600 181.050 619.050 ;
        RECT 202.950 618.600 205.050 619.050 ;
        RECT 88.950 617.400 205.050 618.600 ;
        RECT 88.950 616.950 91.050 617.400 ;
        RECT 178.950 616.950 181.050 617.400 ;
        RECT 202.950 616.950 205.050 617.400 ;
        RECT 226.950 618.600 229.050 619.050 ;
        RECT 280.950 618.600 283.050 619.050 ;
        RECT 226.950 617.400 283.050 618.600 ;
        RECT 226.950 616.950 229.050 617.400 ;
        RECT 280.950 616.950 283.050 617.400 ;
        RECT 298.950 618.600 301.050 619.050 ;
        RECT 371.400 618.600 372.600 620.400 ;
        RECT 421.950 619.950 424.050 620.400 ;
        RECT 527.400 620.400 703.050 621.600 ;
        RECT 298.950 617.400 372.600 618.600 ;
        RECT 463.950 618.600 466.050 619.050 ;
        RECT 527.400 618.600 528.600 620.400 ;
        RECT 700.950 619.950 703.050 620.400 ;
        RECT 715.950 621.600 718.050 622.050 ;
        RECT 724.950 621.600 727.050 622.050 ;
        RECT 715.950 620.400 727.050 621.600 ;
        RECT 715.950 619.950 718.050 620.400 ;
        RECT 724.950 619.950 727.050 620.400 ;
        RECT 763.950 621.600 766.050 622.050 ;
        RECT 781.950 621.600 784.050 622.050 ;
        RECT 763.950 620.400 784.050 621.600 ;
        RECT 763.950 619.950 766.050 620.400 ;
        RECT 781.950 619.950 784.050 620.400 ;
        RECT 892.950 621.600 895.050 622.050 ;
        RECT 916.950 621.600 919.050 622.050 ;
        RECT 892.950 620.400 919.050 621.600 ;
        RECT 892.950 619.950 895.050 620.400 ;
        RECT 916.950 619.950 919.050 620.400 ;
        RECT 463.950 617.400 528.600 618.600 ;
        RECT 571.950 618.600 574.050 619.050 ;
        RECT 649.950 618.600 652.050 619.050 ;
        RECT 571.950 617.400 652.050 618.600 ;
        RECT 298.950 616.950 301.050 617.400 ;
        RECT 463.950 616.950 466.050 617.400 ;
        RECT 571.950 616.950 574.050 617.400 ;
        RECT 649.950 616.950 652.050 617.400 ;
        RECT 874.950 618.600 877.050 619.050 ;
        RECT 874.950 617.400 882.600 618.600 ;
        RECT 874.950 616.950 877.050 617.400 ;
        RECT 106.950 615.600 109.050 616.050 ;
        RECT 163.950 615.600 166.050 616.050 ;
        RECT 172.950 615.600 175.050 616.050 ;
        RECT 106.950 614.400 175.050 615.600 ;
        RECT 106.950 613.950 109.050 614.400 ;
        RECT 163.950 613.950 166.050 614.400 ;
        RECT 172.950 613.950 175.050 614.400 ;
        RECT 295.950 615.600 298.050 616.050 ;
        RECT 325.950 615.600 328.050 616.050 ;
        RECT 295.950 614.400 328.050 615.600 ;
        RECT 295.950 613.950 298.050 614.400 ;
        RECT 325.950 613.950 328.050 614.400 ;
        RECT 412.950 615.600 415.050 616.050 ;
        RECT 433.950 615.600 436.050 616.050 ;
        RECT 412.950 614.400 436.050 615.600 ;
        RECT 412.950 613.950 415.050 614.400 ;
        RECT 433.950 613.950 436.050 614.400 ;
        RECT 535.950 615.600 538.050 616.050 ;
        RECT 565.950 615.600 568.050 616.050 ;
        RECT 535.950 614.400 568.050 615.600 ;
        RECT 535.950 613.950 538.050 614.400 ;
        RECT 565.950 613.950 568.050 614.400 ;
        RECT 577.950 615.600 580.050 616.050 ;
        RECT 628.950 615.600 631.050 616.050 ;
        RECT 577.950 614.400 631.050 615.600 ;
        RECT 577.950 613.950 580.050 614.400 ;
        RECT 628.950 613.950 631.050 614.400 ;
        RECT 715.950 615.600 718.050 616.050 ;
        RECT 757.950 615.600 760.050 616.050 ;
        RECT 715.950 614.400 760.050 615.600 ;
        RECT 715.950 613.950 718.050 614.400 ;
        RECT 757.950 613.950 760.050 614.400 ;
        RECT 817.950 615.600 820.050 616.050 ;
        RECT 841.950 615.600 844.050 616.050 ;
        RECT 817.950 614.400 844.050 615.600 ;
        RECT 817.950 613.950 820.050 614.400 ;
        RECT 841.950 613.950 844.050 614.400 ;
        RECT 850.950 615.600 853.050 616.050 ;
        RECT 871.950 615.600 874.050 616.050 ;
        RECT 850.950 614.400 874.050 615.600 ;
        RECT 881.400 615.600 882.600 617.400 ;
        RECT 916.950 615.600 919.050 616.050 ;
        RECT 881.400 614.400 919.050 615.600 ;
        RECT 850.950 613.950 853.050 614.400 ;
        RECT 871.950 613.950 874.050 614.400 ;
        RECT 916.950 613.950 919.050 614.400 ;
        RECT 928.950 613.950 934.050 616.050 ;
        RECT 7.950 612.600 10.050 613.050 ;
        RECT 28.950 612.600 31.050 613.050 ;
        RECT 7.950 611.400 31.050 612.600 ;
        RECT 7.950 610.950 10.050 611.400 ;
        RECT 28.950 610.950 31.050 611.400 ;
        RECT 115.950 612.600 118.050 612.900 ;
        RECT 145.950 612.600 148.050 613.050 ;
        RECT 187.950 612.600 190.050 613.050 ;
        RECT 115.950 611.400 190.050 612.600 ;
        RECT 115.950 610.800 118.050 611.400 ;
        RECT 145.950 610.950 148.050 611.400 ;
        RECT 187.950 610.950 190.050 611.400 ;
        RECT 205.950 612.600 208.050 613.050 ;
        RECT 214.950 612.600 217.050 613.050 ;
        RECT 205.950 611.400 217.050 612.600 ;
        RECT 205.950 610.950 208.050 611.400 ;
        RECT 214.950 610.950 217.050 611.400 ;
        RECT 220.950 612.600 223.050 613.050 ;
        RECT 229.950 612.600 232.050 613.050 ;
        RECT 220.950 611.400 232.050 612.600 ;
        RECT 220.950 610.950 223.050 611.400 ;
        RECT 229.950 610.950 232.050 611.400 ;
        RECT 244.950 612.600 247.050 613.050 ;
        RECT 271.950 612.600 274.050 613.050 ;
        RECT 316.950 612.600 319.050 613.050 ;
        RECT 244.950 611.400 274.050 612.600 ;
        RECT 244.950 610.950 247.050 611.400 ;
        RECT 271.950 610.950 274.050 611.400 ;
        RECT 308.400 611.400 319.050 612.600 ;
        RECT 31.950 609.600 34.050 610.050 ;
        RECT 40.950 609.600 43.050 610.050 ;
        RECT 31.950 608.400 43.050 609.600 ;
        RECT 31.950 607.950 34.050 608.400 ;
        RECT 40.950 607.950 43.050 608.400 ;
        RECT 22.950 606.750 25.050 607.200 ;
        RECT 28.950 606.750 31.050 607.200 ;
        RECT 22.950 605.550 31.050 606.750 ;
        RECT 22.950 605.100 25.050 605.550 ;
        RECT 28.950 605.100 31.050 605.550 ;
        RECT 46.950 606.750 49.050 607.200 ;
        RECT 52.950 606.750 55.050 607.200 ;
        RECT 46.950 605.550 55.050 606.750 ;
        RECT 46.950 605.100 49.050 605.550 ;
        RECT 52.950 605.100 55.050 605.550 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 64.950 606.600 67.050 607.200 ;
        RECT 85.950 606.600 88.050 607.200 ;
        RECT 64.950 605.400 88.050 606.600 ;
        RECT 64.950 605.100 67.050 605.400 ;
        RECT 85.950 605.100 88.050 605.400 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 169.950 605.100 172.050 607.200 ;
        RECT 184.950 606.600 187.050 610.050 ;
        RECT 274.950 609.600 277.050 610.050 ;
        RECT 283.950 609.600 286.050 610.050 ;
        RECT 274.950 608.400 286.050 609.600 ;
        RECT 274.950 607.950 277.050 608.400 ;
        RECT 283.950 607.950 286.050 608.400 ;
        RECT 292.950 609.600 295.050 610.050 ;
        RECT 308.400 609.600 309.600 611.400 ;
        RECT 316.950 610.950 319.050 611.400 ;
        RECT 397.950 612.600 400.050 613.050 ;
        RECT 409.950 612.600 412.050 613.050 ;
        RECT 417.000 612.600 421.050 613.050 ;
        RECT 397.950 611.400 412.050 612.600 ;
        RECT 397.950 610.950 400.050 611.400 ;
        RECT 409.950 610.950 412.050 611.400 ;
        RECT 416.400 610.950 421.050 612.600 ;
        RECT 427.950 612.600 430.050 613.050 ;
        RECT 457.950 612.600 460.050 613.050 ;
        RECT 427.950 611.400 460.050 612.600 ;
        RECT 427.950 610.950 430.050 611.400 ;
        RECT 457.950 610.950 460.050 611.400 ;
        RECT 568.950 612.600 571.050 613.050 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 568.950 611.400 598.050 612.600 ;
        RECT 568.950 610.950 571.050 611.400 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 670.950 612.600 673.050 613.050 ;
        RECT 679.950 612.600 682.050 613.050 ;
        RECT 670.950 611.400 682.050 612.600 ;
        RECT 670.950 610.950 673.050 611.400 ;
        RECT 679.950 610.950 682.050 611.400 ;
        RECT 697.950 612.600 700.050 613.050 ;
        RECT 712.950 612.600 715.050 613.050 ;
        RECT 859.950 612.600 862.050 613.050 ;
        RECT 697.950 611.400 715.050 612.600 ;
        RECT 697.950 610.950 700.050 611.400 ;
        RECT 712.950 610.950 715.050 611.400 ;
        RECT 806.400 611.400 862.050 612.600 ;
        RECT 292.950 608.400 309.600 609.600 ;
        RECT 292.950 607.950 295.050 608.400 ;
        RECT 193.950 606.600 196.050 607.200 ;
        RECT 184.950 606.000 196.050 606.600 ;
        RECT 185.400 605.400 196.050 606.000 ;
        RECT 193.950 605.100 196.050 605.400 ;
        RECT 199.950 606.600 202.050 607.200 ;
        RECT 211.950 606.600 214.050 607.200 ;
        RECT 226.950 606.600 229.050 607.200 ;
        RECT 244.950 606.600 247.050 607.200 ;
        RECT 199.950 605.400 214.050 606.600 ;
        RECT 199.950 605.100 202.050 605.400 ;
        RECT 211.950 605.100 214.050 605.400 ;
        RECT 215.400 605.400 247.050 606.600 ;
        RECT 19.950 600.600 22.050 601.050 ;
        RECT 28.950 600.600 31.050 601.050 ;
        RECT 19.950 599.400 31.050 600.600 ;
        RECT 59.400 600.600 60.600 604.950 ;
        RECT 93.000 603.600 97.050 604.050 ;
        RECT 92.400 603.000 97.050 603.600 ;
        RECT 91.950 601.950 97.050 603.000 ;
        RECT 61.950 600.600 64.050 600.900 ;
        RECT 59.400 599.400 64.050 600.600 ;
        RECT 19.950 598.950 22.050 599.400 ;
        RECT 28.950 598.950 31.050 599.400 ;
        RECT 61.950 598.800 64.050 599.400 ;
        RECT 91.950 598.950 94.050 601.950 ;
        RECT 143.400 601.050 144.600 604.950 ;
        RECT 170.400 603.600 171.600 605.100 ;
        RECT 215.400 603.600 216.600 605.400 ;
        RECT 226.950 605.100 229.050 605.400 ;
        RECT 244.950 605.100 247.050 605.400 ;
        RECT 250.950 605.100 253.050 607.200 ;
        RECT 259.950 606.750 262.050 607.200 ;
        RECT 265.950 606.750 268.050 607.200 ;
        RECT 259.950 605.550 268.050 606.750 ;
        RECT 259.950 605.100 262.050 605.550 ;
        RECT 265.950 605.100 268.050 605.550 ;
        RECT 292.950 605.100 295.050 607.200 ;
        RECT 298.950 605.100 301.050 607.200 ;
        RECT 310.950 606.600 313.050 607.200 ;
        RECT 328.950 606.600 331.050 607.050 ;
        RECT 310.950 605.400 331.050 606.600 ;
        RECT 310.950 605.100 313.050 605.400 ;
        RECT 170.400 602.400 216.600 603.600 ;
        RECT 142.950 598.950 145.050 601.050 ;
        RECT 172.950 600.450 175.050 600.900 ;
        RECT 178.800 600.450 180.900 601.050 ;
        RECT 215.400 600.900 216.600 602.400 ;
        RECT 251.400 601.050 252.600 605.100 ;
        RECT 172.950 599.250 180.900 600.450 ;
        RECT 172.950 598.800 175.050 599.250 ;
        RECT 178.800 598.950 180.900 599.250 ;
        RECT 181.950 600.450 184.050 600.900 ;
        RECT 190.950 600.450 193.050 600.900 ;
        RECT 181.950 599.250 193.050 600.450 ;
        RECT 181.950 598.800 184.050 599.250 ;
        RECT 190.950 598.800 193.050 599.250 ;
        RECT 214.950 598.800 217.050 600.900 ;
        RECT 251.400 599.400 256.050 601.050 ;
        RECT 252.000 598.950 256.050 599.400 ;
        RECT 268.950 600.450 271.050 600.900 ;
        RECT 277.950 600.450 280.050 600.900 ;
        RECT 268.950 599.250 280.050 600.450 ;
        RECT 268.950 598.800 271.050 599.250 ;
        RECT 277.950 598.800 280.050 599.250 ;
        RECT 286.950 600.600 289.050 601.050 ;
        RECT 293.400 600.600 294.600 605.100 ;
        RECT 286.950 599.400 294.600 600.600 ;
        RECT 299.400 600.600 300.600 605.100 ;
        RECT 311.400 603.600 312.600 605.100 ;
        RECT 328.950 604.950 331.050 605.400 ;
        RECT 334.950 605.100 337.050 607.200 ;
        RECT 355.950 605.100 358.050 607.200 ;
        RECT 373.950 605.100 376.050 607.200 ;
        RECT 385.950 606.600 388.050 607.050 ;
        RECT 391.950 606.600 394.050 607.050 ;
        RECT 400.950 606.600 403.050 607.050 ;
        RECT 385.950 605.400 394.050 606.600 ;
        RECT 311.400 602.400 318.600 603.600 ;
        RECT 313.950 600.600 316.050 600.900 ;
        RECT 299.400 599.400 316.050 600.600 ;
        RECT 317.400 600.600 318.600 602.400 ;
        RECT 335.400 601.050 336.600 605.100 ;
        RECT 317.400 599.400 321.600 600.600 ;
        RECT 286.950 598.950 289.050 599.400 ;
        RECT 313.950 598.800 316.050 599.400 ;
        RECT 97.950 597.600 100.050 598.050 ;
        RECT 103.950 597.600 106.050 598.050 ;
        RECT 109.950 597.600 112.050 598.050 ;
        RECT 97.950 596.400 112.050 597.600 ;
        RECT 97.950 595.950 100.050 596.400 ;
        RECT 103.950 595.950 106.050 596.400 ;
        RECT 109.950 595.950 112.050 596.400 ;
        RECT 139.950 597.600 142.050 598.050 ;
        RECT 145.950 597.600 148.050 598.050 ;
        RECT 139.950 596.400 148.050 597.600 ;
        RECT 139.950 595.950 142.050 596.400 ;
        RECT 145.950 595.950 148.050 596.400 ;
        RECT 52.950 594.600 55.050 595.050 ;
        RECT 64.950 594.600 67.050 595.050 ;
        RECT 52.950 593.400 67.050 594.600 ;
        RECT 52.950 592.950 55.050 593.400 ;
        RECT 64.950 592.950 67.050 593.400 ;
        RECT 127.950 594.600 130.050 595.050 ;
        RECT 148.950 594.600 151.050 595.050 ;
        RECT 127.950 593.400 151.050 594.600 ;
        RECT 151.950 594.600 154.050 598.050 ;
        RECT 235.950 597.600 238.050 598.050 ;
        RECT 316.950 597.600 319.050 598.050 ;
        RECT 235.950 596.400 319.050 597.600 ;
        RECT 320.400 597.600 321.600 599.400 ;
        RECT 325.950 600.450 328.050 601.050 ;
        RECT 331.950 600.450 334.050 600.900 ;
        RECT 325.950 599.250 334.050 600.450 ;
        RECT 335.400 599.400 340.050 601.050 ;
        RECT 356.400 600.600 357.600 605.100 ;
        RECT 374.400 603.600 375.600 605.100 ;
        RECT 385.950 604.950 388.050 605.400 ;
        RECT 391.950 604.950 394.050 605.400 ;
        RECT 395.400 605.400 403.050 606.600 ;
        RECT 382.950 603.600 385.050 603.900 ;
        RECT 374.400 602.400 385.050 603.600 ;
        RECT 382.950 601.800 385.050 602.400 ;
        RECT 395.400 600.900 396.600 605.400 ;
        RECT 400.950 604.950 403.050 605.400 ;
        RECT 370.950 600.600 373.050 600.900 ;
        RECT 388.950 600.600 391.050 600.900 ;
        RECT 356.400 599.400 373.050 600.600 ;
        RECT 325.950 598.950 328.050 599.250 ;
        RECT 331.950 598.800 334.050 599.250 ;
        RECT 336.000 598.950 340.050 599.400 ;
        RECT 370.950 598.800 373.050 599.400 ;
        RECT 377.400 599.400 391.050 600.600 ;
        RECT 325.950 597.600 328.050 597.900 ;
        RECT 320.400 596.400 328.050 597.600 ;
        RECT 235.950 595.950 238.050 596.400 ;
        RECT 316.950 595.950 319.050 596.400 ;
        RECT 325.950 595.800 328.050 596.400 ;
        RECT 346.950 597.600 349.050 598.050 ;
        RECT 377.400 597.600 378.600 599.400 ;
        RECT 388.950 598.800 391.050 599.400 ;
        RECT 394.950 598.800 397.050 600.900 ;
        RECT 346.950 596.400 357.600 597.600 ;
        RECT 346.950 595.950 349.050 596.400 ;
        RECT 166.950 594.600 169.050 595.050 ;
        RECT 151.950 594.000 169.050 594.600 ;
        RECT 152.400 593.400 169.050 594.000 ;
        RECT 127.950 592.950 130.050 593.400 ;
        RECT 148.950 592.950 151.050 593.400 ;
        RECT 166.950 592.950 169.050 593.400 ;
        RECT 232.950 594.600 235.050 595.050 ;
        RECT 241.950 594.600 244.050 595.050 ;
        RECT 232.950 593.400 244.050 594.600 ;
        RECT 232.950 592.950 235.050 593.400 ;
        RECT 241.950 592.950 244.050 593.400 ;
        RECT 274.950 594.600 277.050 595.050 ;
        RECT 280.950 594.600 283.050 595.050 ;
        RECT 289.950 594.600 292.050 595.050 ;
        RECT 274.950 593.400 292.050 594.600 ;
        RECT 274.950 592.950 277.050 593.400 ;
        RECT 280.950 592.950 283.050 593.400 ;
        RECT 289.950 592.950 292.050 593.400 ;
        RECT 295.950 594.600 298.050 595.050 ;
        RECT 304.950 594.600 307.050 595.050 ;
        RECT 295.950 593.400 307.050 594.600 ;
        RECT 295.950 592.950 298.050 593.400 ;
        RECT 304.950 592.950 307.050 593.400 ;
        RECT 340.950 594.600 343.050 595.050 ;
        RECT 352.950 594.600 355.050 595.050 ;
        RECT 340.950 593.400 355.050 594.600 ;
        RECT 356.400 594.600 357.600 596.400 ;
        RECT 374.400 596.400 378.600 597.600 ;
        RECT 397.950 597.600 400.050 598.050 ;
        RECT 416.400 597.600 417.600 610.950 ;
        RECT 806.400 610.050 807.600 611.400 ;
        RECT 859.950 610.950 862.050 611.400 ;
        RECT 424.950 609.600 427.050 610.050 ;
        RECT 419.400 608.400 427.050 609.600 ;
        RECT 419.400 600.600 420.600 608.400 ;
        RECT 424.950 607.950 427.050 608.400 ;
        RECT 454.950 607.950 457.050 610.050 ;
        RECT 544.950 609.600 547.050 610.050 ;
        RECT 562.950 609.600 565.050 610.050 ;
        RECT 544.950 608.400 565.050 609.600 ;
        RECT 544.950 607.950 547.050 608.400 ;
        RECT 562.950 607.950 565.050 608.400 ;
        RECT 739.950 609.600 742.050 610.050 ;
        RECT 745.950 609.600 748.050 610.050 ;
        RECT 739.950 608.400 748.050 609.600 ;
        RECT 739.950 607.950 742.050 608.400 ;
        RECT 745.950 607.950 748.050 608.400 ;
        RECT 769.950 609.600 772.050 610.050 ;
        RECT 778.950 609.600 781.050 610.050 ;
        RECT 769.950 608.400 781.050 609.600 ;
        RECT 769.950 607.950 772.050 608.400 ;
        RECT 778.950 607.950 781.050 608.400 ;
        RECT 802.950 608.400 807.600 610.050 ;
        RECT 841.950 609.600 844.050 610.050 ;
        RECT 865.950 609.600 868.050 610.050 ;
        RECT 841.950 608.400 868.050 609.600 ;
        RECT 802.950 607.950 807.000 608.400 ;
        RECT 841.950 607.950 844.050 608.400 ;
        RECT 865.950 607.950 868.050 608.400 ;
        RECT 901.950 609.600 904.050 610.050 ;
        RECT 910.950 609.600 913.050 610.050 ;
        RECT 901.950 608.400 913.050 609.600 ;
        RECT 901.950 607.950 904.050 608.400 ;
        RECT 910.950 607.950 913.050 608.400 ;
        RECT 934.950 609.600 939.000 610.050 ;
        RECT 934.950 607.950 939.600 609.600 ;
        RECT 421.950 605.100 424.050 607.200 ;
        RECT 439.950 606.750 442.050 607.200 ;
        RECT 445.950 606.750 448.050 607.200 ;
        RECT 439.950 605.550 448.050 606.750 ;
        RECT 439.950 605.100 442.050 605.550 ;
        RECT 445.950 605.100 448.050 605.550 ;
        RECT 422.400 603.600 423.600 605.100 ;
        RECT 455.400 603.600 456.600 607.950 ;
        RECT 499.950 606.600 502.050 607.050 ;
        RECT 532.950 606.600 535.050 607.050 ;
        RECT 499.950 605.400 535.050 606.600 ;
        RECT 499.950 604.950 502.050 605.400 ;
        RECT 532.950 604.950 535.050 605.400 ;
        RECT 544.950 605.100 547.050 607.200 ;
        RECT 550.950 606.750 553.050 607.200 ;
        RECT 556.950 606.750 559.050 607.200 ;
        RECT 550.950 605.550 559.050 606.750 ;
        RECT 598.950 606.600 601.050 607.050 ;
        RECT 550.950 605.100 553.050 605.550 ;
        RECT 556.950 605.100 559.050 605.550 ;
        RECT 572.400 605.400 601.050 606.600 ;
        RECT 466.950 603.600 469.050 604.050 ;
        RECT 545.400 603.600 546.600 605.100 ;
        RECT 422.400 602.400 429.600 603.600 ;
        RECT 455.400 602.400 469.050 603.600 ;
        RECT 539.400 603.000 546.600 603.600 ;
        RECT 424.950 600.600 427.050 601.050 ;
        RECT 419.400 599.400 427.050 600.600 ;
        RECT 428.400 600.600 429.600 602.400 ;
        RECT 466.950 601.950 469.050 602.400 ;
        RECT 538.950 602.400 546.600 603.000 ;
        RECT 436.950 600.600 439.050 600.900 ;
        RECT 428.400 599.400 439.050 600.600 ;
        RECT 424.950 598.950 427.050 599.400 ;
        RECT 436.950 598.800 439.050 599.400 ;
        RECT 448.950 600.600 451.050 601.050 ;
        RECT 472.950 600.600 475.050 601.050 ;
        RECT 448.950 599.400 475.050 600.600 ;
        RECT 448.950 598.950 451.050 599.400 ;
        RECT 472.950 598.950 475.050 599.400 ;
        RECT 538.950 598.950 541.050 602.400 ;
        RECT 572.400 601.050 573.600 605.400 ;
        RECT 598.950 604.950 601.050 605.400 ;
        RECT 637.950 606.750 640.050 607.200 ;
        RECT 652.950 606.750 655.050 607.200 ;
        RECT 637.950 605.550 655.050 606.750 ;
        RECT 637.950 605.100 640.050 605.550 ;
        RECT 652.950 605.100 655.050 605.550 ;
        RECT 658.950 606.750 661.050 606.900 ;
        RECT 673.950 606.750 676.050 607.200 ;
        RECT 658.950 605.550 676.050 606.750 ;
        RECT 658.950 604.800 661.050 605.550 ;
        RECT 673.950 605.100 676.050 605.550 ;
        RECT 727.950 606.750 730.050 607.200 ;
        RECT 733.950 606.750 736.050 607.200 ;
        RECT 727.950 605.550 736.050 606.750 ;
        RECT 727.950 605.100 730.050 605.550 ;
        RECT 733.950 605.100 736.050 605.550 ;
        RECT 748.950 606.600 751.050 607.050 ;
        RECT 763.950 606.600 766.050 607.050 ;
        RECT 748.950 605.400 766.050 606.600 ;
        RECT 748.950 604.950 751.050 605.400 ;
        RECT 763.950 604.950 766.050 605.400 ;
        RECT 577.950 603.600 580.050 604.050 ;
        RECT 595.950 603.600 598.050 604.050 ;
        RECT 781.950 603.600 784.050 607.050 ;
        RECT 790.950 606.600 793.050 607.200 ;
        RECT 577.950 602.400 598.050 603.600 ;
        RECT 577.950 601.950 580.050 602.400 ;
        RECT 595.950 601.950 598.050 602.400 ;
        RECT 779.400 603.000 784.050 603.600 ;
        RECT 785.400 605.400 793.050 606.600 ;
        RECT 779.400 602.400 783.600 603.000 ;
        RECT 556.950 600.600 559.050 601.050 ;
        RECT 565.950 600.600 568.050 600.900 ;
        RECT 556.950 599.400 568.050 600.600 ;
        RECT 556.950 598.950 559.050 599.400 ;
        RECT 565.950 598.800 568.050 599.400 ;
        RECT 571.950 598.950 574.050 601.050 ;
        RECT 622.950 600.600 625.050 601.050 ;
        RECT 634.950 600.600 637.050 601.050 ;
        RECT 640.950 600.600 643.050 601.050 ;
        RECT 622.950 599.400 643.050 600.600 ;
        RECT 622.950 598.950 625.050 599.400 ;
        RECT 634.950 598.950 637.050 599.400 ;
        RECT 640.950 598.950 643.050 599.400 ;
        RECT 664.950 600.450 667.050 600.900 ;
        RECT 670.950 600.450 673.050 600.900 ;
        RECT 664.950 599.250 673.050 600.450 ;
        RECT 664.950 598.800 667.050 599.250 ;
        RECT 670.950 598.800 673.050 599.250 ;
        RECT 679.950 600.450 682.050 600.900 ;
        RECT 694.950 600.450 697.050 600.900 ;
        RECT 679.950 599.250 697.050 600.450 ;
        RECT 679.950 598.800 682.050 599.250 ;
        RECT 694.950 598.800 697.050 599.250 ;
        RECT 700.950 600.600 703.050 601.050 ;
        RECT 712.950 600.600 715.050 600.900 ;
        RECT 700.950 599.400 715.050 600.600 ;
        RECT 700.950 598.950 703.050 599.400 ;
        RECT 712.950 598.800 715.050 599.400 ;
        RECT 724.950 600.450 727.050 600.900 ;
        RECT 754.950 600.450 757.050 600.900 ;
        RECT 724.950 599.250 757.050 600.450 ;
        RECT 724.950 598.800 727.050 599.250 ;
        RECT 754.950 598.800 757.050 599.250 ;
        RECT 769.950 600.600 772.050 601.050 ;
        RECT 779.400 600.600 780.600 602.400 ;
        RECT 785.400 601.050 786.600 605.400 ;
        RECT 790.950 605.100 793.050 605.400 ;
        RECT 805.950 606.600 808.050 607.050 ;
        RECT 820.950 606.750 823.050 607.200 ;
        RECT 826.950 606.750 829.050 607.200 ;
        RECT 805.950 605.400 816.600 606.600 ;
        RECT 805.950 604.950 808.050 605.400 ;
        RECT 799.950 603.600 802.050 604.050 ;
        RECT 799.950 602.400 813.600 603.600 ;
        RECT 799.950 601.950 802.050 602.400 ;
        RECT 769.950 599.400 780.600 600.600 ;
        RECT 781.950 599.400 786.600 601.050 ;
        RECT 769.950 598.950 772.050 599.400 ;
        RECT 781.950 598.950 786.000 599.400 ;
        RECT 397.950 596.400 417.600 597.600 ;
        RECT 475.950 597.600 478.050 598.050 ;
        RECT 514.950 597.600 517.050 598.050 ;
        RECT 475.950 596.400 517.050 597.600 ;
        RECT 374.400 594.600 375.600 596.400 ;
        RECT 397.950 595.950 400.050 596.400 ;
        RECT 475.950 595.950 478.050 596.400 ;
        RECT 514.950 595.950 517.050 596.400 ;
        RECT 541.950 597.600 544.050 598.050 ;
        RECT 583.950 597.600 586.050 598.050 ;
        RECT 541.950 596.400 586.050 597.600 ;
        RECT 541.950 595.950 544.050 596.400 ;
        RECT 583.950 595.950 586.050 596.400 ;
        RECT 718.950 597.600 721.050 598.050 ;
        RECT 730.950 597.600 733.050 598.050 ;
        RECT 718.950 596.400 733.050 597.600 ;
        RECT 718.950 595.950 721.050 596.400 ;
        RECT 730.950 595.950 733.050 596.400 ;
        RECT 745.950 597.600 748.050 598.050 ;
        RECT 793.950 597.600 796.050 598.050 ;
        RECT 745.950 596.400 796.050 597.600 ;
        RECT 812.400 597.600 813.600 602.400 ;
        RECT 815.400 600.600 816.600 605.400 ;
        RECT 820.950 605.550 829.050 606.750 ;
        RECT 820.950 605.100 823.050 605.550 ;
        RECT 826.950 605.100 829.050 605.550 ;
        RECT 835.950 605.100 838.050 607.200 ;
        RECT 853.950 605.100 856.050 607.200 ;
        RECT 871.950 606.750 874.050 607.200 ;
        RECT 889.950 606.750 892.050 607.200 ;
        RECT 871.950 606.600 892.050 606.750 ;
        RECT 895.800 606.600 897.900 607.050 ;
        RECT 871.950 605.550 897.900 606.600 ;
        RECT 871.950 605.100 874.050 605.550 ;
        RECT 889.950 605.400 897.900 605.550 ;
        RECT 889.950 605.100 892.050 605.400 ;
        RECT 817.950 600.600 820.050 600.900 ;
        RECT 815.400 599.400 820.050 600.600 ;
        RECT 817.950 598.800 820.050 599.400 ;
        RECT 823.950 600.600 826.050 601.050 ;
        RECT 836.400 600.600 837.600 605.100 ;
        RECT 823.950 599.400 837.600 600.600 ;
        RECT 844.950 600.600 847.050 601.050 ;
        RECT 854.400 600.600 855.600 605.100 ;
        RECT 895.800 604.950 897.900 605.400 ;
        RECT 898.950 604.950 901.050 607.050 ;
        RECT 925.950 605.100 928.050 607.200 ;
        RECT 931.950 605.100 934.050 607.200 ;
        RECT 899.400 601.050 900.600 604.950 ;
        RECT 844.950 599.400 855.600 600.600 ;
        RECT 823.950 598.950 826.050 599.400 ;
        RECT 844.950 598.950 847.050 599.400 ;
        RECT 898.950 598.950 901.050 601.050 ;
        RECT 926.400 600.600 927.600 605.100 ;
        RECT 917.400 599.400 927.600 600.600 ;
        RECT 932.400 601.050 933.600 605.100 ;
        RECT 932.400 599.400 937.050 601.050 ;
        RECT 838.950 597.600 841.050 598.050 ;
        RECT 862.950 597.600 865.050 598.050 ;
        RECT 812.400 596.400 865.050 597.600 ;
        RECT 745.950 595.950 748.050 596.400 ;
        RECT 793.950 595.950 796.050 596.400 ;
        RECT 838.950 595.950 841.050 596.400 ;
        RECT 862.950 595.950 865.050 596.400 ;
        RECT 910.950 597.600 913.050 598.050 ;
        RECT 917.400 597.600 918.600 599.400 ;
        RECT 933.000 598.950 937.050 599.400 ;
        RECT 910.950 596.400 918.600 597.600 ;
        RECT 910.950 595.950 913.050 596.400 ;
        RECT 356.400 593.400 375.600 594.600 ;
        RECT 403.950 594.600 406.050 594.900 ;
        RECT 412.800 594.600 414.900 595.050 ;
        RECT 403.950 593.400 414.900 594.600 ;
        RECT 340.950 592.950 343.050 593.400 ;
        RECT 352.950 592.950 355.050 593.400 ;
        RECT 403.950 592.800 406.050 593.400 ;
        RECT 412.800 592.950 414.900 593.400 ;
        RECT 415.950 594.600 418.050 595.050 ;
        RECT 427.950 594.600 430.050 595.050 ;
        RECT 415.950 593.400 430.050 594.600 ;
        RECT 415.950 592.950 418.050 593.400 ;
        RECT 427.950 592.950 430.050 593.400 ;
        RECT 436.950 594.600 439.050 595.050 ;
        RECT 451.950 594.600 454.050 595.050 ;
        RECT 436.950 593.400 454.050 594.600 ;
        RECT 436.950 592.950 439.050 593.400 ;
        RECT 451.950 592.950 454.050 593.400 ;
        RECT 463.950 594.600 466.050 595.050 ;
        RECT 514.950 594.600 517.050 594.900 ;
        RECT 535.950 594.600 538.050 595.050 ;
        RECT 463.950 593.400 538.050 594.600 ;
        RECT 463.950 592.950 466.050 593.400 ;
        RECT 514.950 592.800 517.050 593.400 ;
        RECT 535.950 592.950 538.050 593.400 ;
        RECT 541.950 594.600 544.050 594.900 ;
        RECT 643.950 594.600 646.050 595.050 ;
        RECT 676.950 594.600 679.050 595.050 ;
        RECT 541.950 593.400 585.600 594.600 ;
        RECT 541.950 592.800 544.050 593.400 ;
        RECT 13.950 591.600 16.050 592.050 ;
        RECT 43.950 591.600 46.050 592.050 ;
        RECT 13.950 590.400 46.050 591.600 ;
        RECT 13.950 589.950 16.050 590.400 ;
        RECT 43.950 589.950 46.050 590.400 ;
        RECT 55.950 591.600 58.050 592.050 ;
        RECT 79.950 591.600 82.050 592.050 ;
        RECT 55.950 590.400 82.050 591.600 ;
        RECT 55.950 589.950 58.050 590.400 ;
        RECT 79.950 589.950 82.050 590.400 ;
        RECT 88.950 591.600 91.050 592.050 ;
        RECT 109.950 591.600 112.050 592.050 ;
        RECT 88.950 590.400 112.050 591.600 ;
        RECT 88.950 589.950 91.050 590.400 ;
        RECT 109.950 589.950 112.050 590.400 ;
        RECT 121.950 591.600 124.050 592.050 ;
        RECT 163.950 591.600 166.050 592.050 ;
        RECT 121.950 590.400 166.050 591.600 ;
        RECT 121.950 589.950 124.050 590.400 ;
        RECT 163.950 589.950 166.050 590.400 ;
        RECT 172.950 591.600 175.050 592.050 ;
        RECT 178.950 591.600 181.050 592.050 ;
        RECT 172.950 590.400 181.050 591.600 ;
        RECT 172.950 589.950 175.050 590.400 ;
        RECT 178.950 589.950 181.050 590.400 ;
        RECT 253.950 591.600 256.050 592.050 ;
        RECT 280.800 591.600 282.900 591.900 ;
        RECT 253.950 590.400 282.900 591.600 ;
        RECT 253.950 589.950 256.050 590.400 ;
        RECT 280.800 589.800 282.900 590.400 ;
        RECT 283.950 591.600 286.050 592.050 ;
        RECT 331.950 591.600 334.050 592.050 ;
        RECT 283.950 590.400 334.050 591.600 ;
        RECT 283.950 589.950 286.050 590.400 ;
        RECT 331.950 589.950 334.050 590.400 ;
        RECT 349.950 591.600 352.050 592.050 ;
        RECT 376.950 591.600 379.050 592.050 ;
        RECT 349.950 590.400 379.050 591.600 ;
        RECT 349.950 589.950 352.050 590.400 ;
        RECT 376.950 589.950 379.050 590.400 ;
        RECT 430.950 591.600 433.050 592.050 ;
        RECT 445.950 591.600 448.050 592.050 ;
        RECT 430.950 590.400 448.050 591.600 ;
        RECT 430.950 589.950 433.050 590.400 ;
        RECT 445.950 589.950 448.050 590.400 ;
        RECT 463.950 591.600 466.050 591.900 ;
        RECT 517.950 591.600 520.050 592.050 ;
        RECT 463.950 590.400 520.050 591.600 ;
        RECT 463.950 589.800 466.050 590.400 ;
        RECT 517.950 589.950 520.050 590.400 ;
        RECT 532.950 591.600 535.050 592.050 ;
        RECT 547.950 591.600 550.050 592.050 ;
        RECT 532.950 590.400 550.050 591.600 ;
        RECT 532.950 589.950 535.050 590.400 ;
        RECT 547.950 589.950 550.050 590.400 ;
        RECT 61.950 588.600 64.050 589.050 ;
        RECT 106.950 588.600 109.050 589.050 ;
        RECT 190.950 588.600 193.050 589.050 ;
        RECT 205.950 588.600 208.050 589.050 ;
        RECT 391.950 588.600 394.050 589.050 ;
        RECT 61.950 587.400 109.050 588.600 ;
        RECT 61.950 586.950 64.050 587.400 ;
        RECT 106.950 586.950 109.050 587.400 ;
        RECT 110.400 587.400 180.600 588.600 ;
        RECT 64.950 585.600 67.050 586.050 ;
        RECT 110.400 585.600 111.600 587.400 ;
        RECT 64.950 584.400 111.600 585.600 ;
        RECT 124.950 585.600 127.050 586.050 ;
        RECT 136.950 585.600 139.050 586.050 ;
        RECT 124.950 584.400 139.050 585.600 ;
        RECT 64.950 583.950 67.050 584.400 ;
        RECT 124.950 583.950 127.050 584.400 ;
        RECT 136.950 583.950 139.050 584.400 ;
        RECT 142.950 585.600 145.050 586.050 ;
        RECT 179.400 585.600 180.600 587.400 ;
        RECT 190.950 587.400 208.050 588.600 ;
        RECT 190.950 586.950 193.050 587.400 ;
        RECT 205.950 586.950 208.050 587.400 ;
        RECT 212.400 587.400 394.050 588.600 ;
        RECT 212.400 585.600 213.600 587.400 ;
        RECT 391.950 586.950 394.050 587.400 ;
        RECT 469.950 588.600 472.050 589.050 ;
        RECT 481.950 588.600 484.050 589.050 ;
        RECT 469.950 587.400 484.050 588.600 ;
        RECT 469.950 586.950 472.050 587.400 ;
        RECT 481.950 586.950 484.050 587.400 ;
        RECT 493.950 588.600 496.050 589.050 ;
        RECT 574.950 588.600 577.050 589.050 ;
        RECT 493.950 587.400 577.050 588.600 ;
        RECT 584.400 588.600 585.600 593.400 ;
        RECT 643.950 593.400 679.050 594.600 ;
        RECT 643.950 592.950 646.050 593.400 ;
        RECT 676.950 592.950 679.050 593.400 ;
        RECT 736.950 594.600 739.050 595.050 ;
        RECT 763.950 594.600 766.050 595.050 ;
        RECT 736.950 593.400 766.050 594.600 ;
        RECT 736.950 592.950 739.050 593.400 ;
        RECT 763.950 592.950 766.050 593.400 ;
        RECT 799.950 594.600 802.050 595.050 ;
        RECT 814.950 594.600 817.050 595.050 ;
        RECT 799.950 593.400 817.050 594.600 ;
        RECT 799.950 592.950 802.050 593.400 ;
        RECT 814.950 592.950 817.050 593.400 ;
        RECT 856.950 594.600 859.050 595.050 ;
        RECT 862.950 594.600 865.050 594.900 ;
        RECT 856.950 593.400 865.050 594.600 ;
        RECT 856.950 592.950 859.050 593.400 ;
        RECT 862.950 592.800 865.050 593.400 ;
        RECT 919.950 594.600 922.050 595.050 ;
        RECT 931.950 594.600 934.050 595.050 ;
        RECT 919.950 593.400 934.050 594.600 ;
        RECT 919.950 592.950 922.050 593.400 ;
        RECT 931.950 592.950 934.050 593.400 ;
        RECT 745.950 591.600 748.050 592.050 ;
        RECT 832.950 591.600 835.050 592.050 ;
        RECT 745.950 590.400 835.050 591.600 ;
        RECT 745.950 589.950 748.050 590.400 ;
        RECT 832.950 589.950 835.050 590.400 ;
        RECT 895.950 591.600 898.050 592.050 ;
        RECT 934.950 591.600 937.050 592.050 ;
        RECT 895.950 590.400 937.050 591.600 ;
        RECT 895.950 589.950 898.050 590.400 ;
        RECT 934.950 589.950 937.050 590.400 ;
        RECT 938.400 589.050 939.600 607.950 ;
        RECT 604.950 588.600 607.050 589.050 ;
        RECT 584.400 587.400 607.050 588.600 ;
        RECT 493.950 586.950 496.050 587.400 ;
        RECT 574.950 586.950 577.050 587.400 ;
        RECT 604.950 586.950 607.050 587.400 ;
        RECT 652.950 588.600 655.050 589.050 ;
        RECT 898.950 588.600 901.050 589.050 ;
        RECT 922.950 588.600 925.050 589.050 ;
        RECT 936.000 588.900 939.600 589.050 ;
        RECT 652.950 587.400 867.600 588.600 ;
        RECT 652.950 586.950 655.050 587.400 ;
        RECT 142.950 584.400 177.600 585.600 ;
        RECT 179.400 584.400 213.600 585.600 ;
        RECT 286.950 585.600 289.050 586.050 ;
        RECT 295.950 585.600 298.050 586.050 ;
        RECT 286.950 584.400 298.050 585.600 ;
        RECT 142.950 583.950 145.050 584.400 ;
        RECT 28.950 582.600 31.050 583.050 ;
        RECT 58.950 582.600 61.050 583.050 ;
        RECT 28.950 581.400 61.050 582.600 ;
        RECT 28.950 580.950 31.050 581.400 ;
        RECT 58.950 580.950 61.050 581.400 ;
        RECT 106.950 582.600 109.050 583.050 ;
        RECT 121.950 582.600 124.050 583.050 ;
        RECT 106.950 581.400 124.050 582.600 ;
        RECT 106.950 580.950 109.050 581.400 ;
        RECT 121.950 580.950 124.050 581.400 ;
        RECT 157.950 582.600 160.050 583.050 ;
        RECT 169.950 582.600 172.050 583.050 ;
        RECT 157.950 581.400 172.050 582.600 ;
        RECT 176.400 582.600 177.600 584.400 ;
        RECT 286.950 583.950 289.050 584.400 ;
        RECT 295.950 583.950 298.050 584.400 ;
        RECT 391.950 585.600 394.050 585.900 ;
        RECT 397.950 585.600 400.050 586.050 ;
        RECT 391.950 584.400 400.050 585.600 ;
        RECT 391.950 583.800 394.050 584.400 ;
        RECT 397.950 583.950 400.050 584.400 ;
        RECT 409.950 585.600 412.050 586.050 ;
        RECT 418.950 585.600 421.050 586.050 ;
        RECT 409.950 584.400 421.050 585.600 ;
        RECT 409.950 583.950 412.050 584.400 ;
        RECT 418.950 583.950 421.050 584.400 ;
        RECT 466.950 585.600 469.050 586.050 ;
        RECT 487.950 585.600 490.050 586.050 ;
        RECT 466.950 584.400 490.050 585.600 ;
        RECT 466.950 583.950 469.050 584.400 ;
        RECT 487.950 583.950 490.050 584.400 ;
        RECT 517.950 585.600 520.050 586.050 ;
        RECT 541.950 585.600 544.050 586.050 ;
        RECT 517.950 584.400 544.050 585.600 ;
        RECT 517.950 583.950 520.050 584.400 ;
        RECT 541.950 583.950 544.050 584.400 ;
        RECT 553.950 585.600 556.050 586.050 ;
        RECT 565.950 585.600 568.050 586.050 ;
        RECT 553.950 584.400 568.050 585.600 ;
        RECT 553.950 583.950 556.050 584.400 ;
        RECT 565.950 583.950 568.050 584.400 ;
        RECT 619.950 585.600 622.050 586.050 ;
        RECT 625.950 585.600 628.050 586.050 ;
        RECT 619.950 584.400 628.050 585.600 ;
        RECT 619.950 583.950 622.050 584.400 ;
        RECT 625.950 583.950 628.050 584.400 ;
        RECT 760.950 585.600 763.050 586.050 ;
        RECT 775.950 585.600 778.050 586.050 ;
        RECT 760.950 584.400 778.050 585.600 ;
        RECT 866.400 585.600 867.600 587.400 ;
        RECT 898.950 587.400 925.050 588.600 ;
        RECT 898.950 586.950 901.050 587.400 ;
        RECT 922.950 586.950 925.050 587.400 ;
        RECT 934.950 587.400 939.600 588.900 ;
        RECT 934.950 586.950 939.000 587.400 ;
        RECT 934.950 586.800 937.050 586.950 ;
        RECT 871.950 585.600 874.050 586.050 ;
        RECT 910.950 585.600 913.050 586.050 ;
        RECT 866.400 584.400 874.050 585.600 ;
        RECT 760.950 583.950 763.050 584.400 ;
        RECT 775.950 583.950 778.050 584.400 ;
        RECT 871.950 583.950 874.050 584.400 ;
        RECT 884.400 584.400 913.050 585.600 ;
        RECT 884.400 583.050 885.600 584.400 ;
        RECT 910.950 583.950 913.050 584.400 ;
        RECT 205.950 582.600 208.050 583.050 ;
        RECT 176.400 581.400 208.050 582.600 ;
        RECT 157.950 580.950 160.050 581.400 ;
        RECT 169.950 580.950 172.050 581.400 ;
        RECT 205.950 580.950 208.050 581.400 ;
        RECT 346.950 582.600 349.050 583.050 ;
        RECT 355.950 582.600 358.050 583.050 ;
        RECT 346.950 581.400 358.050 582.600 ;
        RECT 346.950 580.950 349.050 581.400 ;
        RECT 355.950 580.950 358.050 581.400 ;
        RECT 415.950 582.600 418.050 583.050 ;
        RECT 502.950 582.600 505.050 583.050 ;
        RECT 415.950 581.400 505.050 582.600 ;
        RECT 415.950 580.950 418.050 581.400 ;
        RECT 502.950 580.950 505.050 581.400 ;
        RECT 604.950 582.600 607.050 583.050 ;
        RECT 649.950 582.600 652.050 583.050 ;
        RECT 604.950 581.400 652.050 582.600 ;
        RECT 604.950 580.950 607.050 581.400 ;
        RECT 649.950 580.950 652.050 581.400 ;
        RECT 877.950 582.600 880.050 583.050 ;
        RECT 883.950 582.600 886.050 583.050 ;
        RECT 877.950 581.400 886.050 582.600 ;
        RECT 877.950 580.950 880.050 581.400 ;
        RECT 883.950 580.950 886.050 581.400 ;
        RECT 127.950 579.600 130.050 580.050 ;
        RECT 142.950 579.600 145.050 580.050 ;
        RECT 127.950 578.400 145.050 579.600 ;
        RECT 127.950 577.950 130.050 578.400 ;
        RECT 142.950 577.950 145.050 578.400 ;
        RECT 154.950 579.600 157.050 580.050 ;
        RECT 178.950 579.600 181.050 580.050 ;
        RECT 154.950 578.400 181.050 579.600 ;
        RECT 154.950 577.950 157.050 578.400 ;
        RECT 178.950 577.950 181.050 578.400 ;
        RECT 214.950 579.600 217.050 580.050 ;
        RECT 223.950 579.600 226.050 580.050 ;
        RECT 214.950 578.400 226.050 579.600 ;
        RECT 214.950 577.950 217.050 578.400 ;
        RECT 223.950 577.950 226.050 578.400 ;
        RECT 343.950 579.600 346.050 580.050 ;
        RECT 358.950 579.600 361.050 580.050 ;
        RECT 343.950 578.400 361.050 579.600 ;
        RECT 343.950 577.950 346.050 578.400 ;
        RECT 358.950 577.950 361.050 578.400 ;
        RECT 385.950 579.600 388.050 580.050 ;
        RECT 409.950 579.600 412.050 580.050 ;
        RECT 385.950 578.400 412.050 579.600 ;
        RECT 385.950 577.950 388.050 578.400 ;
        RECT 409.950 577.950 412.050 578.400 ;
        RECT 526.950 579.600 529.050 580.050 ;
        RECT 553.950 579.600 556.050 580.050 ;
        RECT 526.950 578.400 556.050 579.600 ;
        RECT 526.950 577.950 529.050 578.400 ;
        RECT 553.950 577.950 556.050 578.400 ;
        RECT 613.950 579.600 616.050 580.050 ;
        RECT 631.950 579.600 634.050 580.050 ;
        RECT 613.950 578.400 634.050 579.600 ;
        RECT 613.950 577.950 616.050 578.400 ;
        RECT 631.950 577.950 634.050 578.400 ;
        RECT 718.950 579.600 721.050 580.050 ;
        RECT 733.950 579.600 736.050 580.050 ;
        RECT 718.950 578.400 736.050 579.600 ;
        RECT 718.950 577.950 721.050 578.400 ;
        RECT 733.950 577.950 736.050 578.400 ;
        RECT 790.950 579.600 793.050 580.050 ;
        RECT 802.950 579.600 805.050 580.050 ;
        RECT 790.950 578.400 805.050 579.600 ;
        RECT 790.950 577.950 793.050 578.400 ;
        RECT 802.950 577.950 805.050 578.400 ;
        RECT 847.950 579.600 850.050 580.050 ;
        RECT 853.950 579.600 856.050 580.050 ;
        RECT 847.950 578.400 856.050 579.600 ;
        RECT 847.950 577.950 850.050 578.400 ;
        RECT 853.950 577.950 856.050 578.400 ;
        RECT 58.950 576.600 61.050 577.050 ;
        RECT 82.950 576.600 85.050 577.050 ;
        RECT 88.950 576.600 91.050 577.050 ;
        RECT 58.950 575.400 66.600 576.600 ;
        RECT 58.950 574.950 61.050 575.400 ;
        RECT 16.950 572.100 19.050 574.200 ;
        RECT 34.950 573.600 37.050 574.200 ;
        RECT 43.950 573.600 46.050 574.050 ;
        RECT 34.950 572.400 46.050 573.600 ;
        RECT 34.950 572.100 37.050 572.400 ;
        RECT 17.400 570.600 18.600 572.100 ;
        RECT 43.950 571.950 46.050 572.400 ;
        RECT 52.950 573.750 55.050 574.200 ;
        RECT 61.950 573.750 64.050 574.200 ;
        RECT 52.950 572.550 64.050 573.750 ;
        RECT 52.950 572.100 55.050 572.550 ;
        RECT 61.950 572.100 64.050 572.550 ;
        RECT 17.400 570.000 27.600 570.600 ;
        RECT 17.400 569.400 28.050 570.000 ;
        RECT 25.950 565.950 28.050 569.400 ;
        RECT 65.400 567.600 66.600 575.400 ;
        RECT 82.950 575.400 91.050 576.600 ;
        RECT 82.950 574.950 85.050 575.400 ;
        RECT 88.950 574.950 91.050 575.400 ;
        RECT 103.950 576.600 106.050 577.050 ;
        RECT 151.950 576.600 154.050 577.050 ;
        RECT 103.950 575.400 154.050 576.600 ;
        RECT 103.950 574.950 106.050 575.400 ;
        RECT 151.950 574.950 154.050 575.400 ;
        RECT 211.950 576.600 214.050 577.050 ;
        RECT 220.950 576.600 223.050 577.200 ;
        RECT 211.950 575.400 223.050 576.600 ;
        RECT 211.950 574.950 214.050 575.400 ;
        RECT 220.950 575.100 223.050 575.400 ;
        RECT 283.950 576.600 286.050 577.050 ;
        RECT 298.950 576.600 301.050 577.050 ;
        RECT 319.950 576.600 322.050 577.050 ;
        RECT 283.950 575.400 322.050 576.600 ;
        RECT 283.950 574.950 286.050 575.400 ;
        RECT 298.950 574.950 301.050 575.400 ;
        RECT 319.950 574.950 322.050 575.400 ;
        RECT 415.950 574.950 418.050 577.050 ;
        RECT 478.950 576.600 481.050 577.050 ;
        RECT 484.950 576.600 487.050 577.050 ;
        RECT 478.950 575.400 487.050 576.600 ;
        RECT 478.950 574.950 481.050 575.400 ;
        RECT 484.950 574.950 487.050 575.400 ;
        RECT 79.950 572.100 82.050 574.200 ;
        RECT 91.950 573.600 94.050 574.050 ;
        RECT 115.950 573.600 118.050 574.200 ;
        RECT 127.950 573.600 130.050 574.050 ;
        RECT 91.950 572.400 114.600 573.600 ;
        RECT 80.400 570.600 81.600 572.100 ;
        RECT 91.950 571.950 94.050 572.400 ;
        RECT 80.400 570.000 87.600 570.600 ;
        RECT 80.400 569.400 88.050 570.000 ;
        RECT 70.950 567.600 73.050 567.900 ;
        RECT 65.400 566.400 73.050 567.600 ;
        RECT 70.950 565.800 73.050 566.400 ;
        RECT 85.950 565.950 88.050 569.400 ;
        RECT 113.400 567.900 114.600 572.400 ;
        RECT 115.950 572.400 130.050 573.600 ;
        RECT 115.950 572.100 118.050 572.400 ;
        RECT 127.950 571.950 130.050 572.400 ;
        RECT 133.950 572.100 136.050 574.200 ;
        RECT 139.950 573.600 142.050 574.200 ;
        RECT 148.950 573.600 151.050 574.050 ;
        RECT 139.950 572.400 151.050 573.600 ;
        RECT 139.950 572.100 142.050 572.400 ;
        RECT 94.950 567.600 97.050 567.900 ;
        RECT 94.950 567.000 102.600 567.600 ;
        RECT 94.950 566.400 103.050 567.000 ;
        RECT 94.950 565.800 97.050 566.400 ;
        RECT 22.950 564.600 25.050 565.050 ;
        RECT 31.950 564.600 34.050 565.050 ;
        RECT 22.950 563.400 34.050 564.600 ;
        RECT 22.950 562.950 25.050 563.400 ;
        RECT 31.950 562.950 34.050 563.400 ;
        RECT 49.950 564.600 52.050 565.050 ;
        RECT 88.950 564.600 91.050 565.050 ;
        RECT 49.950 563.400 91.050 564.600 ;
        RECT 49.950 562.950 52.050 563.400 ;
        RECT 88.950 562.950 91.050 563.400 ;
        RECT 100.950 564.600 103.050 566.400 ;
        RECT 112.950 565.800 115.050 567.900 ;
        RECT 134.400 564.600 135.600 572.100 ;
        RECT 148.950 571.950 151.050 572.400 ;
        RECT 157.950 572.100 160.050 574.200 ;
        RECT 136.950 567.450 139.050 567.900 ;
        RECT 142.950 567.450 145.050 567.900 ;
        RECT 136.950 566.250 145.050 567.450 ;
        RECT 136.950 565.800 139.050 566.250 ;
        RECT 142.950 565.800 145.050 566.250 ;
        RECT 148.950 567.600 151.050 568.050 ;
        RECT 158.400 567.600 159.600 572.100 ;
        RECT 163.950 571.950 166.050 574.050 ;
        RECT 193.950 573.600 196.050 574.050 ;
        RECT 199.950 573.600 202.050 574.200 ;
        RECT 193.950 572.400 202.050 573.600 ;
        RECT 193.950 571.950 196.050 572.400 ;
        RECT 199.950 572.100 202.050 572.400 ;
        RECT 220.950 571.950 223.050 574.050 ;
        RECT 310.950 573.600 313.050 574.200 ;
        RECT 337.950 573.600 340.050 574.200 ;
        RECT 352.950 573.600 355.050 574.200 ;
        RECT 310.950 572.400 330.600 573.600 ;
        RECT 310.950 572.100 313.050 572.400 ;
        RECT 164.400 568.050 165.600 571.950 ;
        RECT 148.950 566.400 159.600 567.600 ;
        RECT 148.950 565.950 151.050 566.400 ;
        RECT 163.950 565.950 166.050 568.050 ;
        RECT 172.950 567.600 175.050 568.050 ;
        RECT 208.950 567.600 211.050 567.900 ;
        RECT 172.950 567.450 211.050 567.600 ;
        RECT 217.950 567.450 220.050 567.900 ;
        RECT 172.950 566.400 220.050 567.450 ;
        RECT 172.950 565.950 175.050 566.400 ;
        RECT 208.950 566.250 220.050 566.400 ;
        RECT 208.950 565.800 211.050 566.250 ;
        RECT 217.950 565.800 220.050 566.250 ;
        RECT 221.400 565.050 222.600 571.950 ;
        RECT 226.950 567.600 229.050 567.900 ;
        RECT 235.950 567.600 238.050 571.050 ;
        RECT 280.950 570.600 283.050 571.050 ;
        RECT 292.950 570.600 295.050 571.200 ;
        RECT 280.950 569.400 295.050 570.600 ;
        RECT 280.950 568.950 283.050 569.400 ;
        RECT 292.950 569.100 295.050 569.400 ;
        RECT 226.950 567.000 238.050 567.600 ;
        RECT 256.950 567.600 259.050 568.050 ;
        RECT 277.950 567.600 280.050 568.050 ;
        RECT 226.950 566.400 237.600 567.000 ;
        RECT 256.950 566.400 280.050 567.600 ;
        RECT 226.950 565.800 229.050 566.400 ;
        RECT 256.950 565.950 259.050 566.400 ;
        RECT 277.950 565.950 280.050 566.400 ;
        RECT 301.950 567.600 304.050 568.050 ;
        RECT 329.400 567.900 330.600 572.400 ;
        RECT 337.950 572.400 355.050 573.600 ;
        RECT 337.950 572.100 340.050 572.400 ;
        RECT 352.950 572.100 355.050 572.400 ;
        RECT 367.950 573.600 370.050 574.050 ;
        RECT 376.950 573.600 379.050 574.200 ;
        RECT 367.950 572.400 379.050 573.600 ;
        RECT 367.950 571.950 370.050 572.400 ;
        RECT 376.950 572.100 379.050 572.400 ;
        RECT 397.950 573.600 400.050 574.200 ;
        RECT 403.950 573.750 406.050 574.200 ;
        RECT 412.950 573.750 415.050 574.200 ;
        RECT 397.950 572.400 402.600 573.600 ;
        RECT 397.950 572.100 400.050 572.400 ;
        RECT 307.950 567.600 310.050 567.900 ;
        RECT 301.950 566.400 310.050 567.600 ;
        RECT 301.950 565.950 304.050 566.400 ;
        RECT 307.950 565.800 310.050 566.400 ;
        RECT 328.950 565.800 331.050 567.900 ;
        RECT 361.950 567.450 364.050 567.900 ;
        RECT 367.950 567.450 370.050 567.900 ;
        RECT 361.950 566.250 370.050 567.450 ;
        RECT 361.950 565.800 364.050 566.250 ;
        RECT 367.950 565.800 370.050 566.250 ;
        RECT 382.950 567.600 385.050 568.050 ;
        RECT 388.950 567.600 391.050 568.050 ;
        RECT 382.950 566.400 391.050 567.600 ;
        RECT 401.400 567.600 402.600 572.400 ;
        RECT 403.950 572.550 415.050 573.750 ;
        RECT 403.950 572.100 406.050 572.550 ;
        RECT 412.950 572.100 415.050 572.550 ;
        RECT 409.950 567.600 412.050 568.050 ;
        RECT 416.400 567.900 417.600 574.950 ;
        RECT 418.950 572.100 421.050 574.200 ;
        RECT 401.400 566.400 412.050 567.600 ;
        RECT 382.950 565.950 385.050 566.400 ;
        RECT 388.950 565.950 391.050 566.400 ;
        RECT 409.950 565.950 412.050 566.400 ;
        RECT 415.950 565.800 418.050 567.900 ;
        RECT 419.400 565.050 420.600 572.100 ;
        RECT 424.950 571.950 427.050 574.050 ;
        RECT 496.950 573.750 499.050 574.200 ;
        RECT 505.950 573.750 508.050 574.200 ;
        RECT 496.950 572.550 508.050 573.750 ;
        RECT 496.950 572.100 499.050 572.550 ;
        RECT 505.950 572.100 508.050 572.550 ;
        RECT 520.950 573.600 523.050 574.050 ;
        RECT 532.950 573.600 535.050 574.200 ;
        RECT 520.950 572.400 535.050 573.600 ;
        RECT 544.950 573.600 547.050 577.050 ;
        RECT 580.950 576.600 583.050 577.050 ;
        RECT 592.950 576.600 595.050 577.050 ;
        RECT 580.950 575.400 595.050 576.600 ;
        RECT 580.950 574.950 583.050 575.400 ;
        RECT 592.950 574.950 595.050 575.400 ;
        RECT 601.950 576.600 604.050 577.050 ;
        RECT 616.950 576.600 619.050 577.050 ;
        RECT 601.950 575.400 619.050 576.600 ;
        RECT 601.950 574.950 604.050 575.400 ;
        RECT 616.950 574.950 619.050 575.400 ;
        RECT 646.950 576.600 649.050 577.050 ;
        RECT 670.950 576.600 673.050 577.050 ;
        RECT 646.950 575.400 673.050 576.600 ;
        RECT 646.950 574.950 649.050 575.400 ;
        RECT 670.950 574.950 673.050 575.400 ;
        RECT 688.950 576.600 691.050 577.050 ;
        RECT 694.950 576.600 697.050 577.050 ;
        RECT 739.950 576.600 742.050 577.050 ;
        RECT 688.950 575.400 697.050 576.600 ;
        RECT 688.950 574.950 691.050 575.400 ;
        RECT 694.950 574.950 697.050 575.400 ;
        RECT 731.400 575.400 742.050 576.600 ;
        RECT 550.950 573.600 553.050 574.200 ;
        RECT 619.950 573.600 622.050 574.050 ;
        RECT 544.950 573.000 553.050 573.600 ;
        RECT 545.400 572.400 553.050 573.000 ;
        RECT 520.950 571.950 523.050 572.400 ;
        RECT 532.950 572.100 535.050 572.400 ;
        RECT 550.950 572.100 553.050 572.400 ;
        RECT 563.400 572.400 622.050 573.600 ;
        RECT 100.950 563.400 135.600 564.600 ;
        RECT 169.950 564.600 172.050 565.050 ;
        RECT 205.950 564.600 208.050 565.050 ;
        RECT 169.950 563.400 208.050 564.600 ;
        RECT 100.950 562.950 103.050 563.400 ;
        RECT 169.950 562.950 172.050 563.400 ;
        RECT 205.950 562.950 208.050 563.400 ;
        RECT 220.950 562.950 223.050 565.050 ;
        RECT 226.950 564.450 229.050 564.900 ;
        RECT 232.950 564.450 235.050 564.900 ;
        RECT 226.950 563.250 235.050 564.450 ;
        RECT 226.950 562.800 229.050 563.250 ;
        RECT 232.950 562.800 235.050 563.250 ;
        RECT 313.950 564.600 316.050 565.050 ;
        RECT 334.950 564.600 337.050 565.050 ;
        RECT 394.950 564.600 397.050 565.050 ;
        RECT 313.950 563.400 397.050 564.600 ;
        RECT 313.950 562.950 316.050 563.400 ;
        RECT 334.950 562.950 337.050 563.400 ;
        RECT 394.950 562.950 397.050 563.400 ;
        RECT 418.950 562.950 421.050 565.050 ;
        RECT 425.400 564.600 426.600 571.950 ;
        RECT 430.950 570.600 433.050 571.050 ;
        RECT 430.950 569.400 456.600 570.600 ;
        RECT 430.950 568.950 433.050 569.400 ;
        RECT 455.400 565.050 456.600 569.400 ;
        RECT 478.950 569.100 481.050 571.200 ;
        RECT 563.400 571.050 564.600 572.400 ;
        RECT 619.950 571.950 622.050 572.400 ;
        RECT 625.950 571.950 628.050 574.050 ;
        RECT 631.950 573.600 634.050 574.200 ;
        RECT 631.950 572.400 645.600 573.600 ;
        RECT 631.950 572.100 634.050 572.400 ;
        RECT 479.400 565.050 480.600 569.100 ;
        RECT 484.950 568.950 487.050 571.050 ;
        RECT 559.950 569.400 564.600 571.050 ;
        RECT 580.950 570.600 583.050 570.900 ;
        RECT 601.950 570.600 604.050 571.050 ;
        RECT 566.400 569.400 604.050 570.600 ;
        RECT 559.950 568.950 564.000 569.400 ;
        RECT 485.400 565.050 486.600 568.950 ;
        RECT 499.950 567.450 502.050 567.900 ;
        RECT 529.950 567.450 532.050 567.900 ;
        RECT 499.950 566.250 532.050 567.450 ;
        RECT 499.950 565.800 502.050 566.250 ;
        RECT 529.950 565.800 532.050 566.250 ;
        RECT 547.950 567.600 550.050 567.900 ;
        RECT 566.400 567.600 567.600 569.400 ;
        RECT 580.950 568.800 583.050 569.400 ;
        RECT 601.950 568.950 604.050 569.400 ;
        RECT 547.950 566.400 567.600 567.600 ;
        RECT 568.950 567.600 571.050 567.900 ;
        RECT 589.950 567.600 592.050 567.900 ;
        RECT 568.950 566.400 592.050 567.600 ;
        RECT 547.950 565.800 550.050 566.400 ;
        RECT 568.950 565.800 571.050 566.400 ;
        RECT 589.950 565.800 592.050 566.400 ;
        RECT 598.950 567.450 601.050 567.900 ;
        RECT 604.950 567.450 607.050 568.050 ;
        RECT 610.950 567.450 613.050 567.900 ;
        RECT 598.950 566.250 613.050 567.450 ;
        RECT 598.950 565.800 601.050 566.250 ;
        RECT 604.950 565.950 607.050 566.250 ;
        RECT 610.950 565.800 613.050 566.250 ;
        RECT 619.950 567.600 622.050 568.050 ;
        RECT 626.400 567.600 627.600 571.950 ;
        RECT 644.400 567.900 645.600 572.400 ;
        RECT 664.950 571.950 667.050 574.050 ;
        RECT 676.950 572.100 679.050 574.200 ;
        RECT 709.950 573.750 712.050 574.200 ;
        RECT 724.950 573.750 727.050 574.200 ;
        RECT 709.950 572.550 727.050 573.750 ;
        RECT 709.950 572.100 712.050 572.550 ;
        RECT 724.950 572.100 727.050 572.550 ;
        RECT 619.950 566.400 627.600 567.600 ;
        RECT 619.950 565.950 622.050 566.400 ;
        RECT 643.950 565.800 646.050 567.900 ;
        RECT 430.950 564.600 433.050 565.050 ;
        RECT 425.400 563.400 433.050 564.600 ;
        RECT 430.950 562.950 433.050 563.400 ;
        RECT 451.950 563.400 456.600 565.050 ;
        RECT 475.950 563.400 480.600 565.050 ;
        RECT 451.950 562.950 456.000 563.400 ;
        RECT 475.950 562.950 480.000 563.400 ;
        RECT 484.950 562.950 487.050 565.050 ;
        RECT 665.400 564.600 666.600 571.950 ;
        RECT 670.950 564.600 673.050 565.050 ;
        RECT 665.400 563.400 673.050 564.600 ;
        RECT 670.950 562.950 673.050 563.400 ;
        RECT 677.400 562.050 678.600 572.100 ;
        RECT 682.950 570.600 685.050 571.050 ;
        RECT 700.950 570.600 703.050 571.050 ;
        RECT 682.950 569.400 703.050 570.600 ;
        RECT 682.950 568.950 685.050 569.400 ;
        RECT 700.950 568.950 703.050 569.400 ;
        RECT 712.950 567.600 715.050 567.900 ;
        RECT 721.950 567.600 724.050 568.050 ;
        RECT 731.400 567.900 732.600 575.400 ;
        RECT 739.950 574.950 742.050 575.400 ;
        RECT 748.800 576.000 750.900 577.050 ;
        RECT 751.950 576.600 754.050 577.050 ;
        RECT 787.950 576.600 790.050 577.050 ;
        RECT 796.950 576.600 799.050 577.050 ;
        RECT 883.950 576.600 886.050 577.050 ;
        RECT 748.800 574.950 751.050 576.000 ;
        RECT 751.950 575.400 799.050 576.600 ;
        RECT 751.950 574.950 754.050 575.400 ;
        RECT 787.950 574.950 790.050 575.400 ;
        RECT 796.950 574.950 799.050 575.400 ;
        RECT 878.400 575.400 886.050 576.600 ;
        RECT 748.950 573.600 751.050 574.950 ;
        RECT 772.950 573.600 775.050 574.200 ;
        RECT 778.950 573.600 781.050 574.200 ;
        RECT 737.400 572.400 775.050 573.600 ;
        RECT 737.400 567.900 738.600 572.400 ;
        RECT 772.950 572.100 775.050 572.400 ;
        RECT 776.400 572.400 781.050 573.600 ;
        RECT 776.400 570.600 777.600 572.400 ;
        RECT 778.950 572.100 781.050 572.400 ;
        RECT 793.950 573.600 796.050 574.050 ;
        RECT 793.950 572.400 801.600 573.600 ;
        RECT 793.950 571.950 796.050 572.400 ;
        RECT 755.400 569.400 777.600 570.600 ;
        RECT 755.400 567.900 756.600 569.400 ;
        RECT 800.400 567.900 801.600 572.400 ;
        RECT 802.950 572.100 805.050 574.200 ;
        RECT 803.400 570.600 804.600 572.100 ;
        RECT 817.950 571.950 820.050 574.050 ;
        RECT 832.950 573.750 835.050 574.200 ;
        RECT 838.950 573.750 841.050 574.200 ;
        RECT 832.950 572.550 841.050 573.750 ;
        RECT 832.950 572.100 835.050 572.550 ;
        RECT 838.950 572.100 841.050 572.550 ;
        RECT 868.950 573.750 871.050 574.200 ;
        RECT 874.950 573.750 877.050 574.200 ;
        RECT 868.950 572.550 877.050 573.750 ;
        RECT 868.950 572.100 871.050 572.550 ;
        RECT 874.950 572.100 877.050 572.550 ;
        RECT 803.400 569.400 807.600 570.600 ;
        RECT 806.400 568.050 807.600 569.400 ;
        RECT 818.400 568.050 819.600 571.950 ;
        RECT 878.400 570.600 879.600 575.400 ;
        RECT 883.950 574.950 886.050 575.400 ;
        RECT 901.950 574.950 904.050 577.050 ;
        RECT 880.950 571.950 883.050 574.050 ;
        RECT 875.400 569.400 879.600 570.600 ;
        RECT 712.950 566.400 724.050 567.600 ;
        RECT 712.950 565.800 715.050 566.400 ;
        RECT 721.950 565.950 724.050 566.400 ;
        RECT 730.950 565.800 733.050 567.900 ;
        RECT 736.950 565.800 739.050 567.900 ;
        RECT 754.950 565.800 757.050 567.900 ;
        RECT 781.950 567.450 784.050 567.900 ;
        RECT 787.950 567.450 790.050 567.900 ;
        RECT 781.950 566.250 790.050 567.450 ;
        RECT 781.950 565.800 784.050 566.250 ;
        RECT 787.950 565.800 790.050 566.250 ;
        RECT 799.950 565.800 802.050 567.900 ;
        RECT 806.400 566.400 811.050 568.050 ;
        RECT 807.000 565.950 811.050 566.400 ;
        RECT 817.950 565.950 820.050 568.050 ;
        RECT 871.950 567.600 874.050 567.900 ;
        RECT 875.400 567.600 876.600 569.400 ;
        RECT 881.400 568.050 882.600 571.950 ;
        RECT 902.400 570.600 903.600 574.950 ;
        RECT 907.950 573.600 910.050 574.050 ;
        RECT 913.950 573.600 916.050 574.050 ;
        RECT 919.950 573.600 922.050 574.050 ;
        RECT 907.950 572.400 922.050 573.600 ;
        RECT 907.950 571.950 910.050 572.400 ;
        RECT 913.950 571.950 916.050 572.400 ;
        RECT 919.950 571.950 922.050 572.400 ;
        RECT 922.950 570.600 925.050 571.050 ;
        RECT 899.400 570.000 903.600 570.600 ;
        RECT 914.400 570.000 925.050 570.600 ;
        RECT 898.950 569.400 903.600 570.000 ;
        RECT 913.950 569.400 925.050 570.000 ;
        RECT 871.950 566.400 876.600 567.600 ;
        RECT 871.950 565.800 874.050 566.400 ;
        RECT 880.950 565.950 883.050 568.050 ;
        RECT 898.950 565.950 901.050 569.400 ;
        RECT 913.950 565.950 916.050 569.400 ;
        RECT 922.950 568.950 925.050 569.400 ;
        RECT 754.950 564.600 757.050 564.750 ;
        RECT 763.950 564.600 766.050 565.050 ;
        RECT 754.950 563.400 766.050 564.600 ;
        RECT 754.950 562.650 757.050 563.400 ;
        RECT 763.950 562.950 766.050 563.400 ;
        RECT 904.950 564.600 907.050 565.050 ;
        RECT 916.950 564.600 919.050 565.050 ;
        RECT 904.950 563.400 919.050 564.600 ;
        RECT 904.950 562.950 907.050 563.400 ;
        RECT 916.950 562.950 919.050 563.400 ;
        RECT 37.950 561.600 40.050 562.050 ;
        RECT 73.950 561.600 76.050 561.900 ;
        RECT 37.950 560.400 76.050 561.600 ;
        RECT 37.950 559.950 40.050 560.400 ;
        RECT 73.950 559.800 76.050 560.400 ;
        RECT 94.950 561.600 97.050 562.050 ;
        RECT 112.950 561.600 115.050 562.050 ;
        RECT 94.950 560.400 115.050 561.600 ;
        RECT 94.950 559.950 97.050 560.400 ;
        RECT 112.950 559.950 115.050 560.400 ;
        RECT 127.950 561.600 130.050 562.050 ;
        RECT 139.950 561.600 142.050 562.050 ;
        RECT 127.950 560.400 142.050 561.600 ;
        RECT 127.950 559.950 130.050 560.400 ;
        RECT 139.950 559.950 142.050 560.400 ;
        RECT 166.950 561.600 169.050 562.050 ;
        RECT 223.950 561.600 226.050 562.050 ;
        RECT 166.950 560.400 226.050 561.600 ;
        RECT 166.950 559.950 169.050 560.400 ;
        RECT 223.950 559.950 226.050 560.400 ;
        RECT 325.950 561.600 328.050 562.050 ;
        RECT 403.950 561.600 406.050 562.050 ;
        RECT 448.950 561.600 451.050 562.050 ;
        RECT 325.950 560.400 406.050 561.600 ;
        RECT 325.950 559.950 328.050 560.400 ;
        RECT 403.950 559.950 406.050 560.400 ;
        RECT 437.400 560.400 451.050 561.600 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 112.950 558.600 115.050 558.900 ;
        RECT 88.950 557.400 115.050 558.600 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 112.950 556.800 115.050 557.400 ;
        RECT 118.950 558.600 121.050 559.050 ;
        RECT 124.950 558.600 127.050 559.050 ;
        RECT 154.950 558.600 157.050 559.050 ;
        RECT 118.950 557.400 157.050 558.600 ;
        RECT 118.950 556.950 121.050 557.400 ;
        RECT 124.950 556.950 127.050 557.400 ;
        RECT 154.950 556.950 157.050 557.400 ;
        RECT 181.950 558.600 184.050 559.050 ;
        RECT 214.950 558.600 217.050 559.050 ;
        RECT 319.950 558.600 322.050 559.050 ;
        RECT 418.950 558.600 421.050 559.050 ;
        RECT 437.400 558.600 438.600 560.400 ;
        RECT 448.950 559.950 451.050 560.400 ;
        RECT 472.950 561.600 475.050 562.050 ;
        RECT 487.950 561.600 490.050 562.050 ;
        RECT 472.950 560.400 490.050 561.600 ;
        RECT 472.950 559.950 475.050 560.400 ;
        RECT 487.950 559.950 490.050 560.400 ;
        RECT 529.950 561.600 532.050 562.050 ;
        RECT 541.950 561.600 544.050 562.050 ;
        RECT 553.950 561.600 556.050 562.050 ;
        RECT 529.950 560.400 556.050 561.600 ;
        RECT 529.950 559.950 532.050 560.400 ;
        RECT 541.950 559.950 544.050 560.400 ;
        RECT 553.950 559.950 556.050 560.400 ;
        RECT 610.950 561.600 613.050 562.050 ;
        RECT 643.950 561.600 646.050 562.050 ;
        RECT 675.000 561.900 678.600 562.050 ;
        RECT 610.950 560.400 646.050 561.600 ;
        RECT 610.950 559.950 613.050 560.400 ;
        RECT 643.950 559.950 646.050 560.400 ;
        RECT 673.950 560.400 678.600 561.900 ;
        RECT 844.950 561.600 847.050 562.050 ;
        RECT 877.950 561.600 880.050 562.050 ;
        RECT 844.950 560.400 880.050 561.600 ;
        RECT 673.950 559.950 678.000 560.400 ;
        RECT 844.950 559.950 847.050 560.400 ;
        RECT 877.950 559.950 880.050 560.400 ;
        RECT 673.950 559.800 676.050 559.950 ;
        RECT 181.950 557.400 217.050 558.600 ;
        RECT 181.950 556.950 184.050 557.400 ;
        RECT 214.950 556.950 217.050 557.400 ;
        RECT 239.400 557.400 312.600 558.600 ;
        RECT 25.950 555.600 28.050 556.050 ;
        RECT 67.950 555.600 70.050 556.050 ;
        RECT 25.950 554.400 70.050 555.600 ;
        RECT 25.950 553.950 28.050 554.400 ;
        RECT 67.950 553.950 70.050 554.400 ;
        RECT 97.950 555.600 100.050 556.050 ;
        RECT 136.950 555.600 139.050 556.050 ;
        RECT 97.950 554.400 139.050 555.600 ;
        RECT 97.950 553.950 100.050 554.400 ;
        RECT 136.950 553.950 139.050 554.400 ;
        RECT 217.950 555.600 220.050 556.050 ;
        RECT 235.950 555.600 238.050 556.050 ;
        RECT 239.400 555.600 240.600 557.400 ;
        RECT 217.950 554.400 240.600 555.600 ;
        RECT 311.400 555.600 312.600 557.400 ;
        RECT 319.950 557.400 417.600 558.600 ;
        RECT 319.950 556.950 322.050 557.400 ;
        RECT 340.950 555.600 343.050 556.050 ;
        RECT 311.400 554.400 343.050 555.600 ;
        RECT 217.950 553.950 220.050 554.400 ;
        RECT 235.950 553.950 238.050 554.400 ;
        RECT 340.950 553.950 343.050 554.400 ;
        RECT 346.950 555.600 349.050 556.050 ;
        RECT 379.950 555.600 382.050 556.050 ;
        RECT 346.950 554.400 382.050 555.600 ;
        RECT 416.400 555.600 417.600 557.400 ;
        RECT 418.950 557.400 438.600 558.600 ;
        RECT 502.950 558.600 505.050 559.050 ;
        RECT 568.950 558.600 571.050 559.050 ;
        RECT 502.950 557.400 571.050 558.600 ;
        RECT 418.950 556.950 421.050 557.400 ;
        RECT 502.950 556.950 505.050 557.400 ;
        RECT 568.950 556.950 571.050 557.400 ;
        RECT 580.950 558.600 583.050 559.050 ;
        RECT 592.950 558.600 595.050 559.050 ;
        RECT 580.950 557.400 595.050 558.600 ;
        RECT 580.950 556.950 583.050 557.400 ;
        RECT 592.950 556.950 595.050 557.400 ;
        RECT 646.950 558.600 649.050 559.050 ;
        RECT 661.950 558.600 664.050 559.050 ;
        RECT 667.950 558.600 670.050 559.050 ;
        RECT 646.950 557.400 670.050 558.600 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 661.950 556.950 664.050 557.400 ;
        RECT 667.950 556.950 670.050 557.400 ;
        RECT 724.950 558.600 727.050 559.050 ;
        RECT 814.950 558.600 817.050 559.050 ;
        RECT 898.950 558.600 901.050 559.050 ;
        RECT 928.950 558.600 931.050 559.050 ;
        RECT 724.950 557.400 813.600 558.600 ;
        RECT 724.950 556.950 727.050 557.400 ;
        RECT 427.950 555.600 430.050 556.050 ;
        RECT 416.400 554.400 430.050 555.600 ;
        RECT 346.950 553.950 349.050 554.400 ;
        RECT 379.950 553.950 382.050 554.400 ;
        RECT 427.950 553.950 430.050 554.400 ;
        RECT 490.950 555.600 493.050 556.050 ;
        RECT 532.950 555.600 535.050 556.050 ;
        RECT 490.950 554.400 535.050 555.600 ;
        RECT 490.950 553.950 493.050 554.400 ;
        RECT 532.950 553.950 535.050 554.400 ;
        RECT 568.950 555.600 571.050 555.900 ;
        RECT 622.950 555.600 625.050 556.050 ;
        RECT 727.950 555.600 730.050 556.050 ;
        RECT 568.950 554.400 625.050 555.600 ;
        RECT 568.950 553.800 571.050 554.400 ;
        RECT 622.950 553.950 625.050 554.400 ;
        RECT 629.400 554.400 730.050 555.600 ;
        RECT 629.400 553.050 630.600 554.400 ;
        RECT 727.950 553.950 730.050 554.400 ;
        RECT 769.950 555.600 772.050 556.050 ;
        RECT 778.950 555.600 781.050 556.050 ;
        RECT 769.950 554.400 781.050 555.600 ;
        RECT 812.400 555.600 813.600 557.400 ;
        RECT 814.950 557.400 931.050 558.600 ;
        RECT 814.950 556.950 817.050 557.400 ;
        RECT 898.950 556.950 901.050 557.400 ;
        RECT 928.950 556.950 931.050 557.400 ;
        RECT 844.800 555.600 846.900 556.050 ;
        RECT 812.400 554.400 846.900 555.600 ;
        RECT 769.950 553.950 772.050 554.400 ;
        RECT 778.950 553.950 781.050 554.400 ;
        RECT 844.800 553.950 846.900 554.400 ;
        RECT 847.950 555.600 850.050 556.050 ;
        RECT 856.950 555.600 859.050 556.050 ;
        RECT 886.950 555.600 889.050 556.050 ;
        RECT 847.950 554.400 889.050 555.600 ;
        RECT 847.950 553.950 850.050 554.400 ;
        RECT 856.950 553.950 859.050 554.400 ;
        RECT 886.950 553.950 889.050 554.400 ;
        RECT 70.950 552.600 73.050 553.050 ;
        RECT 88.950 552.600 91.050 553.050 ;
        RECT 70.950 551.400 91.050 552.600 ;
        RECT 70.950 550.950 73.050 551.400 ;
        RECT 88.950 550.950 91.050 551.400 ;
        RECT 100.950 552.600 103.050 553.050 ;
        RECT 148.950 552.600 151.050 553.050 ;
        RECT 100.950 551.400 151.050 552.600 ;
        RECT 100.950 550.950 103.050 551.400 ;
        RECT 148.950 550.950 151.050 551.400 ;
        RECT 205.950 552.600 208.050 553.050 ;
        RECT 232.950 552.600 235.050 553.050 ;
        RECT 205.950 551.400 235.050 552.600 ;
        RECT 205.950 550.950 208.050 551.400 ;
        RECT 232.950 550.950 235.050 551.400 ;
        RECT 253.950 552.600 256.050 553.050 ;
        RECT 295.950 552.600 298.050 553.050 ;
        RECT 253.950 551.400 298.050 552.600 ;
        RECT 253.950 550.950 256.050 551.400 ;
        RECT 295.950 550.950 298.050 551.400 ;
        RECT 307.950 552.600 310.050 553.050 ;
        RECT 367.950 552.600 370.050 553.050 ;
        RECT 307.950 551.400 370.050 552.600 ;
        RECT 307.950 550.950 310.050 551.400 ;
        RECT 367.950 550.950 370.050 551.400 ;
        RECT 409.950 552.600 412.050 553.050 ;
        RECT 421.950 552.600 424.050 553.050 ;
        RECT 409.950 551.400 424.050 552.600 ;
        RECT 409.950 550.950 412.050 551.400 ;
        RECT 421.950 550.950 424.050 551.400 ;
        RECT 433.950 552.600 436.050 553.050 ;
        RECT 493.950 552.600 496.050 553.050 ;
        RECT 433.950 551.400 496.050 552.600 ;
        RECT 433.950 550.950 436.050 551.400 ;
        RECT 493.950 550.950 496.050 551.400 ;
        RECT 571.950 552.600 574.050 553.050 ;
        RECT 619.950 552.600 622.050 553.050 ;
        RECT 571.950 551.400 622.050 552.600 ;
        RECT 571.950 550.950 574.050 551.400 ;
        RECT 619.950 550.950 622.050 551.400 ;
        RECT 625.950 551.400 630.600 553.050 ;
        RECT 694.950 552.600 697.050 553.050 ;
        RECT 715.950 552.600 718.050 553.050 ;
        RECT 694.950 551.400 718.050 552.600 ;
        RECT 625.950 550.950 630.000 551.400 ;
        RECT 694.950 550.950 697.050 551.400 ;
        RECT 715.950 550.950 718.050 551.400 ;
        RECT 748.950 552.600 751.050 553.050 ;
        RECT 775.950 552.600 778.050 553.050 ;
        RECT 748.950 551.400 778.050 552.600 ;
        RECT 748.950 550.950 751.050 551.400 ;
        RECT 775.950 550.950 778.050 551.400 ;
        RECT 805.950 552.600 808.050 553.050 ;
        RECT 826.950 552.600 829.050 553.050 ;
        RECT 805.950 551.400 829.050 552.600 ;
        RECT 805.950 550.950 808.050 551.400 ;
        RECT 826.950 550.950 829.050 551.400 ;
        RECT 910.950 552.600 913.050 553.050 ;
        RECT 934.950 552.600 937.050 553.050 ;
        RECT 910.950 551.400 937.050 552.600 ;
        RECT 910.950 550.950 913.050 551.400 ;
        RECT 934.950 550.950 937.050 551.400 ;
        RECT 13.950 549.600 16.050 550.050 ;
        RECT 19.950 549.600 22.050 550.050 ;
        RECT 13.950 548.400 22.050 549.600 ;
        RECT 13.950 547.950 16.050 548.400 ;
        RECT 19.950 547.950 22.050 548.400 ;
        RECT 106.950 549.600 109.050 550.050 ;
        RECT 142.950 549.600 145.050 550.050 ;
        RECT 169.950 549.600 172.050 550.050 ;
        RECT 106.950 548.400 135.600 549.600 ;
        RECT 106.950 547.950 109.050 548.400 ;
        RECT 28.950 546.600 31.050 547.050 ;
        RECT 43.800 546.600 45.900 547.050 ;
        RECT 28.950 545.400 45.900 546.600 ;
        RECT 28.950 544.950 31.050 545.400 ;
        RECT 43.800 544.950 45.900 545.400 ;
        RECT 46.950 546.600 49.050 547.050 ;
        RECT 58.950 546.600 61.050 547.050 ;
        RECT 46.950 545.400 61.050 546.600 ;
        RECT 46.950 544.950 49.050 545.400 ;
        RECT 58.950 544.950 61.050 545.400 ;
        RECT 64.950 546.600 67.050 547.050 ;
        RECT 91.950 546.600 94.050 547.050 ;
        RECT 64.950 545.400 94.050 546.600 ;
        RECT 64.950 544.950 67.050 545.400 ;
        RECT 91.950 544.950 94.050 545.400 ;
        RECT 112.950 546.600 115.050 547.050 ;
        RECT 130.950 546.600 133.050 547.050 ;
        RECT 112.950 545.400 133.050 546.600 ;
        RECT 134.400 546.600 135.600 548.400 ;
        RECT 142.950 548.400 172.050 549.600 ;
        RECT 142.950 547.950 145.050 548.400 ;
        RECT 169.950 547.950 172.050 548.400 ;
        RECT 208.950 549.600 211.050 550.050 ;
        RECT 214.950 549.600 217.050 550.050 ;
        RECT 208.950 548.400 217.050 549.600 ;
        RECT 208.950 547.950 211.050 548.400 ;
        RECT 214.950 547.950 217.050 548.400 ;
        RECT 220.950 549.600 223.050 550.050 ;
        RECT 238.950 549.600 241.050 550.050 ;
        RECT 220.950 548.400 241.050 549.600 ;
        RECT 220.950 547.950 223.050 548.400 ;
        RECT 238.950 547.950 241.050 548.400 ;
        RECT 301.950 549.600 304.050 550.050 ;
        RECT 355.800 549.600 357.900 550.050 ;
        RECT 301.950 548.400 357.900 549.600 ;
        RECT 301.950 547.950 304.050 548.400 ;
        RECT 355.800 547.950 357.900 548.400 ;
        RECT 358.950 549.600 361.050 550.050 ;
        RECT 364.950 549.600 367.050 550.050 ;
        RECT 358.950 548.400 367.050 549.600 ;
        RECT 358.950 547.950 361.050 548.400 ;
        RECT 364.950 547.950 367.050 548.400 ;
        RECT 448.950 549.600 451.050 550.050 ;
        RECT 484.950 549.600 487.050 550.050 ;
        RECT 448.950 548.400 487.050 549.600 ;
        RECT 448.950 547.950 451.050 548.400 ;
        RECT 484.950 547.950 487.050 548.400 ;
        RECT 508.950 549.600 511.050 550.050 ;
        RECT 559.950 549.600 562.050 550.050 ;
        RECT 508.950 548.400 562.050 549.600 ;
        RECT 508.950 547.950 511.050 548.400 ;
        RECT 559.950 547.950 562.050 548.400 ;
        RECT 565.950 549.600 568.050 550.050 ;
        RECT 676.950 549.600 679.050 550.050 ;
        RECT 724.950 549.600 727.050 550.050 ;
        RECT 565.950 548.400 576.600 549.600 ;
        RECT 565.950 547.950 568.050 548.400 ;
        RECT 151.950 546.600 154.050 547.050 ;
        RECT 134.400 545.400 154.050 546.600 ;
        RECT 112.950 544.950 115.050 545.400 ;
        RECT 130.950 544.950 133.050 545.400 ;
        RECT 151.950 544.950 154.050 545.400 ;
        RECT 175.950 546.600 178.050 547.050 ;
        RECT 190.950 546.600 193.050 547.050 ;
        RECT 175.950 545.400 193.050 546.600 ;
        RECT 175.950 544.950 178.050 545.400 ;
        RECT 190.950 544.950 193.050 545.400 ;
        RECT 220.950 546.600 223.050 546.900 ;
        RECT 241.950 546.600 244.050 547.050 ;
        RECT 388.950 546.600 391.050 547.050 ;
        RECT 436.950 546.600 439.050 547.050 ;
        RECT 220.950 545.400 439.050 546.600 ;
        RECT 220.950 544.800 223.050 545.400 ;
        RECT 241.950 544.950 244.050 545.400 ;
        RECT 388.950 544.950 391.050 545.400 ;
        RECT 436.950 544.950 439.050 545.400 ;
        RECT 454.950 546.600 457.050 547.050 ;
        RECT 475.950 546.600 478.050 547.050 ;
        RECT 454.950 545.400 478.050 546.600 ;
        RECT 454.950 544.950 457.050 545.400 ;
        RECT 475.950 544.950 478.050 545.400 ;
        RECT 481.950 546.600 484.050 547.050 ;
        RECT 520.950 546.600 523.050 547.050 ;
        RECT 550.950 546.600 553.050 547.050 ;
        RECT 481.950 545.400 507.600 546.600 ;
        RECT 481.950 544.950 484.050 545.400 ;
        RECT 506.400 544.050 507.600 545.400 ;
        RECT 520.950 545.400 553.050 546.600 ;
        RECT 575.400 546.600 576.600 548.400 ;
        RECT 676.950 548.400 727.050 549.600 ;
        RECT 676.950 547.950 679.050 548.400 ;
        RECT 724.950 547.950 727.050 548.400 ;
        RECT 784.950 549.600 787.050 550.050 ;
        RECT 817.950 549.600 820.050 550.050 ;
        RECT 784.950 548.400 820.050 549.600 ;
        RECT 784.950 547.950 787.050 548.400 ;
        RECT 817.950 547.950 820.050 548.400 ;
        RECT 829.950 549.600 832.050 550.050 ;
        RECT 871.950 549.600 874.050 550.050 ;
        RECT 829.950 548.400 874.050 549.600 ;
        RECT 829.950 547.950 832.050 548.400 ;
        RECT 871.950 547.950 874.050 548.400 ;
        RECT 883.950 549.600 886.050 550.050 ;
        RECT 892.950 549.600 895.050 550.050 ;
        RECT 883.950 548.400 895.050 549.600 ;
        RECT 883.950 547.950 886.050 548.400 ;
        RECT 892.950 547.950 895.050 548.400 ;
        RECT 613.950 546.600 616.050 547.050 ;
        RECT 575.400 545.400 616.050 546.600 ;
        RECT 520.950 544.950 523.050 545.400 ;
        RECT 550.950 544.950 553.050 545.400 ;
        RECT 613.950 544.950 616.050 545.400 ;
        RECT 832.950 546.600 835.050 547.050 ;
        RECT 850.950 546.600 853.050 547.050 ;
        RECT 877.950 546.600 880.050 547.050 ;
        RECT 895.950 546.600 898.050 547.050 ;
        RECT 832.950 545.400 898.050 546.600 ;
        RECT 832.950 544.950 835.050 545.400 ;
        RECT 850.950 544.950 853.050 545.400 ;
        RECT 877.950 544.950 880.050 545.400 ;
        RECT 895.950 544.950 898.050 545.400 ;
        RECT 13.950 543.600 16.050 544.050 ;
        RECT 97.950 543.600 100.050 544.050 ;
        RECT 13.950 542.400 100.050 543.600 ;
        RECT 13.950 541.950 16.050 542.400 ;
        RECT 97.950 541.950 100.050 542.400 ;
        RECT 136.950 543.600 139.050 544.050 ;
        RECT 217.950 543.600 220.050 544.050 ;
        RECT 136.950 542.400 220.050 543.600 ;
        RECT 136.950 541.950 139.050 542.400 ;
        RECT 217.950 541.950 220.050 542.400 ;
        RECT 223.950 543.600 226.050 544.050 ;
        RECT 271.950 543.600 274.050 544.050 ;
        RECT 223.950 542.400 274.050 543.600 ;
        RECT 223.950 541.950 226.050 542.400 ;
        RECT 271.950 541.950 274.050 542.400 ;
        RECT 337.950 543.600 340.050 544.050 ;
        RECT 343.950 543.600 346.050 544.050 ;
        RECT 337.950 542.400 346.050 543.600 ;
        RECT 337.950 541.950 340.050 542.400 ;
        RECT 343.950 541.950 346.050 542.400 ;
        RECT 361.950 543.600 364.050 544.050 ;
        RECT 409.950 543.600 412.050 544.050 ;
        RECT 433.950 543.600 436.050 544.050 ;
        RECT 496.950 543.600 499.050 544.050 ;
        RECT 361.950 542.400 412.050 543.600 ;
        RECT 361.950 541.950 364.050 542.400 ;
        RECT 409.950 541.950 412.050 542.400 ;
        RECT 425.400 542.400 436.050 543.600 ;
        RECT 88.950 540.600 91.050 541.050 ;
        RECT 127.950 540.600 130.050 541.050 ;
        RECT 88.950 539.400 130.050 540.600 ;
        RECT 88.950 538.950 91.050 539.400 ;
        RECT 127.950 538.950 130.050 539.400 ;
        RECT 163.950 540.600 166.050 541.050 ;
        RECT 199.950 540.600 202.050 541.050 ;
        RECT 163.950 539.400 202.050 540.600 ;
        RECT 163.950 538.950 166.050 539.400 ;
        RECT 199.950 538.950 202.050 539.400 ;
        RECT 367.950 540.600 370.050 541.050 ;
        RECT 425.400 540.600 426.600 542.400 ;
        RECT 433.950 541.950 436.050 542.400 ;
        RECT 473.400 542.400 499.050 543.600 ;
        RECT 367.950 539.400 426.600 540.600 ;
        RECT 451.950 540.600 454.050 541.050 ;
        RECT 473.400 540.600 474.600 542.400 ;
        RECT 496.950 541.950 499.050 542.400 ;
        RECT 505.950 543.600 508.050 544.050 ;
        RECT 511.950 543.600 514.050 544.050 ;
        RECT 505.950 542.400 514.050 543.600 ;
        RECT 505.950 541.950 508.050 542.400 ;
        RECT 511.950 541.950 514.050 542.400 ;
        RECT 628.950 543.600 631.050 544.050 ;
        RECT 694.950 543.600 697.050 544.050 ;
        RECT 628.950 542.400 697.050 543.600 ;
        RECT 628.950 541.950 631.050 542.400 ;
        RECT 694.950 541.950 697.050 542.400 ;
        RECT 700.950 543.600 703.050 544.050 ;
        RECT 835.950 543.600 838.050 544.050 ;
        RECT 700.950 542.400 838.050 543.600 ;
        RECT 700.950 541.950 703.050 542.400 ;
        RECT 835.950 541.950 838.050 542.400 ;
        RECT 451.950 539.400 474.600 540.600 ;
        RECT 475.950 540.600 478.050 541.050 ;
        RECT 508.950 540.600 511.050 541.050 ;
        RECT 475.950 539.400 511.050 540.600 ;
        RECT 367.950 538.950 370.050 539.400 ;
        RECT 451.950 538.950 454.050 539.400 ;
        RECT 475.950 538.950 478.050 539.400 ;
        RECT 508.950 538.950 511.050 539.400 ;
        RECT 532.950 540.600 535.050 541.050 ;
        RECT 565.950 540.600 568.050 541.050 ;
        RECT 532.950 539.400 568.050 540.600 ;
        RECT 532.950 538.950 535.050 539.400 ;
        RECT 565.950 538.950 568.050 539.400 ;
        RECT 619.950 540.600 622.050 541.050 ;
        RECT 658.950 540.600 661.050 541.050 ;
        RECT 619.950 539.400 661.050 540.600 ;
        RECT 619.950 538.950 622.050 539.400 ;
        RECT 658.950 538.950 661.050 539.400 ;
        RECT 703.950 540.600 706.050 541.050 ;
        RECT 751.950 540.600 754.050 541.050 ;
        RECT 703.950 539.400 754.050 540.600 ;
        RECT 703.950 538.950 706.050 539.400 ;
        RECT 751.950 538.950 754.050 539.400 ;
        RECT 766.950 540.600 769.050 541.050 ;
        RECT 823.950 540.600 826.050 541.050 ;
        RECT 766.950 539.400 826.050 540.600 ;
        RECT 766.950 538.950 769.050 539.400 ;
        RECT 823.950 538.950 826.050 539.400 ;
        RECT 865.950 540.600 868.050 541.050 ;
        RECT 883.950 540.600 886.050 541.050 ;
        RECT 865.950 539.400 886.050 540.600 ;
        RECT 865.950 538.950 868.050 539.400 ;
        RECT 883.950 538.950 886.050 539.400 ;
        RECT 82.950 537.600 85.050 538.050 ;
        RECT 106.950 537.600 109.050 538.050 ;
        RECT 82.950 536.400 109.050 537.600 ;
        RECT 82.950 535.950 85.050 536.400 ;
        RECT 106.950 535.950 109.050 536.400 ;
        RECT 118.950 537.600 121.050 538.050 ;
        RECT 145.950 537.600 148.050 538.050 ;
        RECT 118.950 536.400 148.050 537.600 ;
        RECT 118.950 535.950 121.050 536.400 ;
        RECT 145.950 535.950 148.050 536.400 ;
        RECT 238.950 537.600 241.050 538.050 ;
        RECT 280.950 537.600 283.050 538.050 ;
        RECT 238.950 536.400 283.050 537.600 ;
        RECT 238.950 535.950 241.050 536.400 ;
        RECT 280.950 535.950 283.050 536.400 ;
        RECT 406.950 537.600 409.050 538.050 ;
        RECT 418.950 537.600 421.050 538.050 ;
        RECT 436.800 537.600 438.900 538.050 ;
        RECT 406.950 536.400 438.900 537.600 ;
        RECT 406.950 535.950 409.050 536.400 ;
        RECT 418.950 535.950 421.050 536.400 ;
        RECT 436.800 535.950 438.900 536.400 ;
        RECT 439.950 537.600 442.050 538.050 ;
        RECT 490.800 537.600 492.900 538.050 ;
        RECT 495.000 537.600 499.050 538.050 ;
        RECT 499.950 537.600 502.050 538.050 ;
        RECT 439.950 536.400 492.900 537.600 ;
        RECT 494.400 536.400 502.050 537.600 ;
        RECT 439.950 535.950 442.050 536.400 ;
        RECT 490.800 535.950 492.900 536.400 ;
        RECT 495.000 535.950 499.050 536.400 ;
        RECT 499.950 535.950 502.050 536.400 ;
        RECT 601.950 537.600 604.050 538.050 ;
        RECT 700.950 537.600 703.050 538.050 ;
        RECT 601.950 536.400 703.050 537.600 ;
        RECT 601.950 535.950 604.050 536.400 ;
        RECT 700.950 535.950 703.050 536.400 ;
        RECT 727.950 537.600 730.050 538.050 ;
        RECT 784.950 537.600 787.050 538.050 ;
        RECT 727.950 536.400 787.050 537.600 ;
        RECT 727.950 535.950 730.050 536.400 ;
        RECT 784.950 535.950 787.050 536.400 ;
        RECT 7.950 534.600 10.050 535.050 ;
        RECT 127.950 534.600 130.050 535.050 ;
        RECT 187.950 534.600 190.050 535.050 ;
        RECT 217.950 534.600 220.050 535.050 ;
        RECT 268.950 534.600 271.050 535.050 ;
        RECT 7.950 533.400 48.600 534.600 ;
        RECT 7.950 532.950 10.050 533.400 ;
        RECT 1.800 529.950 3.900 532.050 ;
        RECT 4.950 530.100 7.050 532.200 ;
        RECT 47.400 532.050 48.600 533.400 ;
        RECT 127.950 533.400 220.050 534.600 ;
        RECT 127.950 532.950 130.050 533.400 ;
        RECT 187.950 532.950 190.050 533.400 ;
        RECT 217.950 532.950 220.050 533.400 ;
        RECT 242.400 533.400 271.050 534.600 ;
        RECT 47.400 530.400 52.050 532.050 ;
        RECT 2.400 526.050 3.600 529.950 ;
        RECT 5.400 526.050 6.600 530.100 ;
        RECT 48.000 529.950 52.050 530.400 ;
        RECT 61.950 529.950 64.050 532.050 ;
        RECT 103.950 531.600 106.050 532.050 ;
        RECT 127.950 531.600 130.050 531.900 ;
        RECT 103.950 530.400 130.050 531.600 ;
        RECT 103.950 529.950 106.050 530.400 ;
        RECT 62.400 526.050 63.600 529.950 ;
        RECT 127.950 529.800 130.050 530.400 ;
        RECT 157.950 531.600 160.050 532.050 ;
        RECT 178.950 531.600 181.050 532.050 ;
        RECT 157.950 530.400 181.050 531.600 ;
        RECT 157.950 529.950 160.050 530.400 ;
        RECT 178.950 529.950 181.050 530.400 ;
        RECT 190.950 529.950 193.050 532.050 ;
        RECT 242.400 531.600 243.600 533.400 ;
        RECT 268.950 532.950 271.050 533.400 ;
        RECT 277.950 534.600 280.050 535.050 ;
        RECT 361.950 534.600 364.050 535.050 ;
        RECT 277.950 533.400 364.050 534.600 ;
        RECT 277.950 532.950 280.050 533.400 ;
        RECT 361.950 532.950 364.050 533.400 ;
        RECT 409.950 534.600 412.050 535.050 ;
        RECT 598.950 534.600 601.050 535.050 ;
        RECT 409.950 533.400 601.050 534.600 ;
        RECT 409.950 532.950 412.050 533.400 ;
        RECT 598.950 532.950 601.050 533.400 ;
        RECT 628.950 534.600 631.050 535.050 ;
        RECT 646.950 534.600 649.050 535.050 ;
        RECT 628.950 533.400 649.050 534.600 ;
        RECT 628.950 532.950 631.050 533.400 ;
        RECT 646.950 532.950 649.050 533.400 ;
        RECT 655.950 534.600 658.050 535.050 ;
        RECT 718.950 534.600 721.050 535.050 ;
        RECT 655.950 533.400 721.050 534.600 ;
        RECT 655.950 532.950 658.050 533.400 ;
        RECT 718.950 532.950 721.050 533.400 ;
        RECT 847.950 534.600 850.050 535.050 ;
        RECT 853.950 534.600 856.050 535.050 ;
        RECT 847.950 533.400 856.050 534.600 ;
        RECT 847.950 532.950 850.050 533.400 ;
        RECT 853.950 532.950 856.050 533.400 ;
        RECT 898.950 534.600 901.050 535.050 ;
        RECT 922.950 534.600 925.050 535.050 ;
        RECT 898.950 533.400 925.050 534.600 ;
        RECT 898.950 532.950 901.050 533.400 ;
        RECT 922.950 532.950 925.050 533.400 ;
        RECT 224.400 530.400 243.600 531.600 ;
        RECT 244.950 531.600 247.050 532.050 ;
        RECT 262.950 531.600 265.050 532.050 ;
        RECT 244.950 530.400 265.050 531.600 ;
        RECT 67.950 528.600 70.050 529.050 ;
        RECT 79.950 528.600 82.050 529.200 ;
        RECT 67.950 527.400 82.050 528.600 ;
        RECT 67.950 526.950 70.050 527.400 ;
        RECT 79.950 527.100 82.050 527.400 ;
        RECT 85.950 528.600 88.050 529.200 ;
        RECT 97.950 528.600 100.050 529.050 ;
        RECT 109.950 528.600 112.050 529.200 ;
        RECT 85.950 527.400 100.050 528.600 ;
        RECT 85.950 527.100 88.050 527.400 ;
        RECT 97.950 526.950 100.050 527.400 ;
        RECT 101.400 527.400 112.050 528.600 ;
        RECT 1.950 523.950 4.050 526.050 ;
        RECT 5.400 524.400 10.050 526.050 ;
        RECT 6.000 523.950 10.050 524.400 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 55.950 522.600 58.050 523.050 ;
        RECT 64.950 522.600 67.050 523.050 ;
        RECT 55.950 521.400 67.050 522.600 ;
        RECT 55.950 520.950 58.050 521.400 ;
        RECT 64.950 520.950 67.050 521.400 ;
        RECT 70.950 522.600 73.050 523.050 ;
        RECT 82.950 522.600 85.050 522.900 ;
        RECT 70.950 521.400 85.050 522.600 ;
        RECT 70.950 520.950 73.050 521.400 ;
        RECT 82.950 520.800 85.050 521.400 ;
        RECT 88.950 522.600 91.050 522.900 ;
        RECT 101.400 522.600 102.600 527.400 ;
        RECT 109.950 527.100 112.050 527.400 ;
        RECT 133.950 528.600 136.050 529.200 ;
        RECT 142.950 528.750 145.050 529.200 ;
        RECT 151.950 528.750 154.050 529.200 ;
        RECT 142.950 528.600 154.050 528.750 ;
        RECT 160.950 528.600 163.050 529.050 ;
        RECT 133.950 527.550 154.050 528.600 ;
        RECT 133.950 527.400 145.050 527.550 ;
        RECT 133.950 527.100 136.050 527.400 ;
        RECT 142.950 527.100 145.050 527.400 ;
        RECT 151.950 527.100 154.050 527.550 ;
        RECT 155.400 527.400 163.050 528.600 ;
        RECT 155.400 525.600 156.600 527.400 ;
        RECT 160.950 526.950 163.050 527.400 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 116.400 525.000 156.600 525.600 ;
        RECT 88.950 521.400 102.600 522.600 ;
        RECT 115.950 524.400 156.600 525.000 ;
        RECT 88.950 520.800 91.050 521.400 ;
        RECT 115.950 520.950 118.050 524.400 ;
        RECT 182.400 523.050 183.600 526.950 ;
        RECT 121.950 522.600 124.050 523.050 ;
        RECT 148.950 522.600 151.050 522.900 ;
        RECT 121.950 521.400 151.050 522.600 ;
        RECT 121.950 520.950 124.050 521.400 ;
        RECT 148.950 520.800 151.050 521.400 ;
        RECT 163.950 522.450 166.050 523.050 ;
        RECT 172.950 522.450 175.050 522.900 ;
        RECT 163.950 521.250 175.050 522.450 ;
        RECT 163.950 520.950 166.050 521.250 ;
        RECT 172.950 520.800 175.050 521.250 ;
        RECT 181.950 520.950 184.050 523.050 ;
        RECT 191.400 522.900 192.600 529.950 ;
        RECT 193.950 527.100 196.050 529.200 ;
        RECT 194.400 523.050 195.600 527.100 ;
        RECT 202.950 526.950 205.050 529.050 ;
        RECT 208.950 528.600 211.050 529.200 ;
        RECT 224.400 528.600 225.600 530.400 ;
        RECT 244.950 529.950 247.050 530.400 ;
        RECT 262.950 529.950 265.050 530.400 ;
        RECT 295.950 531.750 298.050 532.200 ;
        RECT 313.800 531.750 315.900 532.200 ;
        RECT 295.950 530.550 315.900 531.750 ;
        RECT 295.950 530.100 298.050 530.550 ;
        RECT 313.800 530.100 315.900 530.550 ;
        RECT 400.950 531.600 403.050 532.050 ;
        RECT 421.950 531.600 424.050 532.050 ;
        RECT 439.950 531.600 442.050 532.050 ;
        RECT 400.950 530.400 442.050 531.600 ;
        RECT 400.950 529.950 403.050 530.400 ;
        RECT 421.950 529.950 424.050 530.400 ;
        RECT 439.950 529.950 442.050 530.400 ;
        RECT 505.950 530.100 508.050 532.200 ;
        RECT 811.950 532.050 814.050 532.200 ;
        RECT 574.950 531.600 577.050 532.050 ;
        RECT 583.950 531.600 586.050 532.050 ;
        RECT 625.950 531.600 628.050 532.050 ;
        RECT 574.950 530.400 586.050 531.600 ;
        RECT 208.950 527.400 225.600 528.600 ;
        RECT 226.950 528.600 229.050 529.200 ;
        RECT 232.950 528.600 235.050 529.050 ;
        RECT 256.950 528.600 259.050 529.050 ;
        RECT 226.950 527.400 231.600 528.600 ;
        RECT 208.950 527.100 211.050 527.400 ;
        RECT 203.400 523.050 204.600 526.950 ;
        RECT 190.950 520.800 193.050 522.900 ;
        RECT 194.400 521.400 199.050 523.050 ;
        RECT 195.000 520.950 199.050 521.400 ;
        RECT 202.950 520.950 205.050 523.050 ;
        RECT 221.400 522.600 222.600 527.400 ;
        RECT 226.950 527.100 229.050 527.400 ;
        RECT 230.400 525.600 231.600 527.400 ;
        RECT 232.950 527.400 259.050 528.600 ;
        RECT 232.950 526.950 235.050 527.400 ;
        RECT 256.950 526.950 259.050 527.400 ;
        RECT 271.950 528.600 274.050 529.050 ;
        RECT 283.950 528.600 286.050 529.200 ;
        RECT 292.950 528.600 295.050 529.050 ;
        RECT 397.950 528.600 400.050 529.200 ;
        RECT 271.950 527.400 295.050 528.600 ;
        RECT 311.400 528.000 400.050 528.600 ;
        RECT 271.950 526.950 274.050 527.400 ;
        RECT 283.950 527.100 286.050 527.400 ;
        RECT 292.950 526.950 295.050 527.400 ;
        RECT 310.950 527.400 400.050 528.000 ;
        RECT 230.400 525.000 234.600 525.600 ;
        RECT 230.400 524.400 235.050 525.000 ;
        RECT 223.950 522.600 226.050 522.900 ;
        RECT 221.400 521.400 226.050 522.600 ;
        RECT 223.950 520.800 226.050 521.400 ;
        RECT 232.950 520.950 235.050 524.400 ;
        RECT 310.950 523.950 313.050 527.400 ;
        RECT 397.950 527.100 400.050 527.400 ;
        RECT 442.950 528.750 445.050 529.200 ;
        RECT 466.950 528.750 469.050 529.200 ;
        RECT 442.950 527.550 469.050 528.750 ;
        RECT 442.950 527.100 445.050 527.550 ;
        RECT 466.950 527.100 469.050 527.550 ;
        RECT 484.950 528.750 487.050 529.200 ;
        RECT 493.950 528.750 496.050 529.200 ;
        RECT 484.950 527.550 496.050 528.750 ;
        RECT 484.950 527.100 487.050 527.550 ;
        RECT 493.950 527.100 496.050 527.550 ;
        RECT 403.950 525.600 406.050 526.050 ;
        RECT 403.950 524.400 423.600 525.600 ;
        RECT 403.950 523.950 406.050 524.400 ;
        RECT 265.950 522.600 268.050 522.900 ;
        RECT 289.950 522.600 292.050 522.900 ;
        RECT 307.950 522.600 310.050 522.900 ;
        RECT 265.950 521.400 310.050 522.600 ;
        RECT 422.400 522.600 423.600 524.400 ;
        RECT 506.400 523.050 507.600 530.100 ;
        RECT 574.950 529.950 577.050 530.400 ;
        RECT 583.950 529.950 586.050 530.400 ;
        RECT 587.400 530.400 628.050 531.600 ;
        RECT 529.950 528.600 532.050 529.050 ;
        RECT 550.950 528.600 553.050 529.050 ;
        RECT 571.950 528.600 574.050 529.050 ;
        RECT 529.950 527.400 553.050 528.600 ;
        RECT 554.400 528.000 574.050 528.600 ;
        RECT 529.950 526.950 532.050 527.400 ;
        RECT 550.950 526.950 553.050 527.400 ;
        RECT 553.950 527.400 574.050 528.000 ;
        RECT 553.950 523.950 556.050 527.400 ;
        RECT 571.950 526.950 574.050 527.400 ;
        RECT 577.950 528.600 580.050 529.050 ;
        RECT 587.400 528.600 588.600 530.400 ;
        RECT 625.950 529.950 628.050 530.400 ;
        RECT 652.950 531.600 655.050 532.050 ;
        RECT 691.950 531.600 694.050 532.050 ;
        RECT 652.950 530.400 694.050 531.600 ;
        RECT 652.950 529.950 655.050 530.400 ;
        RECT 691.950 529.950 694.050 530.400 ;
        RECT 733.950 531.600 736.050 532.050 ;
        RECT 757.950 531.600 760.050 532.050 ;
        RECT 733.950 530.400 760.050 531.600 ;
        RECT 733.950 529.950 736.050 530.400 ;
        RECT 757.950 529.950 760.050 530.400 ;
        RECT 766.950 531.600 769.050 532.050 ;
        RECT 790.950 531.600 793.050 532.050 ;
        RECT 802.950 531.600 805.050 532.050 ;
        RECT 810.000 531.600 814.050 532.050 ;
        RECT 871.800 531.600 873.900 532.050 ;
        RECT 766.950 530.400 805.050 531.600 ;
        RECT 766.950 529.950 769.050 530.400 ;
        RECT 790.950 529.950 793.050 530.400 ;
        RECT 802.950 529.950 805.050 530.400 ;
        RECT 809.400 530.100 814.050 531.600 ;
        RECT 860.400 530.400 873.900 531.600 ;
        RECT 809.400 529.950 813.000 530.100 ;
        RECT 577.950 527.400 588.600 528.600 ;
        RECT 631.950 528.750 634.050 529.200 ;
        RECT 640.950 528.750 643.050 529.200 ;
        RECT 631.950 527.550 643.050 528.750 ;
        RECT 577.950 526.950 580.050 527.400 ;
        RECT 631.950 527.100 634.050 527.550 ;
        RECT 640.950 527.100 643.050 527.550 ;
        RECT 664.950 528.600 667.050 529.200 ;
        RECT 679.950 528.600 682.050 529.050 ;
        RECT 693.000 528.600 697.050 529.050 ;
        RECT 664.950 527.400 682.050 528.600 ;
        RECT 664.950 527.100 667.050 527.400 ;
        RECT 439.950 522.600 442.050 522.900 ;
        RECT 496.950 522.600 499.050 522.900 ;
        RECT 422.400 521.400 442.050 522.600 ;
        RECT 265.950 520.800 268.050 521.400 ;
        RECT 289.950 520.800 292.050 521.400 ;
        RECT 307.950 520.800 310.050 521.400 ;
        RECT 439.950 520.800 442.050 521.400 ;
        RECT 485.400 521.400 499.050 522.600 ;
        RECT 506.400 521.400 511.050 523.050 ;
        RECT 118.950 519.600 121.050 520.050 ;
        RECT 160.950 519.600 163.050 520.050 ;
        RECT 118.950 518.400 163.050 519.600 ;
        RECT 118.950 517.950 121.050 518.400 ;
        RECT 160.950 517.950 163.050 518.400 ;
        RECT 199.950 519.600 202.050 520.050 ;
        RECT 208.950 519.600 211.050 520.050 ;
        RECT 229.950 519.600 232.050 520.050 ;
        RECT 241.950 519.600 244.050 520.050 ;
        RECT 199.950 518.400 244.050 519.600 ;
        RECT 199.950 517.950 202.050 518.400 ;
        RECT 208.950 517.950 211.050 518.400 ;
        RECT 229.950 517.950 232.050 518.400 ;
        RECT 241.950 517.950 244.050 518.400 ;
        RECT 361.950 519.600 364.050 520.050 ;
        RECT 418.950 519.600 421.050 520.050 ;
        RECT 361.950 518.400 421.050 519.600 ;
        RECT 361.950 517.950 364.050 518.400 ;
        RECT 418.950 517.950 421.050 518.400 ;
        RECT 427.950 519.600 430.050 520.050 ;
        RECT 433.950 519.600 436.050 520.050 ;
        RECT 427.950 518.400 436.050 519.600 ;
        RECT 427.950 517.950 430.050 518.400 ;
        RECT 433.950 517.950 436.050 518.400 ;
        RECT 466.950 519.600 469.050 520.050 ;
        RECT 485.400 519.600 486.600 521.400 ;
        RECT 496.950 520.800 499.050 521.400 ;
        RECT 507.000 520.950 511.050 521.400 ;
        RECT 571.950 522.450 574.050 522.900 ;
        RECT 580.950 522.450 583.050 522.900 ;
        RECT 613.950 522.600 616.050 523.050 ;
        RECT 571.950 521.250 583.050 522.450 ;
        RECT 571.950 520.800 574.050 521.250 ;
        RECT 580.950 520.800 583.050 521.250 ;
        RECT 590.400 521.400 616.050 522.600 ;
        RECT 590.400 520.050 591.600 521.400 ;
        RECT 613.950 520.950 616.050 521.400 ;
        RECT 643.950 522.600 646.050 522.900 ;
        RECT 658.950 522.600 661.050 523.050 ;
        RECT 643.950 521.400 661.050 522.600 ;
        RECT 665.400 522.600 666.600 527.100 ;
        RECT 679.950 526.950 682.050 527.400 ;
        RECT 692.400 526.950 697.050 528.600 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 712.950 528.600 715.050 529.200 ;
        RECT 739.800 528.600 741.900 529.200 ;
        RECT 712.950 527.400 741.900 528.600 ;
        RECT 712.950 527.100 715.050 527.400 ;
        RECT 739.800 527.100 741.900 527.400 ;
        RECT 742.950 528.750 745.050 529.200 ;
        RECT 787.950 528.750 790.050 529.200 ;
        RECT 742.950 527.550 790.050 528.750 ;
        RECT 742.950 527.100 745.050 527.550 ;
        RECT 787.950 527.100 790.050 527.550 ;
        RECT 793.950 527.100 796.050 529.200 ;
        RECT 798.000 528.600 802.050 529.050 ;
        RECT 679.950 522.600 682.050 523.050 ;
        RECT 665.400 521.400 682.050 522.600 ;
        RECT 643.950 520.800 646.050 521.400 ;
        RECT 658.950 520.950 661.050 521.400 ;
        RECT 679.950 520.950 682.050 521.400 ;
        RECT 688.950 522.600 691.050 522.900 ;
        RECT 692.400 522.600 693.600 526.950 ;
        RECT 704.400 523.050 705.600 526.950 ;
        RECT 721.950 525.600 724.050 526.050 ;
        RECT 754.950 525.600 757.050 526.050 ;
        RECT 721.950 524.400 735.600 525.600 ;
        RECT 721.950 523.950 724.050 524.400 ;
        RECT 688.950 521.400 693.600 522.600 ;
        RECT 688.950 520.800 691.050 521.400 ;
        RECT 703.950 520.950 706.050 523.050 ;
        RECT 709.950 522.600 712.050 522.900 ;
        RECT 718.950 522.600 721.050 523.050 ;
        RECT 709.950 521.400 721.050 522.600 ;
        RECT 709.950 520.800 712.050 521.400 ;
        RECT 718.950 520.950 721.050 521.400 ;
        RECT 734.400 520.050 735.600 524.400 ;
        RECT 754.950 524.400 777.600 525.600 ;
        RECT 754.950 523.950 757.050 524.400 ;
        RECT 763.950 522.450 766.050 522.900 ;
        RECT 769.950 522.450 772.050 522.900 ;
        RECT 763.950 521.250 772.050 522.450 ;
        RECT 776.400 522.600 777.600 524.400 ;
        RECT 790.950 522.600 793.050 522.900 ;
        RECT 776.400 521.400 793.050 522.600 ;
        RECT 763.950 520.800 766.050 521.250 ;
        RECT 769.950 520.800 772.050 521.250 ;
        RECT 790.950 520.800 793.050 521.400 ;
        RECT 466.950 518.400 486.600 519.600 ;
        RECT 559.950 519.600 562.050 520.050 ;
        RECT 577.950 519.600 580.050 520.050 ;
        RECT 559.950 518.400 580.050 519.600 ;
        RECT 466.950 517.950 469.050 518.400 ;
        RECT 559.950 517.950 562.050 518.400 ;
        RECT 577.950 517.950 580.050 518.400 ;
        RECT 586.950 518.400 591.600 520.050 ;
        RECT 595.950 519.600 598.050 520.050 ;
        RECT 601.950 519.600 604.050 520.050 ;
        RECT 595.950 518.400 604.050 519.600 ;
        RECT 586.950 517.950 591.000 518.400 ;
        RECT 595.950 517.950 598.050 518.400 ;
        RECT 601.950 517.950 604.050 518.400 ;
        RECT 661.950 519.600 664.050 520.050 ;
        RECT 673.950 519.600 676.050 520.050 ;
        RECT 661.950 518.400 676.050 519.600 ;
        RECT 661.950 517.950 664.050 518.400 ;
        RECT 673.950 517.950 676.050 518.400 ;
        RECT 733.950 517.950 736.050 520.050 ;
        RECT 745.950 519.600 748.050 520.050 ;
        RECT 772.950 519.600 775.050 520.050 ;
        RECT 745.950 518.400 775.050 519.600 ;
        RECT 745.950 517.950 748.050 518.400 ;
        RECT 772.950 517.950 775.050 518.400 ;
        RECT 61.950 516.600 64.050 517.050 ;
        RECT 70.950 516.600 73.050 517.050 ;
        RECT 61.950 515.400 73.050 516.600 ;
        RECT 61.950 514.950 64.050 515.400 ;
        RECT 70.950 514.950 73.050 515.400 ;
        RECT 97.950 516.600 100.050 517.050 ;
        RECT 109.950 516.600 112.050 517.050 ;
        RECT 97.950 515.400 112.050 516.600 ;
        RECT 97.950 514.950 100.050 515.400 ;
        RECT 109.950 514.950 112.050 515.400 ;
        RECT 124.950 516.600 127.050 517.050 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 124.950 515.400 133.050 516.600 ;
        RECT 124.950 514.950 127.050 515.400 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 136.950 516.600 139.050 517.050 ;
        RECT 154.950 516.600 157.050 517.050 ;
        RECT 136.950 515.400 157.050 516.600 ;
        RECT 136.950 514.950 139.050 515.400 ;
        RECT 154.950 514.950 157.050 515.400 ;
        RECT 220.950 516.600 223.050 517.050 ;
        RECT 226.950 516.600 229.050 517.050 ;
        RECT 220.950 515.400 229.050 516.600 ;
        RECT 220.950 514.950 223.050 515.400 ;
        RECT 226.950 514.950 229.050 515.400 ;
        RECT 253.950 516.600 256.050 517.050 ;
        RECT 271.950 516.600 274.050 517.050 ;
        RECT 253.950 515.400 274.050 516.600 ;
        RECT 253.950 514.950 256.050 515.400 ;
        RECT 271.950 514.950 274.050 515.400 ;
        RECT 280.950 516.600 283.050 517.050 ;
        RECT 415.950 516.600 418.050 517.050 ;
        RECT 280.950 515.400 418.050 516.600 ;
        RECT 280.950 514.950 283.050 515.400 ;
        RECT 415.950 514.950 418.050 515.400 ;
        RECT 487.950 516.600 490.050 517.050 ;
        RECT 496.950 516.600 499.050 517.050 ;
        RECT 487.950 515.400 499.050 516.600 ;
        RECT 487.950 514.950 490.050 515.400 ;
        RECT 496.950 514.950 499.050 515.400 ;
        RECT 595.950 516.600 598.050 516.900 ;
        RECT 616.950 516.600 619.050 517.050 ;
        RECT 595.950 515.400 619.050 516.600 ;
        RECT 110.400 513.600 111.600 514.950 ;
        RECT 595.950 514.800 598.050 515.400 ;
        RECT 616.950 514.950 619.050 515.400 ;
        RECT 700.950 516.600 703.050 517.050 ;
        RECT 709.950 516.600 712.050 517.050 ;
        RECT 700.950 515.400 712.050 516.600 ;
        RECT 700.950 514.950 703.050 515.400 ;
        RECT 709.950 514.950 712.050 515.400 ;
        RECT 769.950 516.600 772.050 517.050 ;
        RECT 794.400 516.600 795.600 527.100 ;
        RECT 797.400 526.950 802.050 528.600 ;
        RECT 797.400 519.600 798.600 526.950 ;
        RECT 809.400 523.050 810.600 529.950 ;
        RECT 811.950 526.950 814.050 529.050 ;
        RECT 826.950 526.950 829.050 529.050 ;
        RECT 835.950 528.750 838.050 529.200 ;
        RECT 841.950 528.750 844.050 529.050 ;
        RECT 844.950 528.750 847.050 529.200 ;
        RECT 835.950 527.550 847.050 528.750 ;
        RECT 835.950 527.100 838.050 527.550 ;
        RECT 841.950 526.950 844.050 527.550 ;
        RECT 844.950 527.100 847.050 527.550 ;
        RECT 805.950 521.400 810.600 523.050 ;
        RECT 805.950 520.950 810.000 521.400 ;
        RECT 812.400 519.600 813.600 526.950 ;
        RECT 814.950 522.600 817.050 522.900 ;
        RECT 827.400 522.600 828.600 526.950 ;
        RECT 814.950 521.400 828.600 522.600 ;
        RECT 850.950 522.600 853.050 523.050 ;
        RECT 860.400 522.600 861.600 530.400 ;
        RECT 871.800 529.950 873.900 530.400 ;
        RECT 874.950 531.600 877.050 532.050 ;
        RECT 883.950 531.600 886.050 532.050 ;
        RECT 874.950 530.400 886.050 531.600 ;
        RECT 874.950 529.950 877.050 530.400 ;
        RECT 883.950 529.950 886.050 530.400 ;
        RECT 862.950 528.600 865.050 529.200 ;
        RECT 883.950 528.600 886.050 529.200 ;
        RECT 862.950 527.400 886.050 528.600 ;
        RECT 862.950 527.100 865.050 527.400 ;
        RECT 883.950 527.100 886.050 527.400 ;
        RECT 904.950 528.750 907.050 529.200 ;
        RECT 910.950 528.750 913.050 528.900 ;
        RECT 904.950 527.550 913.050 528.750 ;
        RECT 904.950 527.100 907.050 527.550 ;
        RECT 910.950 526.800 913.050 527.550 ;
        RECT 916.950 525.600 919.050 529.050 ;
        RECT 928.950 527.100 931.050 529.200 ;
        RECT 850.950 521.400 861.600 522.600 ;
        RECT 878.400 525.000 919.050 525.600 ;
        RECT 878.400 524.400 918.600 525.000 ;
        RECT 814.950 520.800 817.050 521.400 ;
        RECT 850.950 520.950 853.050 521.400 ;
        RECT 797.400 518.400 813.600 519.600 ;
        RECT 826.950 519.600 829.050 520.050 ;
        RECT 832.950 519.600 835.050 520.050 ;
        RECT 826.950 518.400 835.050 519.600 ;
        RECT 826.950 517.950 829.050 518.400 ;
        RECT 832.950 517.950 835.050 518.400 ;
        RECT 862.950 519.600 865.050 520.050 ;
        RECT 878.400 519.600 879.600 524.400 ;
        RECT 880.950 522.450 883.050 522.900 ;
        RECT 889.950 522.450 892.050 522.900 ;
        RECT 880.950 521.250 892.050 522.450 ;
        RECT 880.950 520.800 883.050 521.250 ;
        RECT 889.950 520.800 892.050 521.250 ;
        RECT 929.400 520.050 930.600 527.100 ;
        RECT 862.950 518.400 879.600 519.600 ;
        RECT 862.950 517.950 865.050 518.400 ;
        RECT 928.950 517.950 931.050 520.050 ;
        RECT 808.950 516.600 811.050 517.050 ;
        RECT 769.950 515.400 811.050 516.600 ;
        RECT 769.950 514.950 772.050 515.400 ;
        RECT 808.950 514.950 811.050 515.400 ;
        RECT 859.950 516.600 862.050 517.050 ;
        RECT 868.950 516.600 871.050 517.050 ;
        RECT 919.950 516.600 922.050 517.050 ;
        RECT 859.950 515.400 922.050 516.600 ;
        RECT 859.950 514.950 862.050 515.400 ;
        RECT 868.950 514.950 871.050 515.400 ;
        RECT 919.950 514.950 922.050 515.400 ;
        RECT 166.950 513.600 169.050 514.050 ;
        RECT 110.400 512.400 169.050 513.600 ;
        RECT 166.950 511.950 169.050 512.400 ;
        RECT 178.950 513.600 181.050 514.050 ;
        RECT 199.950 513.600 202.050 514.050 ;
        RECT 247.950 513.600 250.050 514.050 ;
        RECT 367.950 513.600 370.050 514.050 ;
        RECT 178.950 512.400 250.050 513.600 ;
        RECT 178.950 511.950 181.050 512.400 ;
        RECT 199.950 511.950 202.050 512.400 ;
        RECT 247.950 511.950 250.050 512.400 ;
        RECT 362.400 512.400 370.050 513.600 ;
        RECT 13.950 510.600 16.050 511.050 ;
        RECT 19.950 510.600 22.050 511.050 ;
        RECT 13.950 509.400 22.050 510.600 ;
        RECT 13.950 508.950 16.050 509.400 ;
        RECT 19.950 508.950 22.050 509.400 ;
        RECT 28.950 510.600 31.050 511.050 ;
        RECT 58.950 510.600 61.050 511.050 ;
        RECT 28.950 509.400 61.050 510.600 ;
        RECT 28.950 508.950 31.050 509.400 ;
        RECT 58.950 508.950 61.050 509.400 ;
        RECT 64.950 510.600 67.050 511.050 ;
        RECT 76.950 510.600 79.050 511.050 ;
        RECT 64.950 509.400 79.050 510.600 ;
        RECT 64.950 508.950 67.050 509.400 ;
        RECT 76.950 508.950 79.050 509.400 ;
        RECT 88.950 510.600 91.050 511.050 ;
        RECT 205.950 510.600 208.050 511.050 ;
        RECT 88.950 509.400 208.050 510.600 ;
        RECT 88.950 508.950 91.050 509.400 ;
        RECT 205.950 508.950 208.050 509.400 ;
        RECT 349.950 510.600 352.050 511.050 ;
        RECT 362.400 510.600 363.600 512.400 ;
        RECT 367.950 511.950 370.050 512.400 ;
        RECT 373.950 513.600 376.050 514.050 ;
        RECT 388.950 513.600 391.050 514.050 ;
        RECT 373.950 512.400 391.050 513.600 ;
        RECT 373.950 511.950 376.050 512.400 ;
        RECT 388.950 511.950 391.050 512.400 ;
        RECT 412.950 513.600 415.050 514.050 ;
        RECT 475.950 513.600 478.050 514.050 ;
        RECT 412.950 512.400 478.050 513.600 ;
        RECT 412.950 511.950 415.050 512.400 ;
        RECT 475.950 511.950 478.050 512.400 ;
        RECT 568.950 513.600 571.050 514.050 ;
        RECT 580.950 513.600 583.050 514.050 ;
        RECT 607.950 513.600 610.050 514.050 ;
        RECT 625.950 513.600 628.050 514.050 ;
        RECT 568.950 512.400 610.050 513.600 ;
        RECT 568.950 511.950 571.050 512.400 ;
        RECT 580.950 511.950 583.050 512.400 ;
        RECT 607.950 511.950 610.050 512.400 ;
        RECT 620.400 512.400 628.050 513.600 ;
        RECT 349.950 509.400 363.600 510.600 ;
        RECT 418.950 510.600 421.050 511.050 ;
        RECT 454.950 510.600 457.050 511.050 ;
        RECT 418.950 509.400 457.050 510.600 ;
        RECT 349.950 508.950 352.050 509.400 ;
        RECT 418.950 508.950 421.050 509.400 ;
        RECT 454.950 508.950 457.050 509.400 ;
        RECT 484.950 510.600 487.050 511.050 ;
        RECT 535.950 510.600 538.050 511.050 ;
        RECT 559.950 510.600 562.050 511.050 ;
        RECT 484.950 509.400 562.050 510.600 ;
        RECT 484.950 508.950 487.050 509.400 ;
        RECT 535.950 508.950 538.050 509.400 ;
        RECT 559.950 508.950 562.050 509.400 ;
        RECT 577.950 510.600 580.050 511.050 ;
        RECT 592.950 510.600 595.050 511.050 ;
        RECT 620.400 510.600 621.600 512.400 ;
        RECT 625.950 511.950 628.050 512.400 ;
        RECT 676.950 513.600 679.050 514.050 ;
        RECT 682.950 513.600 685.050 514.050 ;
        RECT 676.950 512.400 685.050 513.600 ;
        RECT 676.950 511.950 679.050 512.400 ;
        RECT 682.950 511.950 685.050 512.400 ;
        RECT 703.950 513.600 706.050 514.050 ;
        RECT 715.950 513.600 718.050 514.050 ;
        RECT 703.950 512.400 718.050 513.600 ;
        RECT 703.950 511.950 706.050 512.400 ;
        RECT 715.950 511.950 718.050 512.400 ;
        RECT 814.950 513.600 817.050 514.050 ;
        RECT 844.950 513.600 847.050 514.050 ;
        RECT 895.950 513.600 898.050 514.050 ;
        RECT 814.950 512.400 828.600 513.600 ;
        RECT 814.950 511.950 817.050 512.400 ;
        RECT 577.950 509.400 621.600 510.600 ;
        RECT 622.950 510.600 625.050 511.050 ;
        RECT 631.950 510.600 634.050 511.050 ;
        RECT 655.800 510.600 657.900 511.050 ;
        RECT 622.950 509.400 634.050 510.600 ;
        RECT 577.950 508.950 580.050 509.400 ;
        RECT 592.950 508.950 595.050 509.400 ;
        RECT 622.950 508.950 625.050 509.400 ;
        RECT 631.950 508.950 634.050 509.400 ;
        RECT 635.400 509.400 657.900 510.600 ;
        RECT 49.950 507.600 52.050 508.050 ;
        RECT 14.400 506.400 52.050 507.600 ;
        RECT 14.400 505.050 15.600 506.400 ;
        RECT 49.950 505.950 52.050 506.400 ;
        RECT 124.950 507.600 127.050 508.050 ;
        RECT 139.800 507.600 141.900 508.050 ;
        RECT 124.950 506.400 141.900 507.600 ;
        RECT 124.950 505.950 127.050 506.400 ;
        RECT 139.800 505.950 141.900 506.400 ;
        RECT 142.950 507.600 145.050 508.050 ;
        RECT 169.950 507.600 172.050 508.050 ;
        RECT 142.950 506.400 172.050 507.600 ;
        RECT 142.950 505.950 145.050 506.400 ;
        RECT 169.950 505.950 172.050 506.400 ;
        RECT 298.950 507.600 301.050 508.050 ;
        RECT 304.950 507.600 307.050 508.050 ;
        RECT 364.950 507.600 367.050 508.050 ;
        RECT 298.950 506.400 367.050 507.600 ;
        RECT 298.950 505.950 301.050 506.400 ;
        RECT 304.950 505.950 307.050 506.400 ;
        RECT 364.950 505.950 367.050 506.400 ;
        RECT 427.950 507.600 430.050 508.050 ;
        RECT 451.950 507.600 454.050 508.050 ;
        RECT 427.950 506.400 454.050 507.600 ;
        RECT 427.950 505.950 430.050 506.400 ;
        RECT 451.950 505.950 454.050 506.400 ;
        RECT 457.950 507.600 460.050 508.050 ;
        RECT 463.950 507.600 466.050 508.050 ;
        RECT 457.950 506.400 466.050 507.600 ;
        RECT 457.950 505.950 460.050 506.400 ;
        RECT 463.950 505.950 466.050 506.400 ;
        RECT 529.950 507.600 532.050 508.050 ;
        RECT 574.950 507.600 577.050 508.050 ;
        RECT 529.950 506.400 577.050 507.600 ;
        RECT 529.950 505.950 532.050 506.400 ;
        RECT 574.950 505.950 577.050 506.400 ;
        RECT 598.950 507.600 601.050 508.050 ;
        RECT 635.400 507.600 636.600 509.400 ;
        RECT 655.800 508.950 657.900 509.400 ;
        RECT 658.950 510.600 661.050 511.050 ;
        RECT 691.950 510.600 694.050 511.050 ;
        RECT 697.950 510.600 700.050 511.050 ;
        RECT 658.950 509.400 690.600 510.600 ;
        RECT 658.950 508.950 661.050 509.400 ;
        RECT 598.950 506.400 636.600 507.600 ;
        RECT 649.950 507.600 652.050 508.050 ;
        RECT 689.400 507.600 690.600 509.400 ;
        RECT 691.950 509.400 700.050 510.600 ;
        RECT 691.950 508.950 694.050 509.400 ;
        RECT 697.950 508.950 700.050 509.400 ;
        RECT 745.950 510.600 748.050 511.050 ;
        RECT 760.950 510.600 763.050 511.050 ;
        RECT 745.950 509.400 763.050 510.600 ;
        RECT 827.400 510.600 828.600 512.400 ;
        RECT 844.950 512.400 898.050 513.600 ;
        RECT 844.950 511.950 847.050 512.400 ;
        RECT 895.950 511.950 898.050 512.400 ;
        RECT 916.950 513.600 919.050 514.050 ;
        RECT 925.950 513.600 928.050 514.050 ;
        RECT 916.950 512.400 928.050 513.600 ;
        RECT 916.950 511.950 919.050 512.400 ;
        RECT 925.950 511.950 928.050 512.400 ;
        RECT 853.950 510.600 856.050 511.050 ;
        RECT 827.400 509.400 856.050 510.600 ;
        RECT 745.950 508.950 748.050 509.400 ;
        RECT 760.950 508.950 763.050 509.400 ;
        RECT 853.950 508.950 856.050 509.400 ;
        RECT 901.950 510.600 904.050 511.050 ;
        RECT 928.950 510.600 931.050 511.050 ;
        RECT 901.950 509.400 931.050 510.600 ;
        RECT 901.950 508.950 904.050 509.400 ;
        RECT 928.950 508.950 931.050 509.400 ;
        RECT 694.950 507.600 697.050 508.050 ;
        RECT 649.950 506.400 672.600 507.600 ;
        RECT 689.400 506.400 697.050 507.600 ;
        RECT 598.950 505.950 601.050 506.400 ;
        RECT 649.950 505.950 652.050 506.400 ;
        RECT 10.950 503.400 15.600 505.050 ;
        RECT 94.950 504.600 97.050 505.050 ;
        RECT 106.950 504.600 109.050 505.050 ;
        RECT 94.950 503.400 109.050 504.600 ;
        RECT 10.950 502.950 15.000 503.400 ;
        RECT 94.950 502.950 97.050 503.400 ;
        RECT 106.950 502.950 109.050 503.400 ;
        RECT 172.950 504.600 175.050 505.050 ;
        RECT 229.950 504.600 232.050 505.050 ;
        RECT 172.950 503.400 232.050 504.600 ;
        RECT 172.950 502.950 175.050 503.400 ;
        RECT 229.950 502.950 232.050 503.400 ;
        RECT 307.950 504.600 310.050 505.050 ;
        RECT 412.950 504.600 415.050 505.050 ;
        RECT 307.950 503.400 415.050 504.600 ;
        RECT 307.950 502.950 310.050 503.400 ;
        RECT 412.950 502.950 415.050 503.400 ;
        RECT 433.950 504.600 436.050 505.050 ;
        RECT 439.950 504.600 442.050 505.050 ;
        RECT 433.950 503.400 442.050 504.600 ;
        RECT 433.950 502.950 436.050 503.400 ;
        RECT 439.950 502.950 442.050 503.400 ;
        RECT 574.950 504.600 577.050 504.900 ;
        RECT 580.950 504.600 583.050 505.050 ;
        RECT 574.950 503.400 583.050 504.600 ;
        RECT 574.950 502.800 577.050 503.400 ;
        RECT 580.950 502.950 583.050 503.400 ;
        RECT 586.950 504.600 589.050 505.050 ;
        RECT 592.950 504.600 595.050 505.050 ;
        RECT 586.950 503.400 595.050 504.600 ;
        RECT 586.950 502.950 589.050 503.400 ;
        RECT 592.950 502.950 595.050 503.400 ;
        RECT 652.950 504.600 655.050 505.050 ;
        RECT 667.950 504.600 670.050 505.050 ;
        RECT 652.950 503.400 670.050 504.600 ;
        RECT 671.400 504.600 672.600 506.400 ;
        RECT 694.950 505.950 697.050 506.400 ;
        RECT 730.950 507.600 733.050 508.050 ;
        RECT 739.950 507.600 742.050 508.050 ;
        RECT 796.950 507.600 799.050 508.050 ;
        RECT 730.950 506.400 742.050 507.600 ;
        RECT 730.950 505.950 733.050 506.400 ;
        RECT 739.950 505.950 742.050 506.400 ;
        RECT 758.400 506.400 799.050 507.600 ;
        RECT 697.950 504.600 700.050 505.050 ;
        RECT 671.400 503.400 700.050 504.600 ;
        RECT 652.950 502.950 655.050 503.400 ;
        RECT 667.950 502.950 670.050 503.400 ;
        RECT 697.950 502.950 700.050 503.400 ;
        RECT 703.950 504.600 706.050 505.050 ;
        RECT 721.950 504.600 724.050 505.050 ;
        RECT 703.950 503.400 724.050 504.600 ;
        RECT 703.950 502.950 706.050 503.400 ;
        RECT 721.950 502.950 724.050 503.400 ;
        RECT 727.950 504.600 730.050 505.050 ;
        RECT 758.400 504.600 759.600 506.400 ;
        RECT 796.950 505.950 799.050 506.400 ;
        RECT 823.950 507.600 826.050 508.050 ;
        RECT 859.950 507.600 862.050 508.050 ;
        RECT 823.950 506.400 862.050 507.600 ;
        RECT 823.950 505.950 826.050 506.400 ;
        RECT 859.950 505.950 862.050 506.400 ;
        RECT 910.950 507.600 913.050 508.050 ;
        RECT 922.950 507.600 925.050 508.050 ;
        RECT 910.950 506.400 925.050 507.600 ;
        RECT 910.950 505.950 913.050 506.400 ;
        RECT 922.950 505.950 925.050 506.400 ;
        RECT 805.950 504.600 808.050 505.050 ;
        RECT 727.950 503.400 759.600 504.600 ;
        RECT 761.400 503.400 808.050 504.600 ;
        RECT 727.950 502.950 730.050 503.400 ;
        RECT 761.400 502.050 762.600 503.400 ;
        RECT 805.950 502.950 808.050 503.400 ;
        RECT 826.950 504.600 829.050 505.050 ;
        RECT 868.950 504.600 871.050 505.050 ;
        RECT 826.950 503.400 871.050 504.600 ;
        RECT 826.950 502.950 829.050 503.400 ;
        RECT 868.950 502.950 871.050 503.400 ;
        RECT 886.950 504.600 889.050 505.050 ;
        RECT 901.950 504.600 904.050 505.050 ;
        RECT 886.950 503.400 904.050 504.600 ;
        RECT 886.950 502.950 889.050 503.400 ;
        RECT 901.950 502.950 904.050 503.400 ;
        RECT 175.950 501.600 178.050 502.050 ;
        RECT 181.950 501.600 184.050 502.050 ;
        RECT 277.950 501.600 280.050 502.050 ;
        RECT 175.950 500.400 184.050 501.600 ;
        RECT 175.950 499.950 178.050 500.400 ;
        RECT 181.950 499.950 184.050 500.400 ;
        RECT 236.400 500.400 280.050 501.600 ;
        RECT 112.950 498.600 115.050 499.050 ;
        RECT 172.950 498.600 175.050 499.050 ;
        RECT 112.950 497.400 175.050 498.600 ;
        RECT 112.950 496.950 115.050 497.400 ;
        RECT 172.950 496.950 175.050 497.400 ;
        RECT 196.950 498.600 199.050 499.050 ;
        RECT 236.400 498.600 237.600 500.400 ;
        RECT 277.950 499.950 280.050 500.400 ;
        RECT 322.950 501.600 325.050 502.050 ;
        RECT 343.950 501.600 346.050 502.050 ;
        RECT 322.950 500.400 346.050 501.600 ;
        RECT 322.950 499.950 325.050 500.400 ;
        RECT 343.950 499.950 346.050 500.400 ;
        RECT 367.950 501.600 370.050 502.050 ;
        RECT 403.950 501.600 406.050 502.050 ;
        RECT 367.950 500.400 406.050 501.600 ;
        RECT 367.950 499.950 370.050 500.400 ;
        RECT 403.950 499.950 406.050 500.400 ;
        RECT 415.950 501.600 418.050 502.050 ;
        RECT 427.950 501.600 430.050 502.050 ;
        RECT 415.950 500.400 430.050 501.600 ;
        RECT 415.950 499.950 418.050 500.400 ;
        RECT 427.950 499.950 430.050 500.400 ;
        RECT 433.950 501.600 436.050 501.900 ;
        RECT 460.950 501.600 463.050 502.050 ;
        RECT 433.950 500.400 463.050 501.600 ;
        RECT 433.950 499.800 436.050 500.400 ;
        RECT 460.950 499.950 463.050 500.400 ;
        RECT 589.950 501.600 592.050 502.050 ;
        RECT 664.950 501.600 667.050 502.050 ;
        RECT 760.950 501.600 763.050 502.050 ;
        RECT 589.950 500.400 763.050 501.600 ;
        RECT 589.950 499.950 592.050 500.400 ;
        RECT 664.950 499.950 667.050 500.400 ;
        RECT 760.950 499.950 763.050 500.400 ;
        RECT 811.950 501.600 814.050 502.050 ;
        RECT 832.950 501.600 835.050 502.050 ;
        RECT 850.800 501.600 852.900 502.050 ;
        RECT 811.950 500.400 852.900 501.600 ;
        RECT 811.950 499.950 814.050 500.400 ;
        RECT 832.950 499.950 835.050 500.400 ;
        RECT 850.800 499.950 852.900 500.400 ;
        RECT 853.950 501.600 856.050 502.050 ;
        RECT 865.950 501.600 868.050 502.050 ;
        RECT 853.950 500.400 868.050 501.600 ;
        RECT 853.950 499.950 856.050 500.400 ;
        RECT 865.950 499.950 868.050 500.400 ;
        RECT 934.950 501.600 939.000 502.050 ;
        RECT 934.950 499.950 939.600 501.600 ;
        RECT 523.950 498.600 526.050 499.050 ;
        RECT 196.950 497.400 237.600 498.600 ;
        RECT 497.400 497.400 526.050 498.600 ;
        RECT 196.950 496.950 199.050 497.400 ;
        RECT 4.950 495.600 7.050 496.050 ;
        RECT 19.950 495.600 22.050 496.200 ;
        RECT 4.950 494.400 22.050 495.600 ;
        RECT 4.950 493.950 7.050 494.400 ;
        RECT 19.950 494.100 22.050 494.400 ;
        RECT 28.950 492.600 31.050 493.050 ;
        RECT 46.800 492.600 48.900 493.050 ;
        RECT 28.950 491.400 48.900 492.600 ;
        RECT 28.950 490.950 31.050 491.400 ;
        RECT 46.800 490.950 48.900 491.400 ;
        RECT 49.950 492.600 52.050 492.900 ;
        RECT 70.950 492.600 73.050 496.050 ;
        RECT 88.950 495.750 91.050 496.200 ;
        RECT 103.950 495.750 106.050 496.200 ;
        RECT 88.950 494.550 106.050 495.750 ;
        RECT 114.000 495.600 118.050 496.050 ;
        RECT 88.950 494.100 91.050 494.550 ;
        RECT 103.950 494.100 106.050 494.550 ;
        RECT 49.950 492.000 73.050 492.600 ;
        RECT 113.400 493.950 118.050 495.600 ;
        RECT 124.950 495.600 129.000 496.050 ;
        RECT 187.950 495.600 192.000 496.050 ;
        RECT 124.950 493.950 129.600 495.600 ;
        RECT 187.950 493.950 192.600 495.600 ;
        RECT 49.950 491.400 72.600 492.000 ;
        RECT 49.950 490.800 52.050 491.400 ;
        RECT 113.400 487.050 114.600 493.950 ;
        RECT 128.400 492.600 129.600 493.950 ;
        RECT 139.950 492.600 142.050 492.900 ;
        RECT 128.400 491.400 142.050 492.600 ;
        RECT 139.950 490.800 142.050 491.400 ;
        RECT 166.950 491.100 169.050 493.200 ;
        RECT 175.950 491.100 178.050 493.200 ;
        RECT 124.950 489.600 127.050 490.050 ;
        RECT 167.400 489.600 168.600 491.100 ;
        RECT 176.400 489.600 177.600 491.100 ;
        RECT 124.950 488.400 168.600 489.600 ;
        RECT 173.400 489.000 177.600 489.600 ;
        RECT 172.950 488.400 177.600 489.000 ;
        RECT 124.950 487.950 127.050 488.400 ;
        RECT 7.950 486.600 10.050 487.050 ;
        RECT 13.950 486.600 16.050 487.050 ;
        RECT 34.950 486.600 37.050 487.050 ;
        RECT 82.950 486.600 85.050 487.050 ;
        RECT 7.950 485.400 85.050 486.600 ;
        RECT 7.950 484.950 10.050 485.400 ;
        RECT 13.950 484.950 16.050 485.400 ;
        RECT 34.950 484.950 37.050 485.400 ;
        RECT 82.950 484.950 85.050 485.400 ;
        RECT 112.950 484.950 115.050 487.050 ;
        RECT 172.950 484.950 175.050 488.400 ;
        RECT 191.400 487.050 192.600 493.950 ;
        RECT 226.950 492.600 229.050 496.050 ;
        RECT 244.950 495.600 247.050 496.200 ;
        RECT 262.950 495.600 265.050 496.200 ;
        RECT 221.400 492.000 229.050 492.600 ;
        RECT 236.400 494.400 247.050 495.600 ;
        RECT 221.400 491.400 228.600 492.000 ;
        RECT 196.950 489.600 199.050 489.900 ;
        RECT 221.400 489.600 222.600 491.400 ;
        RECT 236.400 490.050 237.600 494.400 ;
        RECT 244.950 494.100 247.050 494.400 ;
        RECT 248.400 494.400 265.050 495.600 ;
        RECT 196.950 488.400 222.600 489.600 ;
        RECT 223.950 489.450 226.050 489.900 ;
        RECT 229.950 489.450 232.050 489.900 ;
        RECT 196.950 487.800 199.050 488.400 ;
        RECT 223.950 488.250 232.050 489.450 ;
        RECT 223.950 487.800 226.050 488.250 ;
        RECT 229.950 487.800 232.050 488.250 ;
        RECT 235.950 487.950 238.050 490.050 ;
        RECT 248.400 489.900 249.600 494.400 ;
        RECT 262.950 494.100 265.050 494.400 ;
        RECT 364.950 495.750 367.050 496.200 ;
        RECT 376.950 495.750 379.050 496.200 ;
        RECT 364.950 494.550 379.050 495.750 ;
        RECT 364.950 494.100 367.050 494.550 ;
        RECT 376.950 494.100 379.050 494.550 ;
        RECT 382.950 495.600 385.050 496.050 ;
        RECT 403.950 495.600 406.050 496.050 ;
        RECT 382.950 494.400 406.050 495.600 ;
        RECT 382.950 493.950 385.050 494.400 ;
        RECT 403.950 493.950 406.050 494.400 ;
        RECT 412.950 495.600 415.050 496.200 ;
        RECT 424.950 495.600 427.050 496.050 ;
        RECT 412.950 494.400 427.050 495.600 ;
        RECT 412.950 494.100 415.050 494.400 ;
        RECT 424.950 493.950 427.050 494.400 ;
        RECT 292.950 492.600 295.050 493.050 ;
        RECT 260.400 491.400 295.050 492.600 ;
        RECT 260.400 489.900 261.600 491.400 ;
        RECT 292.950 490.950 295.050 491.400 ;
        RECT 247.950 487.800 250.050 489.900 ;
        RECT 259.950 487.800 262.050 489.900 ;
        RECT 283.950 489.600 286.050 489.900 ;
        RECT 295.950 489.600 298.050 490.050 ;
        RECT 283.950 488.400 298.050 489.600 ;
        RECT 283.950 487.800 286.050 488.400 ;
        RECT 295.950 487.950 298.050 488.400 ;
        RECT 355.950 489.600 358.050 489.900 ;
        RECT 361.950 489.600 364.050 490.050 ;
        RECT 457.950 489.600 460.050 493.050 ;
        RECT 481.950 492.600 484.050 492.900 ;
        RECT 497.400 492.600 498.600 497.400 ;
        RECT 523.950 496.950 526.050 497.400 ;
        RECT 628.950 498.600 631.050 499.050 ;
        RECT 634.950 498.600 637.050 499.050 ;
        RECT 685.950 498.600 688.050 499.050 ;
        RECT 628.950 497.400 688.050 498.600 ;
        RECT 628.950 496.950 631.050 497.400 ;
        RECT 634.950 496.950 637.050 497.400 ;
        RECT 685.950 496.950 688.050 497.400 ;
        RECT 724.950 498.600 727.050 499.050 ;
        RECT 736.950 498.600 739.050 499.050 ;
        RECT 724.950 497.400 739.050 498.600 ;
        RECT 724.950 496.950 727.050 497.400 ;
        RECT 736.950 496.950 739.050 497.400 ;
        RECT 751.950 498.600 754.050 499.050 ;
        RECT 757.950 498.600 760.050 499.050 ;
        RECT 751.950 497.400 760.050 498.600 ;
        RECT 751.950 496.950 754.050 497.400 ;
        RECT 757.950 496.950 760.050 497.400 ;
        RECT 781.950 498.600 784.050 499.050 ;
        RECT 793.950 498.600 796.050 499.050 ;
        RECT 781.950 497.400 796.050 498.600 ;
        RECT 781.950 496.950 784.050 497.400 ;
        RECT 793.950 496.950 796.050 497.400 ;
        RECT 547.950 495.600 550.050 496.200 ;
        RECT 481.950 491.400 498.600 492.600 ;
        RECT 521.400 494.400 550.050 495.600 ;
        RECT 481.950 490.800 484.050 491.400 ;
        RECT 521.400 489.900 522.600 494.400 ;
        RECT 547.950 494.100 550.050 494.400 ;
        RECT 562.950 495.600 565.050 496.200 ;
        RECT 568.950 495.600 571.050 496.050 ;
        RECT 562.950 494.400 571.050 495.600 ;
        RECT 562.950 494.100 565.050 494.400 ;
        RECT 568.950 493.950 571.050 494.400 ;
        RECT 577.950 495.600 580.050 496.050 ;
        RECT 586.950 495.600 589.050 496.200 ;
        RECT 577.950 494.400 589.050 495.600 ;
        RECT 577.950 493.950 580.050 494.400 ;
        RECT 586.950 494.100 589.050 494.400 ;
        RECT 604.950 495.600 607.050 496.200 ;
        RECT 619.950 495.600 622.050 496.050 ;
        RECT 604.950 494.400 622.050 495.600 ;
        RECT 604.950 494.100 607.050 494.400 ;
        RECT 619.950 493.950 622.050 494.400 ;
        RECT 625.950 495.600 628.050 496.050 ;
        RECT 658.950 495.600 661.050 496.050 ;
        RECT 625.950 494.400 661.050 495.600 ;
        RECT 625.950 493.950 628.050 494.400 ;
        RECT 658.950 493.950 661.050 494.400 ;
        RECT 670.950 495.750 673.050 496.200 ;
        RECT 703.950 495.750 706.050 496.200 ;
        RECT 670.950 494.550 706.050 495.750 ;
        RECT 670.950 494.100 673.050 494.550 ;
        RECT 569.400 490.050 570.600 493.950 ;
        RECT 355.950 488.400 364.050 489.600 ;
        RECT 355.950 487.800 358.050 488.400 ;
        RECT 361.950 487.950 364.050 488.400 ;
        RECT 455.400 489.000 460.050 489.600 ;
        RECT 455.400 488.400 459.600 489.000 ;
        RECT 191.400 485.400 196.050 487.050 ;
        RECT 192.000 484.950 196.050 485.400 ;
        RECT 199.950 486.600 202.050 487.050 ;
        RECT 205.950 486.600 208.050 487.050 ;
        RECT 217.950 486.600 220.050 487.050 ;
        RECT 199.950 485.400 220.050 486.600 ;
        RECT 199.950 484.950 202.050 485.400 ;
        RECT 205.950 484.950 208.050 485.400 ;
        RECT 217.950 484.950 220.050 485.400 ;
        RECT 241.950 486.600 244.050 487.050 ;
        RECT 259.950 486.600 262.050 487.050 ;
        RECT 241.950 485.400 262.050 486.600 ;
        RECT 241.950 484.950 244.050 485.400 ;
        RECT 259.950 484.950 262.050 485.400 ;
        RECT 298.950 486.600 301.050 487.050 ;
        RECT 304.950 486.600 307.050 487.050 ;
        RECT 298.950 485.400 307.050 486.600 ;
        RECT 298.950 484.950 301.050 485.400 ;
        RECT 304.950 484.950 307.050 485.400 ;
        RECT 343.950 486.600 346.050 487.050 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 409.950 486.600 412.050 487.050 ;
        RECT 343.950 485.400 412.050 486.600 ;
        RECT 343.950 484.950 346.050 485.400 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 409.950 484.950 412.050 485.400 ;
        RECT 424.950 486.600 427.050 487.050 ;
        RECT 455.400 486.600 456.600 488.400 ;
        RECT 520.950 487.800 523.050 489.900 ;
        RECT 526.950 489.600 529.050 489.900 ;
        RECT 544.950 489.600 547.050 489.900 ;
        RECT 526.950 488.400 547.050 489.600 ;
        RECT 526.950 487.800 529.050 488.400 ;
        RECT 544.950 487.800 547.050 488.400 ;
        RECT 568.950 487.950 571.050 490.050 ;
        RECT 580.950 487.800 583.050 489.900 ;
        RECT 595.950 489.600 598.050 490.050 ;
        RECT 695.400 489.900 696.600 494.550 ;
        RECT 703.950 494.100 706.050 494.550 ;
        RECT 709.950 495.600 712.050 496.200 ;
        RECT 733.950 495.600 736.050 496.050 ;
        RECT 709.950 494.400 714.600 495.600 ;
        RECT 709.950 494.100 712.050 494.400 ;
        RECT 713.400 490.050 714.600 494.400 ;
        RECT 733.950 494.400 741.600 495.600 ;
        RECT 733.950 493.950 736.050 494.400 ;
        RECT 740.400 490.050 741.600 494.400 ;
        RECT 745.950 494.100 748.050 496.200 ;
        RECT 760.950 495.600 765.000 496.050 ;
        RECT 766.950 495.750 769.050 496.200 ;
        RECT 775.950 495.750 778.050 496.200 ;
        RECT 616.950 489.600 619.050 489.900 ;
        RECT 595.950 489.450 619.050 489.600 ;
        RECT 646.950 489.450 649.050 489.900 ;
        RECT 595.950 488.400 649.050 489.450 ;
        RECT 595.950 487.950 598.050 488.400 ;
        RECT 616.950 488.250 649.050 488.400 ;
        RECT 616.950 487.800 619.050 488.250 ;
        RECT 646.950 487.800 649.050 488.250 ;
        RECT 658.950 489.450 661.050 489.900 ;
        RECT 667.950 489.450 670.050 489.900 ;
        RECT 658.950 488.250 670.050 489.450 ;
        RECT 658.950 487.800 661.050 488.250 ;
        RECT 667.950 487.800 670.050 488.250 ;
        RECT 694.950 487.800 697.050 489.900 ;
        RECT 712.950 487.950 715.050 490.050 ;
        RECT 730.950 489.450 733.050 489.900 ;
        RECT 736.800 489.450 738.900 489.900 ;
        RECT 730.950 488.250 738.900 489.450 ;
        RECT 730.950 487.800 733.050 488.250 ;
        RECT 736.800 487.800 738.900 488.250 ;
        RECT 739.950 487.950 742.050 490.050 ;
        RECT 746.400 489.600 747.600 494.100 ;
        RECT 760.950 493.950 765.600 495.600 ;
        RECT 766.950 494.550 778.050 495.750 ;
        RECT 766.950 494.100 769.050 494.550 ;
        RECT 775.950 494.100 778.050 494.550 ;
        RECT 784.950 495.600 787.050 496.200 ;
        RECT 826.950 495.600 829.050 496.050 ;
        RECT 838.950 495.600 841.050 496.200 ;
        RECT 843.000 495.600 847.050 496.050 ;
        RECT 849.000 495.600 853.050 496.050 ;
        RECT 784.950 495.000 801.600 495.600 ;
        RECT 784.950 494.400 802.050 495.000 ;
        RECT 784.950 494.100 787.050 494.400 ;
        RECT 754.950 489.600 757.050 490.050 ;
        RECT 764.400 489.900 765.600 493.950 ;
        RECT 799.950 490.800 802.050 494.400 ;
        RECT 826.950 494.400 841.050 495.600 ;
        RECT 826.950 493.950 829.050 494.400 ;
        RECT 838.950 494.100 841.050 494.400 ;
        RECT 842.400 493.950 847.050 495.600 ;
        RECT 848.400 493.950 853.050 495.600 ;
        RECT 856.950 494.100 859.050 496.200 ;
        RECT 868.950 495.600 871.050 496.050 ;
        RECT 874.950 495.600 877.050 496.050 ;
        RECT 868.950 494.400 877.050 495.600 ;
        RECT 842.400 492.600 843.600 493.950 ;
        RECT 836.400 491.400 843.600 492.600 ;
        RECT 746.400 488.400 757.050 489.600 ;
        RECT 754.950 487.950 757.050 488.400 ;
        RECT 763.950 489.600 766.050 489.900 ;
        RECT 772.950 489.600 775.050 490.050 ;
        RECT 836.400 489.900 837.600 491.400 ;
        RECT 848.400 490.050 849.600 493.950 ;
        RECT 763.950 488.400 775.050 489.600 ;
        RECT 763.950 487.800 766.050 488.400 ;
        RECT 772.950 487.950 775.050 488.400 ;
        RECT 787.950 489.600 790.050 489.900 ;
        RECT 796.950 489.600 799.050 489.900 ;
        RECT 787.950 489.450 799.050 489.600 ;
        RECT 802.950 489.450 805.050 489.900 ;
        RECT 787.950 488.400 805.050 489.450 ;
        RECT 787.950 487.800 790.050 488.400 ;
        RECT 796.950 488.250 805.050 488.400 ;
        RECT 796.950 487.800 799.050 488.250 ;
        RECT 802.950 487.800 805.050 488.250 ;
        RECT 835.950 487.800 838.050 489.900 ;
        RECT 844.950 488.400 849.600 490.050 ;
        RECT 844.950 487.950 849.000 488.400 ;
        RECT 424.950 485.400 456.600 486.600 ;
        RECT 505.950 486.450 508.050 486.900 ;
        RECT 511.950 486.450 514.050 486.900 ;
        RECT 581.400 486.600 582.600 487.800 ;
        RECT 857.400 487.050 858.600 494.100 ;
        RECT 868.950 493.950 871.050 494.400 ;
        RECT 874.950 493.950 877.050 494.400 ;
        RECT 880.950 494.100 883.050 496.200 ;
        RECT 907.950 495.600 910.050 496.200 ;
        RECT 919.950 495.750 922.050 496.200 ;
        RECT 934.950 495.750 937.050 496.200 ;
        RECT 919.950 495.600 937.050 495.750 ;
        RECT 907.950 494.550 937.050 495.600 ;
        RECT 907.950 494.400 922.050 494.550 ;
        RECT 907.950 494.100 910.050 494.400 ;
        RECT 919.950 494.100 922.050 494.400 ;
        RECT 934.950 494.100 937.050 494.550 ;
        RECT 859.950 489.600 862.050 489.900 ;
        RECT 881.400 489.600 882.600 494.100 ;
        RECT 938.400 492.600 939.600 499.950 ;
        RECT 932.400 492.000 939.600 492.600 ;
        RECT 859.950 488.400 882.600 489.600 ;
        RECT 931.950 491.400 939.600 492.000 ;
        RECT 859.950 487.800 862.050 488.400 ;
        RECT 931.950 487.950 934.050 491.400 ;
        RECT 424.950 484.950 427.050 485.400 ;
        RECT 505.950 485.250 514.050 486.450 ;
        RECT 83.400 483.600 84.600 484.950 ;
        RECT 505.950 484.800 508.050 485.250 ;
        RECT 511.950 484.800 514.050 485.250 ;
        RECT 578.400 485.400 582.600 486.600 ;
        RECT 586.950 486.600 589.050 487.050 ;
        RECT 592.950 486.600 595.050 487.050 ;
        RECT 586.950 485.400 595.050 486.600 ;
        RECT 115.950 483.600 118.050 484.050 ;
        RECT 496.950 483.600 499.050 484.050 ;
        RECT 541.950 483.600 544.050 484.050 ;
        RECT 83.400 482.400 118.050 483.600 ;
        RECT 115.950 481.950 118.050 482.400 ;
        RECT 341.400 482.400 544.050 483.600 ;
        RECT 97.950 480.600 100.050 481.050 ;
        RECT 265.950 480.600 268.050 481.050 ;
        RECT 341.400 480.600 342.600 482.400 ;
        RECT 496.950 481.950 499.050 482.400 ;
        RECT 541.950 481.950 544.050 482.400 ;
        RECT 550.950 483.600 553.050 484.050 ;
        RECT 578.400 483.600 579.600 485.400 ;
        RECT 586.950 484.950 589.050 485.400 ;
        RECT 592.950 484.950 595.050 485.400 ;
        RECT 679.950 486.600 682.050 487.050 ;
        RECT 703.950 486.600 706.050 487.050 ;
        RECT 679.950 485.400 706.050 486.600 ;
        RECT 679.950 484.950 682.050 485.400 ;
        RECT 703.950 484.950 706.050 485.400 ;
        RECT 823.950 486.600 826.050 487.050 ;
        RECT 823.950 485.400 834.600 486.600 ;
        RECT 823.950 484.950 826.050 485.400 ;
        RECT 550.950 482.400 579.600 483.600 ;
        RECT 589.950 483.600 592.050 484.050 ;
        RECT 613.950 483.600 616.050 484.050 ;
        RECT 622.950 483.600 625.050 484.050 ;
        RECT 589.950 482.400 625.050 483.600 ;
        RECT 550.950 481.950 553.050 482.400 ;
        RECT 589.950 481.950 592.050 482.400 ;
        RECT 613.950 481.950 616.050 482.400 ;
        RECT 622.950 481.950 625.050 482.400 ;
        RECT 682.950 483.600 685.050 484.050 ;
        RECT 700.950 483.600 703.050 484.050 ;
        RECT 724.950 483.600 727.050 484.050 ;
        RECT 682.950 482.400 727.050 483.600 ;
        RECT 682.950 481.950 685.050 482.400 ;
        RECT 700.950 481.950 703.050 482.400 ;
        RECT 724.950 481.950 727.050 482.400 ;
        RECT 763.950 483.600 766.050 483.900 ;
        RECT 775.950 483.600 778.050 484.050 ;
        RECT 763.950 482.400 778.050 483.600 ;
        RECT 833.400 483.600 834.600 485.400 ;
        RECT 856.950 484.950 859.050 487.050 ;
        RECT 841.950 483.600 844.050 484.050 ;
        RECT 833.400 482.400 844.050 483.600 ;
        RECT 763.950 481.800 766.050 482.400 ;
        RECT 775.950 481.950 778.050 482.400 ;
        RECT 841.950 481.950 844.050 482.400 ;
        RECT 904.950 483.600 907.050 483.900 ;
        RECT 934.950 483.600 937.050 484.050 ;
        RECT 904.950 482.400 937.050 483.600 ;
        RECT 904.950 481.800 907.050 482.400 ;
        RECT 934.950 481.950 937.050 482.400 ;
        RECT 97.950 479.400 114.600 480.600 ;
        RECT 97.950 478.950 100.050 479.400 ;
        RECT 73.950 477.600 76.050 478.050 ;
        RECT 79.950 477.600 82.050 478.050 ;
        RECT 73.950 476.400 82.050 477.600 ;
        RECT 113.400 477.600 114.600 479.400 ;
        RECT 265.950 479.400 342.600 480.600 ;
        RECT 397.950 480.600 400.050 481.050 ;
        RECT 415.950 480.600 418.050 481.050 ;
        RECT 436.950 480.600 439.050 481.050 ;
        RECT 397.950 479.400 439.050 480.600 ;
        RECT 265.950 478.950 268.050 479.400 ;
        RECT 397.950 478.950 400.050 479.400 ;
        RECT 415.950 478.950 418.050 479.400 ;
        RECT 436.950 478.950 439.050 479.400 ;
        RECT 547.950 480.600 550.050 481.050 ;
        RECT 652.950 480.600 655.050 481.050 ;
        RECT 547.950 479.400 655.050 480.600 ;
        RECT 547.950 478.950 550.050 479.400 ;
        RECT 652.950 478.950 655.050 479.400 ;
        RECT 781.950 480.600 784.050 481.050 ;
        RECT 820.950 480.600 823.050 481.050 ;
        RECT 781.950 479.400 823.050 480.600 ;
        RECT 781.950 478.950 784.050 479.400 ;
        RECT 820.950 478.950 823.050 479.400 ;
        RECT 859.950 480.600 862.050 481.050 ;
        RECT 895.950 480.600 898.050 481.050 ;
        RECT 859.950 479.400 898.050 480.600 ;
        RECT 859.950 478.950 862.050 479.400 ;
        RECT 895.950 478.950 898.050 479.400 ;
        RECT 139.950 477.600 142.050 478.050 ;
        RECT 113.400 476.400 142.050 477.600 ;
        RECT 73.950 475.950 76.050 476.400 ;
        RECT 79.950 475.950 82.050 476.400 ;
        RECT 139.950 475.950 142.050 476.400 ;
        RECT 172.950 477.600 175.050 478.050 ;
        RECT 199.950 477.600 202.050 478.050 ;
        RECT 172.950 476.400 202.050 477.600 ;
        RECT 172.950 475.950 175.050 476.400 ;
        RECT 199.950 475.950 202.050 476.400 ;
        RECT 334.950 477.600 337.050 478.050 ;
        RECT 358.950 477.600 361.050 478.050 ;
        RECT 334.950 476.400 361.050 477.600 ;
        RECT 334.950 475.950 337.050 476.400 ;
        RECT 358.950 475.950 361.050 476.400 ;
        RECT 379.950 477.600 382.050 478.050 ;
        RECT 433.800 477.600 435.900 478.050 ;
        RECT 379.950 476.400 435.900 477.600 ;
        RECT 437.400 477.600 438.600 478.950 ;
        RECT 526.950 477.600 529.050 478.050 ;
        RECT 437.400 476.400 529.050 477.600 ;
        RECT 379.950 475.950 382.050 476.400 ;
        RECT 433.800 475.950 435.900 476.400 ;
        RECT 526.950 475.950 529.050 476.400 ;
        RECT 565.950 477.600 568.050 478.050 ;
        RECT 607.950 477.600 610.050 478.050 ;
        RECT 565.950 476.400 610.050 477.600 ;
        RECT 565.950 475.950 568.050 476.400 ;
        RECT 607.950 475.950 610.050 476.400 ;
        RECT 667.950 477.600 670.050 478.050 ;
        RECT 712.950 477.600 715.050 478.050 ;
        RECT 742.950 477.600 745.050 478.050 ;
        RECT 769.950 477.600 772.050 478.050 ;
        RECT 667.950 476.400 711.600 477.600 ;
        RECT 667.950 475.950 670.050 476.400 ;
        RECT 142.950 474.600 145.050 475.050 ;
        RECT 169.950 474.600 172.050 475.050 ;
        RECT 142.950 473.400 172.050 474.600 ;
        RECT 142.950 472.950 145.050 473.400 ;
        RECT 169.950 472.950 172.050 473.400 ;
        RECT 181.950 474.600 184.050 475.050 ;
        RECT 187.950 474.600 190.050 475.050 ;
        RECT 181.950 473.400 190.050 474.600 ;
        RECT 181.950 472.950 184.050 473.400 ;
        RECT 187.950 472.950 190.050 473.400 ;
        RECT 394.950 474.600 397.050 475.050 ;
        RECT 400.950 474.600 403.050 475.050 ;
        RECT 394.950 473.400 403.050 474.600 ;
        RECT 394.950 472.950 397.050 473.400 ;
        RECT 400.950 472.950 403.050 473.400 ;
        RECT 451.950 474.600 454.050 475.050 ;
        RECT 514.950 474.600 517.050 475.050 ;
        RECT 577.950 474.600 580.050 475.050 ;
        RECT 451.950 473.400 517.050 474.600 ;
        RECT 451.950 472.950 454.050 473.400 ;
        RECT 514.950 472.950 517.050 473.400 ;
        RECT 539.400 473.400 580.050 474.600 ;
        RECT 115.950 471.600 118.050 472.050 ;
        RECT 133.950 471.600 136.050 472.050 ;
        RECT 115.950 470.400 136.050 471.600 ;
        RECT 115.950 469.950 118.050 470.400 ;
        RECT 133.950 469.950 136.050 470.400 ;
        RECT 271.950 471.600 274.050 472.050 ;
        RECT 283.950 471.600 286.050 472.050 ;
        RECT 271.950 470.400 286.050 471.600 ;
        RECT 271.950 469.950 274.050 470.400 ;
        RECT 283.950 469.950 286.050 470.400 ;
        RECT 388.950 471.600 391.050 472.050 ;
        RECT 539.400 471.600 540.600 473.400 ;
        RECT 577.950 472.950 580.050 473.400 ;
        RECT 613.950 474.600 616.050 475.050 ;
        RECT 658.950 474.600 661.050 475.050 ;
        RECT 679.950 474.600 682.050 475.050 ;
        RECT 613.950 473.400 682.050 474.600 ;
        RECT 710.400 474.600 711.600 476.400 ;
        RECT 712.950 476.400 772.050 477.600 ;
        RECT 712.950 475.950 715.050 476.400 ;
        RECT 742.950 475.950 745.050 476.400 ;
        RECT 769.950 475.950 772.050 476.400 ;
        RECT 826.950 477.600 829.050 478.050 ;
        RECT 871.950 477.600 874.050 478.050 ;
        RECT 826.950 476.400 874.050 477.600 ;
        RECT 826.950 475.950 829.050 476.400 ;
        RECT 871.950 475.950 874.050 476.400 ;
        RECT 883.950 477.600 886.050 478.050 ;
        RECT 928.950 477.600 931.050 478.050 ;
        RECT 883.950 476.400 931.050 477.600 ;
        RECT 883.950 475.950 886.050 476.400 ;
        RECT 928.950 475.950 931.050 476.400 ;
        RECT 781.950 474.600 784.050 475.050 ;
        RECT 820.950 474.600 823.050 475.050 ;
        RECT 710.400 473.400 784.050 474.600 ;
        RECT 613.950 472.950 616.050 473.400 ;
        RECT 658.950 472.950 661.050 473.400 ;
        RECT 679.950 472.950 682.050 473.400 ;
        RECT 781.950 472.950 784.050 473.400 ;
        RECT 788.400 473.400 823.050 474.600 ;
        RECT 649.950 471.600 652.050 472.050 ;
        RECT 688.950 471.600 691.050 472.050 ;
        RECT 694.950 471.600 697.050 472.050 ;
        RECT 388.950 470.400 540.600 471.600 ;
        RECT 617.400 470.400 652.050 471.600 ;
        RECT 388.950 469.950 391.050 470.400 ;
        RECT 37.950 468.600 40.050 469.050 ;
        RECT 49.950 468.600 52.050 469.050 ;
        RECT 37.950 467.400 52.050 468.600 ;
        RECT 37.950 466.950 40.050 467.400 ;
        RECT 49.950 466.950 52.050 467.400 ;
        RECT 73.950 468.600 76.050 469.050 ;
        RECT 124.950 468.600 127.050 469.050 ;
        RECT 73.950 467.400 127.050 468.600 ;
        RECT 73.950 466.950 76.050 467.400 ;
        RECT 124.950 466.950 127.050 467.400 ;
        RECT 136.950 468.600 139.050 469.050 ;
        RECT 211.950 468.600 214.050 469.050 ;
        RECT 136.950 467.400 214.050 468.600 ;
        RECT 136.950 466.950 139.050 467.400 ;
        RECT 211.950 466.950 214.050 467.400 ;
        RECT 217.950 468.600 220.050 469.050 ;
        RECT 265.950 468.600 268.050 469.050 ;
        RECT 217.950 467.400 268.050 468.600 ;
        RECT 217.950 466.950 220.050 467.400 ;
        RECT 265.950 466.950 268.050 467.400 ;
        RECT 310.950 468.600 313.050 469.050 ;
        RECT 316.950 468.600 319.050 469.050 ;
        RECT 310.950 467.400 319.050 468.600 ;
        RECT 310.950 466.950 313.050 467.400 ;
        RECT 316.950 466.950 319.050 467.400 ;
        RECT 349.950 468.600 352.050 469.050 ;
        RECT 421.950 468.600 424.050 469.050 ;
        RECT 442.950 468.600 445.050 469.050 ;
        RECT 349.950 467.400 372.600 468.600 ;
        RECT 349.950 466.950 352.050 467.400 ;
        RECT 100.950 465.600 103.050 466.050 ;
        RECT 106.950 465.600 109.050 466.050 ;
        RECT 100.950 464.400 109.050 465.600 ;
        RECT 100.950 463.950 103.050 464.400 ;
        RECT 106.950 463.950 109.050 464.400 ;
        RECT 181.950 465.600 184.050 466.050 ;
        RECT 193.950 465.600 196.050 466.050 ;
        RECT 181.950 464.400 196.050 465.600 ;
        RECT 181.950 463.950 184.050 464.400 ;
        RECT 193.950 463.950 196.050 464.400 ;
        RECT 232.950 465.600 235.050 466.050 ;
        RECT 238.950 465.600 241.050 466.050 ;
        RECT 232.950 464.400 241.050 465.600 ;
        RECT 232.950 463.950 235.050 464.400 ;
        RECT 238.950 463.950 241.050 464.400 ;
        RECT 253.950 465.600 256.050 466.050 ;
        RECT 259.950 465.600 262.050 466.050 ;
        RECT 253.950 464.400 262.050 465.600 ;
        RECT 371.400 465.600 372.600 467.400 ;
        RECT 421.950 467.400 445.050 468.600 ;
        RECT 421.950 466.950 424.050 467.400 ;
        RECT 442.950 466.950 445.050 467.400 ;
        RECT 478.950 468.600 481.050 469.050 ;
        RECT 532.950 468.600 535.050 469.050 ;
        RECT 571.950 468.600 574.050 469.050 ;
        RECT 478.950 467.400 535.050 468.600 ;
        RECT 478.950 466.950 481.050 467.400 ;
        RECT 532.950 466.950 535.050 467.400 ;
        RECT 539.400 467.400 574.050 468.600 ;
        RECT 539.400 466.050 540.600 467.400 ;
        RECT 571.950 466.950 574.050 467.400 ;
        RECT 577.950 468.600 580.050 469.050 ;
        RECT 617.400 468.600 618.600 470.400 ;
        RECT 649.950 469.950 652.050 470.400 ;
        RECT 677.400 470.400 697.050 471.600 ;
        RECT 577.950 467.400 618.600 468.600 ;
        RECT 619.950 468.600 622.050 469.050 ;
        RECT 677.400 468.600 678.600 470.400 ;
        RECT 688.950 469.950 691.050 470.400 ;
        RECT 694.950 469.950 697.050 470.400 ;
        RECT 715.950 471.600 718.050 472.050 ;
        RECT 745.950 471.600 748.050 472.050 ;
        RECT 715.950 470.400 748.050 471.600 ;
        RECT 715.950 469.950 718.050 470.400 ;
        RECT 745.950 469.950 748.050 470.400 ;
        RECT 766.950 471.600 769.050 472.050 ;
        RECT 788.400 471.600 789.600 473.400 ;
        RECT 820.950 472.950 823.050 473.400 ;
        RECT 847.950 474.600 850.050 475.050 ;
        RECT 868.950 474.600 871.050 475.050 ;
        RECT 847.950 473.400 871.050 474.600 ;
        RECT 847.950 472.950 850.050 473.400 ;
        RECT 868.950 472.950 871.050 473.400 ;
        RECT 766.950 470.400 789.600 471.600 ;
        RECT 811.950 471.600 814.050 472.050 ;
        RECT 883.950 471.600 886.050 472.050 ;
        RECT 811.950 470.400 886.050 471.600 ;
        RECT 766.950 469.950 769.050 470.400 ;
        RECT 811.950 469.950 814.050 470.400 ;
        RECT 883.950 469.950 886.050 470.400 ;
        RECT 619.950 467.400 678.600 468.600 ;
        RECT 679.950 468.600 682.050 469.050 ;
        RECT 757.800 468.600 759.900 469.050 ;
        RECT 679.950 467.400 759.900 468.600 ;
        RECT 577.950 466.950 580.050 467.400 ;
        RECT 619.950 466.950 622.050 467.400 ;
        RECT 679.950 466.950 682.050 467.400 ;
        RECT 757.800 466.950 759.900 467.400 ;
        RECT 760.950 468.600 763.050 469.050 ;
        RECT 844.950 468.600 847.050 469.050 ;
        RECT 760.950 467.400 847.050 468.600 ;
        RECT 760.950 466.950 763.050 467.400 ;
        RECT 844.950 466.950 847.050 467.400 ;
        RECT 886.950 468.600 889.050 469.050 ;
        RECT 913.950 468.600 916.050 469.050 ;
        RECT 886.950 467.400 916.050 468.600 ;
        RECT 886.950 466.950 889.050 467.400 ;
        RECT 913.950 466.950 916.050 467.400 ;
        RECT 412.950 465.600 415.050 466.050 ;
        RECT 371.400 464.400 415.050 465.600 ;
        RECT 253.950 463.950 256.050 464.400 ;
        RECT 259.950 463.950 262.050 464.400 ;
        RECT 412.950 463.950 415.050 464.400 ;
        RECT 424.950 465.600 427.050 466.050 ;
        RECT 538.950 465.600 541.050 466.050 ;
        RECT 424.950 464.400 541.050 465.600 ;
        RECT 424.950 463.950 427.050 464.400 ;
        RECT 538.950 463.950 541.050 464.400 ;
        RECT 631.950 465.600 634.050 466.050 ;
        RECT 667.950 465.600 670.050 466.050 ;
        RECT 631.950 464.400 670.050 465.600 ;
        RECT 631.950 463.950 634.050 464.400 ;
        RECT 667.950 463.950 670.050 464.400 ;
        RECT 808.950 465.600 811.050 466.050 ;
        RECT 832.950 465.600 835.050 466.050 ;
        RECT 808.950 464.400 835.050 465.600 ;
        RECT 808.950 463.950 811.050 464.400 ;
        RECT 832.950 463.950 835.050 464.400 ;
        RECT 856.950 465.600 859.050 466.050 ;
        RECT 865.950 465.600 868.050 466.050 ;
        RECT 877.950 465.600 880.050 466.050 ;
        RECT 910.950 465.600 913.050 466.050 ;
        RECT 856.950 464.400 913.050 465.600 ;
        RECT 856.950 463.950 859.050 464.400 ;
        RECT 865.950 463.950 868.050 464.400 ;
        RECT 877.950 463.950 880.050 464.400 ;
        RECT 910.950 463.950 913.050 464.400 ;
        RECT 130.950 462.600 133.050 463.050 ;
        RECT 196.950 462.600 199.050 463.050 ;
        RECT 130.950 461.400 199.050 462.600 ;
        RECT 130.950 460.950 133.050 461.400 ;
        RECT 196.950 460.950 199.050 461.400 ;
        RECT 235.950 462.600 238.050 463.050 ;
        RECT 367.950 462.600 370.050 463.050 ;
        RECT 235.950 461.400 243.600 462.600 ;
        RECT 235.950 460.950 238.050 461.400 ;
        RECT 10.950 459.600 13.050 460.050 ;
        RECT 28.950 459.600 31.050 460.050 ;
        RECT 10.950 458.400 31.050 459.600 ;
        RECT 10.950 457.950 13.050 458.400 ;
        RECT 28.950 457.950 31.050 458.400 ;
        RECT 127.950 459.600 130.050 460.050 ;
        RECT 184.950 459.600 187.050 460.050 ;
        RECT 127.950 458.400 187.050 459.600 ;
        RECT 127.950 457.950 130.050 458.400 ;
        RECT 184.950 457.950 187.050 458.400 ;
        RECT 242.400 457.050 243.600 461.400 ;
        RECT 362.400 461.400 370.050 462.600 ;
        RECT 362.400 457.050 363.600 461.400 ;
        RECT 367.950 460.950 370.050 461.400 ;
        RECT 517.950 462.600 520.050 463.050 ;
        RECT 544.800 462.600 546.900 463.050 ;
        RECT 517.950 461.400 546.900 462.600 ;
        RECT 517.950 460.950 520.050 461.400 ;
        RECT 544.800 460.950 546.900 461.400 ;
        RECT 547.950 462.600 550.050 463.050 ;
        RECT 583.950 462.600 586.050 463.050 ;
        RECT 616.950 462.600 619.050 463.050 ;
        RECT 667.950 462.600 670.050 462.900 ;
        RECT 547.950 461.400 619.050 462.600 ;
        RECT 547.950 460.950 550.050 461.400 ;
        RECT 583.950 460.950 586.050 461.400 ;
        RECT 616.950 460.950 619.050 461.400 ;
        RECT 635.400 461.400 670.050 462.600 ;
        RECT 409.950 459.600 412.050 460.050 ;
        RECT 478.950 459.600 481.050 460.050 ;
        RECT 502.950 459.600 505.050 460.050 ;
        RECT 409.950 458.400 481.050 459.600 ;
        RECT 409.950 457.950 412.050 458.400 ;
        RECT 478.950 457.950 481.050 458.400 ;
        RECT 482.400 458.400 505.050 459.600 ;
        RECT 139.950 456.600 144.000 457.050 ;
        RECT 139.950 454.950 144.600 456.600 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 262.950 456.600 265.050 457.050 ;
        RECT 271.950 456.600 274.050 457.050 ;
        RECT 325.950 456.600 328.050 457.050 ;
        RECT 340.950 456.600 343.050 457.050 ;
        RECT 262.950 455.400 343.050 456.600 ;
        RECT 262.950 454.950 265.050 455.400 ;
        RECT 271.950 454.950 274.050 455.400 ;
        RECT 325.950 454.950 328.050 455.400 ;
        RECT 340.950 454.950 343.050 455.400 ;
        RECT 361.950 454.950 364.050 457.050 ;
        RECT 412.950 456.600 415.050 457.050 ;
        RECT 482.400 456.600 483.600 458.400 ;
        RECT 502.950 457.950 505.050 458.400 ;
        RECT 532.950 459.600 535.050 460.050 ;
        RECT 550.950 459.600 553.050 460.050 ;
        RECT 635.400 459.600 636.600 461.400 ;
        RECT 667.950 460.800 670.050 461.400 ;
        RECT 736.950 462.600 739.050 463.050 ;
        RECT 769.950 462.600 772.050 463.050 ;
        RECT 736.950 461.400 772.050 462.600 ;
        RECT 736.950 460.950 739.050 461.400 ;
        RECT 769.950 460.950 772.050 461.400 ;
        RECT 778.950 462.600 781.050 463.050 ;
        RECT 853.950 462.600 856.050 463.050 ;
        RECT 778.950 461.400 856.050 462.600 ;
        RECT 778.950 460.950 781.050 461.400 ;
        RECT 853.950 460.950 856.050 461.400 ;
        RECT 532.950 458.400 636.600 459.600 ;
        RECT 640.950 459.600 643.050 460.050 ;
        RECT 649.950 459.600 652.050 460.050 ;
        RECT 640.950 458.400 652.050 459.600 ;
        RECT 532.950 457.950 535.050 458.400 ;
        RECT 550.950 457.950 553.050 458.400 ;
        RECT 640.950 457.950 643.050 458.400 ;
        RECT 649.950 457.950 652.050 458.400 ;
        RECT 691.950 459.600 694.050 460.050 ;
        RECT 721.950 459.600 724.050 460.050 ;
        RECT 691.950 458.400 724.050 459.600 ;
        RECT 691.950 457.950 694.050 458.400 ;
        RECT 721.950 457.950 724.050 458.400 ;
        RECT 790.950 459.600 793.050 460.050 ;
        RECT 805.950 459.600 808.050 460.050 ;
        RECT 790.950 458.400 808.050 459.600 ;
        RECT 790.950 457.950 793.050 458.400 ;
        RECT 805.950 457.950 808.050 458.400 ;
        RECT 859.950 459.600 862.050 460.050 ;
        RECT 868.950 459.600 871.050 460.050 ;
        RECT 898.950 459.600 901.050 460.050 ;
        RECT 859.950 458.400 871.050 459.600 ;
        RECT 859.950 457.950 862.050 458.400 ;
        RECT 868.950 457.950 871.050 458.400 ;
        RECT 893.400 458.400 901.050 459.600 ;
        RECT 412.950 455.400 483.600 456.600 ;
        RECT 523.950 456.600 526.050 457.050 ;
        RECT 553.950 456.600 556.050 457.050 ;
        RECT 613.950 456.600 616.050 457.050 ;
        RECT 523.950 455.400 556.050 456.600 ;
        RECT 412.950 454.950 415.050 455.400 ;
        RECT 523.950 454.950 526.050 455.400 ;
        RECT 553.950 454.950 556.050 455.400 ;
        RECT 608.400 455.400 616.050 456.600 ;
        RECT 130.950 451.950 133.050 454.050 ;
        RECT 136.950 451.950 139.050 454.050 ;
        RECT 143.400 453.600 144.600 454.950 ;
        RECT 157.950 453.600 160.050 454.050 ;
        RECT 143.400 452.400 160.050 453.600 ;
        RECT 157.950 451.950 160.050 452.400 ;
        RECT 181.950 451.950 184.050 454.050 ;
        RECT 190.950 453.600 193.050 454.050 ;
        RECT 196.950 453.600 199.050 454.050 ;
        RECT 190.950 452.400 199.050 453.600 ;
        RECT 190.950 451.950 193.050 452.400 ;
        RECT 196.950 451.950 199.050 452.400 ;
        RECT 259.950 451.950 262.050 454.050 ;
        RECT 268.950 451.950 271.050 454.050 ;
        RECT 487.950 453.750 490.050 454.200 ;
        RECT 505.950 453.750 508.050 454.200 ;
        RECT 487.950 452.550 508.050 453.750 ;
        RECT 601.950 453.600 604.050 454.050 ;
        RECT 487.950 452.100 490.050 452.550 ;
        RECT 505.950 452.100 508.050 452.550 ;
        RECT 575.400 452.400 604.050 453.600 ;
        RECT 4.950 450.750 7.050 451.200 ;
        RECT 13.950 450.750 16.050 451.200 ;
        RECT 4.950 449.550 16.050 450.750 ;
        RECT 4.950 449.100 7.050 449.550 ;
        RECT 13.950 449.100 16.050 449.550 ;
        RECT 100.950 450.600 103.050 451.200 ;
        RECT 112.950 450.600 115.050 451.050 ;
        RECT 121.950 450.600 124.050 451.200 ;
        RECT 100.950 449.400 124.050 450.600 ;
        RECT 100.950 449.100 103.050 449.400 ;
        RECT 112.950 448.950 115.050 449.400 ;
        RECT 121.950 449.100 124.050 449.400 ;
        RECT 58.950 447.600 61.050 448.200 ;
        RECT 58.950 446.400 81.600 447.600 ;
        RECT 58.950 446.100 61.050 446.400 ;
        RECT 16.950 444.450 19.050 444.900 ;
        RECT 22.950 444.450 25.050 444.900 ;
        RECT 16.950 443.250 25.050 444.450 ;
        RECT 80.400 444.600 81.600 446.400 ;
        RECT 131.400 445.050 132.600 451.950 ;
        RECT 137.400 445.050 138.600 451.950 ;
        RECT 182.400 448.050 183.600 451.950 ;
        RECT 238.950 450.600 241.050 451.050 ;
        RECT 238.950 449.400 258.600 450.600 ;
        RECT 238.950 448.950 241.050 449.400 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 202.950 447.450 205.050 447.900 ;
        RECT 217.950 447.450 220.050 447.900 ;
        RECT 202.950 446.250 220.050 447.450 ;
        RECT 103.950 444.600 106.050 444.900 ;
        RECT 124.950 444.600 127.050 444.900 ;
        RECT 80.400 443.400 106.050 444.600 ;
        RECT 119.400 444.000 127.050 444.600 ;
        RECT 16.950 442.800 19.050 443.250 ;
        RECT 22.950 442.800 25.050 443.250 ;
        RECT 103.950 442.800 106.050 443.400 ;
        RECT 118.950 443.400 127.050 444.000 ;
        RECT 118.950 439.950 121.050 443.400 ;
        RECT 124.950 442.800 127.050 443.400 ;
        RECT 130.800 442.950 132.900 445.050 ;
        RECT 133.950 443.400 138.600 445.050 ;
        RECT 133.950 442.950 138.000 443.400 ;
        RECT 139.950 441.600 142.050 442.050 ;
        RECT 155.400 441.600 156.600 445.950 ;
        RECT 202.950 445.800 205.050 446.250 ;
        RECT 217.950 445.800 220.050 446.250 ;
        RECT 257.400 444.600 258.600 449.400 ;
        RECT 260.400 448.050 261.600 451.950 ;
        RECT 269.400 448.050 270.600 451.950 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 268.950 445.950 271.050 448.050 ;
        RECT 280.950 447.600 283.050 448.050 ;
        RECT 295.950 447.600 298.050 448.200 ;
        RECT 280.950 446.400 298.050 447.600 ;
        RECT 280.950 445.950 283.050 446.400 ;
        RECT 295.950 446.100 298.050 446.400 ;
        RECT 343.950 447.600 346.050 448.050 ;
        RECT 364.950 447.600 367.050 451.050 ;
        RECT 511.950 450.600 514.050 451.200 ;
        RECT 547.950 450.600 550.050 451.200 ;
        RECT 511.950 449.400 550.050 450.600 ;
        RECT 511.950 449.100 514.050 449.400 ;
        RECT 547.950 449.100 550.050 449.400 ;
        RECT 556.950 450.600 559.050 451.200 ;
        RECT 575.400 450.600 576.600 452.400 ;
        RECT 601.950 451.950 604.050 452.400 ;
        RECT 556.950 449.400 576.600 450.600 ;
        RECT 577.950 450.600 580.050 451.050 ;
        RECT 577.950 449.400 600.600 450.600 ;
        RECT 556.950 449.100 559.050 449.400 ;
        RECT 577.950 448.950 580.050 449.400 ;
        RECT 388.950 447.600 391.050 448.050 ;
        RECT 343.950 446.400 391.050 447.600 ;
        RECT 343.950 445.950 346.050 446.400 ;
        RECT 388.950 445.950 391.050 446.400 ;
        RECT 400.950 447.450 403.050 447.900 ;
        RECT 433.950 447.450 436.050 447.900 ;
        RECT 400.950 446.250 436.050 447.450 ;
        RECT 400.950 445.800 403.050 446.250 ;
        RECT 433.950 445.800 436.050 446.250 ;
        RECT 274.950 444.600 277.050 445.050 ;
        RECT 257.400 443.400 277.050 444.600 ;
        RECT 274.950 442.950 277.050 443.400 ;
        RECT 331.950 444.600 334.050 445.050 ;
        RECT 340.950 444.600 343.050 445.050 ;
        RECT 526.950 444.600 529.050 444.900 ;
        RECT 331.950 443.400 343.050 444.600 ;
        RECT 331.950 442.950 334.050 443.400 ;
        RECT 340.950 442.950 343.050 443.400 ;
        RECT 515.400 443.400 529.050 444.600 ;
        RECT 515.400 442.050 516.600 443.400 ;
        RECT 526.950 442.800 529.050 443.400 ;
        RECT 544.950 444.450 547.050 444.900 ;
        RECT 553.950 444.450 556.050 444.900 ;
        RECT 544.950 443.250 556.050 444.450 ;
        RECT 544.950 442.800 547.050 443.250 ;
        RECT 553.950 442.800 556.050 443.250 ;
        RECT 571.950 444.600 574.050 444.900 ;
        RECT 592.950 444.600 595.050 444.900 ;
        RECT 571.950 443.400 595.050 444.600 ;
        RECT 571.950 442.800 574.050 443.400 ;
        RECT 592.950 442.800 595.050 443.400 ;
        RECT 599.400 442.050 600.600 449.400 ;
        RECT 604.950 448.950 607.050 451.050 ;
        RECT 605.400 445.050 606.600 448.950 ;
        RECT 604.950 442.950 607.050 445.050 ;
        RECT 608.400 442.050 609.600 455.400 ;
        RECT 613.950 454.950 616.050 455.400 ;
        RECT 637.950 456.600 640.050 457.050 ;
        RECT 676.950 456.600 679.050 457.050 ;
        RECT 637.950 455.400 679.050 456.600 ;
        RECT 637.950 454.950 640.050 455.400 ;
        RECT 676.950 454.950 679.050 455.400 ;
        RECT 697.950 456.600 700.050 457.050 ;
        RECT 706.950 456.600 709.050 457.050 ;
        RECT 697.950 455.400 709.050 456.600 ;
        RECT 697.950 454.950 700.050 455.400 ;
        RECT 706.950 454.950 709.050 455.400 ;
        RECT 739.950 456.600 742.050 457.050 ;
        RECT 748.950 456.600 751.050 457.050 ;
        RECT 739.950 455.400 751.050 456.600 ;
        RECT 739.950 454.950 742.050 455.400 ;
        RECT 748.950 454.950 751.050 455.400 ;
        RECT 760.950 456.600 763.050 457.050 ;
        RECT 775.950 456.600 778.050 457.050 ;
        RECT 760.950 455.400 778.050 456.600 ;
        RECT 760.950 454.950 763.050 455.400 ;
        RECT 775.950 454.950 778.050 455.400 ;
        RECT 781.950 456.600 784.050 457.050 ;
        RECT 793.950 456.600 796.050 457.050 ;
        RECT 781.950 455.400 796.050 456.600 ;
        RECT 781.950 454.950 784.050 455.400 ;
        RECT 793.950 454.950 796.050 455.400 ;
        RECT 853.950 456.600 856.050 457.050 ;
        RECT 893.400 456.600 894.600 458.400 ;
        RECT 898.950 457.950 901.050 458.400 ;
        RECT 853.950 455.400 894.600 456.600 ;
        RECT 895.950 456.600 898.050 457.050 ;
        RECT 895.950 455.400 921.600 456.600 ;
        RECT 853.950 454.950 856.050 455.400 ;
        RECT 895.950 454.950 898.050 455.400 ;
        RECT 682.950 453.600 685.050 454.050 ;
        RECT 665.400 452.400 685.050 453.600 ;
        RECT 613.950 449.100 616.050 451.200 ;
        RECT 619.950 450.600 622.050 451.200 ;
        RECT 631.950 450.750 634.050 451.200 ;
        RECT 646.950 450.750 649.050 451.200 ;
        RECT 665.400 451.050 666.600 452.400 ;
        RECT 682.950 451.950 685.050 452.400 ;
        RECT 694.950 453.600 697.050 453.900 ;
        RECT 727.950 453.600 730.050 454.050 ;
        RECT 694.950 452.400 730.050 453.600 ;
        RECT 694.950 451.800 697.050 452.400 ;
        RECT 727.950 451.950 730.050 452.400 ;
        RECT 757.950 453.600 760.050 454.050 ;
        RECT 772.950 453.600 775.050 454.050 ;
        RECT 757.950 452.400 775.050 453.600 ;
        RECT 757.950 451.950 760.050 452.400 ;
        RECT 772.950 451.950 775.050 452.400 ;
        RECT 787.950 453.600 790.050 454.050 ;
        RECT 814.950 453.600 817.050 454.050 ;
        RECT 787.950 452.400 817.050 453.600 ;
        RECT 787.950 451.950 790.050 452.400 ;
        RECT 814.950 451.950 817.050 452.400 ;
        RECT 853.950 453.600 856.050 453.900 ;
        RECT 883.950 453.600 886.050 454.050 ;
        RECT 853.950 452.400 886.050 453.600 ;
        RECT 853.950 451.800 856.050 452.400 ;
        RECT 883.950 451.950 886.050 452.400 ;
        RECT 631.950 450.600 649.050 450.750 ;
        RECT 619.950 449.550 649.050 450.600 ;
        RECT 619.950 449.400 634.050 449.550 ;
        RECT 619.950 449.100 622.050 449.400 ;
        RECT 631.950 449.100 634.050 449.400 ;
        RECT 646.950 449.100 649.050 449.550 ;
        RECT 614.400 447.600 615.600 449.100 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 673.950 450.600 676.050 451.050 ;
        RECT 688.950 450.600 691.050 451.200 ;
        RECT 673.950 449.400 691.050 450.600 ;
        RECT 673.950 448.950 676.050 449.400 ;
        RECT 688.950 449.100 691.050 449.400 ;
        RECT 703.950 449.100 706.050 451.200 ;
        RECT 709.950 450.750 712.050 451.200 ;
        RECT 715.950 450.750 718.050 451.200 ;
        RECT 709.950 449.550 718.050 450.750 ;
        RECT 745.950 450.600 748.050 451.200 ;
        RECT 709.950 449.100 712.050 449.550 ;
        RECT 715.950 449.100 718.050 449.550 ;
        RECT 719.400 449.400 748.050 450.600 ;
        RECT 625.950 447.600 628.050 448.050 ;
        RECT 691.950 447.600 694.050 448.050 ;
        RECT 614.400 447.000 624.600 447.600 ;
        RECT 614.400 446.400 625.050 447.000 ;
        RECT 622.950 442.950 625.050 446.400 ;
        RECT 625.950 446.400 694.050 447.600 ;
        RECT 625.950 445.950 628.050 446.400 ;
        RECT 691.950 445.950 694.050 446.400 ;
        RECT 646.950 444.600 649.050 445.050 ;
        RECT 661.950 444.600 664.050 444.900 ;
        RECT 646.950 443.400 664.050 444.600 ;
        RECT 646.950 442.950 649.050 443.400 ;
        RECT 661.950 442.800 664.050 443.400 ;
        RECT 667.950 444.600 670.050 445.050 ;
        RECT 667.950 444.000 684.600 444.600 ;
        RECT 691.950 444.450 694.050 444.900 ;
        RECT 700.950 444.450 703.050 444.900 ;
        RECT 667.950 443.400 685.050 444.000 ;
        RECT 667.950 442.950 670.050 443.400 ;
        RECT 139.950 440.400 156.600 441.600 ;
        RECT 193.950 441.600 196.050 442.050 ;
        RECT 208.950 441.600 211.050 442.050 ;
        RECT 322.950 441.600 325.050 442.050 ;
        RECT 193.950 440.400 211.050 441.600 ;
        RECT 139.950 439.950 142.050 440.400 ;
        RECT 193.950 439.950 196.050 440.400 ;
        RECT 208.950 439.950 211.050 440.400 ;
        RECT 278.400 440.400 325.050 441.600 ;
        RECT 214.950 438.600 217.050 439.050 ;
        RECT 278.400 438.600 279.600 440.400 ;
        RECT 322.950 439.950 325.050 440.400 ;
        RECT 430.950 441.600 433.050 442.050 ;
        RECT 514.950 441.600 517.050 442.050 ;
        RECT 556.950 441.600 559.050 442.050 ;
        RECT 430.950 440.400 517.050 441.600 ;
        RECT 430.950 439.950 433.050 440.400 ;
        RECT 514.950 439.950 517.050 440.400 ;
        RECT 530.400 440.400 559.050 441.600 ;
        RECT 214.950 437.400 279.600 438.600 ;
        RECT 433.950 438.600 436.050 439.050 ;
        RECT 484.950 438.600 487.050 439.050 ;
        RECT 433.950 437.400 487.050 438.600 ;
        RECT 214.950 436.950 217.050 437.400 ;
        RECT 433.950 436.950 436.050 437.400 ;
        RECT 484.950 436.950 487.050 437.400 ;
        RECT 502.950 438.600 505.050 439.050 ;
        RECT 530.400 438.600 531.600 440.400 ;
        RECT 556.950 439.950 559.050 440.400 ;
        RECT 595.950 440.400 600.600 442.050 ;
        RECT 595.950 439.950 600.000 440.400 ;
        RECT 607.950 439.950 610.050 442.050 ;
        RECT 664.950 441.600 667.050 442.050 ;
        RECT 670.950 441.600 673.050 442.050 ;
        RECT 664.950 440.400 673.050 441.600 ;
        RECT 664.950 439.950 667.050 440.400 ;
        RECT 670.950 439.950 673.050 440.400 ;
        RECT 682.950 439.950 685.050 443.400 ;
        RECT 691.950 443.250 703.050 444.450 ;
        RECT 691.950 442.800 694.050 443.250 ;
        RECT 700.950 442.800 703.050 443.250 ;
        RECT 704.400 441.600 705.600 449.100 ;
        RECT 719.400 445.050 720.600 449.400 ;
        RECT 745.950 449.100 748.050 449.400 ;
        RECT 778.950 448.950 781.050 451.050 ;
        RECT 784.950 450.750 787.050 451.200 ;
        RECT 790.950 450.750 793.050 451.200 ;
        RECT 784.950 449.550 793.050 450.750 ;
        RECT 784.950 449.100 787.050 449.550 ;
        RECT 790.950 449.100 793.050 449.550 ;
        RECT 799.950 450.600 802.050 451.200 ;
        RECT 811.950 450.600 814.050 451.050 ;
        RECT 838.950 450.600 841.050 451.200 ;
        RECT 799.950 449.400 814.050 450.600 ;
        RECT 799.950 449.100 802.050 449.400 ;
        RECT 811.950 448.950 814.050 449.400 ;
        RECT 824.400 449.400 841.050 450.600 ;
        RECT 718.950 442.950 721.050 445.050 ;
        RECT 730.950 444.600 733.050 444.900 ;
        RECT 736.950 444.600 739.050 445.050 ;
        RECT 730.950 443.400 739.050 444.600 ;
        RECT 730.950 442.800 733.050 443.400 ;
        RECT 736.950 442.950 739.050 443.400 ;
        RECT 751.950 444.450 754.050 444.900 ;
        RECT 757.950 444.450 760.050 444.900 ;
        RECT 751.950 443.250 760.050 444.450 ;
        RECT 751.950 442.800 754.050 443.250 ;
        RECT 757.950 442.800 760.050 443.250 ;
        RECT 772.950 444.600 775.050 444.900 ;
        RECT 779.400 444.600 780.600 448.950 ;
        RECT 824.400 447.600 825.600 449.400 ;
        RECT 838.950 449.100 841.050 449.400 ;
        RECT 850.950 448.950 853.050 451.050 ;
        RECT 865.950 448.950 868.050 451.050 ;
        RECT 904.950 449.100 907.050 451.200 ;
        RECT 920.400 450.600 921.600 455.400 ;
        RECT 925.950 454.950 928.050 457.050 ;
        RECT 922.950 450.600 925.050 451.050 ;
        RECT 920.400 449.400 925.050 450.600 ;
        RECT 772.950 443.400 780.600 444.600 ;
        RECT 809.400 446.400 825.600 447.600 ;
        RECT 772.950 442.800 775.050 443.400 ;
        RECT 721.950 441.600 724.050 442.050 ;
        RECT 704.400 440.400 724.050 441.600 ;
        RECT 721.950 439.950 724.050 440.400 ;
        RECT 799.950 441.600 802.050 442.050 ;
        RECT 809.400 441.600 810.600 446.400 ;
        RECT 851.400 445.050 852.600 448.950 ;
        RECT 826.950 444.450 829.050 444.900 ;
        RECT 835.950 444.450 838.050 444.900 ;
        RECT 826.950 443.250 838.050 444.450 ;
        RECT 826.950 442.800 829.050 443.250 ;
        RECT 835.950 442.800 838.050 443.250 ;
        RECT 850.950 442.950 853.050 445.050 ;
        RECT 862.950 444.600 865.050 444.900 ;
        RECT 866.400 444.600 867.600 448.950 ;
        RECT 905.400 447.600 906.600 449.100 ;
        RECT 922.950 448.950 925.050 449.400 ;
        RECT 902.400 446.400 906.600 447.600 ;
        RECT 862.950 443.400 867.600 444.600 ;
        RECT 886.950 444.600 889.050 444.900 ;
        RECT 902.400 444.600 903.600 446.400 ;
        RECT 926.400 444.900 927.600 454.950 ;
        RECT 934.950 448.950 937.050 451.050 ;
        RECT 935.400 445.050 936.600 448.950 ;
        RECT 886.950 443.400 903.600 444.600 ;
        RECT 862.950 442.800 865.050 443.400 ;
        RECT 886.950 442.800 889.050 443.400 ;
        RECT 925.950 442.800 928.050 444.900 ;
        RECT 934.950 442.950 937.050 445.050 ;
        RECT 799.950 440.400 810.600 441.600 ;
        RECT 817.950 441.600 820.050 442.050 ;
        RECT 874.950 441.600 877.050 442.050 ;
        RECT 817.950 440.400 877.050 441.600 ;
        RECT 799.950 439.950 802.050 440.400 ;
        RECT 817.950 439.950 820.050 440.400 ;
        RECT 874.950 439.950 877.050 440.400 ;
        RECT 502.950 437.400 531.600 438.600 ;
        RECT 592.950 438.600 595.050 439.050 ;
        RECT 625.800 438.600 627.900 439.050 ;
        RECT 592.950 437.400 627.900 438.600 ;
        RECT 502.950 436.950 505.050 437.400 ;
        RECT 592.950 436.950 595.050 437.400 ;
        RECT 625.800 436.950 627.900 437.400 ;
        RECT 628.950 438.600 631.050 438.900 ;
        RECT 652.950 438.600 655.050 439.050 ;
        RECT 628.950 437.400 655.050 438.600 ;
        RECT 628.950 436.800 631.050 437.400 ;
        RECT 652.950 436.950 655.050 437.400 ;
        RECT 673.950 438.600 676.050 439.050 ;
        RECT 715.950 438.600 718.050 439.050 ;
        RECT 673.950 437.400 718.050 438.600 ;
        RECT 673.950 436.950 676.050 437.400 ;
        RECT 715.950 436.950 718.050 437.400 ;
        RECT 730.950 438.600 733.050 439.050 ;
        RECT 784.950 438.600 787.050 439.050 ;
        RECT 823.950 438.600 826.050 439.050 ;
        RECT 730.950 437.400 787.050 438.600 ;
        RECT 730.950 436.950 733.050 437.400 ;
        RECT 784.950 436.950 787.050 437.400 ;
        RECT 812.400 437.400 826.050 438.600 ;
        RECT 4.950 435.600 7.050 436.050 ;
        RECT 97.950 435.600 100.050 436.050 ;
        RECT 343.950 435.600 346.050 436.050 ;
        RECT 4.950 434.400 100.050 435.600 ;
        RECT 305.400 435.000 346.050 435.600 ;
        RECT 4.950 433.950 7.050 434.400 ;
        RECT 97.950 433.950 100.050 434.400 ;
        RECT 304.950 434.400 346.050 435.000 ;
        RECT 31.950 432.600 34.050 433.050 ;
        RECT 43.950 432.600 46.050 433.050 ;
        RECT 73.950 432.600 76.050 433.050 ;
        RECT 31.950 431.400 76.050 432.600 ;
        RECT 31.950 430.950 34.050 431.400 ;
        RECT 43.950 430.950 46.050 431.400 ;
        RECT 73.950 430.950 76.050 431.400 ;
        RECT 184.950 432.600 187.050 433.050 ;
        RECT 214.950 432.600 217.050 433.050 ;
        RECT 184.950 431.400 217.050 432.600 ;
        RECT 184.950 430.950 187.050 431.400 ;
        RECT 214.950 430.950 217.050 431.400 ;
        RECT 304.950 430.950 307.050 434.400 ;
        RECT 343.950 433.950 346.050 434.400 ;
        RECT 499.950 435.600 502.050 436.050 ;
        RECT 535.950 435.600 538.050 436.050 ;
        RECT 499.950 434.400 538.050 435.600 ;
        RECT 499.950 433.950 502.050 434.400 ;
        RECT 535.950 433.950 538.050 434.400 ;
        RECT 568.950 435.600 571.050 436.050 ;
        RECT 598.950 435.600 601.050 436.050 ;
        RECT 568.950 434.400 601.050 435.600 ;
        RECT 568.950 433.950 571.050 434.400 ;
        RECT 598.950 433.950 601.050 434.400 ;
        RECT 643.950 435.600 646.050 436.050 ;
        RECT 649.950 435.600 652.050 436.050 ;
        RECT 643.950 434.400 652.050 435.600 ;
        RECT 643.950 433.950 646.050 434.400 ;
        RECT 649.950 433.950 652.050 434.400 ;
        RECT 658.950 435.600 661.050 436.050 ;
        RECT 667.950 435.600 670.050 436.050 ;
        RECT 658.950 434.400 670.050 435.600 ;
        RECT 658.950 433.950 661.050 434.400 ;
        RECT 667.950 433.950 670.050 434.400 ;
        RECT 694.950 435.600 697.050 436.050 ;
        RECT 706.950 435.600 709.050 436.050 ;
        RECT 694.950 434.400 709.050 435.600 ;
        RECT 694.950 433.950 697.050 434.400 ;
        RECT 706.950 433.950 709.050 434.400 ;
        RECT 715.950 435.600 718.050 435.900 ;
        RECT 724.950 435.600 727.050 436.050 ;
        RECT 796.950 435.600 799.050 436.050 ;
        RECT 715.950 434.400 727.050 435.600 ;
        RECT 715.950 433.800 718.050 434.400 ;
        RECT 724.950 433.950 727.050 434.400 ;
        RECT 767.400 434.400 799.050 435.600 ;
        RECT 382.950 432.600 385.050 433.050 ;
        RECT 391.950 432.600 394.050 433.050 ;
        RECT 436.950 432.600 439.050 433.050 ;
        RECT 382.950 431.400 439.050 432.600 ;
        RECT 382.950 430.950 385.050 431.400 ;
        RECT 391.950 430.950 394.050 431.400 ;
        RECT 436.950 430.950 439.050 431.400 ;
        RECT 457.950 432.600 460.050 433.050 ;
        RECT 559.950 432.600 562.050 433.050 ;
        RECT 457.950 431.400 562.050 432.600 ;
        RECT 457.950 430.950 460.050 431.400 ;
        RECT 559.950 430.950 562.050 431.400 ;
        RECT 622.950 432.600 625.050 433.050 ;
        RECT 628.950 432.600 631.050 433.050 ;
        RECT 622.950 431.400 631.050 432.600 ;
        RECT 622.950 430.950 625.050 431.400 ;
        RECT 628.950 430.950 631.050 431.400 ;
        RECT 640.950 432.600 643.050 433.050 ;
        RECT 760.950 432.600 763.050 433.050 ;
        RECT 767.400 432.600 768.600 434.400 ;
        RECT 796.950 433.950 799.050 434.400 ;
        RECT 805.950 435.600 808.050 436.050 ;
        RECT 812.400 435.600 813.600 437.400 ;
        RECT 823.950 436.950 826.050 437.400 ;
        RECT 856.950 438.600 859.050 439.050 ;
        RECT 880.950 438.600 883.050 439.050 ;
        RECT 856.950 437.400 883.050 438.600 ;
        RECT 856.950 436.950 859.050 437.400 ;
        RECT 880.950 436.950 883.050 437.400 ;
        RECT 838.950 435.600 841.050 436.050 ;
        RECT 805.950 434.400 813.600 435.600 ;
        RECT 815.400 434.400 841.050 435.600 ;
        RECT 805.950 433.950 808.050 434.400 ;
        RECT 640.950 431.400 768.600 432.600 ;
        RECT 787.950 432.600 790.050 433.050 ;
        RECT 815.400 432.600 816.600 434.400 ;
        RECT 838.950 433.950 841.050 434.400 ;
        RECT 913.950 435.600 916.050 436.050 ;
        RECT 931.950 435.600 934.050 436.050 ;
        RECT 913.950 434.400 934.050 435.600 ;
        RECT 913.950 433.950 916.050 434.400 ;
        RECT 931.950 433.950 934.050 434.400 ;
        RECT 856.950 432.600 859.050 433.050 ;
        RECT 787.950 431.400 816.600 432.600 ;
        RECT 818.400 431.400 859.050 432.600 ;
        RECT 640.950 430.950 643.050 431.400 ;
        RECT 760.950 430.950 763.050 431.400 ;
        RECT 787.950 430.950 790.050 431.400 ;
        RECT 133.950 429.600 136.050 430.050 ;
        RECT 157.950 429.600 160.050 430.050 ;
        RECT 133.950 428.400 160.050 429.600 ;
        RECT 133.950 427.950 136.050 428.400 ;
        RECT 157.950 427.950 160.050 428.400 ;
        RECT 250.950 429.600 253.050 430.050 ;
        RECT 274.950 429.600 277.050 430.050 ;
        RECT 250.950 428.400 277.050 429.600 ;
        RECT 250.950 427.950 253.050 428.400 ;
        RECT 274.950 427.950 277.050 428.400 ;
        RECT 313.950 429.600 316.050 430.050 ;
        RECT 325.950 429.600 328.050 430.050 ;
        RECT 313.950 428.400 328.050 429.600 ;
        RECT 313.950 427.950 316.050 428.400 ;
        RECT 325.950 427.950 328.050 428.400 ;
        RECT 391.950 429.600 394.050 429.900 ;
        RECT 421.950 429.600 424.050 430.050 ;
        RECT 391.950 428.400 424.050 429.600 ;
        RECT 391.950 427.800 394.050 428.400 ;
        RECT 421.950 427.950 424.050 428.400 ;
        RECT 577.950 429.600 580.050 430.050 ;
        RECT 616.950 429.600 619.050 430.050 ;
        RECT 634.950 429.600 637.050 430.050 ;
        RECT 577.950 428.400 637.050 429.600 ;
        RECT 577.950 427.950 580.050 428.400 ;
        RECT 616.950 427.950 619.050 428.400 ;
        RECT 634.950 427.950 637.050 428.400 ;
        RECT 682.950 429.600 685.050 430.050 ;
        RECT 694.950 429.600 697.050 430.050 ;
        RECT 718.950 429.600 721.050 430.050 ;
        RECT 682.950 428.400 693.600 429.600 ;
        RECT 682.950 427.950 685.050 428.400 ;
        RECT 7.950 426.600 10.050 427.050 ;
        RECT 70.950 426.600 73.050 427.050 ;
        RECT 7.950 425.400 73.050 426.600 ;
        RECT 7.950 424.950 10.050 425.400 ;
        RECT 70.950 424.950 73.050 425.400 ;
        RECT 88.950 426.600 91.050 427.050 ;
        RECT 124.950 426.600 127.050 427.050 ;
        RECT 130.950 426.600 133.050 427.050 ;
        RECT 88.950 425.400 133.050 426.600 ;
        RECT 88.950 424.950 91.050 425.400 ;
        RECT 124.950 424.950 127.050 425.400 ;
        RECT 130.950 424.950 133.050 425.400 ;
        RECT 175.950 426.600 178.050 427.050 ;
        RECT 187.950 426.600 190.050 427.050 ;
        RECT 175.950 425.400 190.050 426.600 ;
        RECT 175.950 424.950 178.050 425.400 ;
        RECT 187.950 424.950 190.050 425.400 ;
        RECT 232.950 426.600 235.050 427.050 ;
        RECT 268.950 426.600 271.050 427.050 ;
        RECT 232.950 425.400 271.050 426.600 ;
        RECT 232.950 424.950 235.050 425.400 ;
        RECT 268.950 424.950 271.050 425.400 ;
        RECT 388.950 426.600 391.050 427.050 ;
        RECT 589.950 426.600 592.050 427.050 ;
        RECT 595.950 426.600 598.050 427.050 ;
        RECT 601.950 426.600 604.050 427.050 ;
        RECT 388.950 425.400 429.600 426.600 ;
        RECT 388.950 424.950 391.050 425.400 ;
        RECT 428.400 424.050 429.600 425.400 ;
        RECT 589.950 425.400 604.050 426.600 ;
        RECT 589.950 424.950 592.050 425.400 ;
        RECT 595.950 424.950 598.050 425.400 ;
        RECT 601.950 424.950 604.050 425.400 ;
        RECT 652.950 426.600 655.050 427.050 ;
        RECT 673.950 426.600 676.050 427.050 ;
        RECT 652.950 425.400 676.050 426.600 ;
        RECT 652.950 424.950 655.050 425.400 ;
        RECT 673.950 424.950 676.050 425.400 ;
        RECT 679.950 426.600 682.050 427.050 ;
        RECT 685.950 426.600 688.050 427.050 ;
        RECT 679.950 425.400 688.050 426.600 ;
        RECT 692.400 426.600 693.600 428.400 ;
        RECT 694.950 428.400 721.050 429.600 ;
        RECT 694.950 427.950 697.050 428.400 ;
        RECT 718.950 427.950 721.050 428.400 ;
        RECT 775.950 429.600 778.050 430.050 ;
        RECT 784.950 429.600 787.050 430.050 ;
        RECT 818.400 429.600 819.600 431.400 ;
        RECT 856.950 430.950 859.050 431.400 ;
        RECT 886.950 432.600 889.050 433.050 ;
        RECT 922.950 432.600 925.050 433.050 ;
        RECT 886.950 431.400 925.050 432.600 ;
        RECT 886.950 430.950 889.050 431.400 ;
        RECT 922.950 430.950 925.050 431.400 ;
        RECT 775.950 428.400 819.600 429.600 ;
        RECT 820.950 429.600 823.050 430.050 ;
        RECT 841.950 429.600 844.050 430.050 ;
        RECT 820.950 428.400 844.050 429.600 ;
        RECT 775.950 427.950 778.050 428.400 ;
        RECT 784.950 427.950 787.050 428.400 ;
        RECT 820.950 427.950 823.050 428.400 ;
        RECT 841.950 427.950 844.050 428.400 ;
        RECT 856.950 429.600 859.050 429.900 ;
        RECT 868.950 429.600 871.050 430.050 ;
        RECT 856.950 428.400 871.050 429.600 ;
        RECT 856.950 427.800 859.050 428.400 ;
        RECT 868.950 427.950 871.050 428.400 ;
        RECT 916.950 429.600 919.050 430.050 ;
        RECT 928.950 429.600 931.050 430.050 ;
        RECT 916.950 428.400 931.050 429.600 ;
        RECT 916.950 427.950 919.050 428.400 ;
        RECT 928.950 427.950 931.050 428.400 ;
        RECT 715.950 426.600 718.050 427.050 ;
        RECT 692.400 425.400 718.050 426.600 ;
        RECT 679.950 424.950 682.050 425.400 ;
        RECT 685.950 424.950 688.050 425.400 ;
        RECT 715.950 424.950 718.050 425.400 ;
        RECT 742.950 426.600 745.050 427.050 ;
        RECT 757.800 426.600 759.900 427.050 ;
        RECT 742.950 425.400 759.900 426.600 ;
        RECT 742.950 424.950 745.050 425.400 ;
        RECT 757.800 424.950 759.900 425.400 ;
        RECT 760.950 426.600 763.050 427.050 ;
        RECT 907.950 426.600 910.050 427.050 ;
        RECT 934.950 426.600 937.050 427.050 ;
        RECT 760.950 425.400 840.600 426.600 ;
        RECT 760.950 424.950 763.050 425.400 ;
        RECT 839.400 424.050 840.600 425.400 ;
        RECT 907.950 425.400 937.050 426.600 ;
        RECT 907.950 424.950 910.050 425.400 ;
        RECT 934.950 424.950 937.050 425.400 ;
        RECT 79.950 423.600 82.050 424.050 ;
        RECT 91.950 423.600 94.050 424.050 ;
        RECT 79.950 422.400 94.050 423.600 ;
        RECT 79.950 421.950 82.050 422.400 ;
        RECT 91.950 421.950 94.050 422.400 ;
        RECT 97.950 423.600 100.050 424.050 ;
        RECT 112.950 423.600 115.050 424.050 ;
        RECT 97.950 422.400 115.050 423.600 ;
        RECT 97.950 421.950 100.050 422.400 ;
        RECT 112.950 421.950 115.050 422.400 ;
        RECT 7.950 420.600 10.050 421.050 ;
        RECT 37.950 420.600 40.050 421.050 ;
        RECT 7.950 419.400 40.050 420.600 ;
        RECT 7.950 418.950 10.050 419.400 ;
        RECT 37.950 418.950 40.050 419.400 ;
        RECT 136.950 420.600 139.050 420.900 ;
        RECT 142.950 420.600 145.050 421.050 ;
        RECT 136.950 419.400 145.050 420.600 ;
        RECT 136.950 418.800 139.050 419.400 ;
        RECT 142.950 418.950 145.050 419.400 ;
        RECT 154.950 420.600 157.050 421.050 ;
        RECT 160.950 420.600 163.050 421.050 ;
        RECT 184.950 420.600 187.050 421.050 ;
        RECT 199.950 420.600 202.050 424.050 ;
        RECT 322.950 423.600 325.050 424.050 ;
        RECT 382.950 423.600 385.050 424.050 ;
        RECT 412.950 423.600 415.050 424.050 ;
        RECT 322.950 422.400 385.050 423.600 ;
        RECT 322.950 421.950 325.050 422.400 ;
        RECT 382.950 421.950 385.050 422.400 ;
        RECT 386.400 422.400 415.050 423.600 ;
        RECT 154.950 420.000 202.050 420.600 ;
        RECT 214.950 420.600 217.050 421.050 ;
        RECT 247.950 420.600 250.050 421.050 ;
        RECT 154.950 419.400 201.600 420.000 ;
        RECT 214.950 419.400 250.050 420.600 ;
        RECT 154.950 418.950 157.050 419.400 ;
        RECT 160.950 418.950 163.050 419.400 ;
        RECT 184.950 418.950 187.050 419.400 ;
        RECT 214.950 418.950 217.050 419.400 ;
        RECT 247.950 418.950 250.050 419.400 ;
        RECT 253.950 420.600 256.050 420.900 ;
        RECT 265.950 420.600 268.050 421.050 ;
        RECT 253.950 419.400 268.050 420.600 ;
        RECT 253.950 418.800 256.050 419.400 ;
        RECT 265.950 418.950 268.050 419.400 ;
        RECT 274.950 420.600 277.050 421.050 ;
        RECT 289.950 420.600 292.050 421.050 ;
        RECT 274.950 419.400 292.050 420.600 ;
        RECT 274.950 418.950 277.050 419.400 ;
        RECT 289.950 418.950 292.050 419.400 ;
        RECT 376.950 420.600 379.050 421.050 ;
        RECT 386.400 420.600 387.600 422.400 ;
        RECT 412.950 421.950 415.050 422.400 ;
        RECT 427.950 423.600 430.050 424.050 ;
        RECT 445.950 423.600 448.050 424.050 ;
        RECT 505.950 423.600 508.050 424.050 ;
        RECT 427.950 422.400 508.050 423.600 ;
        RECT 427.950 421.950 430.050 422.400 ;
        RECT 445.950 421.950 448.050 422.400 ;
        RECT 505.950 421.950 508.050 422.400 ;
        RECT 556.950 423.600 559.050 424.050 ;
        RECT 571.950 423.600 574.050 424.050 ;
        RECT 556.950 422.400 574.050 423.600 ;
        RECT 556.950 421.950 559.050 422.400 ;
        RECT 571.950 421.950 574.050 422.400 ;
        RECT 613.950 423.600 616.050 424.050 ;
        RECT 631.950 423.600 634.050 424.050 ;
        RECT 613.950 422.400 634.050 423.600 ;
        RECT 613.950 421.950 616.050 422.400 ;
        RECT 631.950 421.950 634.050 422.400 ;
        RECT 637.950 423.600 640.050 424.050 ;
        RECT 649.950 423.600 652.050 424.050 ;
        RECT 637.950 422.400 652.050 423.600 ;
        RECT 637.950 421.950 640.050 422.400 ;
        RECT 649.950 421.950 652.050 422.400 ;
        RECT 688.950 423.600 691.050 424.050 ;
        RECT 718.950 423.600 721.050 424.050 ;
        RECT 745.950 423.600 748.050 424.050 ;
        RECT 688.950 422.400 748.050 423.600 ;
        RECT 688.950 421.950 691.050 422.400 ;
        RECT 718.950 421.950 721.050 422.400 ;
        RECT 745.950 421.950 748.050 422.400 ;
        RECT 754.950 423.600 757.050 424.050 ;
        RECT 790.950 423.600 793.050 424.050 ;
        RECT 754.950 422.400 793.050 423.600 ;
        RECT 839.400 422.400 844.050 424.050 ;
        RECT 754.950 421.950 757.050 422.400 ;
        RECT 790.950 421.950 793.050 422.400 ;
        RECT 840.000 421.950 844.050 422.400 ;
        RECT 850.950 423.600 853.050 424.050 ;
        RECT 862.950 423.600 865.050 424.050 ;
        RECT 850.950 422.400 865.050 423.600 ;
        RECT 850.950 421.950 853.050 422.400 ;
        RECT 862.950 421.950 865.050 422.400 ;
        RECT 376.950 419.400 387.600 420.600 ;
        RECT 529.950 420.600 532.050 421.050 ;
        RECT 541.950 420.600 544.050 421.050 ;
        RECT 592.950 420.600 595.050 421.050 ;
        RECT 604.950 420.600 607.050 421.050 ;
        RECT 529.950 419.400 579.600 420.600 ;
        RECT 376.950 418.950 379.050 419.400 ;
        RECT 529.950 418.950 532.050 419.400 ;
        RECT 541.950 418.950 544.050 419.400 ;
        RECT 1.950 417.750 4.050 418.200 ;
        RECT 52.950 417.750 55.050 418.200 ;
        RECT 1.950 416.550 55.050 417.750 ;
        RECT 1.950 416.100 4.050 416.550 ;
        RECT 52.950 416.100 55.050 416.550 ;
        RECT 58.950 417.600 61.050 418.200 ;
        RECT 115.950 417.600 118.050 418.050 ;
        RECT 121.800 417.600 123.900 418.050 ;
        RECT 58.950 416.400 63.600 417.600 ;
        RECT 58.950 416.100 61.050 416.400 ;
        RECT 62.400 412.050 63.600 416.400 ;
        RECT 115.950 416.400 123.900 417.600 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 121.800 415.950 123.900 416.400 ;
        RECT 124.950 417.600 127.050 418.050 ;
        RECT 145.950 417.600 148.050 418.200 ;
        RECT 124.950 416.400 148.050 417.600 ;
        RECT 124.950 415.950 127.050 416.400 ;
        RECT 145.950 416.100 148.050 416.400 ;
        RECT 169.950 417.750 172.050 418.200 ;
        RECT 178.950 417.750 181.050 418.200 ;
        RECT 169.950 416.550 181.050 417.750 ;
        RECT 169.950 416.100 172.050 416.550 ;
        RECT 178.950 416.100 181.050 416.550 ;
        RECT 190.950 417.600 193.050 418.200 ;
        RECT 202.950 417.600 205.050 418.050 ;
        RECT 211.950 417.600 214.050 418.200 ;
        RECT 190.950 416.400 201.600 417.600 ;
        RECT 190.950 416.100 193.050 416.400 ;
        RECT 146.400 412.050 147.600 416.100 ;
        RECT 200.400 414.600 201.600 416.400 ;
        RECT 202.950 416.400 214.050 417.600 ;
        RECT 202.950 415.950 205.050 416.400 ;
        RECT 211.950 416.100 214.050 416.400 ;
        RECT 229.950 417.600 232.050 418.050 ;
        RECT 259.950 417.600 262.050 418.050 ;
        RECT 274.800 417.600 276.900 417.900 ;
        RECT 322.950 417.600 325.050 418.200 ;
        RECT 229.950 416.400 276.900 417.600 ;
        RECT 229.950 415.950 232.050 416.400 ;
        RECT 259.950 415.950 262.050 416.400 ;
        RECT 274.800 415.800 276.900 416.400 ;
        RECT 320.400 416.400 325.050 417.600 ;
        RECT 214.950 414.600 217.050 415.050 ;
        RECT 200.400 413.400 217.050 414.600 ;
        RECT 214.950 412.950 217.050 413.400 ;
        RECT 320.400 412.050 321.600 416.400 ;
        RECT 322.950 416.100 325.050 416.400 ;
        RECT 409.950 417.600 412.050 418.200 ;
        RECT 415.950 417.600 418.050 418.050 ;
        RECT 409.950 416.400 418.050 417.600 ;
        RECT 409.950 416.100 412.050 416.400 ;
        RECT 415.950 415.950 418.050 416.400 ;
        RECT 454.950 417.750 457.050 418.200 ;
        RECT 466.950 417.750 469.050 418.200 ;
        RECT 454.950 416.550 469.050 417.750 ;
        RECT 454.950 416.100 457.050 416.550 ;
        RECT 466.950 416.100 469.050 416.550 ;
        RECT 484.950 417.600 487.050 418.200 ;
        RECT 499.950 417.600 502.050 418.200 ;
        RECT 484.950 416.400 502.050 417.600 ;
        RECT 484.950 416.100 487.050 416.400 ;
        RECT 499.950 416.100 502.050 416.400 ;
        RECT 559.950 417.600 562.050 418.200 ;
        RECT 574.950 417.600 577.050 418.050 ;
        RECT 559.950 416.400 577.050 417.600 ;
        RECT 578.400 417.600 579.600 419.400 ;
        RECT 592.950 419.400 607.050 420.600 ;
        RECT 592.950 418.950 595.050 419.400 ;
        RECT 604.950 418.950 607.050 419.400 ;
        RECT 640.950 418.950 643.050 421.050 ;
        RECT 697.950 420.600 700.050 421.050 ;
        RECT 703.950 420.600 706.050 421.050 ;
        RECT 697.950 419.400 706.050 420.600 ;
        RECT 697.950 418.950 700.050 419.400 ;
        RECT 703.950 418.950 706.050 419.400 ;
        RECT 769.950 420.600 772.050 421.050 ;
        RECT 793.950 420.600 796.050 421.050 ;
        RECT 805.950 420.600 808.050 421.050 ;
        RECT 769.950 419.400 808.050 420.600 ;
        RECT 769.950 418.950 772.050 419.400 ;
        RECT 793.950 418.950 796.050 419.400 ;
        RECT 805.950 418.950 808.050 419.400 ;
        RECT 811.950 420.600 814.050 421.050 ;
        RECT 817.950 420.600 820.050 421.050 ;
        RECT 811.950 419.400 820.050 420.600 ;
        RECT 811.950 418.950 814.050 419.400 ;
        RECT 817.950 418.950 820.050 419.400 ;
        RECT 880.950 420.600 883.050 421.050 ;
        RECT 886.950 420.600 889.050 421.050 ;
        RECT 880.950 419.400 889.050 420.600 ;
        RECT 880.950 418.950 883.050 419.400 ;
        RECT 886.950 418.950 889.050 419.400 ;
        RECT 613.950 417.600 616.050 418.050 ;
        RECT 578.400 416.400 616.050 417.600 ;
        RECT 559.950 416.100 562.050 416.400 ;
        RECT 574.950 415.950 577.050 416.400 ;
        RECT 613.950 415.950 616.050 416.400 ;
        RECT 625.950 417.600 628.050 418.200 ;
        RECT 637.950 417.600 640.050 418.050 ;
        RECT 625.950 416.400 640.050 417.600 ;
        RECT 625.950 416.100 628.050 416.400 ;
        RECT 637.950 415.950 640.050 416.400 ;
        RECT 641.400 414.600 642.600 418.950 ;
        RECT 643.950 417.600 646.050 418.200 ;
        RECT 649.950 417.600 652.050 418.050 ;
        RECT 643.950 416.400 652.050 417.600 ;
        RECT 643.950 416.100 646.050 416.400 ;
        RECT 649.950 415.950 652.050 416.400 ;
        RECT 658.950 417.600 661.050 418.050 ;
        RECT 676.950 417.600 679.050 418.050 ;
        RECT 658.950 416.400 679.050 417.600 ;
        RECT 658.950 415.950 661.050 416.400 ;
        RECT 676.950 415.950 679.050 416.400 ;
        RECT 682.950 415.950 685.050 418.050 ;
        RECT 693.000 417.600 697.050 418.050 ;
        RECT 692.400 415.950 697.050 417.600 ;
        RECT 709.950 417.600 712.050 418.200 ;
        RECT 709.950 416.400 726.600 417.600 ;
        RECT 709.950 416.100 712.050 416.400 ;
        RECT 655.950 414.600 658.050 414.900 ;
        RECT 641.400 413.400 658.050 414.600 ;
        RECT 655.950 412.800 658.050 413.400 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 97.950 411.450 100.050 411.900 ;
        RECT 106.950 411.450 109.050 411.900 ;
        RECT 97.950 410.250 109.050 411.450 ;
        RECT 97.950 409.800 100.050 410.250 ;
        RECT 106.950 409.800 109.050 410.250 ;
        RECT 130.950 411.450 133.050 411.900 ;
        RECT 136.950 411.450 139.050 411.900 ;
        RECT 130.950 410.250 139.050 411.450 ;
        RECT 130.950 409.800 133.050 410.250 ;
        RECT 136.950 409.800 139.050 410.250 ;
        RECT 142.950 410.400 147.600 412.050 ;
        RECT 160.950 411.450 163.050 411.900 ;
        RECT 166.950 411.450 169.050 411.900 ;
        RECT 229.950 411.600 232.050 412.050 ;
        RECT 142.950 409.950 147.000 410.400 ;
        RECT 160.950 410.250 169.050 411.450 ;
        RECT 160.950 409.800 163.050 410.250 ;
        RECT 166.950 409.800 169.050 410.250 ;
        RECT 170.400 410.400 232.050 411.600 ;
        RECT 151.950 408.600 154.050 409.050 ;
        RECT 170.400 408.600 171.600 410.400 ;
        RECT 229.950 409.950 232.050 410.400 ;
        RECT 268.950 411.450 271.050 411.900 ;
        RECT 277.950 411.450 280.050 411.900 ;
        RECT 268.950 410.250 280.050 411.450 ;
        RECT 268.950 409.800 271.050 410.250 ;
        RECT 277.950 409.800 280.050 410.250 ;
        RECT 319.950 409.950 322.050 412.050 ;
        RECT 355.950 411.600 358.050 412.050 ;
        RECT 385.950 411.600 388.050 412.050 ;
        RECT 355.950 410.400 388.050 411.600 ;
        RECT 355.950 409.950 358.050 410.400 ;
        RECT 385.950 409.950 388.050 410.400 ;
        RECT 406.950 411.600 409.050 411.900 ;
        RECT 424.950 411.600 427.050 411.900 ;
        RECT 406.950 410.400 427.050 411.600 ;
        RECT 406.950 409.800 409.050 410.400 ;
        RECT 424.950 409.800 427.050 410.400 ;
        RECT 451.950 411.600 454.050 411.900 ;
        RECT 463.950 411.600 466.050 411.900 ;
        RECT 478.950 411.600 481.050 411.900 ;
        RECT 451.950 410.400 481.050 411.600 ;
        RECT 451.950 409.800 454.050 410.400 ;
        RECT 463.950 409.800 466.050 410.400 ;
        RECT 478.950 409.800 481.050 410.400 ;
        RECT 604.950 411.600 607.050 411.900 ;
        RECT 628.950 411.600 631.050 411.900 ;
        RECT 640.950 411.600 643.050 411.900 ;
        RECT 604.950 410.400 643.050 411.600 ;
        RECT 604.950 409.800 607.050 410.400 ;
        RECT 628.950 409.800 631.050 410.400 ;
        RECT 640.950 409.800 643.050 410.400 ;
        RECT 646.950 411.450 649.050 411.900 ;
        RECT 652.950 411.450 655.050 411.900 ;
        RECT 646.950 410.250 655.050 411.450 ;
        RECT 683.400 411.600 684.600 415.950 ;
        RECT 692.400 411.900 693.600 415.950 ;
        RECT 725.400 412.050 726.600 416.400 ;
        RECT 730.950 416.100 733.050 418.200 ;
        RECT 736.950 417.600 739.050 418.050 ;
        RECT 736.950 416.400 744.600 417.600 ;
        RECT 731.400 414.600 732.600 416.100 ;
        RECT 736.950 415.950 739.050 416.400 ;
        RECT 731.400 413.400 741.600 414.600 ;
        RECT 685.950 411.600 688.050 411.900 ;
        RECT 683.400 410.400 688.050 411.600 ;
        RECT 646.950 409.800 649.050 410.250 ;
        RECT 652.950 409.800 655.050 410.250 ;
        RECT 685.950 409.800 688.050 410.400 ;
        RECT 691.950 409.800 694.050 411.900 ;
        RECT 706.950 409.800 709.050 411.900 ;
        RECT 712.950 411.450 715.050 411.900 ;
        RECT 718.950 411.450 721.050 411.900 ;
        RECT 712.950 410.250 721.050 411.450 ;
        RECT 712.950 409.800 715.050 410.250 ;
        RECT 718.950 409.800 721.050 410.250 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 151.950 407.400 171.600 408.600 ;
        RECT 229.950 408.600 232.050 408.900 ;
        RECT 250.950 408.600 253.050 409.050 ;
        RECT 229.950 407.400 253.050 408.600 ;
        RECT 151.950 406.950 154.050 407.400 ;
        RECT 229.950 406.800 232.050 407.400 ;
        RECT 250.950 406.950 253.050 407.400 ;
        RECT 313.950 408.450 316.050 408.900 ;
        RECT 331.950 408.450 334.050 408.900 ;
        RECT 313.950 407.250 334.050 408.450 ;
        RECT 313.950 406.800 316.050 407.250 ;
        RECT 331.950 406.800 334.050 407.250 ;
        RECT 520.950 408.600 523.050 409.050 ;
        RECT 553.950 408.600 556.050 409.050 ;
        RECT 520.950 407.400 556.050 408.600 ;
        RECT 520.950 406.950 523.050 407.400 ;
        RECT 553.950 406.950 556.050 407.400 ;
        RECT 562.950 408.600 565.050 409.050 ;
        RECT 601.950 408.600 604.050 409.050 ;
        RECT 562.950 407.400 604.050 408.600 ;
        RECT 562.950 406.950 565.050 407.400 ;
        RECT 601.950 406.950 604.050 407.400 ;
        RECT 673.950 408.600 676.050 409.050 ;
        RECT 688.950 408.600 691.050 409.050 ;
        RECT 673.950 407.400 691.050 408.600 ;
        RECT 673.950 406.950 676.050 407.400 ;
        RECT 688.950 406.950 691.050 407.400 ;
        RECT 694.950 408.600 697.050 409.050 ;
        RECT 707.400 408.600 708.600 409.800 ;
        RECT 694.950 407.400 708.600 408.600 ;
        RECT 740.400 408.600 741.600 413.400 ;
        RECT 743.400 412.050 744.600 416.400 ;
        RECT 754.950 415.950 757.050 418.050 ;
        RECT 802.950 415.950 805.050 418.050 ;
        RECT 820.950 417.600 823.050 417.900 ;
        RECT 832.950 417.600 835.050 418.200 ;
        RECT 820.950 416.400 835.050 417.600 ;
        RECT 755.400 412.050 756.600 415.950 ;
        RECT 803.400 412.050 804.600 415.950 ;
        RECT 820.950 415.800 823.050 416.400 ;
        RECT 832.950 416.100 835.050 416.400 ;
        RECT 838.950 417.600 841.050 418.200 ;
        RECT 850.950 417.600 853.050 418.200 ;
        RECT 874.950 417.600 877.050 418.200 ;
        RECT 838.950 416.400 853.050 417.600 ;
        RECT 838.950 416.100 841.050 416.400 ;
        RECT 850.950 416.100 853.050 416.400 ;
        RECT 869.400 416.400 877.050 417.600 ;
        RECT 742.950 409.950 745.050 412.050 ;
        RECT 754.950 409.950 757.050 412.050 ;
        RECT 760.950 411.600 763.050 412.050 ;
        RECT 766.950 411.600 769.050 411.900 ;
        RECT 790.950 411.600 793.050 411.900 ;
        RECT 760.950 410.400 793.050 411.600 ;
        RECT 760.950 409.950 763.050 410.400 ;
        RECT 766.950 409.800 769.050 410.400 ;
        RECT 790.950 409.800 793.050 410.400 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 805.950 411.600 808.050 415.050 ;
        RECT 869.400 414.600 870.600 416.400 ;
        RECT 874.950 416.100 877.050 416.400 ;
        RECT 883.950 415.950 886.050 418.050 ;
        RECT 901.950 417.750 904.050 418.200 ;
        RECT 910.950 417.750 913.050 418.200 ;
        RECT 901.950 416.550 913.050 417.750 ;
        RECT 901.950 416.100 904.050 416.550 ;
        RECT 910.950 416.100 913.050 416.550 ;
        RECT 931.950 415.950 934.050 418.050 ;
        RECT 860.400 413.400 870.600 414.600 ;
        RECT 860.400 411.900 861.600 413.400 ;
        RECT 884.400 412.050 885.600 415.950 ;
        RECT 932.400 412.050 933.600 415.950 ;
        RECT 814.950 411.600 817.050 411.900 ;
        RECT 829.950 411.600 832.050 411.900 ;
        RECT 805.950 411.000 832.050 411.600 ;
        RECT 806.400 410.400 832.050 411.000 ;
        RECT 814.950 409.800 817.050 410.400 ;
        RECT 829.950 409.800 832.050 410.400 ;
        RECT 859.950 409.800 862.050 411.900 ;
        RECT 883.950 409.950 886.050 412.050 ;
        RECT 889.950 411.450 892.050 411.900 ;
        RECT 898.950 411.450 901.050 411.900 ;
        RECT 889.950 410.250 901.050 411.450 ;
        RECT 889.950 409.800 892.050 410.250 ;
        RECT 898.950 409.800 901.050 410.250 ;
        RECT 931.950 409.950 934.050 412.050 ;
        RECT 772.950 408.600 775.050 409.050 ;
        RECT 841.950 408.600 844.050 409.050 ;
        RECT 865.950 408.600 868.050 409.050 ;
        RECT 877.950 408.600 880.050 409.050 ;
        RECT 740.400 407.400 880.050 408.600 ;
        RECT 694.950 406.950 697.050 407.400 ;
        RECT 772.950 406.950 775.050 407.400 ;
        RECT 841.950 406.950 844.050 407.400 ;
        RECT 865.950 406.950 868.050 407.400 ;
        RECT 877.950 406.950 880.050 407.400 ;
        RECT 886.950 408.600 889.050 409.050 ;
        RECT 904.950 408.600 907.050 409.050 ;
        RECT 886.950 407.400 907.050 408.600 ;
        RECT 886.950 406.950 889.050 407.400 ;
        RECT 904.950 406.950 907.050 407.400 ;
        RECT 76.950 405.600 79.050 406.050 ;
        RECT 130.950 405.600 133.050 406.050 ;
        RECT 76.950 404.400 133.050 405.600 ;
        RECT 76.950 403.950 79.050 404.400 ;
        RECT 130.950 403.950 133.050 404.400 ;
        RECT 142.950 405.600 145.050 406.050 ;
        RECT 148.950 405.600 151.050 406.050 ;
        RECT 187.950 405.600 190.050 406.050 ;
        RECT 142.950 404.400 190.050 405.600 ;
        RECT 142.950 403.950 145.050 404.400 ;
        RECT 148.950 403.950 151.050 404.400 ;
        RECT 187.950 403.950 190.050 404.400 ;
        RECT 253.950 405.600 256.050 406.050 ;
        RECT 271.950 405.600 274.050 406.050 ;
        RECT 253.950 404.400 274.050 405.600 ;
        RECT 253.950 403.950 256.050 404.400 ;
        RECT 271.950 403.950 274.050 404.400 ;
        RECT 286.950 405.600 289.050 406.050 ;
        RECT 316.950 405.600 319.050 406.050 ;
        RECT 286.950 404.400 319.050 405.600 ;
        RECT 286.950 403.950 289.050 404.400 ;
        RECT 316.950 403.950 319.050 404.400 ;
        RECT 421.950 405.600 424.050 406.050 ;
        RECT 442.950 405.600 445.050 406.050 ;
        RECT 421.950 404.400 445.050 405.600 ;
        RECT 421.950 403.950 424.050 404.400 ;
        RECT 442.950 403.950 445.050 404.400 ;
        RECT 538.950 405.600 541.050 406.050 ;
        RECT 574.950 405.600 577.050 406.050 ;
        RECT 631.950 405.600 634.050 406.050 ;
        RECT 538.950 404.400 549.600 405.600 ;
        RECT 538.950 403.950 541.050 404.400 ;
        RECT 49.950 402.600 52.050 403.050 ;
        RECT 79.950 402.600 82.050 403.050 ;
        RECT 49.950 401.400 82.050 402.600 ;
        RECT 49.950 400.950 52.050 401.400 ;
        RECT 79.950 400.950 82.050 401.400 ;
        RECT 139.950 402.600 142.050 403.050 ;
        RECT 208.950 402.600 211.050 403.050 ;
        RECT 139.950 401.400 211.050 402.600 ;
        RECT 139.950 400.950 142.050 401.400 ;
        RECT 208.950 400.950 211.050 401.400 ;
        RECT 277.950 402.600 280.050 403.050 ;
        RECT 340.950 402.600 343.050 403.050 ;
        RECT 442.950 402.600 445.050 402.900 ;
        RECT 277.950 401.400 445.050 402.600 ;
        RECT 277.950 400.950 280.050 401.400 ;
        RECT 340.950 400.950 343.050 401.400 ;
        RECT 442.950 400.800 445.050 401.400 ;
        RECT 502.950 402.600 505.050 403.050 ;
        RECT 508.950 402.600 511.050 403.050 ;
        RECT 523.950 402.600 526.050 403.050 ;
        RECT 539.400 402.600 540.600 403.950 ;
        RECT 502.950 401.400 540.600 402.600 ;
        RECT 548.400 402.600 549.600 404.400 ;
        RECT 574.950 404.400 634.050 405.600 ;
        RECT 574.950 403.950 577.050 404.400 ;
        RECT 631.950 403.950 634.050 404.400 ;
        RECT 667.950 405.600 670.050 406.050 ;
        RECT 691.950 405.600 694.050 406.050 ;
        RECT 667.950 404.400 694.050 405.600 ;
        RECT 667.950 403.950 670.050 404.400 ;
        RECT 691.950 403.950 694.050 404.400 ;
        RECT 748.950 405.600 751.050 406.050 ;
        RECT 769.950 405.600 772.050 406.050 ;
        RECT 748.950 404.400 772.050 405.600 ;
        RECT 748.950 403.950 751.050 404.400 ;
        RECT 769.950 403.950 772.050 404.400 ;
        RECT 775.950 405.600 778.050 406.050 ;
        RECT 796.950 405.600 799.050 406.050 ;
        RECT 835.950 405.600 838.050 406.050 ;
        RECT 775.950 404.400 838.050 405.600 ;
        RECT 775.950 403.950 778.050 404.400 ;
        RECT 796.950 403.950 799.050 404.400 ;
        RECT 835.950 403.950 838.050 404.400 ;
        RECT 847.950 405.600 850.050 406.050 ;
        RECT 871.950 405.600 874.050 406.050 ;
        RECT 847.950 404.400 874.050 405.600 ;
        RECT 847.950 403.950 850.050 404.400 ;
        RECT 871.950 403.950 874.050 404.400 ;
        RECT 580.950 402.600 583.050 403.050 ;
        RECT 548.400 401.400 583.050 402.600 ;
        RECT 502.950 400.950 505.050 401.400 ;
        RECT 508.950 400.950 511.050 401.400 ;
        RECT 523.950 400.950 526.050 401.400 ;
        RECT 580.950 400.950 583.050 401.400 ;
        RECT 589.950 402.600 592.050 403.050 ;
        RECT 625.950 402.600 628.050 403.050 ;
        RECT 589.950 401.400 628.050 402.600 ;
        RECT 589.950 400.950 592.050 401.400 ;
        RECT 625.950 400.950 628.050 401.400 ;
        RECT 646.950 402.600 649.050 403.050 ;
        RECT 694.950 402.600 697.050 403.050 ;
        RECT 646.950 401.400 697.050 402.600 ;
        RECT 646.950 400.950 649.050 401.400 ;
        RECT 694.950 400.950 697.050 401.400 ;
        RECT 712.950 402.600 715.050 403.050 ;
        RECT 739.950 402.600 742.050 403.050 ;
        RECT 814.800 402.600 816.900 403.050 ;
        RECT 712.950 401.400 742.050 402.600 ;
        RECT 712.950 400.950 715.050 401.400 ;
        RECT 739.950 400.950 742.050 401.400 ;
        RECT 779.400 401.400 816.900 402.600 ;
        RECT 779.400 400.050 780.600 401.400 ;
        RECT 814.800 400.950 816.900 401.400 ;
        RECT 817.950 402.600 820.050 403.050 ;
        RECT 835.950 402.600 838.050 402.900 ;
        RECT 817.950 401.400 838.050 402.600 ;
        RECT 817.950 400.950 820.050 401.400 ;
        RECT 835.950 400.800 838.050 401.400 ;
        RECT 262.950 399.600 265.050 400.050 ;
        RECT 286.950 399.600 289.050 400.050 ;
        RECT 262.950 398.400 289.050 399.600 ;
        RECT 262.950 397.950 265.050 398.400 ;
        RECT 286.950 397.950 289.050 398.400 ;
        RECT 322.950 399.600 325.050 400.050 ;
        RECT 421.950 399.600 424.050 400.050 ;
        RECT 322.950 398.400 424.050 399.600 ;
        RECT 322.950 397.950 325.050 398.400 ;
        RECT 421.950 397.950 424.050 398.400 ;
        RECT 544.950 399.600 547.050 400.050 ;
        RECT 598.950 399.600 601.050 400.050 ;
        RECT 544.950 398.400 601.050 399.600 ;
        RECT 544.950 397.950 547.050 398.400 ;
        RECT 598.950 397.950 601.050 398.400 ;
        RECT 610.950 399.600 613.050 400.050 ;
        RECT 622.950 399.600 625.050 400.050 ;
        RECT 697.950 399.600 700.050 400.050 ;
        RECT 610.950 398.400 625.050 399.600 ;
        RECT 610.950 397.950 613.050 398.400 ;
        RECT 622.950 397.950 625.050 398.400 ;
        RECT 626.400 398.400 700.050 399.600 ;
        RECT 40.950 396.600 43.050 397.050 ;
        RECT 67.950 396.600 70.050 397.050 ;
        RECT 151.950 396.600 154.050 397.050 ;
        RECT 40.950 395.400 154.050 396.600 ;
        RECT 40.950 394.950 43.050 395.400 ;
        RECT 67.950 394.950 70.050 395.400 ;
        RECT 151.950 394.950 154.050 395.400 ;
        RECT 184.950 396.600 187.050 397.050 ;
        RECT 223.950 396.600 226.050 397.050 ;
        RECT 184.950 395.400 226.050 396.600 ;
        RECT 184.950 394.950 187.050 395.400 ;
        RECT 223.950 394.950 226.050 395.400 ;
        RECT 325.950 396.600 328.050 397.050 ;
        RECT 376.950 396.600 379.050 397.050 ;
        RECT 325.950 395.400 379.050 396.600 ;
        RECT 325.950 394.950 328.050 395.400 ;
        RECT 376.950 394.950 379.050 395.400 ;
        RECT 550.950 396.600 553.050 397.050 ;
        RECT 595.950 396.600 598.050 397.050 ;
        RECT 626.400 396.600 627.600 398.400 ;
        RECT 697.950 397.950 700.050 398.400 ;
        RECT 718.950 399.600 721.050 400.050 ;
        RECT 778.950 399.600 781.050 400.050 ;
        RECT 718.950 398.400 781.050 399.600 ;
        RECT 718.950 397.950 721.050 398.400 ;
        RECT 778.950 397.950 781.050 398.400 ;
        RECT 784.950 399.600 787.050 400.050 ;
        RECT 838.950 399.600 841.050 400.050 ;
        RECT 784.950 398.400 841.050 399.600 ;
        RECT 784.950 397.950 787.050 398.400 ;
        RECT 838.950 397.950 841.050 398.400 ;
        RECT 847.950 399.600 850.050 400.050 ;
        RECT 883.950 399.600 886.050 400.050 ;
        RECT 847.950 398.400 886.050 399.600 ;
        RECT 847.950 397.950 850.050 398.400 ;
        RECT 883.950 397.950 886.050 398.400 ;
        RECT 550.950 395.400 627.600 396.600 ;
        RECT 676.950 396.600 679.050 397.050 ;
        RECT 715.950 396.600 718.050 397.050 ;
        RECT 676.950 395.400 718.050 396.600 ;
        RECT 550.950 394.950 553.050 395.400 ;
        RECT 595.950 394.950 598.050 395.400 ;
        RECT 676.950 394.950 679.050 395.400 ;
        RECT 715.950 394.950 718.050 395.400 ;
        RECT 724.950 396.600 727.050 397.050 ;
        RECT 766.950 396.600 769.050 397.050 ;
        RECT 805.950 396.600 808.050 397.050 ;
        RECT 817.800 396.600 819.900 397.050 ;
        RECT 724.950 395.400 769.050 396.600 ;
        RECT 724.950 394.950 727.050 395.400 ;
        RECT 766.950 394.950 769.050 395.400 ;
        RECT 803.400 395.400 819.900 396.600 ;
        RECT 112.950 393.600 115.050 394.050 ;
        RECT 160.950 393.600 163.050 394.050 ;
        RECT 112.950 392.400 163.050 393.600 ;
        RECT 112.950 391.950 115.050 392.400 ;
        RECT 160.950 391.950 163.050 392.400 ;
        RECT 565.950 393.600 568.050 394.050 ;
        RECT 574.950 393.600 577.050 394.050 ;
        RECT 565.950 392.400 577.050 393.600 ;
        RECT 565.950 391.950 568.050 392.400 ;
        RECT 574.950 391.950 577.050 392.400 ;
        RECT 607.950 393.600 610.050 394.050 ;
        RECT 646.950 393.600 649.050 394.050 ;
        RECT 607.950 392.400 649.050 393.600 ;
        RECT 607.950 391.950 610.050 392.400 ;
        RECT 646.950 391.950 649.050 392.400 ;
        RECT 778.950 393.600 781.050 394.050 ;
        RECT 803.400 393.600 804.600 395.400 ;
        RECT 805.950 394.950 808.050 395.400 ;
        RECT 817.800 394.950 819.900 395.400 ;
        RECT 820.950 396.600 823.050 397.050 ;
        RECT 910.950 396.600 913.050 397.050 ;
        RECT 919.950 396.600 922.050 397.050 ;
        RECT 820.950 395.400 922.050 396.600 ;
        RECT 820.950 394.950 823.050 395.400 ;
        RECT 910.950 394.950 913.050 395.400 ;
        RECT 919.950 394.950 922.050 395.400 ;
        RECT 883.950 393.600 886.050 394.050 ;
        RECT 778.950 392.400 804.600 393.600 ;
        RECT 851.400 392.400 886.050 393.600 ;
        RECT 778.950 391.950 781.050 392.400 ;
        RECT 28.950 390.600 31.050 391.050 ;
        RECT 184.950 390.600 187.050 391.050 ;
        RECT 28.950 389.400 187.050 390.600 ;
        RECT 28.950 388.950 31.050 389.400 ;
        RECT 184.950 388.950 187.050 389.400 ;
        RECT 313.950 390.600 316.050 391.050 ;
        RECT 346.950 390.600 349.050 391.050 ;
        RECT 394.950 390.600 397.050 391.050 ;
        RECT 409.950 390.600 412.050 391.050 ;
        RECT 457.950 390.600 460.050 391.050 ;
        RECT 313.950 389.400 460.050 390.600 ;
        RECT 313.950 388.950 316.050 389.400 ;
        RECT 346.950 388.950 349.050 389.400 ;
        RECT 394.950 388.950 397.050 389.400 ;
        RECT 409.950 388.950 412.050 389.400 ;
        RECT 457.950 388.950 460.050 389.400 ;
        RECT 547.950 390.600 550.050 391.050 ;
        RECT 577.950 390.600 580.050 391.050 ;
        RECT 661.950 390.600 664.050 391.050 ;
        RECT 667.950 390.600 670.050 391.050 ;
        RECT 547.950 389.400 670.050 390.600 ;
        RECT 547.950 388.950 550.050 389.400 ;
        RECT 577.950 388.950 580.050 389.400 ;
        RECT 661.950 388.950 664.050 389.400 ;
        RECT 667.950 388.950 670.050 389.400 ;
        RECT 691.950 390.600 694.050 391.050 ;
        RECT 718.950 390.600 721.050 391.050 ;
        RECT 691.950 389.400 721.050 390.600 ;
        RECT 691.950 388.950 694.050 389.400 ;
        RECT 718.950 388.950 721.050 389.400 ;
        RECT 724.950 390.600 727.050 391.050 ;
        RECT 754.950 390.600 757.050 391.050 ;
        RECT 724.950 389.400 757.050 390.600 ;
        RECT 724.950 388.950 727.050 389.400 ;
        RECT 754.950 388.950 757.050 389.400 ;
        RECT 805.950 390.600 808.050 391.050 ;
        RECT 851.400 390.600 852.600 392.400 ;
        RECT 883.950 391.950 886.050 392.400 ;
        RECT 805.950 389.400 852.600 390.600 ;
        RECT 805.950 388.950 808.050 389.400 ;
        RECT 40.950 387.600 43.050 388.050 ;
        RECT 55.950 387.600 58.050 388.050 ;
        RECT 40.950 386.400 58.050 387.600 ;
        RECT 40.950 385.950 43.050 386.400 ;
        RECT 55.950 385.950 58.050 386.400 ;
        RECT 157.950 387.600 160.050 388.050 ;
        RECT 163.950 387.600 166.050 388.050 ;
        RECT 157.950 386.400 166.050 387.600 ;
        RECT 157.950 385.950 160.050 386.400 ;
        RECT 163.950 385.950 166.050 386.400 ;
        RECT 214.950 387.600 217.050 388.050 ;
        RECT 220.950 387.600 223.050 388.050 ;
        RECT 271.950 387.600 274.050 388.050 ;
        RECT 295.950 387.600 298.050 388.050 ;
        RECT 214.950 386.400 298.050 387.600 ;
        RECT 214.950 385.950 217.050 386.400 ;
        RECT 220.950 385.950 223.050 386.400 ;
        RECT 271.950 385.950 274.050 386.400 ;
        RECT 295.950 385.950 298.050 386.400 ;
        RECT 388.950 387.600 391.050 388.050 ;
        RECT 415.950 387.600 418.050 388.050 ;
        RECT 388.950 386.400 418.050 387.600 ;
        RECT 388.950 385.950 391.050 386.400 ;
        RECT 415.950 385.950 418.050 386.400 ;
        RECT 505.950 387.600 508.050 388.050 ;
        RECT 562.950 387.600 565.050 388.050 ;
        RECT 505.950 386.400 565.050 387.600 ;
        RECT 505.950 385.950 508.050 386.400 ;
        RECT 562.950 385.950 565.050 386.400 ;
        RECT 580.950 387.600 583.050 388.050 ;
        RECT 625.950 387.600 628.050 388.050 ;
        RECT 580.950 386.400 628.050 387.600 ;
        RECT 580.950 385.950 583.050 386.400 ;
        RECT 625.950 385.950 628.050 386.400 ;
        RECT 637.950 387.600 640.050 388.050 ;
        RECT 661.950 387.600 664.050 387.900 ;
        RECT 637.950 386.400 664.050 387.600 ;
        RECT 637.950 385.950 640.050 386.400 ;
        RECT 661.950 385.800 664.050 386.400 ;
        RECT 697.950 387.600 700.050 388.050 ;
        RECT 715.950 387.600 718.050 388.050 ;
        RECT 697.950 386.400 718.050 387.600 ;
        RECT 697.950 385.950 700.050 386.400 ;
        RECT 715.950 385.950 718.050 386.400 ;
        RECT 721.950 387.600 724.050 388.050 ;
        RECT 772.950 387.600 775.050 388.050 ;
        RECT 721.950 386.400 775.050 387.600 ;
        RECT 721.950 385.950 724.050 386.400 ;
        RECT 772.950 385.950 775.050 386.400 ;
        RECT 814.950 387.600 817.050 388.050 ;
        RECT 853.950 387.600 856.050 388.050 ;
        RECT 814.950 386.400 856.050 387.600 ;
        RECT 814.950 385.950 817.050 386.400 ;
        RECT 853.950 385.950 856.050 386.400 ;
        RECT 121.950 384.600 124.050 385.050 ;
        RECT 154.950 384.600 157.050 385.050 ;
        RECT 121.950 383.400 157.050 384.600 ;
        RECT 121.950 382.950 124.050 383.400 ;
        RECT 154.950 382.950 157.050 383.400 ;
        RECT 217.950 384.600 220.050 385.050 ;
        RECT 241.950 384.600 244.050 385.050 ;
        RECT 217.950 383.400 244.050 384.600 ;
        RECT 217.950 382.950 220.050 383.400 ;
        RECT 241.950 382.950 244.050 383.400 ;
        RECT 301.950 384.600 304.050 385.050 ;
        RECT 319.950 384.600 322.050 385.050 ;
        RECT 466.950 384.600 469.050 385.050 ;
        RECT 301.950 383.400 469.050 384.600 ;
        RECT 301.950 382.950 304.050 383.400 ;
        RECT 319.950 382.950 322.050 383.400 ;
        RECT 466.950 382.950 469.050 383.400 ;
        RECT 520.950 384.600 523.050 385.050 ;
        RECT 541.950 384.600 544.050 385.050 ;
        RECT 520.950 383.400 544.050 384.600 ;
        RECT 520.950 382.950 523.050 383.400 ;
        RECT 541.950 382.950 544.050 383.400 ;
        RECT 601.950 384.600 604.050 385.050 ;
        RECT 712.950 384.600 715.050 385.050 ;
        RECT 727.950 384.600 730.050 385.050 ;
        RECT 601.950 383.400 730.050 384.600 ;
        RECT 601.950 382.950 604.050 383.400 ;
        RECT 712.950 382.950 715.050 383.400 ;
        RECT 727.950 382.950 730.050 383.400 ;
        RECT 808.950 384.600 811.050 385.050 ;
        RECT 829.950 384.600 832.050 385.050 ;
        RECT 808.950 383.400 832.050 384.600 ;
        RECT 808.950 382.950 811.050 383.400 ;
        RECT 829.950 382.950 832.050 383.400 ;
        RECT 106.950 381.600 109.050 382.050 ;
        RECT 190.950 381.600 193.050 382.050 ;
        RECT 106.950 380.400 193.050 381.600 ;
        RECT 106.950 379.950 109.050 380.400 ;
        RECT 190.950 379.950 193.050 380.400 ;
        RECT 280.950 381.600 283.050 382.050 ;
        RECT 325.950 381.600 328.050 382.050 ;
        RECT 280.950 380.400 328.050 381.600 ;
        RECT 280.950 379.950 283.050 380.400 ;
        RECT 325.950 379.950 328.050 380.400 ;
        RECT 331.950 381.600 334.050 382.050 ;
        RECT 379.950 381.600 382.050 382.050 ;
        RECT 331.950 380.400 382.050 381.600 ;
        RECT 467.400 381.600 468.600 382.950 ;
        RECT 544.950 381.600 547.050 382.050 ;
        RECT 467.400 380.400 547.050 381.600 ;
        RECT 331.950 379.950 334.050 380.400 ;
        RECT 379.950 379.950 382.050 380.400 ;
        RECT 544.950 379.950 547.050 380.400 ;
        RECT 586.950 381.600 589.050 382.050 ;
        RECT 610.950 381.600 613.050 382.050 ;
        RECT 643.950 381.600 646.050 382.050 ;
        RECT 586.950 380.400 646.050 381.600 ;
        RECT 586.950 379.950 589.050 380.400 ;
        RECT 610.950 379.950 613.050 380.400 ;
        RECT 643.950 379.950 646.050 380.400 ;
        RECT 688.950 381.600 691.050 382.050 ;
        RECT 694.950 381.600 697.050 382.050 ;
        RECT 706.950 381.600 709.050 382.050 ;
        RECT 688.950 380.400 709.050 381.600 ;
        RECT 688.950 379.950 691.050 380.400 ;
        RECT 694.950 379.950 697.050 380.400 ;
        RECT 706.950 379.950 709.050 380.400 ;
        RECT 160.950 378.600 163.050 379.050 ;
        RECT 175.950 378.600 178.050 379.050 ;
        RECT 160.950 377.400 178.050 378.600 ;
        RECT 160.950 376.950 163.050 377.400 ;
        RECT 175.950 376.950 178.050 377.400 ;
        RECT 205.950 378.600 208.050 379.050 ;
        RECT 217.950 378.600 220.050 379.050 ;
        RECT 232.950 378.600 235.050 379.050 ;
        RECT 205.950 377.400 235.050 378.600 ;
        RECT 205.950 376.950 208.050 377.400 ;
        RECT 217.950 376.950 220.050 377.400 ;
        RECT 232.950 376.950 235.050 377.400 ;
        RECT 277.950 378.600 280.050 379.050 ;
        RECT 304.950 378.600 307.050 379.050 ;
        RECT 277.950 377.400 307.050 378.600 ;
        RECT 277.950 376.950 280.050 377.400 ;
        RECT 304.950 376.950 307.050 377.400 ;
        RECT 361.950 378.600 364.050 379.050 ;
        RECT 376.950 378.600 379.050 379.050 ;
        RECT 361.950 377.400 379.050 378.600 ;
        RECT 361.950 376.950 364.050 377.400 ;
        RECT 376.950 376.950 379.050 377.400 ;
        RECT 394.950 378.600 397.050 379.050 ;
        RECT 430.950 378.600 433.050 379.050 ;
        RECT 394.950 377.400 433.050 378.600 ;
        RECT 394.950 376.950 397.050 377.400 ;
        RECT 430.950 376.950 433.050 377.400 ;
        RECT 454.950 378.600 457.050 379.050 ;
        RECT 550.950 378.600 553.050 379.050 ;
        RECT 607.950 378.600 610.050 379.050 ;
        RECT 454.950 377.400 553.050 378.600 ;
        RECT 454.950 376.950 457.050 377.400 ;
        RECT 550.950 376.950 553.050 377.400 ;
        RECT 596.400 377.400 610.050 378.600 ;
        RECT 34.950 375.600 37.050 376.050 ;
        RECT 43.950 375.600 46.050 376.050 ;
        RECT 76.950 375.600 79.050 376.050 ;
        RECT 34.950 374.400 79.050 375.600 ;
        RECT 34.950 373.950 37.050 374.400 ;
        RECT 43.950 373.950 46.050 374.400 ;
        RECT 76.950 373.950 79.050 374.400 ;
        RECT 121.950 375.600 124.050 376.050 ;
        RECT 130.950 375.600 133.050 376.200 ;
        RECT 121.950 374.400 133.050 375.600 ;
        RECT 121.950 373.950 124.050 374.400 ;
        RECT 130.950 374.100 133.050 374.400 ;
        RECT 151.950 375.600 154.050 376.050 ;
        RECT 208.950 375.600 211.050 376.050 ;
        RECT 235.950 375.600 238.050 376.050 ;
        RECT 151.950 374.400 171.600 375.600 ;
        RECT 151.950 373.950 154.050 374.400 ;
        RECT 46.950 372.750 49.050 373.200 ;
        RECT 52.950 372.750 55.050 373.200 ;
        RECT 46.950 371.550 55.050 372.750 ;
        RECT 46.950 371.100 49.050 371.550 ;
        RECT 52.950 371.100 55.050 371.550 ;
        RECT 58.950 372.600 61.050 373.200 ;
        RECT 67.950 372.600 72.000 373.050 ;
        RECT 58.950 371.400 66.600 372.600 ;
        RECT 58.950 371.100 61.050 371.400 ;
        RECT 65.400 367.050 66.600 371.400 ;
        RECT 67.950 370.950 72.600 372.600 ;
        RECT 71.400 369.900 72.600 370.950 ;
        RECT 70.950 367.800 73.050 369.900 ;
        RECT 65.400 365.400 70.050 367.050 ;
        RECT 66.000 364.950 70.050 365.400 ;
        RECT 127.950 366.600 130.050 367.050 ;
        RECT 145.950 366.600 148.050 366.900 ;
        RECT 166.800 366.600 168.900 367.050 ;
        RECT 170.400 366.900 171.600 374.400 ;
        RECT 208.950 374.400 238.050 375.600 ;
        RECT 208.950 373.950 211.050 374.400 ;
        RECT 235.950 373.950 238.050 374.400 ;
        RECT 307.950 375.600 310.050 376.050 ;
        RECT 340.950 375.600 343.050 376.050 ;
        RECT 307.950 374.400 343.050 375.600 ;
        RECT 307.950 373.950 310.050 374.400 ;
        RECT 340.950 373.950 343.050 374.400 ;
        RECT 562.950 375.600 565.050 376.050 ;
        RECT 596.400 375.600 597.600 377.400 ;
        RECT 607.950 376.950 610.050 377.400 ;
        RECT 631.950 378.600 634.050 379.050 ;
        RECT 673.950 378.600 676.050 379.050 ;
        RECT 631.950 377.400 676.050 378.600 ;
        RECT 631.950 376.950 634.050 377.400 ;
        RECT 673.950 376.950 676.050 377.400 ;
        RECT 724.950 378.600 727.050 379.050 ;
        RECT 733.950 378.600 736.050 379.050 ;
        RECT 793.950 378.600 796.050 379.050 ;
        RECT 811.950 378.600 814.050 379.050 ;
        RECT 724.950 377.400 814.050 378.600 ;
        RECT 724.950 376.950 727.050 377.400 ;
        RECT 733.950 376.950 736.050 377.400 ;
        RECT 793.950 376.950 796.050 377.400 ;
        RECT 811.950 376.950 814.050 377.400 ;
        RECT 835.950 378.600 838.050 379.050 ;
        RECT 850.950 378.600 853.050 379.050 ;
        RECT 835.950 377.400 853.050 378.600 ;
        RECT 835.950 376.950 838.050 377.400 ;
        RECT 850.950 376.950 853.050 377.400 ;
        RECT 898.950 378.600 901.050 379.050 ;
        RECT 913.950 378.600 916.050 379.050 ;
        RECT 898.950 377.400 916.050 378.600 ;
        RECT 898.950 376.950 901.050 377.400 ;
        RECT 913.950 376.950 916.050 377.400 ;
        RECT 562.950 374.400 597.600 375.600 ;
        RECT 622.950 375.600 625.050 376.050 ;
        RECT 688.950 375.600 691.050 376.050 ;
        RECT 700.950 375.600 703.050 376.050 ;
        RECT 622.950 374.400 630.600 375.600 ;
        RECT 562.950 373.950 565.050 374.400 ;
        RECT 622.950 373.950 625.050 374.400 ;
        RECT 172.950 372.600 175.050 373.200 ;
        RECT 184.950 372.600 187.050 373.200 ;
        RECT 172.950 371.400 187.050 372.600 ;
        RECT 172.950 371.100 175.050 371.400 ;
        RECT 184.950 371.100 187.050 371.400 ;
        RECT 196.950 370.950 199.050 373.050 ;
        RECT 205.950 372.600 208.050 373.050 ;
        RECT 211.950 372.600 214.050 373.200 ;
        RECT 229.950 372.600 232.050 373.200 ;
        RECT 205.950 371.400 214.050 372.600 ;
        RECT 205.950 370.950 208.050 371.400 ;
        RECT 211.950 371.100 214.050 371.400 ;
        RECT 224.400 371.400 232.050 372.600 ;
        RECT 127.950 365.400 148.050 366.600 ;
        RECT 127.950 364.950 130.050 365.400 ;
        RECT 145.950 364.800 148.050 365.400 ;
        RECT 152.400 365.400 168.900 366.600 ;
        RECT 22.950 363.600 25.050 364.050 ;
        RECT 55.950 363.600 58.050 364.050 ;
        RECT 85.950 363.600 88.050 364.050 ;
        RECT 124.950 363.600 127.050 364.050 ;
        RECT 152.400 363.600 153.600 365.400 ;
        RECT 166.800 364.950 168.900 365.400 ;
        RECT 169.950 364.800 172.050 366.900 ;
        RECT 22.950 362.400 153.600 363.600 ;
        RECT 154.950 363.600 157.050 364.050 ;
        RECT 163.950 363.600 166.050 364.050 ;
        RECT 154.950 362.400 166.050 363.600 ;
        RECT 197.400 363.600 198.600 370.950 ;
        RECT 224.400 369.600 225.600 371.400 ;
        RECT 229.950 371.100 232.050 371.400 ;
        RECT 235.950 371.100 238.050 373.200 ;
        RECT 247.950 372.600 250.050 373.200 ;
        RECT 256.950 372.600 259.050 373.050 ;
        RECT 247.950 371.400 259.050 372.600 ;
        RECT 247.950 371.100 250.050 371.400 ;
        RECT 221.400 368.400 225.600 369.600 ;
        RECT 221.400 364.050 222.600 368.400 ;
        RECT 236.400 366.600 237.600 371.100 ;
        RECT 256.950 370.950 259.050 371.400 ;
        RECT 265.950 372.750 268.050 373.200 ;
        RECT 274.950 372.750 277.050 373.200 ;
        RECT 265.950 372.600 277.050 372.750 ;
        RECT 289.950 372.600 292.050 373.200 ;
        RECT 265.950 371.550 292.050 372.600 ;
        RECT 265.950 371.100 268.050 371.550 ;
        RECT 274.950 371.400 292.050 371.550 ;
        RECT 274.950 371.100 277.050 371.400 ;
        RECT 289.950 371.100 292.050 371.400 ;
        RECT 304.950 372.600 307.050 373.050 ;
        RECT 322.950 372.600 325.050 373.050 ;
        RECT 304.950 371.400 325.050 372.600 ;
        RECT 304.950 370.950 307.050 371.400 ;
        RECT 322.950 370.950 325.050 371.400 ;
        RECT 370.950 372.600 373.050 373.200 ;
        RECT 394.800 372.600 396.900 373.200 ;
        RECT 370.950 371.400 396.900 372.600 ;
        RECT 370.950 371.100 373.050 371.400 ;
        RECT 394.800 371.100 396.900 371.400 ;
        RECT 355.950 369.600 358.050 370.050 ;
        RECT 397.950 369.600 400.050 373.050 ;
        RECT 418.950 372.600 421.050 373.200 ;
        RECT 436.950 372.600 439.050 373.200 ;
        RECT 448.950 372.600 451.050 373.200 ;
        RECT 418.950 371.400 451.050 372.600 ;
        RECT 418.950 371.100 421.050 371.400 ;
        RECT 436.950 371.100 439.050 371.400 ;
        RECT 448.950 371.100 451.050 371.400 ;
        RECT 481.950 372.600 484.050 373.200 ;
        RECT 487.950 372.750 490.050 373.200 ;
        RECT 493.950 372.750 496.050 373.200 ;
        RECT 487.950 372.600 496.050 372.750 ;
        RECT 481.950 371.550 496.050 372.600 ;
        RECT 481.950 371.400 490.050 371.550 ;
        RECT 481.950 371.100 484.050 371.400 ;
        RECT 487.950 371.100 490.050 371.400 ;
        RECT 493.950 371.100 496.050 371.550 ;
        RECT 499.950 372.600 502.050 373.200 ;
        RECT 511.950 372.600 514.050 373.200 ;
        RECT 535.950 372.600 538.050 373.200 ;
        RECT 559.950 372.600 562.050 373.050 ;
        RECT 499.950 371.400 538.050 372.600 ;
        RECT 499.950 371.100 502.050 371.400 ;
        RECT 511.950 371.100 514.050 371.400 ;
        RECT 535.950 371.100 538.050 371.400 ;
        RECT 551.400 371.400 562.050 372.600 ;
        RECT 355.950 369.000 400.050 369.600 ;
        RECT 442.950 369.600 445.050 370.050 ;
        RECT 551.400 369.600 552.600 371.400 ;
        RECT 559.950 370.950 562.050 371.400 ;
        RECT 568.950 372.600 571.050 373.050 ;
        RECT 589.950 372.600 592.050 373.050 ;
        RECT 598.950 372.600 601.050 373.050 ;
        RECT 568.950 371.400 588.600 372.600 ;
        RECT 568.950 370.950 571.050 371.400 ;
        RECT 355.950 368.400 399.600 369.000 ;
        RECT 442.950 368.400 552.600 369.600 ;
        RECT 553.950 369.600 556.050 370.050 ;
        RECT 574.950 369.600 577.050 370.050 ;
        RECT 553.950 368.400 577.050 369.600 ;
        RECT 587.400 369.600 588.600 371.400 ;
        RECT 589.950 371.400 601.050 372.600 ;
        RECT 589.950 370.950 592.050 371.400 ;
        RECT 598.950 370.950 601.050 371.400 ;
        RECT 604.950 372.600 607.050 373.200 ;
        RECT 616.950 372.600 619.050 373.050 ;
        RECT 604.950 371.400 619.050 372.600 ;
        RECT 629.400 372.600 630.600 374.400 ;
        RECT 688.950 374.400 703.050 375.600 ;
        RECT 688.950 373.950 691.050 374.400 ;
        RECT 700.950 373.950 703.050 374.400 ;
        RECT 838.950 373.950 841.050 376.050 ;
        RECT 631.950 372.600 634.050 373.050 ;
        RECT 649.950 372.600 652.050 373.200 ;
        RECT 629.400 371.400 652.050 372.600 ;
        RECT 604.950 371.100 607.050 371.400 ;
        RECT 616.950 370.950 619.050 371.400 ;
        RECT 631.950 370.950 634.050 371.400 ;
        RECT 649.950 371.100 652.050 371.400 ;
        RECT 661.950 371.100 664.050 373.200 ;
        RECT 667.950 372.600 670.050 373.200 ;
        RECT 682.950 372.600 685.050 373.200 ;
        RECT 738.000 372.600 742.050 373.050 ;
        RECT 667.950 371.400 685.050 372.600 ;
        RECT 667.950 371.100 670.050 371.400 ;
        RECT 682.950 371.100 685.050 371.400 ;
        RECT 662.400 369.600 663.600 371.100 ;
        RECT 737.400 370.950 742.050 372.600 ;
        RECT 748.950 371.100 751.050 373.200 ;
        RECT 760.950 372.750 763.050 373.200 ;
        RECT 766.950 372.750 769.050 373.200 ;
        RECT 760.950 371.550 769.050 372.750 ;
        RECT 760.950 371.100 763.050 371.550 ;
        RECT 766.950 371.100 769.050 371.550 ;
        RECT 587.400 368.400 594.600 369.600 ;
        RECT 662.400 368.400 690.600 369.600 ;
        RECT 355.950 367.950 358.050 368.400 ;
        RECT 442.950 367.950 445.050 368.400 ;
        RECT 553.950 367.950 556.050 368.400 ;
        RECT 574.950 367.950 577.050 368.400 ;
        RECT 250.950 366.600 253.050 366.900 ;
        RECT 236.400 365.400 253.050 366.600 ;
        RECT 250.950 364.800 253.050 365.400 ;
        RECT 256.950 366.450 259.050 366.900 ;
        RECT 262.950 366.450 265.050 366.900 ;
        RECT 256.950 365.250 265.050 366.450 ;
        RECT 256.950 364.800 259.050 365.250 ;
        RECT 262.950 364.800 265.050 365.250 ;
        RECT 268.950 366.600 271.050 366.900 ;
        RECT 280.950 366.600 283.050 367.050 ;
        RECT 268.950 365.400 283.050 366.600 ;
        RECT 268.950 364.800 271.050 365.400 ;
        RECT 280.950 364.950 283.050 365.400 ;
        RECT 298.950 366.600 301.050 367.050 ;
        RECT 328.950 366.600 331.050 366.900 ;
        RECT 298.950 365.400 331.050 366.600 ;
        RECT 298.950 364.950 301.050 365.400 ;
        RECT 328.950 364.800 331.050 365.400 ;
        RECT 340.950 366.450 343.050 366.900 ;
        RECT 367.950 366.450 370.050 366.900 ;
        RECT 340.950 365.250 370.050 366.450 ;
        RECT 340.950 364.800 343.050 365.250 ;
        RECT 367.950 364.800 370.050 365.250 ;
        RECT 382.950 366.600 385.050 367.050 ;
        RECT 400.950 366.600 403.050 367.050 ;
        RECT 382.950 365.400 403.050 366.600 ;
        RECT 382.950 364.950 385.050 365.400 ;
        RECT 400.950 364.950 403.050 365.400 ;
        RECT 415.950 366.450 418.050 366.900 ;
        RECT 424.950 366.450 427.050 366.900 ;
        RECT 415.950 365.250 427.050 366.450 ;
        RECT 415.950 364.800 418.050 365.250 ;
        RECT 424.950 364.800 427.050 365.250 ;
        RECT 457.950 366.600 460.050 366.900 ;
        RECT 466.950 366.600 469.050 366.900 ;
        RECT 457.950 366.450 469.050 366.600 ;
        RECT 472.950 366.450 475.050 366.900 ;
        RECT 457.950 365.400 475.050 366.450 ;
        RECT 457.950 364.800 460.050 365.400 ;
        RECT 466.950 365.250 475.050 365.400 ;
        RECT 466.950 364.800 469.050 365.250 ;
        RECT 472.950 364.800 475.050 365.250 ;
        RECT 478.950 366.600 481.050 366.900 ;
        RECT 526.950 366.600 529.050 367.050 ;
        RECT 478.950 365.400 529.050 366.600 ;
        RECT 478.950 364.800 481.050 365.400 ;
        RECT 526.950 364.950 529.050 365.400 ;
        RECT 544.950 366.450 547.050 366.900 ;
        RECT 550.950 366.450 553.050 366.900 ;
        RECT 544.950 365.250 553.050 366.450 ;
        RECT 544.950 364.800 547.050 365.250 ;
        RECT 550.950 364.800 553.050 365.250 ;
        RECT 593.400 364.050 594.600 368.400 ;
        RECT 595.950 366.450 598.050 367.050 ;
        RECT 601.950 366.450 604.050 366.900 ;
        RECT 595.950 365.250 604.050 366.450 ;
        RECT 595.950 364.950 598.050 365.250 ;
        RECT 601.950 364.800 604.050 365.250 ;
        RECT 623.400 365.400 648.600 366.600 ;
        RECT 211.950 363.600 214.050 364.050 ;
        RECT 197.400 362.400 214.050 363.600 ;
        RECT 22.950 361.950 25.050 362.400 ;
        RECT 55.950 361.950 58.050 362.400 ;
        RECT 85.950 361.950 88.050 362.400 ;
        RECT 124.950 361.950 127.050 362.400 ;
        RECT 154.950 361.950 157.050 362.400 ;
        RECT 163.950 361.950 166.050 362.400 ;
        RECT 211.950 361.950 214.050 362.400 ;
        RECT 217.950 362.400 222.600 364.050 ;
        RECT 226.950 363.600 229.050 364.050 ;
        RECT 232.950 363.600 235.050 364.050 ;
        RECT 226.950 362.400 235.050 363.600 ;
        RECT 593.400 363.900 597.000 364.050 ;
        RECT 593.400 362.400 598.050 363.900 ;
        RECT 217.950 361.950 222.000 362.400 ;
        RECT 226.950 361.950 229.050 362.400 ;
        RECT 232.950 361.950 235.050 362.400 ;
        RECT 594.000 361.950 598.050 362.400 ;
        RECT 604.950 363.600 607.050 364.050 ;
        RECT 623.400 363.600 624.600 365.400 ;
        RECT 604.950 362.400 624.600 363.600 ;
        RECT 647.400 363.600 648.600 365.400 ;
        RECT 673.950 366.450 676.050 366.900 ;
        RECT 679.950 366.450 682.050 367.050 ;
        RECT 685.950 366.450 688.050 366.900 ;
        RECT 673.950 365.250 688.050 366.450 ;
        RECT 689.400 366.600 690.600 368.400 ;
        RECT 737.400 366.900 738.600 370.950 ;
        RECT 691.950 366.600 694.050 366.900 ;
        RECT 709.950 366.600 712.050 366.900 ;
        RECT 689.400 365.400 712.050 366.600 ;
        RECT 673.950 364.800 676.050 365.250 ;
        RECT 679.950 364.950 682.050 365.250 ;
        RECT 685.950 364.800 688.050 365.250 ;
        RECT 691.950 364.800 694.050 365.400 ;
        RECT 709.950 364.800 712.050 365.400 ;
        RECT 736.950 364.800 739.050 366.900 ;
        RECT 749.400 364.050 750.600 371.100 ;
        RECT 778.950 370.950 781.050 373.050 ;
        RECT 787.950 372.600 790.050 373.200 ;
        RECT 785.400 371.400 790.050 372.600 ;
        RECT 775.950 366.600 778.050 366.900 ;
        RECT 779.400 366.600 780.600 370.950 ;
        RECT 785.400 367.050 786.600 371.400 ;
        RECT 787.950 371.100 790.050 371.400 ;
        RECT 805.950 369.600 808.050 373.050 ;
        RECT 817.950 370.950 820.050 373.050 ;
        RECT 835.950 372.600 838.050 373.200 ;
        RECT 833.400 371.400 838.050 372.600 ;
        RECT 803.400 369.000 808.050 369.600 ;
        RECT 803.400 368.400 807.600 369.000 ;
        RECT 775.950 365.400 780.600 366.600 ;
        RECT 775.950 364.800 778.050 365.400 ;
        RECT 784.950 364.950 787.050 367.050 ;
        RECT 670.950 363.600 673.050 364.050 ;
        RECT 647.400 362.400 673.050 363.600 ;
        RECT 604.950 361.950 607.050 362.400 ;
        RECT 670.950 361.950 673.050 362.400 ;
        RECT 700.950 363.600 703.050 364.050 ;
        RECT 721.950 363.600 724.050 364.050 ;
        RECT 700.950 362.400 724.050 363.600 ;
        RECT 700.950 361.950 703.050 362.400 ;
        RECT 721.950 361.950 724.050 362.400 ;
        RECT 748.950 361.950 751.050 364.050 ;
        RECT 760.950 363.600 763.050 364.050 ;
        RECT 772.950 363.600 775.050 364.050 ;
        RECT 760.950 362.400 775.050 363.600 ;
        RECT 760.950 361.950 763.050 362.400 ;
        RECT 772.950 361.950 775.050 362.400 ;
        RECT 790.950 363.600 793.050 364.050 ;
        RECT 803.400 363.600 804.600 368.400 ;
        RECT 818.400 367.050 819.600 370.950 ;
        RECT 814.950 366.600 817.050 366.900 ;
        RECT 806.400 366.000 817.050 366.600 ;
        RECT 790.950 362.400 804.600 363.600 ;
        RECT 805.950 365.400 817.050 366.000 ;
        RECT 818.400 365.400 823.050 367.050 ;
        RECT 790.950 361.950 793.050 362.400 ;
        RECT 805.950 361.950 808.050 365.400 ;
        RECT 814.950 364.800 817.050 365.400 ;
        RECT 819.000 364.950 823.050 365.400 ;
        RECT 833.400 364.050 834.600 371.400 ;
        RECT 835.950 371.100 838.050 371.400 ;
        RECT 839.400 366.900 840.600 373.950 ;
        RECT 847.950 372.600 850.050 376.050 ;
        RECT 862.950 375.600 865.050 376.050 ;
        RECT 871.950 375.600 874.050 376.050 ;
        RECT 862.950 374.400 874.050 375.600 ;
        RECT 862.950 373.950 865.050 374.400 ;
        RECT 871.950 373.950 874.050 374.400 ;
        RECT 889.950 375.600 892.050 376.050 ;
        RECT 895.950 375.600 898.050 376.050 ;
        RECT 889.950 374.400 898.050 375.600 ;
        RECT 889.950 373.950 892.050 374.400 ;
        RECT 895.950 373.950 898.050 374.400 ;
        RECT 845.400 372.000 850.050 372.600 ;
        RECT 853.950 372.600 858.000 373.050 ;
        RECT 883.950 372.600 886.050 373.200 ;
        RECT 904.950 372.600 907.050 373.200 ;
        RECT 845.400 371.400 849.600 372.000 ;
        RECT 845.400 367.050 846.600 371.400 ;
        RECT 853.950 370.950 858.600 372.600 ;
        RECT 883.950 371.400 907.050 372.600 ;
        RECT 883.950 371.100 886.050 371.400 ;
        RECT 904.950 371.100 907.050 371.400 ;
        RECT 838.950 364.800 841.050 366.900 ;
        RECT 844.950 364.950 847.050 367.050 ;
        RECT 857.400 366.900 858.600 370.950 ;
        RECT 856.950 364.800 859.050 366.900 ;
        RECT 862.950 366.600 865.050 366.900 ;
        RECT 895.950 366.600 898.050 367.050 ;
        RECT 862.950 365.400 898.050 366.600 ;
        RECT 862.950 364.800 865.050 365.400 ;
        RECT 895.950 364.950 898.050 365.400 ;
        RECT 833.400 362.400 838.050 364.050 ;
        RECT 834.000 361.950 838.050 362.400 ;
        RECT 874.950 363.600 877.050 364.050 ;
        RECT 883.950 363.600 886.050 364.050 ;
        RECT 874.950 362.400 886.050 363.600 ;
        RECT 874.950 361.950 877.050 362.400 ;
        RECT 883.950 361.950 886.050 362.400 ;
        RECT 595.950 361.800 598.050 361.950 ;
        RECT 223.950 360.600 226.050 361.050 ;
        RECT 286.800 360.600 288.900 361.050 ;
        RECT 223.950 359.400 288.900 360.600 ;
        RECT 223.950 358.950 226.050 359.400 ;
        RECT 286.800 358.950 288.900 359.400 ;
        RECT 289.950 360.600 292.050 361.050 ;
        RECT 310.950 360.600 313.050 361.050 ;
        RECT 289.950 359.400 313.050 360.600 ;
        RECT 289.950 358.950 292.050 359.400 ;
        RECT 310.950 358.950 313.050 359.400 ;
        RECT 316.950 360.600 319.050 361.050 ;
        RECT 349.950 360.600 352.050 361.050 ;
        RECT 385.950 360.600 388.050 361.050 ;
        RECT 316.950 359.400 388.050 360.600 ;
        RECT 316.950 358.950 319.050 359.400 ;
        RECT 349.950 358.950 352.050 359.400 ;
        RECT 385.950 358.950 388.050 359.400 ;
        RECT 391.950 360.600 394.050 361.050 ;
        RECT 406.950 360.600 409.050 361.050 ;
        RECT 391.950 359.400 409.050 360.600 ;
        RECT 391.950 358.950 394.050 359.400 ;
        RECT 406.950 358.950 409.050 359.400 ;
        RECT 514.950 360.600 517.050 361.050 ;
        RECT 547.950 360.600 550.050 361.050 ;
        RECT 703.950 360.600 706.050 361.050 ;
        RECT 901.950 360.600 904.050 361.050 ;
        RECT 514.950 359.400 550.050 360.600 ;
        RECT 514.950 358.950 517.050 359.400 ;
        RECT 547.950 358.950 550.050 359.400 ;
        RECT 578.400 359.400 706.050 360.600 ;
        RECT 130.950 357.600 133.050 358.050 ;
        RECT 205.950 357.600 208.050 358.050 ;
        RECT 130.950 356.400 208.050 357.600 ;
        RECT 130.950 355.950 133.050 356.400 ;
        RECT 205.950 355.950 208.050 356.400 ;
        RECT 211.950 357.600 214.050 358.050 ;
        RECT 298.950 357.600 301.050 358.050 ;
        RECT 211.950 356.400 301.050 357.600 ;
        RECT 211.950 355.950 214.050 356.400 ;
        RECT 298.950 355.950 301.050 356.400 ;
        RECT 373.950 357.600 376.050 358.050 ;
        RECT 415.950 357.600 418.050 358.050 ;
        RECT 373.950 356.400 418.050 357.600 ;
        RECT 373.950 355.950 376.050 356.400 ;
        RECT 415.950 355.950 418.050 356.400 ;
        RECT 463.950 357.600 466.050 358.050 ;
        RECT 550.950 357.600 553.050 358.050 ;
        RECT 463.950 356.400 553.050 357.600 ;
        RECT 463.950 355.950 466.050 356.400 ;
        RECT 550.950 355.950 553.050 356.400 ;
        RECT 571.950 357.600 574.050 358.050 ;
        RECT 578.400 357.600 579.600 359.400 ;
        RECT 703.950 358.950 706.050 359.400 ;
        RECT 764.400 359.400 771.600 360.600 ;
        RECT 571.950 356.400 579.600 357.600 ;
        RECT 589.950 357.600 592.050 358.050 ;
        RECT 604.950 357.600 607.050 358.050 ;
        RECT 589.950 356.400 607.050 357.600 ;
        RECT 571.950 355.950 574.050 356.400 ;
        RECT 589.950 355.950 592.050 356.400 ;
        RECT 604.950 355.950 607.050 356.400 ;
        RECT 748.950 357.600 751.050 358.050 ;
        RECT 764.400 357.600 765.600 359.400 ;
        RECT 748.950 356.400 765.600 357.600 ;
        RECT 770.400 357.600 771.600 359.400 ;
        RECT 901.950 359.400 918.600 360.600 ;
        RECT 901.950 358.950 904.050 359.400 ;
        RECT 787.950 357.600 790.050 358.050 ;
        RECT 770.400 356.400 790.050 357.600 ;
        RECT 748.950 355.950 751.050 356.400 ;
        RECT 787.950 355.950 790.050 356.400 ;
        RECT 838.950 357.600 841.050 358.050 ;
        RECT 871.950 357.600 874.050 358.050 ;
        RECT 838.950 356.400 874.050 357.600 ;
        RECT 917.400 357.600 918.600 359.400 ;
        RECT 925.950 357.600 928.050 358.050 ;
        RECT 917.400 356.400 928.050 357.600 ;
        RECT 838.950 355.950 841.050 356.400 ;
        RECT 871.950 355.950 874.050 356.400 ;
        RECT 925.950 355.950 928.050 356.400 ;
        RECT 28.950 354.600 31.050 355.050 ;
        RECT 112.950 354.600 115.050 355.050 ;
        RECT 28.950 353.400 115.050 354.600 ;
        RECT 28.950 352.950 31.050 353.400 ;
        RECT 112.950 352.950 115.050 353.400 ;
        RECT 166.950 354.600 169.050 355.050 ;
        RECT 187.950 354.600 190.050 355.050 ;
        RECT 166.950 353.400 190.050 354.600 ;
        RECT 166.950 352.950 169.050 353.400 ;
        RECT 187.950 352.950 190.050 353.400 ;
        RECT 253.950 354.600 256.050 355.050 ;
        RECT 259.950 354.600 262.050 355.050 ;
        RECT 277.950 354.600 280.050 355.050 ;
        RECT 253.950 353.400 280.050 354.600 ;
        RECT 253.950 352.950 256.050 353.400 ;
        RECT 259.950 352.950 262.050 353.400 ;
        RECT 277.950 352.950 280.050 353.400 ;
        RECT 325.950 354.600 328.050 355.050 ;
        RECT 340.950 354.600 343.050 355.050 ;
        RECT 374.400 354.600 375.600 355.950 ;
        RECT 325.950 353.400 375.600 354.600 ;
        RECT 532.950 354.600 535.050 355.050 ;
        RECT 541.950 354.600 544.050 355.050 ;
        RECT 532.950 353.400 544.050 354.600 ;
        RECT 325.950 352.950 328.050 353.400 ;
        RECT 340.950 352.950 343.050 353.400 ;
        RECT 532.950 352.950 535.050 353.400 ;
        RECT 541.950 352.950 544.050 353.400 ;
        RECT 556.950 354.600 559.050 355.050 ;
        RECT 562.950 354.600 565.050 355.050 ;
        RECT 556.950 353.400 565.050 354.600 ;
        RECT 556.950 352.950 559.050 353.400 ;
        RECT 562.950 352.950 565.050 353.400 ;
        RECT 607.950 354.600 610.050 355.050 ;
        RECT 613.950 354.600 616.050 355.050 ;
        RECT 607.950 353.400 616.050 354.600 ;
        RECT 607.950 352.950 610.050 353.400 ;
        RECT 613.950 352.950 616.050 353.400 ;
        RECT 622.950 354.600 625.050 355.050 ;
        RECT 640.950 354.600 643.050 355.050 ;
        RECT 649.950 354.600 652.050 355.050 ;
        RECT 622.950 353.400 652.050 354.600 ;
        RECT 622.950 352.950 625.050 353.400 ;
        RECT 640.950 352.950 643.050 353.400 ;
        RECT 649.950 352.950 652.050 353.400 ;
        RECT 664.950 354.600 667.050 355.050 ;
        RECT 700.950 354.600 703.050 355.050 ;
        RECT 718.800 354.600 720.900 355.050 ;
        RECT 664.950 353.400 720.900 354.600 ;
        RECT 664.950 352.950 667.050 353.400 ;
        RECT 700.950 352.950 703.050 353.400 ;
        RECT 718.800 352.950 720.900 353.400 ;
        RECT 721.950 354.600 724.050 355.050 ;
        RECT 766.950 354.600 769.050 355.050 ;
        RECT 796.950 354.600 799.050 355.050 ;
        RECT 808.950 354.600 811.050 355.050 ;
        RECT 721.950 353.400 811.050 354.600 ;
        RECT 721.950 352.950 724.050 353.400 ;
        RECT 766.950 352.950 769.050 353.400 ;
        RECT 796.950 352.950 799.050 353.400 ;
        RECT 808.950 352.950 811.050 353.400 ;
        RECT 814.950 354.600 817.050 355.050 ;
        RECT 853.950 354.600 856.050 355.050 ;
        RECT 814.950 353.400 856.050 354.600 ;
        RECT 814.950 352.950 817.050 353.400 ;
        RECT 853.950 352.950 856.050 353.400 ;
        RECT 865.950 354.600 868.050 355.050 ;
        RECT 886.950 354.600 889.050 355.050 ;
        RECT 907.950 354.600 910.050 355.050 ;
        RECT 865.950 353.400 910.050 354.600 ;
        RECT 865.950 352.950 868.050 353.400 ;
        RECT 886.950 352.950 889.050 353.400 ;
        RECT 907.950 352.950 910.050 353.400 ;
        RECT 208.950 351.600 211.050 352.050 ;
        RECT 229.950 351.600 232.050 352.050 ;
        RECT 208.950 350.400 232.050 351.600 ;
        RECT 208.950 349.950 211.050 350.400 ;
        RECT 229.950 349.950 232.050 350.400 ;
        RECT 268.950 351.600 271.050 352.050 ;
        RECT 292.950 351.600 295.050 352.050 ;
        RECT 268.950 350.400 295.050 351.600 ;
        RECT 268.950 349.950 271.050 350.400 ;
        RECT 292.950 349.950 295.050 350.400 ;
        RECT 334.950 351.600 337.050 352.050 ;
        RECT 352.950 351.600 355.050 352.050 ;
        RECT 334.950 350.400 355.050 351.600 ;
        RECT 334.950 349.950 337.050 350.400 ;
        RECT 352.950 349.950 355.050 350.400 ;
        RECT 523.950 351.600 526.050 352.050 ;
        RECT 544.950 351.600 547.050 352.050 ;
        RECT 523.950 350.400 547.050 351.600 ;
        RECT 523.950 349.950 526.050 350.400 ;
        RECT 544.950 349.950 547.050 350.400 ;
        RECT 610.950 351.600 613.050 352.050 ;
        RECT 718.950 351.600 721.050 351.900 ;
        RECT 751.950 351.600 754.050 352.050 ;
        RECT 769.950 351.600 772.050 352.050 ;
        RECT 784.950 351.600 787.050 352.050 ;
        RECT 610.950 350.400 787.050 351.600 ;
        RECT 610.950 349.950 613.050 350.400 ;
        RECT 718.950 349.800 721.050 350.400 ;
        RECT 751.950 349.950 754.050 350.400 ;
        RECT 769.950 349.950 772.050 350.400 ;
        RECT 784.950 349.950 787.050 350.400 ;
        RECT 847.950 351.600 850.050 352.050 ;
        RECT 862.950 351.600 865.050 352.050 ;
        RECT 847.950 350.400 865.050 351.600 ;
        RECT 847.950 349.950 850.050 350.400 ;
        RECT 862.950 349.950 865.050 350.400 ;
        RECT 868.950 351.600 871.050 352.050 ;
        RECT 874.950 351.600 877.050 352.050 ;
        RECT 880.950 351.600 883.050 352.050 ;
        RECT 868.950 350.400 883.050 351.600 ;
        RECT 868.950 349.950 871.050 350.400 ;
        RECT 874.950 349.950 877.050 350.400 ;
        RECT 880.950 349.950 883.050 350.400 ;
        RECT 913.950 351.600 916.050 352.050 ;
        RECT 931.950 351.600 934.050 352.050 ;
        RECT 913.950 350.400 934.050 351.600 ;
        RECT 913.950 349.950 916.050 350.400 ;
        RECT 931.950 349.950 934.050 350.400 ;
        RECT 61.950 348.600 64.050 349.050 ;
        RECT 127.950 348.600 130.050 349.050 ;
        RECT 61.950 347.400 130.050 348.600 ;
        RECT 61.950 346.950 64.050 347.400 ;
        RECT 127.950 346.950 130.050 347.400 ;
        RECT 145.950 348.600 148.050 349.050 ;
        RECT 151.950 348.600 154.050 349.050 ;
        RECT 166.950 348.600 169.050 349.050 ;
        RECT 145.950 347.400 169.050 348.600 ;
        RECT 145.950 346.950 148.050 347.400 ;
        RECT 151.950 346.950 154.050 347.400 ;
        RECT 166.950 346.950 169.050 347.400 ;
        RECT 199.950 348.600 202.050 349.050 ;
        RECT 226.950 348.600 229.050 349.050 ;
        RECT 199.950 347.400 229.050 348.600 ;
        RECT 199.950 346.950 202.050 347.400 ;
        RECT 226.950 346.950 229.050 347.400 ;
        RECT 232.950 348.600 235.050 349.050 ;
        RECT 280.950 348.600 283.050 349.050 ;
        RECT 232.950 347.400 283.050 348.600 ;
        RECT 232.950 346.950 235.050 347.400 ;
        RECT 280.950 346.950 283.050 347.400 ;
        RECT 427.950 348.600 430.050 349.050 ;
        RECT 451.950 348.600 454.050 349.050 ;
        RECT 427.950 347.400 454.050 348.600 ;
        RECT 427.950 346.950 430.050 347.400 ;
        RECT 451.950 346.950 454.050 347.400 ;
        RECT 547.950 348.600 550.050 349.050 ;
        RECT 553.950 348.600 556.050 349.050 ;
        RECT 562.950 348.600 565.050 349.050 ;
        RECT 547.950 347.400 565.050 348.600 ;
        RECT 547.950 346.950 550.050 347.400 ;
        RECT 553.950 346.950 556.050 347.400 ;
        RECT 562.950 346.950 565.050 347.400 ;
        RECT 646.950 348.600 649.050 349.050 ;
        RECT 658.950 348.600 661.050 349.050 ;
        RECT 646.950 347.400 661.050 348.600 ;
        RECT 646.950 346.950 649.050 347.400 ;
        RECT 658.950 346.950 661.050 347.400 ;
        RECT 673.950 348.600 676.050 349.050 ;
        RECT 712.950 348.600 715.050 349.050 ;
        RECT 727.950 348.600 730.050 349.050 ;
        RECT 673.950 347.400 715.050 348.600 ;
        RECT 673.950 346.950 676.050 347.400 ;
        RECT 712.950 346.950 715.050 347.400 ;
        RECT 722.400 347.400 730.050 348.600 ;
        RECT 67.950 345.600 70.050 346.050 ;
        RECT 76.950 345.600 79.050 346.050 ;
        RECT 67.950 344.400 79.050 345.600 ;
        RECT 67.950 343.950 70.050 344.400 ;
        RECT 76.950 343.950 79.050 344.400 ;
        RECT 151.950 345.600 154.050 345.900 ;
        RECT 160.950 345.600 163.050 346.050 ;
        RECT 151.950 344.400 163.050 345.600 ;
        RECT 151.950 343.800 154.050 344.400 ;
        RECT 160.950 343.950 163.050 344.400 ;
        RECT 190.950 345.600 193.050 346.050 ;
        RECT 217.950 345.600 220.050 346.050 ;
        RECT 190.950 344.400 220.050 345.600 ;
        RECT 190.950 343.950 193.050 344.400 ;
        RECT 217.950 343.950 220.050 344.400 ;
        RECT 274.950 345.600 277.050 346.050 ;
        RECT 301.950 345.600 304.050 346.050 ;
        RECT 274.950 344.400 304.050 345.600 ;
        RECT 274.950 343.950 277.050 344.400 ;
        RECT 301.950 343.950 304.050 344.400 ;
        RECT 397.950 345.600 400.050 346.050 ;
        RECT 424.950 345.600 427.050 346.050 ;
        RECT 397.950 344.400 427.050 345.600 ;
        RECT 397.950 343.950 400.050 344.400 ;
        RECT 424.950 343.950 427.050 344.400 ;
        RECT 454.950 345.600 457.050 346.050 ;
        RECT 472.950 345.600 475.050 346.050 ;
        RECT 454.950 344.400 475.050 345.600 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 472.950 343.950 475.050 344.400 ;
        RECT 487.950 345.600 490.050 346.050 ;
        RECT 496.800 345.600 498.900 346.050 ;
        RECT 487.950 344.400 498.900 345.600 ;
        RECT 487.950 343.950 490.050 344.400 ;
        RECT 496.800 343.950 498.900 344.400 ;
        RECT 499.950 345.600 502.050 346.050 ;
        RECT 517.950 345.600 520.050 346.050 ;
        RECT 499.950 344.400 520.050 345.600 ;
        RECT 499.950 343.950 502.050 344.400 ;
        RECT 517.950 343.950 520.050 344.400 ;
        RECT 526.950 345.600 529.050 346.050 ;
        RECT 538.950 345.600 541.050 346.050 ;
        RECT 526.950 344.400 541.050 345.600 ;
        RECT 526.950 343.950 529.050 344.400 ;
        RECT 538.950 343.950 541.050 344.400 ;
        RECT 574.950 345.600 577.050 346.050 ;
        RECT 589.950 345.600 592.050 346.050 ;
        RECT 574.950 344.400 592.050 345.600 ;
        RECT 574.950 343.950 577.050 344.400 ;
        RECT 589.950 343.950 592.050 344.400 ;
        RECT 598.950 345.600 601.050 346.050 ;
        RECT 616.800 345.600 618.900 346.050 ;
        RECT 598.950 344.400 618.900 345.600 ;
        RECT 598.950 343.950 601.050 344.400 ;
        RECT 616.800 343.950 618.900 344.400 ;
        RECT 619.950 345.600 622.050 346.050 ;
        RECT 634.950 345.600 637.050 346.050 ;
        RECT 619.950 344.400 637.050 345.600 ;
        RECT 619.950 343.950 622.050 344.400 ;
        RECT 634.950 343.950 637.050 344.400 ;
        RECT 646.950 345.600 649.050 345.900 ;
        RECT 655.950 345.600 658.050 346.050 ;
        RECT 722.400 345.600 723.600 347.400 ;
        RECT 727.950 346.950 730.050 347.400 ;
        RECT 787.950 348.600 790.050 349.050 ;
        RECT 820.950 348.600 823.050 349.050 ;
        RECT 787.950 347.400 823.050 348.600 ;
        RECT 787.950 346.950 790.050 347.400 ;
        RECT 820.950 346.950 823.050 347.400 ;
        RECT 841.950 348.600 844.050 349.050 ;
        RECT 847.950 348.600 850.050 348.900 ;
        RECT 910.950 348.600 913.050 349.050 ;
        RECT 841.950 347.400 913.050 348.600 ;
        RECT 841.950 346.950 844.050 347.400 ;
        RECT 847.950 346.800 850.050 347.400 ;
        RECT 646.950 344.400 658.050 345.600 ;
        RECT 646.950 343.800 649.050 344.400 ;
        RECT 655.950 343.950 658.050 344.400 ;
        RECT 716.400 344.400 723.600 345.600 ;
        RECT 850.950 345.600 853.050 346.050 ;
        RECT 859.950 345.600 862.050 346.050 ;
        RECT 850.950 344.400 862.050 345.600 ;
        RECT 112.950 342.600 115.050 343.050 ;
        RECT 175.950 342.600 178.050 343.050 ;
        RECT 250.950 342.600 253.050 343.050 ;
        RECT 112.950 341.400 156.600 342.600 ;
        RECT 112.950 340.950 115.050 341.400 ;
        RECT 37.950 339.600 40.050 340.050 ;
        RECT 70.950 339.600 73.050 340.050 ;
        RECT 37.950 338.400 73.050 339.600 ;
        RECT 37.950 337.950 40.050 338.400 ;
        RECT 70.950 337.950 73.050 338.400 ;
        RECT 121.950 339.600 124.050 340.050 ;
        RECT 127.950 339.600 130.050 340.050 ;
        RECT 150.000 339.600 154.050 340.050 ;
        RECT 121.950 338.400 130.050 339.600 ;
        RECT 121.950 337.950 124.050 338.400 ;
        RECT 127.950 337.950 130.050 338.400 ;
        RECT 149.400 337.950 154.050 339.600 ;
        RECT 155.400 339.600 156.600 341.400 ;
        RECT 175.950 341.400 253.050 342.600 ;
        RECT 175.950 340.950 178.050 341.400 ;
        RECT 250.950 340.950 253.050 341.400 ;
        RECT 433.950 342.600 436.050 343.050 ;
        RECT 442.950 342.600 445.050 343.050 ;
        RECT 433.950 341.400 445.050 342.600 ;
        RECT 433.950 340.950 436.050 341.400 ;
        RECT 442.950 340.950 445.050 341.400 ;
        RECT 448.950 342.600 451.050 343.050 ;
        RECT 526.950 342.600 529.050 342.900 ;
        RECT 448.950 341.400 529.050 342.600 ;
        RECT 448.950 340.950 451.050 341.400 ;
        RECT 526.950 340.800 529.050 341.400 ;
        RECT 535.950 340.950 538.050 343.050 ;
        RECT 541.950 342.600 544.050 343.050 ;
        RECT 556.950 342.600 559.050 343.050 ;
        RECT 583.950 342.600 586.050 343.050 ;
        RECT 541.950 341.400 586.050 342.600 ;
        RECT 541.950 340.950 544.050 341.400 ;
        RECT 556.950 340.950 559.050 341.400 ;
        RECT 583.950 340.950 586.050 341.400 ;
        RECT 595.950 342.600 598.050 343.050 ;
        RECT 640.950 342.600 643.050 343.050 ;
        RECT 595.950 341.400 643.050 342.600 ;
        RECT 595.950 340.950 598.050 341.400 ;
        RECT 640.950 340.950 643.050 341.400 ;
        RECT 649.950 342.600 652.050 343.050 ;
        RECT 706.950 342.600 709.050 343.050 ;
        RECT 716.400 342.600 717.600 344.400 ;
        RECT 850.950 343.950 853.050 344.400 ;
        RECT 859.950 343.950 862.050 344.400 ;
        RECT 883.950 343.800 886.050 347.400 ;
        RECT 910.950 346.950 913.050 347.400 ;
        RECT 898.950 345.600 901.050 346.050 ;
        RECT 907.950 345.600 910.050 346.050 ;
        RECT 898.950 344.400 910.050 345.600 ;
        RECT 898.950 343.950 901.050 344.400 ;
        RECT 907.950 343.950 910.050 344.400 ;
        RECT 919.950 345.600 922.050 346.050 ;
        RECT 931.950 345.600 934.050 346.050 ;
        RECT 919.950 344.400 934.050 345.600 ;
        RECT 919.950 343.950 922.050 344.400 ;
        RECT 931.950 343.950 934.050 344.400 ;
        RECT 649.950 341.400 709.050 342.600 ;
        RECT 649.950 340.950 652.050 341.400 ;
        RECT 706.950 340.950 709.050 341.400 ;
        RECT 713.400 341.400 717.600 342.600 ;
        RECT 724.950 342.600 727.050 343.050 ;
        RECT 736.950 342.600 739.050 343.050 ;
        RECT 724.950 341.400 739.050 342.600 ;
        RECT 160.950 339.600 163.050 340.200 ;
        RECT 155.400 338.400 163.050 339.600 ;
        RECT 160.950 338.100 163.050 338.400 ;
        RECT 166.950 339.750 169.050 340.200 ;
        RECT 178.950 339.750 181.050 340.200 ;
        RECT 166.950 338.550 181.050 339.750 ;
        RECT 166.950 338.100 169.050 338.550 ;
        RECT 178.950 338.100 181.050 338.550 ;
        RECT 184.950 339.600 187.050 340.200 ;
        RECT 196.950 339.600 199.050 340.050 ;
        RECT 184.950 338.400 199.050 339.600 ;
        RECT 184.950 338.100 187.050 338.400 ;
        RECT 196.950 337.950 199.050 338.400 ;
        RECT 202.950 339.600 205.050 340.050 ;
        RECT 217.950 339.600 220.050 340.050 ;
        RECT 202.950 338.400 220.050 339.600 ;
        RECT 202.950 337.950 205.050 338.400 ;
        RECT 217.950 337.950 220.050 338.400 ;
        RECT 235.950 339.600 238.050 340.050 ;
        RECT 241.950 339.600 244.050 340.200 ;
        RECT 235.950 338.400 244.050 339.600 ;
        RECT 235.950 337.950 238.050 338.400 ;
        RECT 241.950 338.100 244.050 338.400 ;
        RECT 298.950 339.600 301.050 340.200 ;
        RECT 307.950 339.600 310.050 340.050 ;
        RECT 319.950 339.600 322.050 340.200 ;
        RECT 324.000 339.600 328.050 340.050 ;
        RECT 298.950 338.400 310.050 339.600 ;
        RECT 298.950 338.100 301.050 338.400 ;
        RECT 307.950 337.950 310.050 338.400 ;
        RECT 314.400 338.400 322.050 339.600 ;
        RECT 61.950 336.600 64.050 337.200 ;
        RECT 67.950 336.600 70.050 337.050 ;
        RECT 61.950 335.400 70.050 336.600 ;
        RECT 61.950 335.100 64.050 335.400 ;
        RECT 67.950 334.950 70.050 335.400 ;
        RECT 76.950 336.450 79.050 336.900 ;
        RECT 97.950 336.450 100.050 336.900 ;
        RECT 76.950 335.250 100.050 336.450 ;
        RECT 76.950 334.800 79.050 335.250 ;
        RECT 97.950 334.800 100.050 335.250 ;
        RECT 124.950 336.600 127.050 337.050 ;
        RECT 124.950 335.400 141.600 336.600 ;
        RECT 124.950 334.950 127.050 335.400 ;
        RECT 46.950 333.600 49.050 334.050 ;
        RECT 52.950 333.600 55.050 333.900 ;
        RECT 46.950 332.400 55.050 333.600 ;
        RECT 140.400 333.600 141.600 335.400 ;
        RECT 149.400 333.900 150.600 337.950 ;
        RECT 314.400 334.050 315.600 338.400 ;
        RECT 319.950 338.100 322.050 338.400 ;
        RECT 323.400 337.950 328.050 339.600 ;
        RECT 331.950 339.600 334.050 340.050 ;
        RECT 346.950 339.600 349.050 340.200 ;
        RECT 367.950 339.600 370.050 340.200 ;
        RECT 331.950 338.400 370.050 339.600 ;
        RECT 331.950 337.950 334.050 338.400 ;
        RECT 346.950 338.100 349.050 338.400 ;
        RECT 367.950 338.100 370.050 338.400 ;
        RECT 388.950 338.100 391.050 340.200 ;
        RECT 406.950 339.600 409.050 340.200 ;
        RECT 412.950 339.600 415.050 340.200 ;
        RECT 418.950 339.600 421.050 340.050 ;
        RECT 406.950 338.400 411.600 339.600 ;
        RECT 406.950 338.100 409.050 338.400 ;
        RECT 142.950 333.600 145.050 333.900 ;
        RECT 140.400 332.400 145.050 333.600 ;
        RECT 46.950 331.950 49.050 332.400 ;
        RECT 52.950 331.800 55.050 332.400 ;
        RECT 142.950 331.800 145.050 332.400 ;
        RECT 148.950 331.800 151.050 333.900 ;
        RECT 157.950 333.450 160.050 333.900 ;
        RECT 163.950 333.450 166.050 333.900 ;
        RECT 157.950 332.250 166.050 333.450 ;
        RECT 157.950 331.800 160.050 332.250 ;
        RECT 163.950 331.800 166.050 332.250 ;
        RECT 274.950 333.600 277.050 333.900 ;
        RECT 292.950 333.600 295.050 334.050 ;
        RECT 274.950 332.400 295.050 333.600 ;
        RECT 274.950 331.800 277.050 332.400 ;
        RECT 292.950 331.950 295.050 332.400 ;
        RECT 313.950 331.950 316.050 334.050 ;
        RECT 323.400 333.900 324.600 337.950 ;
        RECT 389.400 336.600 390.600 338.100 ;
        RECT 374.400 335.400 390.600 336.600 ;
        RECT 410.400 336.600 411.600 338.400 ;
        RECT 412.950 338.400 421.050 339.600 ;
        RECT 412.950 338.100 415.050 338.400 ;
        RECT 418.950 337.950 421.050 338.400 ;
        RECT 436.950 339.600 439.050 340.050 ;
        RECT 463.950 339.750 466.050 340.200 ;
        RECT 478.950 339.750 481.050 340.200 ;
        RECT 436.950 338.400 447.600 339.600 ;
        RECT 436.950 337.950 439.050 338.400 ;
        RECT 446.400 336.600 447.600 338.400 ;
        RECT 463.950 338.550 481.050 339.750 ;
        RECT 463.950 338.100 466.050 338.550 ;
        RECT 478.950 338.100 481.050 338.550 ;
        RECT 493.950 339.750 496.050 340.200 ;
        RECT 505.950 339.750 508.050 340.200 ;
        RECT 493.950 338.550 508.050 339.750 ;
        RECT 493.950 338.100 496.050 338.550 ;
        RECT 505.950 338.100 508.050 338.550 ;
        RECT 532.950 338.100 535.050 340.200 ;
        RECT 410.400 335.400 426.600 336.600 ;
        RECT 446.400 335.400 465.600 336.600 ;
        RECT 322.950 331.800 325.050 333.900 ;
        RECT 358.950 333.450 361.050 333.900 ;
        RECT 364.950 333.450 367.050 333.900 ;
        RECT 358.950 332.250 367.050 333.450 ;
        RECT 358.950 331.800 361.050 332.250 ;
        RECT 364.950 331.800 367.050 332.250 ;
        RECT 370.950 333.600 373.050 333.900 ;
        RECT 374.400 333.600 375.600 335.400 ;
        RECT 425.400 333.900 426.600 335.400 ;
        RECT 370.950 332.400 375.600 333.600 ;
        RECT 370.950 331.800 373.050 332.400 ;
        RECT 424.950 331.800 427.050 333.900 ;
        RECT 121.950 330.450 124.050 330.900 ;
        RECT 127.950 330.450 130.050 330.900 ;
        RECT 121.950 329.250 130.050 330.450 ;
        RECT 121.950 328.800 124.050 329.250 ;
        RECT 127.950 328.800 130.050 329.250 ;
        RECT 181.950 330.600 184.050 331.050 ;
        RECT 199.950 330.600 202.050 331.050 ;
        RECT 181.950 329.400 202.050 330.600 ;
        RECT 181.950 328.950 184.050 329.400 ;
        RECT 199.950 328.950 202.050 329.400 ;
        RECT 211.950 330.600 214.050 331.050 ;
        RECT 253.950 330.600 256.050 331.050 ;
        RECT 211.950 329.400 256.050 330.600 ;
        RECT 211.950 328.950 214.050 329.400 ;
        RECT 253.950 328.950 256.050 329.400 ;
        RECT 298.950 330.600 301.050 331.050 ;
        RECT 367.950 330.600 370.050 331.050 ;
        RECT 376.950 330.600 379.050 331.050 ;
        RECT 298.950 329.400 306.600 330.600 ;
        RECT 298.950 328.950 301.050 329.400 ;
        RECT 148.950 327.600 151.050 328.050 ;
        RECT 154.950 327.600 157.050 328.050 ;
        RECT 148.950 326.400 157.050 327.600 ;
        RECT 148.950 325.950 151.050 326.400 ;
        RECT 154.950 325.950 157.050 326.400 ;
        RECT 205.950 327.600 208.050 328.050 ;
        RECT 235.950 327.600 238.050 328.050 ;
        RECT 295.950 327.600 298.050 328.050 ;
        RECT 205.950 326.400 298.050 327.600 ;
        RECT 305.400 327.600 306.600 329.400 ;
        RECT 367.950 329.400 379.050 330.600 ;
        RECT 367.950 328.950 370.050 329.400 ;
        RECT 376.950 328.950 379.050 329.400 ;
        RECT 382.950 330.600 385.050 331.050 ;
        RECT 388.950 330.600 391.050 331.050 ;
        RECT 382.950 329.400 391.050 330.600 ;
        RECT 464.400 330.600 465.600 335.400 ;
        RECT 466.950 333.600 469.050 334.050 ;
        RECT 496.950 333.600 499.050 333.900 ;
        RECT 466.950 332.400 499.050 333.600 ;
        RECT 466.950 331.950 469.050 332.400 ;
        RECT 496.950 331.800 499.050 332.400 ;
        RECT 502.950 333.600 505.050 334.050 ;
        RECT 508.950 333.600 511.050 337.050 ;
        RECT 502.950 333.000 511.050 333.600 ;
        RECT 502.950 332.400 510.600 333.000 ;
        RECT 502.950 331.950 505.050 332.400 ;
        RECT 533.400 331.050 534.600 338.100 ;
        RECT 536.400 333.900 537.600 340.950 ;
        RECT 550.950 339.600 555.000 340.050 ;
        RECT 556.950 339.600 559.050 340.200 ;
        RECT 562.950 339.600 565.050 340.200 ;
        RECT 622.950 339.600 625.050 340.050 ;
        RECT 550.950 337.950 555.600 339.600 ;
        RECT 556.950 338.400 561.600 339.600 ;
        RECT 556.950 338.100 559.050 338.400 ;
        RECT 554.400 333.900 555.600 337.950 ;
        RECT 560.400 336.600 561.600 338.400 ;
        RECT 562.950 338.400 582.600 339.600 ;
        RECT 562.950 338.100 565.050 338.400 ;
        RECT 560.400 335.400 564.600 336.600 ;
        RECT 535.950 331.800 538.050 333.900 ;
        RECT 553.950 331.800 556.050 333.900 ;
        RECT 563.400 333.600 564.600 335.400 ;
        RECT 568.950 333.600 571.050 334.050 ;
        RECT 581.400 333.900 582.600 338.400 ;
        RECT 617.400 338.400 625.050 339.600 ;
        RECT 617.400 334.050 618.600 338.400 ;
        RECT 622.950 337.950 625.050 338.400 ;
        RECT 637.950 337.950 640.050 340.050 ;
        RECT 667.950 338.100 670.050 340.200 ;
        RECT 682.950 339.600 685.050 340.050 ;
        RECT 691.950 339.600 694.050 340.200 ;
        RECT 703.950 339.600 706.050 340.050 ;
        RECT 682.950 338.400 694.050 339.600 ;
        RECT 638.400 334.050 639.600 337.950 ;
        RECT 563.400 332.400 571.050 333.600 ;
        RECT 568.950 331.950 571.050 332.400 ;
        RECT 580.950 331.800 583.050 333.900 ;
        RECT 616.950 331.950 619.050 334.050 ;
        RECT 637.950 331.950 640.050 334.050 ;
        RECT 649.950 333.600 652.050 333.900 ;
        RECT 668.400 333.600 669.600 338.100 ;
        RECT 682.950 337.950 685.050 338.400 ;
        RECT 691.950 338.100 694.050 338.400 ;
        RECT 695.400 338.400 706.050 339.600 ;
        RECT 695.400 333.900 696.600 338.400 ;
        RECT 703.950 337.950 706.050 338.400 ;
        RECT 713.400 334.050 714.600 341.400 ;
        RECT 724.950 340.950 727.050 341.400 ;
        RECT 736.950 340.950 739.050 341.400 ;
        RECT 718.950 339.600 723.000 340.050 ;
        RECT 742.950 339.600 745.050 340.200 ;
        RECT 754.950 339.600 757.050 343.050 ;
        RECT 775.950 342.600 778.050 343.050 ;
        RECT 781.950 342.600 784.050 343.050 ;
        RECT 775.950 341.400 784.050 342.600 ;
        RECT 775.950 340.950 778.050 341.400 ;
        RECT 781.950 340.950 784.050 341.400 ;
        RECT 796.950 342.600 799.050 343.050 ;
        RECT 802.950 342.600 805.050 343.050 ;
        RECT 796.950 341.400 805.050 342.600 ;
        RECT 796.950 340.950 799.050 341.400 ;
        RECT 802.950 340.950 805.050 341.400 ;
        RECT 817.950 342.600 820.050 343.050 ;
        RECT 823.950 342.600 826.050 343.050 ;
        RECT 841.950 342.600 844.050 343.050 ;
        RECT 916.950 342.600 919.050 343.050 ;
        RECT 817.950 341.400 826.050 342.600 ;
        RECT 817.950 340.950 820.050 341.400 ;
        RECT 823.950 340.950 826.050 341.400 ;
        RECT 827.400 341.400 844.050 342.600 ;
        RECT 718.950 337.950 723.600 339.600 ;
        RECT 742.950 339.000 757.050 339.600 ;
        RECT 790.950 339.600 793.050 340.200 ;
        RECT 805.950 339.600 808.050 340.200 ;
        RECT 827.400 339.600 828.600 341.400 ;
        RECT 841.950 340.950 844.050 341.400 ;
        RECT 851.400 341.400 924.600 342.600 ;
        RECT 742.950 338.400 756.600 339.000 ;
        RECT 790.950 338.400 801.600 339.600 ;
        RECT 742.950 338.100 745.050 338.400 ;
        RECT 790.950 338.100 793.050 338.400 ;
        RECT 722.400 336.600 723.600 337.950 ;
        RECT 800.400 336.600 801.600 338.400 ;
        RECT 805.950 338.400 828.600 339.600 ;
        RECT 805.950 338.100 808.050 338.400 ;
        RECT 829.950 338.100 832.050 340.200 ;
        RECT 820.950 336.600 823.050 337.050 ;
        RECT 830.400 336.600 831.600 338.100 ;
        RECT 722.400 335.400 726.600 336.600 ;
        RECT 800.400 335.400 804.600 336.600 ;
        RECT 649.950 332.400 669.600 333.600 ;
        RECT 679.950 333.450 682.050 333.900 ;
        RECT 688.950 333.450 691.050 333.900 ;
        RECT 649.950 331.800 652.050 332.400 ;
        RECT 679.950 332.250 691.050 333.450 ;
        RECT 679.950 331.800 682.050 332.250 ;
        RECT 688.950 331.800 691.050 332.250 ;
        RECT 694.950 331.800 697.050 333.900 ;
        RECT 712.950 331.950 715.050 334.050 ;
        RECT 725.400 333.900 726.600 335.400 ;
        RECT 724.950 331.800 727.050 333.900 ;
        RECT 736.950 333.450 739.050 333.900 ;
        RECT 745.950 333.450 748.050 333.900 ;
        RECT 736.950 332.250 748.050 333.450 ;
        RECT 736.950 331.800 739.050 332.250 ;
        RECT 745.950 331.800 748.050 332.250 ;
        RECT 751.950 333.600 754.050 333.900 ;
        RECT 763.950 333.600 766.050 333.900 ;
        RECT 772.950 333.600 775.050 334.050 ;
        RECT 781.950 333.600 784.050 333.900 ;
        RECT 751.950 332.400 784.050 333.600 ;
        RECT 803.400 333.600 804.600 335.400 ;
        RECT 820.950 335.400 831.600 336.600 ;
        RECT 820.950 334.950 823.050 335.400 ;
        RECT 844.950 333.600 847.050 334.050 ;
        RECT 851.400 333.900 852.600 341.400 ;
        RECT 859.950 339.600 862.050 340.050 ;
        RECT 883.950 339.600 886.050 340.050 ;
        RECT 859.950 338.400 870.600 339.600 ;
        RECT 859.950 337.950 862.050 338.400 ;
        RECT 803.400 332.400 847.050 333.600 ;
        RECT 751.950 331.800 754.050 332.400 ;
        RECT 763.950 331.800 766.050 332.400 ;
        RECT 772.950 331.950 775.050 332.400 ;
        RECT 781.950 331.800 784.050 332.400 ;
        RECT 844.950 331.950 847.050 332.400 ;
        RECT 850.950 331.800 853.050 333.900 ;
        RECT 475.950 330.600 478.050 331.050 ;
        RECT 464.400 329.400 478.050 330.600 ;
        RECT 382.950 328.950 385.050 329.400 ;
        RECT 388.950 328.950 391.050 329.400 ;
        RECT 475.950 328.950 478.050 329.400 ;
        RECT 532.950 328.950 535.050 331.050 ;
        RECT 658.950 330.600 661.050 331.050 ;
        RECT 670.950 330.600 673.050 331.050 ;
        RECT 658.950 329.400 673.050 330.600 ;
        RECT 869.400 330.600 870.600 338.400 ;
        RECT 872.400 338.400 886.050 339.600 ;
        RECT 872.400 333.900 873.600 338.400 ;
        RECT 883.950 337.950 886.050 338.400 ;
        RECT 889.950 337.950 892.050 340.050 ;
        RECT 895.950 338.100 898.050 340.200 ;
        RECT 890.400 334.050 891.600 337.950 ;
        RECT 871.950 331.800 874.050 333.900 ;
        RECT 889.950 331.950 892.050 334.050 ;
        RECT 896.400 331.050 897.600 338.100 ;
        RECT 899.400 333.900 900.600 341.400 ;
        RECT 916.950 340.950 919.050 341.400 ;
        RECT 901.950 338.100 904.050 340.200 ;
        RECT 902.400 336.600 903.600 338.100 ;
        RECT 902.400 336.000 906.600 336.600 ;
        RECT 902.400 335.400 907.050 336.000 ;
        RECT 898.950 331.800 901.050 333.900 ;
        RECT 904.950 331.950 907.050 335.400 ;
        RECT 923.400 333.900 924.600 341.400 ;
        RECT 910.950 333.450 913.050 333.900 ;
        RECT 916.950 333.450 919.050 333.900 ;
        RECT 910.950 332.250 919.050 333.450 ;
        RECT 910.950 331.800 913.050 332.250 ;
        RECT 916.950 331.800 919.050 332.250 ;
        RECT 922.950 331.800 925.050 333.900 ;
        RECT 877.950 330.600 880.050 331.050 ;
        RECT 869.400 329.400 880.050 330.600 ;
        RECT 658.950 328.950 661.050 329.400 ;
        RECT 670.950 328.950 673.050 329.400 ;
        RECT 877.950 328.950 880.050 329.400 ;
        RECT 895.950 328.950 898.050 331.050 ;
        RECT 316.950 327.600 319.050 328.050 ;
        RECT 328.950 327.600 331.050 328.050 ;
        RECT 305.400 326.400 331.050 327.600 ;
        RECT 205.950 325.950 208.050 326.400 ;
        RECT 235.950 325.950 238.050 326.400 ;
        RECT 295.950 325.950 298.050 326.400 ;
        RECT 316.950 325.950 319.050 326.400 ;
        RECT 328.950 325.950 331.050 326.400 ;
        RECT 361.950 327.600 364.050 328.050 ;
        RECT 376.950 327.600 379.050 327.900 ;
        RECT 361.950 326.400 379.050 327.600 ;
        RECT 361.950 325.950 364.050 326.400 ;
        RECT 376.950 325.800 379.050 326.400 ;
        RECT 403.950 327.600 406.050 328.050 ;
        RECT 430.950 327.600 433.050 328.050 ;
        RECT 403.950 326.400 433.050 327.600 ;
        RECT 403.950 325.950 406.050 326.400 ;
        RECT 430.950 325.950 433.050 326.400 ;
        RECT 583.950 327.600 586.050 328.050 ;
        RECT 592.950 327.600 595.050 328.050 ;
        RECT 583.950 326.400 595.050 327.600 ;
        RECT 583.950 325.950 586.050 326.400 ;
        RECT 592.950 325.950 595.050 326.400 ;
        RECT 613.950 327.600 616.050 328.050 ;
        RECT 628.950 327.600 631.050 328.050 ;
        RECT 613.950 326.400 631.050 327.600 ;
        RECT 613.950 325.950 616.050 326.400 ;
        RECT 628.950 325.950 631.050 326.400 ;
        RECT 646.950 327.600 649.050 328.050 ;
        RECT 652.950 327.600 655.050 328.050 ;
        RECT 646.950 326.400 655.050 327.600 ;
        RECT 646.950 325.950 649.050 326.400 ;
        RECT 652.950 325.950 655.050 326.400 ;
        RECT 658.950 327.600 661.050 327.900 ;
        RECT 664.950 327.600 667.050 328.050 ;
        RECT 658.950 326.400 667.050 327.600 ;
        RECT 658.950 325.800 661.050 326.400 ;
        RECT 664.950 325.950 667.050 326.400 ;
        RECT 688.950 327.600 691.050 328.050 ;
        RECT 694.950 327.600 697.050 328.050 ;
        RECT 688.950 326.400 697.050 327.600 ;
        RECT 688.950 325.950 691.050 326.400 ;
        RECT 694.950 325.950 697.050 326.400 ;
        RECT 715.950 327.600 718.050 328.050 ;
        RECT 730.950 327.600 733.050 328.050 ;
        RECT 787.950 327.600 790.050 328.050 ;
        RECT 715.950 326.400 790.050 327.600 ;
        RECT 715.950 325.950 718.050 326.400 ;
        RECT 730.950 325.950 733.050 326.400 ;
        RECT 787.950 325.950 790.050 326.400 ;
        RECT 844.950 327.600 847.050 328.050 ;
        RECT 865.950 327.600 868.050 328.050 ;
        RECT 844.950 326.400 868.050 327.600 ;
        RECT 844.950 325.950 847.050 326.400 ;
        RECT 865.950 325.950 868.050 326.400 ;
        RECT 40.950 324.600 43.050 325.050 ;
        RECT 58.950 324.600 61.050 325.050 ;
        RECT 40.950 323.400 61.050 324.600 ;
        RECT 40.950 322.950 43.050 323.400 ;
        RECT 58.950 322.950 61.050 323.400 ;
        RECT 169.950 324.600 172.050 325.050 ;
        RECT 196.950 324.600 199.050 325.050 ;
        RECT 169.950 323.400 199.050 324.600 ;
        RECT 169.950 322.950 172.050 323.400 ;
        RECT 196.950 322.950 199.050 323.400 ;
        RECT 205.950 324.600 208.050 324.900 ;
        RECT 280.950 324.600 283.050 325.050 ;
        RECT 205.950 323.400 283.050 324.600 ;
        RECT 205.950 322.800 208.050 323.400 ;
        RECT 280.950 322.950 283.050 323.400 ;
        RECT 301.950 324.600 304.050 325.050 ;
        RECT 331.950 324.600 334.050 325.050 ;
        RECT 301.950 323.400 334.050 324.600 ;
        RECT 301.950 322.950 304.050 323.400 ;
        RECT 331.950 322.950 334.050 323.400 ;
        RECT 355.950 324.600 358.050 325.050 ;
        RECT 397.950 324.600 400.050 325.050 ;
        RECT 355.950 323.400 400.050 324.600 ;
        RECT 355.950 322.950 358.050 323.400 ;
        RECT 397.950 322.950 400.050 323.400 ;
        RECT 415.950 324.600 418.050 325.050 ;
        RECT 535.950 324.600 538.050 325.050 ;
        RECT 415.950 323.400 538.050 324.600 ;
        RECT 415.950 322.950 418.050 323.400 ;
        RECT 535.950 322.950 538.050 323.400 ;
        RECT 550.950 324.600 553.050 325.050 ;
        RECT 559.800 324.600 561.900 325.050 ;
        RECT 550.950 323.400 561.900 324.600 ;
        RECT 550.950 322.950 553.050 323.400 ;
        RECT 559.800 322.950 561.900 323.400 ;
        RECT 562.950 324.600 565.050 325.050 ;
        RECT 595.950 324.600 598.050 325.050 ;
        RECT 604.950 324.600 607.050 325.050 ;
        RECT 562.950 323.400 607.050 324.600 ;
        RECT 562.950 322.950 565.050 323.400 ;
        RECT 595.950 322.950 598.050 323.400 ;
        RECT 604.950 322.950 607.050 323.400 ;
        RECT 613.950 324.600 616.050 324.900 ;
        RECT 655.950 324.600 658.050 325.050 ;
        RECT 676.950 324.600 679.050 325.050 ;
        RECT 613.950 323.400 679.050 324.600 ;
        RECT 613.950 322.800 616.050 323.400 ;
        RECT 655.950 322.950 658.050 323.400 ;
        RECT 676.950 322.950 679.050 323.400 ;
        RECT 685.950 324.600 688.050 325.050 ;
        RECT 709.950 324.600 712.050 325.050 ;
        RECT 685.950 323.400 712.050 324.600 ;
        RECT 685.950 322.950 688.050 323.400 ;
        RECT 709.950 322.950 712.050 323.400 ;
        RECT 835.950 324.600 838.050 325.050 ;
        RECT 904.950 324.600 907.050 325.050 ;
        RECT 835.950 323.400 907.050 324.600 ;
        RECT 835.950 322.950 838.050 323.400 ;
        RECT 904.950 322.950 907.050 323.400 ;
        RECT 214.950 321.600 217.050 322.050 ;
        RECT 244.950 321.600 247.050 322.050 ;
        RECT 214.950 320.400 247.050 321.600 ;
        RECT 214.950 319.950 217.050 320.400 ;
        RECT 244.950 319.950 247.050 320.400 ;
        RECT 259.950 321.600 262.050 322.050 ;
        RECT 271.950 321.600 274.050 322.050 ;
        RECT 298.950 321.600 301.050 322.050 ;
        RECT 259.950 320.400 274.050 321.600 ;
        RECT 259.950 319.950 262.050 320.400 ;
        RECT 271.950 319.950 274.050 320.400 ;
        RECT 284.400 320.400 301.050 321.600 ;
        RECT 250.950 318.600 253.050 319.050 ;
        RECT 284.400 318.600 285.600 320.400 ;
        RECT 298.950 319.950 301.050 320.400 ;
        RECT 304.950 321.600 307.050 322.050 ;
        RECT 325.950 321.600 328.050 322.050 ;
        RECT 304.950 320.400 328.050 321.600 ;
        RECT 304.950 319.950 307.050 320.400 ;
        RECT 325.950 319.950 328.050 320.400 ;
        RECT 337.950 321.600 340.050 322.050 ;
        RECT 688.800 321.600 690.900 321.900 ;
        RECT 337.950 320.400 690.900 321.600 ;
        RECT 337.950 319.950 340.050 320.400 ;
        RECT 688.800 319.800 690.900 320.400 ;
        RECT 691.950 321.600 694.050 322.050 ;
        RECT 700.950 321.600 703.050 322.050 ;
        RECT 691.950 320.400 703.050 321.600 ;
        RECT 691.950 319.950 694.050 320.400 ;
        RECT 700.950 319.950 703.050 320.400 ;
        RECT 718.950 321.600 721.050 322.050 ;
        RECT 802.950 321.600 805.050 322.050 ;
        RECT 820.950 321.600 823.050 322.050 ;
        RECT 718.950 320.400 823.050 321.600 ;
        RECT 718.950 319.950 721.050 320.400 ;
        RECT 802.950 319.950 805.050 320.400 ;
        RECT 820.950 319.950 823.050 320.400 ;
        RECT 250.950 317.400 285.600 318.600 ;
        RECT 304.950 318.600 307.050 318.900 ;
        RECT 325.950 318.600 328.050 318.900 ;
        RECT 304.950 317.400 328.050 318.600 ;
        RECT 250.950 316.950 253.050 317.400 ;
        RECT 304.950 316.800 307.050 317.400 ;
        RECT 325.950 316.800 328.050 317.400 ;
        RECT 418.950 318.600 421.050 319.050 ;
        RECT 451.950 318.600 454.050 319.050 ;
        RECT 418.950 317.400 454.050 318.600 ;
        RECT 418.950 316.950 421.050 317.400 ;
        RECT 451.950 316.950 454.050 317.400 ;
        RECT 466.950 318.600 469.050 319.050 ;
        RECT 529.950 318.600 532.050 319.050 ;
        RECT 466.950 317.400 532.050 318.600 ;
        RECT 466.950 316.950 469.050 317.400 ;
        RECT 529.950 316.950 532.050 317.400 ;
        RECT 553.950 318.600 556.050 319.050 ;
        RECT 583.950 318.600 586.050 319.050 ;
        RECT 553.950 317.400 586.050 318.600 ;
        RECT 553.950 316.950 556.050 317.400 ;
        RECT 583.950 316.950 586.050 317.400 ;
        RECT 589.950 318.600 592.050 319.050 ;
        RECT 616.800 318.600 618.900 319.050 ;
        RECT 589.950 317.400 618.900 318.600 ;
        RECT 589.950 316.950 592.050 317.400 ;
        RECT 616.800 316.950 618.900 317.400 ;
        RECT 619.950 318.600 622.050 319.050 ;
        RECT 694.950 318.600 697.050 319.050 ;
        RECT 619.950 317.400 697.050 318.600 ;
        RECT 619.950 316.950 622.050 317.400 ;
        RECT 694.950 316.950 697.050 317.400 ;
        RECT 703.950 318.600 706.050 319.050 ;
        RECT 808.950 318.600 811.050 319.050 ;
        RECT 703.950 317.400 811.050 318.600 ;
        RECT 703.950 316.950 706.050 317.400 ;
        RECT 808.950 316.950 811.050 317.400 ;
        RECT 178.950 315.600 181.050 316.050 ;
        RECT 220.950 315.600 223.050 316.050 ;
        RECT 178.950 314.400 223.050 315.600 ;
        RECT 178.950 313.950 181.050 314.400 ;
        RECT 220.950 313.950 223.050 314.400 ;
        RECT 295.950 315.600 298.050 316.050 ;
        RECT 316.950 315.600 319.050 316.050 ;
        RECT 295.950 314.400 319.050 315.600 ;
        RECT 295.950 313.950 298.050 314.400 ;
        RECT 316.950 313.950 319.050 314.400 ;
        RECT 328.950 315.600 331.050 316.050 ;
        RECT 352.950 315.600 355.050 316.050 ;
        RECT 367.950 315.600 370.050 316.050 ;
        RECT 328.950 314.400 370.050 315.600 ;
        RECT 328.950 313.950 331.050 314.400 ;
        RECT 352.950 313.950 355.050 314.400 ;
        RECT 367.950 313.950 370.050 314.400 ;
        RECT 547.950 315.600 550.050 316.050 ;
        RECT 562.950 315.600 565.050 316.050 ;
        RECT 547.950 314.400 565.050 315.600 ;
        RECT 547.950 313.950 550.050 314.400 ;
        RECT 562.950 313.950 565.050 314.400 ;
        RECT 586.950 315.600 589.050 316.050 ;
        RECT 613.950 315.600 616.050 316.050 ;
        RECT 586.950 314.400 616.050 315.600 ;
        RECT 586.950 313.950 589.050 314.400 ;
        RECT 613.950 313.950 616.050 314.400 ;
        RECT 628.950 315.600 631.050 316.050 ;
        RECT 679.950 315.600 682.050 316.050 ;
        RECT 754.950 315.600 757.050 316.050 ;
        RECT 628.950 314.400 682.050 315.600 ;
        RECT 628.950 313.950 631.050 314.400 ;
        RECT 679.950 313.950 682.050 314.400 ;
        RECT 707.400 314.400 757.050 315.600 ;
        RECT 187.950 312.600 190.050 313.050 ;
        RECT 301.950 312.600 304.050 313.050 ;
        RECT 187.950 311.400 304.050 312.600 ;
        RECT 187.950 310.950 190.050 311.400 ;
        RECT 301.950 310.950 304.050 311.400 ;
        RECT 370.950 312.600 373.050 313.050 ;
        RECT 418.950 312.600 421.050 313.050 ;
        RECT 370.950 311.400 421.050 312.600 ;
        RECT 370.950 310.950 373.050 311.400 ;
        RECT 418.950 310.950 421.050 311.400 ;
        RECT 442.950 312.600 445.050 313.050 ;
        RECT 511.950 312.600 514.050 313.050 ;
        RECT 442.950 311.400 514.050 312.600 ;
        RECT 442.950 310.950 445.050 311.400 ;
        RECT 511.950 310.950 514.050 311.400 ;
        RECT 529.950 312.600 532.050 313.050 ;
        RECT 574.950 312.600 577.050 313.050 ;
        RECT 529.950 311.400 577.050 312.600 ;
        RECT 529.950 310.950 532.050 311.400 ;
        RECT 574.950 310.950 577.050 311.400 ;
        RECT 628.950 312.600 631.050 312.900 ;
        RECT 640.950 312.600 643.050 313.050 ;
        RECT 628.950 311.400 643.050 312.600 ;
        RECT 628.950 310.800 631.050 311.400 ;
        RECT 640.950 310.950 643.050 311.400 ;
        RECT 700.950 312.600 703.050 313.050 ;
        RECT 707.400 312.600 708.600 314.400 ;
        RECT 754.950 313.950 757.050 314.400 ;
        RECT 700.950 311.400 708.600 312.600 ;
        RECT 775.950 312.600 778.050 313.050 ;
        RECT 817.950 312.600 820.050 313.050 ;
        RECT 775.950 311.400 820.050 312.600 ;
        RECT 700.950 310.950 703.050 311.400 ;
        RECT 775.950 310.950 778.050 311.400 ;
        RECT 817.950 310.950 820.050 311.400 ;
        RECT 838.950 312.600 841.050 313.050 ;
        RECT 874.950 312.600 877.050 313.050 ;
        RECT 838.950 311.400 877.050 312.600 ;
        RECT 838.950 310.950 841.050 311.400 ;
        RECT 874.950 310.950 877.050 311.400 ;
        RECT 49.950 309.600 52.050 310.050 ;
        RECT 67.950 309.600 70.050 310.050 ;
        RECT 49.950 308.400 70.050 309.600 ;
        RECT 49.950 307.950 52.050 308.400 ;
        RECT 67.950 307.950 70.050 308.400 ;
        RECT 217.950 309.600 220.050 310.050 ;
        RECT 238.950 309.600 241.050 310.050 ;
        RECT 217.950 308.400 241.050 309.600 ;
        RECT 217.950 307.950 220.050 308.400 ;
        RECT 238.950 307.950 241.050 308.400 ;
        RECT 253.950 309.600 256.050 310.050 ;
        RECT 274.950 309.600 277.050 310.050 ;
        RECT 253.950 308.400 277.050 309.600 ;
        RECT 253.950 307.950 256.050 308.400 ;
        RECT 274.950 307.950 277.050 308.400 ;
        RECT 280.950 309.600 283.050 310.050 ;
        RECT 310.950 309.600 313.050 310.050 ;
        RECT 322.800 309.600 324.900 310.050 ;
        RECT 280.950 308.400 324.900 309.600 ;
        RECT 280.950 307.950 283.050 308.400 ;
        RECT 310.950 307.950 313.050 308.400 ;
        RECT 322.800 307.950 324.900 308.400 ;
        RECT 325.950 309.600 328.050 310.050 ;
        RECT 340.950 309.600 343.050 310.050 ;
        RECT 469.950 309.600 472.050 310.050 ;
        RECT 502.950 309.600 505.050 310.050 ;
        RECT 325.950 308.400 441.600 309.600 ;
        RECT 325.950 307.950 328.050 308.400 ;
        RECT 340.950 307.950 343.050 308.400 ;
        RECT 440.400 307.050 441.600 308.400 ;
        RECT 469.950 308.400 505.050 309.600 ;
        RECT 469.950 307.950 472.050 308.400 ;
        RECT 502.950 307.950 505.050 308.400 ;
        RECT 556.950 309.600 559.050 310.050 ;
        RECT 580.950 309.600 583.050 310.050 ;
        RECT 556.950 308.400 583.050 309.600 ;
        RECT 556.950 307.950 559.050 308.400 ;
        RECT 580.950 307.950 583.050 308.400 ;
        RECT 886.950 309.600 889.050 310.050 ;
        RECT 916.950 309.600 919.050 310.050 ;
        RECT 886.950 308.400 919.050 309.600 ;
        RECT 886.950 307.950 889.050 308.400 ;
        RECT 916.950 307.950 919.050 308.400 ;
        RECT 163.950 306.600 166.050 307.050 ;
        RECT 172.950 306.600 175.050 307.050 ;
        RECT 163.950 305.400 175.050 306.600 ;
        RECT 163.950 304.950 166.050 305.400 ;
        RECT 172.950 304.950 175.050 305.400 ;
        RECT 268.950 306.600 271.050 307.050 ;
        RECT 286.950 306.600 289.050 307.050 ;
        RECT 268.950 305.400 289.050 306.600 ;
        RECT 268.950 304.950 271.050 305.400 ;
        RECT 286.950 304.950 289.050 305.400 ;
        RECT 292.950 306.600 295.050 307.050 ;
        RECT 301.950 306.600 304.050 307.050 ;
        RECT 292.950 305.400 304.050 306.600 ;
        RECT 292.950 304.950 295.050 305.400 ;
        RECT 301.950 304.950 304.050 305.400 ;
        RECT 307.950 306.600 310.050 307.050 ;
        RECT 370.950 306.600 373.050 307.050 ;
        RECT 307.950 305.400 373.050 306.600 ;
        RECT 307.950 304.950 310.050 305.400 ;
        RECT 370.950 304.950 373.050 305.400 ;
        RECT 439.950 306.600 442.050 307.050 ;
        RECT 451.950 306.600 454.050 307.050 ;
        RECT 457.950 306.600 460.050 307.050 ;
        RECT 439.950 305.400 460.050 306.600 ;
        RECT 439.950 304.950 442.050 305.400 ;
        RECT 451.950 304.950 454.050 305.400 ;
        RECT 457.950 304.950 460.050 305.400 ;
        RECT 559.950 306.600 562.050 307.050 ;
        RECT 565.950 306.600 568.050 307.050 ;
        RECT 559.950 305.400 568.050 306.600 ;
        RECT 559.950 304.950 562.050 305.400 ;
        RECT 565.950 304.950 568.050 305.400 ;
        RECT 601.950 306.600 604.050 307.050 ;
        RECT 640.950 306.600 643.050 307.050 ;
        RECT 601.950 305.400 643.050 306.600 ;
        RECT 601.950 304.950 604.050 305.400 ;
        RECT 640.950 304.950 643.050 305.400 ;
        RECT 649.950 306.600 652.050 307.050 ;
        RECT 682.950 306.600 685.050 307.050 ;
        RECT 649.950 305.400 685.050 306.600 ;
        RECT 649.950 304.950 652.050 305.400 ;
        RECT 682.950 304.950 685.050 305.400 ;
        RECT 829.950 306.600 832.050 307.050 ;
        RECT 841.950 306.600 844.050 307.050 ;
        RECT 829.950 305.400 844.050 306.600 ;
        RECT 829.950 304.950 832.050 305.400 ;
        RECT 841.950 304.950 844.050 305.400 ;
        RECT 865.950 306.600 868.050 307.050 ;
        RECT 892.950 306.600 895.050 307.050 ;
        RECT 865.950 305.400 895.050 306.600 ;
        RECT 865.950 304.950 868.050 305.400 ;
        RECT 892.950 304.950 895.050 305.400 ;
        RECT 37.950 303.600 40.050 304.050 ;
        RECT 46.950 303.600 49.050 304.050 ;
        RECT 67.950 303.600 70.050 304.050 ;
        RECT 37.950 302.400 70.050 303.600 ;
        RECT 37.950 301.950 40.050 302.400 ;
        RECT 46.950 301.950 49.050 302.400 ;
        RECT 67.950 301.950 70.050 302.400 ;
        RECT 148.950 303.600 151.050 304.050 ;
        RECT 160.950 303.600 163.050 304.050 ;
        RECT 148.950 302.400 163.050 303.600 ;
        RECT 148.950 301.950 151.050 302.400 ;
        RECT 160.950 301.950 163.050 302.400 ;
        RECT 235.950 303.600 238.050 304.050 ;
        RECT 283.950 303.600 286.050 304.050 ;
        RECT 325.800 303.600 327.900 304.050 ;
        RECT 235.950 302.400 270.600 303.600 ;
        RECT 235.950 301.950 238.050 302.400 ;
        RECT 19.950 300.600 22.050 301.050 ;
        RECT 34.950 300.600 37.050 301.050 ;
        RECT 19.950 299.400 37.050 300.600 ;
        RECT 19.950 298.950 22.050 299.400 ;
        RECT 34.950 298.950 37.050 299.400 ;
        RECT 55.950 300.600 58.050 301.050 ;
        RECT 139.950 300.600 142.050 301.050 ;
        RECT 55.950 299.400 142.050 300.600 ;
        RECT 55.950 298.950 58.050 299.400 ;
        RECT 139.950 298.950 142.050 299.400 ;
        RECT 7.950 292.950 10.050 295.050 ;
        RECT 13.950 294.600 16.050 295.200 ;
        RECT 28.950 294.600 31.050 295.200 ;
        RECT 13.950 293.400 31.050 294.600 ;
        RECT 31.950 294.600 34.050 298.050 ;
        RECT 97.950 297.600 100.050 298.050 ;
        RECT 145.950 297.600 148.050 298.050 ;
        RECT 151.950 297.600 154.050 301.050 ;
        RECT 229.950 300.600 232.050 301.050 ;
        RECT 265.950 300.600 268.050 301.050 ;
        RECT 229.950 299.400 268.050 300.600 ;
        RECT 269.400 300.600 270.600 302.400 ;
        RECT 283.950 302.400 327.900 303.600 ;
        RECT 283.950 301.950 286.050 302.400 ;
        RECT 325.800 301.950 327.900 302.400 ;
        RECT 328.950 303.600 331.050 304.050 ;
        RECT 355.950 303.600 358.050 304.050 ;
        RECT 328.950 302.400 358.050 303.600 ;
        RECT 328.950 301.950 331.050 302.400 ;
        RECT 355.950 301.950 358.050 302.400 ;
        RECT 364.950 303.600 367.050 304.050 ;
        RECT 379.950 303.600 382.050 304.050 ;
        RECT 364.950 302.400 382.050 303.600 ;
        RECT 364.950 301.950 367.050 302.400 ;
        RECT 379.950 301.950 382.050 302.400 ;
        RECT 517.950 303.600 520.050 304.050 ;
        RECT 562.950 303.600 565.050 304.050 ;
        RECT 517.950 302.400 565.050 303.600 ;
        RECT 517.950 301.950 520.050 302.400 ;
        RECT 562.950 301.950 565.050 302.400 ;
        RECT 622.950 303.600 625.050 304.050 ;
        RECT 652.950 303.600 655.050 304.050 ;
        RECT 622.950 302.400 655.050 303.600 ;
        RECT 622.950 301.950 625.050 302.400 ;
        RECT 652.950 301.950 655.050 302.400 ;
        RECT 703.950 303.600 706.050 304.050 ;
        RECT 727.950 303.600 730.050 304.050 ;
        RECT 733.950 303.600 736.050 304.050 ;
        RECT 703.950 302.400 736.050 303.600 ;
        RECT 703.950 301.950 706.050 302.400 ;
        RECT 727.950 301.950 730.050 302.400 ;
        RECT 733.950 301.950 736.050 302.400 ;
        RECT 769.950 303.600 772.050 304.050 ;
        RECT 820.950 303.600 823.050 304.050 ;
        RECT 769.950 302.400 823.050 303.600 ;
        RECT 769.950 301.950 772.050 302.400 ;
        RECT 820.950 301.950 823.050 302.400 ;
        RECT 304.950 300.600 307.050 301.050 ;
        RECT 269.400 299.400 307.050 300.600 ;
        RECT 229.950 298.950 232.050 299.400 ;
        RECT 265.950 298.950 268.050 299.400 ;
        RECT 304.950 298.950 307.050 299.400 ;
        RECT 442.950 300.600 445.050 301.050 ;
        RECT 481.950 300.600 484.050 301.050 ;
        RECT 484.950 300.600 487.050 301.050 ;
        RECT 442.950 299.400 487.050 300.600 ;
        RECT 442.950 298.950 445.050 299.400 ;
        RECT 481.950 298.950 484.050 299.400 ;
        RECT 484.950 298.950 487.050 299.400 ;
        RECT 496.950 300.600 499.050 301.050 ;
        RECT 505.950 300.600 508.050 301.050 ;
        RECT 496.950 299.400 508.050 300.600 ;
        RECT 496.950 298.950 499.050 299.400 ;
        RECT 505.950 298.950 508.050 299.400 ;
        RECT 532.950 300.600 535.050 301.050 ;
        RECT 568.950 300.600 571.050 301.050 ;
        RECT 532.950 299.400 571.050 300.600 ;
        RECT 532.950 298.950 535.050 299.400 ;
        RECT 568.950 298.950 571.050 299.400 ;
        RECT 724.950 300.600 727.050 301.050 ;
        RECT 748.950 300.600 751.050 301.050 ;
        RECT 724.950 299.400 751.050 300.600 ;
        RECT 724.950 298.950 727.050 299.400 ;
        RECT 748.950 298.950 751.050 299.400 ;
        RECT 784.950 300.600 787.050 301.050 ;
        RECT 796.950 300.600 799.050 301.050 ;
        RECT 784.950 299.400 799.050 300.600 ;
        RECT 784.950 298.950 787.050 299.400 ;
        RECT 796.950 298.950 799.050 299.400 ;
        RECT 832.950 300.600 835.050 301.050 ;
        RECT 847.950 300.600 850.050 301.050 ;
        RECT 889.950 300.600 892.050 301.050 ;
        RECT 901.950 300.600 904.050 301.050 ;
        RECT 832.950 299.400 850.050 300.600 ;
        RECT 832.950 298.950 835.050 299.400 ;
        RECT 847.950 298.950 850.050 299.400 ;
        RECT 887.400 299.400 904.050 300.600 ;
        RECT 97.950 296.400 148.050 297.600 ;
        RECT 97.950 295.950 100.050 296.400 ;
        RECT 145.950 295.950 148.050 296.400 ;
        RECT 149.400 297.000 154.050 297.600 ;
        RECT 149.400 296.400 153.600 297.000 ;
        RECT 31.950 294.000 39.600 294.600 ;
        RECT 32.400 293.400 39.600 294.000 ;
        RECT 13.950 293.100 16.050 293.400 ;
        RECT 28.950 293.100 31.050 293.400 ;
        RECT 8.400 289.050 9.600 292.950 ;
        RECT 7.950 286.950 10.050 289.050 ;
        RECT 38.400 288.900 39.600 293.400 ;
        RECT 40.950 293.100 43.050 295.200 ;
        RECT 58.950 294.600 61.050 295.050 ;
        RECT 149.400 294.600 150.600 296.400 ;
        RECT 268.950 295.950 271.050 298.050 ;
        RECT 313.950 297.600 316.050 298.050 ;
        RECT 296.400 296.400 316.050 297.600 ;
        RECT 58.950 293.400 69.600 294.600 ;
        RECT 125.400 294.000 150.600 294.600 ;
        RECT 41.400 291.600 42.600 293.100 ;
        RECT 58.950 292.950 61.050 293.400 ;
        RECT 64.950 291.600 67.050 292.050 ;
        RECT 41.400 290.400 67.050 291.600 ;
        RECT 68.400 291.600 69.600 293.400 ;
        RECT 124.950 293.400 150.600 294.000 ;
        RECT 151.950 294.750 154.050 295.200 ;
        RECT 157.950 294.750 160.050 295.200 ;
        RECT 151.950 293.550 160.050 294.750 ;
        RECT 162.000 294.600 166.050 295.050 ;
        RECT 178.950 294.600 181.050 295.050 ;
        RECT 73.950 291.600 76.050 292.050 ;
        RECT 68.400 290.400 76.050 291.600 ;
        RECT 64.950 289.950 67.050 290.400 ;
        RECT 73.950 289.950 76.050 290.400 ;
        RECT 124.950 289.950 127.050 293.400 ;
        RECT 151.950 293.100 154.050 293.550 ;
        RECT 157.950 293.100 160.050 293.550 ;
        RECT 161.400 292.950 166.050 294.600 ;
        RECT 173.400 293.400 181.050 294.600 ;
        RECT 161.400 291.600 162.600 292.950 ;
        RECT 152.400 290.400 162.600 291.600 ;
        RECT 22.950 288.450 25.050 288.900 ;
        RECT 31.950 288.450 34.050 288.900 ;
        RECT 22.950 287.250 34.050 288.450 ;
        RECT 22.950 286.800 25.050 287.250 ;
        RECT 31.950 286.800 34.050 287.250 ;
        RECT 37.950 286.800 40.050 288.900 ;
        RECT 115.950 288.600 118.050 289.050 ;
        RECT 127.950 288.600 130.050 289.050 ;
        RECT 115.950 287.400 130.050 288.600 ;
        RECT 115.950 286.950 118.050 287.400 ;
        RECT 127.950 286.950 130.050 287.400 ;
        RECT 148.950 288.600 151.050 288.900 ;
        RECT 152.400 288.600 153.600 290.400 ;
        RECT 173.400 288.900 174.600 293.400 ;
        RECT 178.950 292.950 181.050 293.400 ;
        RECT 199.950 294.600 202.050 295.050 ;
        RECT 211.950 294.600 214.050 295.200 ;
        RECT 217.950 294.600 220.050 295.050 ;
        RECT 235.950 294.600 238.050 295.050 ;
        RECT 199.950 293.400 216.600 294.600 ;
        RECT 199.950 292.950 202.050 293.400 ;
        RECT 211.950 293.100 214.050 293.400 ;
        RECT 215.400 291.600 216.600 293.400 ;
        RECT 217.950 293.400 238.050 294.600 ;
        RECT 217.950 292.950 220.050 293.400 ;
        RECT 235.950 292.950 238.050 293.400 ;
        RECT 247.950 293.100 250.050 295.200 ;
        RECT 248.400 291.600 249.600 293.100 ;
        RECT 215.400 290.400 249.600 291.600 ;
        RECT 148.950 287.400 153.600 288.600 ;
        RECT 148.950 286.800 151.050 287.400 ;
        RECT 172.950 286.800 175.050 288.900 ;
        RECT 193.950 288.450 196.050 288.900 ;
        RECT 199.950 288.450 202.050 288.900 ;
        RECT 193.950 287.250 202.050 288.450 ;
        RECT 193.950 286.800 196.050 287.250 ;
        RECT 199.950 286.800 202.050 287.250 ;
        RECT 244.950 288.450 247.050 288.900 ;
        RECT 259.950 288.450 262.050 288.900 ;
        RECT 244.950 287.250 262.050 288.450 ;
        RECT 244.950 286.800 247.050 287.250 ;
        RECT 259.950 286.800 262.050 287.250 ;
        RECT 269.400 286.050 270.600 295.950 ;
        RECT 286.950 294.600 289.050 295.050 ;
        RECT 286.950 293.400 294.600 294.600 ;
        RECT 286.950 292.950 289.050 293.400 ;
        RECT 271.950 288.450 274.050 288.900 ;
        RECT 283.950 288.450 286.050 288.900 ;
        RECT 271.950 287.250 286.050 288.450 ;
        RECT 293.400 288.600 294.600 293.400 ;
        RECT 296.400 291.600 297.600 296.400 ;
        RECT 313.950 295.950 316.050 296.400 ;
        RECT 391.950 297.600 394.050 298.050 ;
        RECT 463.950 297.600 466.050 298.050 ;
        RECT 472.950 297.600 475.050 298.050 ;
        RECT 391.950 296.400 475.050 297.600 ;
        RECT 391.950 295.950 394.050 296.400 ;
        RECT 463.950 295.950 466.050 296.400 ;
        RECT 472.950 295.950 475.050 296.400 ;
        RECT 487.950 297.600 490.050 298.050 ;
        RECT 493.950 297.600 496.050 298.050 ;
        RECT 487.950 296.400 496.050 297.600 ;
        RECT 487.950 295.950 490.050 296.400 ;
        RECT 493.950 295.950 496.050 296.400 ;
        RECT 523.950 297.600 526.050 298.050 ;
        RECT 550.950 297.600 553.050 298.050 ;
        RECT 523.950 296.400 553.050 297.600 ;
        RECT 523.950 295.950 526.050 296.400 ;
        RECT 550.950 295.950 553.050 296.400 ;
        RECT 595.950 297.600 600.000 298.050 ;
        RECT 619.950 297.600 622.050 298.050 ;
        RECT 595.950 295.950 600.600 297.600 ;
        RECT 298.950 294.600 301.050 295.200 ;
        RECT 298.950 293.400 306.600 294.600 ;
        RECT 298.950 293.100 301.050 293.400 ;
        RECT 296.400 291.000 303.600 291.600 ;
        RECT 296.400 290.400 304.050 291.000 ;
        RECT 293.400 287.400 297.600 288.600 ;
        RECT 271.950 286.800 274.050 287.250 ;
        RECT 283.950 286.800 286.050 287.250 ;
        RECT 124.950 285.600 127.050 286.050 ;
        RECT 142.950 285.600 145.050 286.050 ;
        RECT 124.950 284.400 145.050 285.600 ;
        RECT 124.950 283.950 127.050 284.400 ;
        RECT 142.950 283.950 145.050 284.400 ;
        RECT 268.950 283.950 271.050 286.050 ;
        RECT 296.400 285.600 297.600 287.400 ;
        RECT 301.950 286.950 304.050 290.400 ;
        RECT 305.400 288.600 306.600 293.400 ;
        RECT 316.950 293.100 319.050 295.200 ;
        RECT 334.950 294.600 337.050 295.200 ;
        RECT 379.950 294.600 382.050 295.200 ;
        RECT 334.950 293.400 382.050 294.600 ;
        RECT 334.950 293.100 337.050 293.400 ;
        RECT 379.950 293.100 382.050 293.400 ;
        RECT 385.950 294.600 388.050 295.200 ;
        RECT 403.950 294.600 406.050 295.200 ;
        RECT 385.950 293.400 406.050 294.600 ;
        RECT 385.950 293.100 388.050 293.400 ;
        RECT 403.950 293.100 406.050 293.400 ;
        RECT 424.950 294.600 427.050 295.200 ;
        RECT 478.950 294.600 481.050 295.200 ;
        RECT 424.950 293.400 481.050 294.600 ;
        RECT 424.950 293.100 427.050 293.400 ;
        RECT 478.950 293.100 481.050 293.400 ;
        RECT 499.950 294.600 502.050 295.050 ;
        RECT 520.950 294.600 523.050 295.050 ;
        RECT 499.950 293.400 523.050 294.600 ;
        RECT 313.950 288.600 316.050 288.900 ;
        RECT 305.400 287.400 316.050 288.600 ;
        RECT 317.400 288.600 318.600 293.100 ;
        RECT 499.950 292.950 502.050 293.400 ;
        RECT 520.950 292.950 523.050 293.400 ;
        RECT 535.950 294.600 538.050 295.200 ;
        RECT 599.400 295.050 600.600 295.950 ;
        RECT 611.400 296.400 622.050 297.600 ;
        RECT 544.950 294.600 547.050 295.050 ;
        RECT 565.800 294.600 567.900 295.050 ;
        RECT 535.950 293.400 543.600 294.600 ;
        RECT 535.950 293.100 538.050 293.400 ;
        RECT 325.950 291.600 330.000 292.050 ;
        RECT 542.400 291.600 543.600 293.400 ;
        RECT 544.950 293.400 567.900 294.600 ;
        RECT 544.950 292.950 547.050 293.400 ;
        RECT 565.800 292.950 567.900 293.400 ;
        RECT 568.950 294.600 571.050 295.050 ;
        RECT 583.950 294.600 586.050 295.050 ;
        RECT 568.950 293.400 586.050 294.600 ;
        RECT 568.950 292.950 571.050 293.400 ;
        RECT 583.950 292.950 586.050 293.400 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 325.950 289.950 330.600 291.600 ;
        RECT 542.400 290.400 567.600 291.600 ;
        RECT 325.950 288.600 328.050 288.900 ;
        RECT 317.400 287.400 328.050 288.600 ;
        RECT 329.400 288.600 330.600 289.950 ;
        RECT 337.950 288.600 340.050 288.900 ;
        RECT 329.400 287.400 340.050 288.600 ;
        RECT 313.950 286.800 316.050 287.400 ;
        RECT 325.950 286.800 328.050 287.400 ;
        RECT 337.950 286.800 340.050 287.400 ;
        RECT 367.950 288.600 370.050 288.900 ;
        RECT 382.950 288.600 385.050 288.900 ;
        RECT 367.950 287.400 385.050 288.600 ;
        RECT 367.950 286.800 370.050 287.400 ;
        RECT 382.950 286.800 385.050 287.400 ;
        RECT 400.950 288.600 403.050 288.900 ;
        RECT 415.950 288.600 418.050 288.900 ;
        RECT 430.950 288.600 433.050 289.050 ;
        RECT 439.950 288.600 442.050 288.900 ;
        RECT 400.950 287.400 442.050 288.600 ;
        RECT 400.950 286.800 403.050 287.400 ;
        RECT 415.950 286.800 418.050 287.400 ;
        RECT 430.950 286.950 433.050 287.400 ;
        RECT 439.950 286.800 442.050 287.400 ;
        RECT 472.950 288.450 475.050 288.900 ;
        RECT 481.950 288.450 484.050 288.900 ;
        RECT 472.950 287.250 484.050 288.450 ;
        RECT 472.950 286.800 475.050 287.250 ;
        RECT 481.950 286.800 484.050 287.250 ;
        RECT 496.950 288.450 499.050 288.900 ;
        RECT 502.950 288.450 505.050 288.900 ;
        RECT 496.950 287.250 505.050 288.450 ;
        RECT 496.950 286.800 499.050 287.250 ;
        RECT 502.950 286.800 505.050 287.250 ;
        RECT 514.950 288.450 517.050 288.900 ;
        RECT 520.950 288.450 523.050 288.900 ;
        RECT 514.950 287.250 523.050 288.450 ;
        RECT 514.950 286.800 517.050 287.250 ;
        RECT 520.950 286.800 523.050 287.250 ;
        RECT 532.950 288.600 535.050 288.900 ;
        RECT 541.950 288.600 544.050 289.050 ;
        RECT 547.950 288.600 550.050 288.900 ;
        RECT 532.950 287.400 550.050 288.600 ;
        RECT 566.400 288.600 567.600 290.400 ;
        RECT 601.950 288.600 604.050 289.050 ;
        RECT 611.400 288.600 612.600 296.400 ;
        RECT 619.950 295.950 622.050 296.400 ;
        RECT 664.950 297.600 667.050 298.050 ;
        RECT 691.950 297.600 694.050 298.050 ;
        RECT 664.950 296.400 694.050 297.600 ;
        RECT 664.950 295.950 667.050 296.400 ;
        RECT 691.950 295.950 694.050 296.400 ;
        RECT 715.950 297.600 718.050 298.050 ;
        RECT 853.950 297.600 856.050 298.050 ;
        RECT 862.950 297.600 865.050 298.050 ;
        RECT 715.950 296.400 726.600 297.600 ;
        RECT 715.950 295.950 718.050 296.400 ;
        RECT 622.950 292.950 625.050 295.050 ;
        RECT 646.950 292.950 649.050 295.050 ;
        RECT 652.950 294.600 657.000 295.050 ;
        RECT 694.950 294.600 697.050 295.200 ;
        RECT 652.950 292.950 657.600 294.600 ;
        RECT 566.400 287.400 579.600 288.600 ;
        RECT 532.950 286.800 535.050 287.400 ;
        RECT 541.950 286.950 544.050 287.400 ;
        RECT 547.950 286.800 550.050 287.400 ;
        RECT 578.400 286.050 579.600 287.400 ;
        RECT 601.950 287.400 612.600 288.600 ;
        RECT 616.950 288.600 619.050 288.900 ;
        RECT 623.400 288.600 624.600 292.950 ;
        RECT 616.950 287.400 624.600 288.600 ;
        RECT 643.950 288.600 646.050 288.900 ;
        RECT 647.400 288.600 648.600 292.950 ;
        RECT 656.400 288.900 657.600 292.950 ;
        RECT 683.400 293.400 697.050 294.600 ;
        RECT 683.400 289.050 684.600 293.400 ;
        RECT 694.950 293.100 697.050 293.400 ;
        RECT 725.400 292.050 726.600 296.400 ;
        RECT 853.950 296.400 865.050 297.600 ;
        RECT 853.950 295.950 856.050 296.400 ;
        RECT 862.950 295.950 865.050 296.400 ;
        RECT 730.950 294.750 733.050 295.200 ;
        RECT 736.950 294.750 739.050 295.200 ;
        RECT 730.950 293.550 739.050 294.750 ;
        RECT 730.950 293.100 733.050 293.550 ;
        RECT 736.950 293.100 739.050 293.550 ;
        RECT 742.950 293.100 745.050 295.200 ;
        RECT 760.950 293.100 763.050 295.200 ;
        RECT 802.950 294.600 805.050 295.200 ;
        RECT 823.950 294.600 826.050 295.200 ;
        RECT 802.950 293.400 826.050 294.600 ;
        RECT 802.950 293.100 805.050 293.400 ;
        RECT 823.950 293.100 826.050 293.400 ;
        RECT 835.950 294.750 838.050 295.200 ;
        RECT 841.950 294.750 844.050 295.200 ;
        RECT 835.950 293.550 844.050 294.750 ;
        RECT 877.950 294.600 880.050 295.050 ;
        RECT 835.950 293.100 838.050 293.550 ;
        RECT 841.950 293.100 844.050 293.550 ;
        RECT 863.400 293.400 880.050 294.600 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 643.950 287.400 648.600 288.600 ;
        RECT 655.950 288.600 658.050 288.900 ;
        RECT 679.800 288.600 681.900 288.900 ;
        RECT 655.950 287.400 681.900 288.600 ;
        RECT 601.950 286.950 604.050 287.400 ;
        RECT 616.950 286.800 619.050 287.400 ;
        RECT 643.950 286.800 646.050 287.400 ;
        RECT 655.950 286.800 658.050 287.400 ;
        RECT 679.800 286.800 681.900 287.400 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 743.400 288.600 744.600 293.100 ;
        RECT 757.950 288.600 760.050 288.900 ;
        RECT 743.400 287.400 760.050 288.600 ;
        RECT 761.400 288.600 762.600 293.100 ;
        RECT 778.950 288.600 781.050 288.900 ;
        RECT 761.400 287.400 781.050 288.600 ;
        RECT 757.950 286.800 760.050 287.400 ;
        RECT 778.950 286.800 781.050 287.400 ;
        RECT 824.400 286.050 825.600 293.100 ;
        RECT 863.400 288.900 864.600 293.400 ;
        RECT 877.950 292.950 880.050 293.400 ;
        RECT 887.400 288.900 888.600 299.400 ;
        RECT 889.950 298.950 892.050 299.400 ;
        RECT 901.950 298.950 904.050 299.400 ;
        RECT 889.950 294.750 892.050 295.200 ;
        RECT 895.950 294.750 898.050 295.200 ;
        RECT 889.950 293.550 898.050 294.750 ;
        RECT 889.950 293.100 892.050 293.550 ;
        RECT 895.950 293.100 898.050 293.550 ;
        RECT 913.950 294.600 916.050 295.050 ;
        RECT 931.950 294.600 934.050 294.900 ;
        RECT 913.950 293.400 934.050 294.600 ;
        RECT 913.950 292.950 916.050 293.400 ;
        RECT 931.950 292.800 934.050 293.400 ;
        RECT 844.950 288.600 847.050 288.900 ;
        RECT 862.950 288.600 865.050 288.900 ;
        RECT 844.950 287.400 865.050 288.600 ;
        RECT 844.950 286.800 847.050 287.400 ;
        RECT 862.950 286.800 865.050 287.400 ;
        RECT 886.950 286.800 889.050 288.900 ;
        RECT 895.950 288.450 898.050 288.900 ;
        RECT 904.950 288.450 907.050 288.900 ;
        RECT 895.950 287.250 907.050 288.450 ;
        RECT 895.950 286.800 898.050 287.250 ;
        RECT 904.950 286.800 907.050 287.250 ;
        RECT 310.950 285.600 313.050 286.050 ;
        RECT 296.400 284.400 313.050 285.600 ;
        RECT 578.400 284.400 583.050 286.050 ;
        RECT 310.950 283.950 313.050 284.400 ;
        RECT 579.000 283.950 583.050 284.400 ;
        RECT 589.950 285.600 592.050 286.050 ;
        RECT 595.950 285.600 598.050 286.050 ;
        RECT 589.950 284.400 598.050 285.600 ;
        RECT 589.950 283.950 592.050 284.400 ;
        RECT 595.950 283.950 598.050 284.400 ;
        RECT 730.950 285.600 733.050 286.050 ;
        RECT 766.950 285.600 769.050 286.050 ;
        RECT 730.950 284.400 769.050 285.600 ;
        RECT 730.950 283.950 733.050 284.400 ;
        RECT 766.950 283.950 769.050 284.400 ;
        RECT 823.950 283.950 826.050 286.050 ;
        RECT 142.950 282.600 145.050 282.900 ;
        RECT 157.950 282.600 160.050 283.050 ;
        RECT 142.950 281.400 160.050 282.600 ;
        RECT 142.950 280.800 145.050 281.400 ;
        RECT 157.950 280.950 160.050 281.400 ;
        RECT 208.950 282.600 211.050 283.050 ;
        RECT 217.950 282.600 220.050 283.050 ;
        RECT 208.950 281.400 220.050 282.600 ;
        RECT 208.950 280.950 211.050 281.400 ;
        RECT 217.950 280.950 220.050 281.400 ;
        RECT 226.950 282.600 229.050 283.050 ;
        RECT 250.950 282.600 253.050 283.050 ;
        RECT 226.950 281.400 253.050 282.600 ;
        RECT 226.950 280.950 229.050 281.400 ;
        RECT 250.950 280.950 253.050 281.400 ;
        RECT 277.950 282.600 280.050 283.050 ;
        RECT 295.950 282.600 298.050 283.050 ;
        RECT 277.950 281.400 298.050 282.600 ;
        RECT 277.950 280.950 280.050 281.400 ;
        RECT 295.950 280.950 298.050 281.400 ;
        RECT 373.950 282.600 376.050 283.050 ;
        RECT 430.950 282.600 433.050 283.050 ;
        RECT 373.950 281.400 433.050 282.600 ;
        RECT 373.950 280.950 376.050 281.400 ;
        RECT 430.950 280.950 433.050 281.400 ;
        RECT 562.950 282.600 565.050 283.050 ;
        RECT 604.950 282.600 607.050 283.050 ;
        RECT 562.950 281.400 607.050 282.600 ;
        RECT 562.950 280.950 565.050 281.400 ;
        RECT 604.950 280.950 607.050 281.400 ;
        RECT 643.950 282.600 646.050 283.050 ;
        RECT 658.950 282.600 661.050 283.050 ;
        RECT 643.950 281.400 661.050 282.600 ;
        RECT 643.950 280.950 646.050 281.400 ;
        RECT 658.950 280.950 661.050 281.400 ;
        RECT 688.950 282.600 691.050 283.050 ;
        RECT 712.950 282.600 715.050 283.050 ;
        RECT 688.950 281.400 715.050 282.600 ;
        RECT 688.950 280.950 691.050 281.400 ;
        RECT 712.950 280.950 715.050 281.400 ;
        RECT 739.950 282.600 742.050 283.050 ;
        RECT 748.950 282.600 751.050 283.050 ;
        RECT 739.950 281.400 751.050 282.600 ;
        RECT 739.950 280.950 742.050 281.400 ;
        RECT 748.950 280.950 751.050 281.400 ;
        RECT 787.950 282.600 790.050 283.050 ;
        RECT 799.950 282.600 802.050 283.050 ;
        RECT 820.950 282.600 823.050 283.050 ;
        RECT 787.950 281.400 823.050 282.600 ;
        RECT 787.950 280.950 790.050 281.400 ;
        RECT 799.950 280.950 802.050 281.400 ;
        RECT 820.950 280.950 823.050 281.400 ;
        RECT 112.950 279.600 115.050 280.050 ;
        RECT 89.400 279.000 115.050 279.600 ;
        RECT 88.950 278.400 115.050 279.000 ;
        RECT 49.950 276.600 52.050 277.050 ;
        RECT 55.950 276.600 58.050 277.050 ;
        RECT 49.950 275.400 58.050 276.600 ;
        RECT 49.950 274.950 52.050 275.400 ;
        RECT 55.950 274.950 58.050 275.400 ;
        RECT 64.950 276.600 67.050 277.050 ;
        RECT 82.950 276.600 85.050 277.050 ;
        RECT 64.950 275.400 85.050 276.600 ;
        RECT 64.950 274.950 67.050 275.400 ;
        RECT 82.950 274.950 85.050 275.400 ;
        RECT 88.950 274.950 91.050 278.400 ;
        RECT 112.950 277.950 115.050 278.400 ;
        RECT 376.950 279.600 379.050 280.050 ;
        RECT 415.950 279.600 418.050 280.050 ;
        RECT 376.950 278.400 418.050 279.600 ;
        RECT 376.950 277.950 379.050 278.400 ;
        RECT 415.950 277.950 418.050 278.400 ;
        RECT 559.950 279.600 562.050 280.050 ;
        RECT 574.950 279.600 577.050 280.050 ;
        RECT 559.950 278.400 577.050 279.600 ;
        RECT 559.950 277.950 562.050 278.400 ;
        RECT 574.950 277.950 577.050 278.400 ;
        RECT 580.950 279.600 583.050 280.050 ;
        RECT 601.950 279.600 604.050 280.050 ;
        RECT 580.950 278.400 604.050 279.600 ;
        RECT 580.950 277.950 583.050 278.400 ;
        RECT 601.950 277.950 604.050 278.400 ;
        RECT 610.950 279.600 613.050 280.050 ;
        RECT 625.950 279.600 628.050 280.050 ;
        RECT 610.950 278.400 628.050 279.600 ;
        RECT 610.950 277.950 613.050 278.400 ;
        RECT 625.950 277.950 628.050 278.400 ;
        RECT 673.950 279.600 676.050 280.050 ;
        RECT 706.950 279.600 709.050 280.050 ;
        RECT 673.950 278.400 709.050 279.600 ;
        RECT 673.950 277.950 676.050 278.400 ;
        RECT 706.950 277.950 709.050 278.400 ;
        RECT 757.950 279.600 760.050 280.050 ;
        RECT 775.950 279.600 778.050 280.050 ;
        RECT 757.950 278.400 778.050 279.600 ;
        RECT 757.950 277.950 760.050 278.400 ;
        RECT 775.950 277.950 778.050 278.400 ;
        RECT 868.950 279.600 871.050 280.050 ;
        RECT 883.950 279.600 886.050 280.050 ;
        RECT 898.950 279.600 901.050 280.050 ;
        RECT 868.950 278.400 901.050 279.600 ;
        RECT 868.950 277.950 871.050 278.400 ;
        RECT 883.950 277.950 886.050 278.400 ;
        RECT 898.950 277.950 901.050 278.400 ;
        RECT 100.950 276.600 103.050 277.050 ;
        RECT 145.950 276.600 148.050 277.050 ;
        RECT 100.950 275.400 148.050 276.600 ;
        RECT 100.950 274.950 103.050 275.400 ;
        RECT 145.950 274.950 148.050 275.400 ;
        RECT 187.950 276.600 190.050 277.050 ;
        RECT 220.950 276.600 223.050 277.050 ;
        RECT 259.950 276.600 262.050 277.050 ;
        RECT 187.950 275.400 262.050 276.600 ;
        RECT 187.950 274.950 190.050 275.400 ;
        RECT 220.950 274.950 223.050 275.400 ;
        RECT 259.950 274.950 262.050 275.400 ;
        RECT 289.950 276.600 292.050 277.050 ;
        RECT 307.950 276.600 310.050 277.050 ;
        RECT 325.950 276.600 328.050 277.050 ;
        RECT 358.950 276.600 361.050 277.050 ;
        RECT 370.950 276.600 373.050 277.050 ;
        RECT 289.950 275.400 357.600 276.600 ;
        RECT 289.950 274.950 292.050 275.400 ;
        RECT 307.950 274.950 310.050 275.400 ;
        RECT 325.950 274.950 328.050 275.400 ;
        RECT 13.950 273.600 16.050 274.050 ;
        RECT 46.950 273.600 49.050 274.050 ;
        RECT 13.950 272.400 49.050 273.600 ;
        RECT 13.950 271.950 16.050 272.400 ;
        RECT 46.950 271.950 49.050 272.400 ;
        RECT 97.950 273.600 100.050 274.050 ;
        RECT 130.950 273.600 133.050 274.050 ;
        RECT 214.950 273.600 217.050 274.050 ;
        RECT 97.950 272.400 133.050 273.600 ;
        RECT 182.400 273.000 217.050 273.600 ;
        RECT 97.950 271.950 100.050 272.400 ;
        RECT 130.950 271.950 133.050 272.400 ;
        RECT 181.950 272.400 217.050 273.000 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 112.950 270.600 115.050 271.050 ;
        RECT 106.950 269.400 115.050 270.600 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 112.950 268.950 115.050 269.400 ;
        RECT 181.950 268.950 184.050 272.400 ;
        RECT 214.950 271.950 217.050 272.400 ;
        RECT 223.950 273.600 226.050 274.050 ;
        RECT 238.950 273.600 241.050 274.050 ;
        RECT 223.950 272.400 241.050 273.600 ;
        RECT 223.950 271.950 226.050 272.400 ;
        RECT 238.950 271.950 241.050 272.400 ;
        RECT 313.950 273.600 316.050 274.050 ;
        RECT 328.950 273.600 331.050 274.050 ;
        RECT 313.950 272.400 331.050 273.600 ;
        RECT 356.400 273.600 357.600 275.400 ;
        RECT 358.950 275.400 373.050 276.600 ;
        RECT 358.950 274.950 361.050 275.400 ;
        RECT 370.950 274.950 373.050 275.400 ;
        RECT 508.950 276.600 511.050 277.050 ;
        RECT 547.950 276.600 550.050 277.050 ;
        RECT 508.950 275.400 550.050 276.600 ;
        RECT 508.950 274.950 511.050 275.400 ;
        RECT 547.950 274.950 550.050 275.400 ;
        RECT 565.950 276.600 568.050 277.050 ;
        RECT 622.950 276.600 625.050 277.050 ;
        RECT 691.950 276.600 694.050 277.050 ;
        RECT 565.950 275.400 694.050 276.600 ;
        RECT 565.950 274.950 568.050 275.400 ;
        RECT 622.950 274.950 625.050 275.400 ;
        RECT 691.950 274.950 694.050 275.400 ;
        RECT 778.950 276.600 781.050 277.050 ;
        RECT 793.950 276.600 796.050 277.050 ;
        RECT 778.950 275.400 796.050 276.600 ;
        RECT 778.950 274.950 781.050 275.400 ;
        RECT 793.950 274.950 796.050 275.400 ;
        RECT 370.950 273.600 373.050 273.900 ;
        RECT 356.400 272.400 373.050 273.600 ;
        RECT 313.950 271.950 316.050 272.400 ;
        RECT 328.950 271.950 331.050 272.400 ;
        RECT 370.950 271.800 373.050 272.400 ;
        RECT 421.950 273.600 424.050 274.050 ;
        RECT 466.950 273.600 469.050 274.050 ;
        RECT 421.950 272.400 469.050 273.600 ;
        RECT 421.950 271.950 424.050 272.400 ;
        RECT 466.950 271.950 469.050 272.400 ;
        RECT 640.950 273.600 643.050 274.050 ;
        RECT 664.950 273.600 667.050 274.050 ;
        RECT 640.950 272.400 667.050 273.600 ;
        RECT 640.950 271.950 643.050 272.400 ;
        RECT 664.950 271.950 667.050 272.400 ;
        RECT 763.950 273.600 766.050 274.050 ;
        RECT 772.950 273.600 775.050 274.050 ;
        RECT 763.950 272.400 775.050 273.600 ;
        RECT 763.950 271.950 766.050 272.400 ;
        RECT 772.950 271.950 775.050 272.400 ;
        RECT 808.950 273.600 811.050 274.050 ;
        RECT 814.950 273.600 817.050 274.050 ;
        RECT 829.950 273.600 832.050 274.050 ;
        RECT 868.950 273.600 871.050 274.050 ;
        RECT 808.950 272.400 871.050 273.600 ;
        RECT 808.950 271.950 811.050 272.400 ;
        RECT 814.950 271.950 817.050 272.400 ;
        RECT 829.950 271.950 832.050 272.400 ;
        RECT 868.950 271.950 871.050 272.400 ;
        RECT 196.950 270.600 199.050 271.050 ;
        RECT 202.950 270.600 205.050 271.050 ;
        RECT 196.950 269.400 205.050 270.600 ;
        RECT 196.950 268.950 199.050 269.400 ;
        RECT 202.950 268.950 205.050 269.400 ;
        RECT 247.950 270.600 250.050 271.050 ;
        RECT 262.950 270.600 265.050 271.050 ;
        RECT 247.950 269.400 265.050 270.600 ;
        RECT 247.950 268.950 250.050 269.400 ;
        RECT 262.950 268.950 265.050 269.400 ;
        RECT 328.950 270.600 331.050 270.900 ;
        RECT 382.950 270.600 385.050 271.050 ;
        RECT 328.950 269.400 385.050 270.600 ;
        RECT 328.950 268.800 331.050 269.400 ;
        RECT 382.950 268.950 385.050 269.400 ;
        RECT 451.950 270.600 454.050 271.050 ;
        RECT 460.950 270.600 463.050 271.050 ;
        RECT 451.950 269.400 463.050 270.600 ;
        RECT 451.950 268.950 454.050 269.400 ;
        RECT 460.950 268.950 463.050 269.400 ;
        RECT 523.950 270.600 526.050 271.050 ;
        RECT 541.950 270.600 544.050 271.050 ;
        RECT 523.950 269.400 544.050 270.600 ;
        RECT 523.950 268.950 526.050 269.400 ;
        RECT 541.950 268.950 544.050 269.400 ;
        RECT 568.950 270.600 571.050 271.050 ;
        RECT 586.950 270.600 589.050 271.050 ;
        RECT 568.950 269.400 589.050 270.600 ;
        RECT 568.950 268.950 571.050 269.400 ;
        RECT 586.950 268.950 589.050 269.400 ;
        RECT 598.950 270.600 601.050 271.050 ;
        RECT 610.950 270.600 613.050 271.050 ;
        RECT 598.950 269.400 613.050 270.600 ;
        RECT 598.950 268.950 601.050 269.400 ;
        RECT 610.950 268.950 613.050 269.400 ;
        RECT 631.950 270.600 634.050 271.050 ;
        RECT 676.950 270.600 679.050 271.050 ;
        RECT 694.950 270.600 697.050 271.050 ;
        RECT 631.950 269.400 697.050 270.600 ;
        RECT 631.950 268.950 634.050 269.400 ;
        RECT 676.950 268.950 679.050 269.400 ;
        RECT 694.950 268.950 697.050 269.400 ;
        RECT 709.950 270.600 712.050 271.050 ;
        RECT 730.950 270.600 733.050 271.050 ;
        RECT 709.950 269.400 733.050 270.600 ;
        RECT 709.950 268.950 712.050 269.400 ;
        RECT 730.950 268.950 733.050 269.400 ;
        RECT 775.950 270.600 778.050 271.050 ;
        RECT 826.950 270.600 829.050 271.050 ;
        RECT 775.950 269.400 829.050 270.600 ;
        RECT 775.950 268.950 778.050 269.400 ;
        RECT 826.950 268.950 829.050 269.400 ;
        RECT 94.950 267.600 97.050 268.050 ;
        RECT 115.950 267.600 118.050 268.050 ;
        RECT 94.950 266.400 118.050 267.600 ;
        RECT 94.950 265.950 97.050 266.400 ;
        RECT 115.950 265.950 118.050 266.400 ;
        RECT 172.950 267.600 175.050 268.050 ;
        RECT 202.950 267.600 205.050 267.900 ;
        RECT 172.950 266.400 205.050 267.600 ;
        RECT 172.950 265.950 175.050 266.400 ;
        RECT 202.950 265.800 205.050 266.400 ;
        RECT 274.950 267.600 277.050 268.050 ;
        RECT 280.950 267.600 283.050 268.050 ;
        RECT 274.950 266.400 283.050 267.600 ;
        RECT 274.950 265.950 277.050 266.400 ;
        RECT 280.950 265.950 283.050 266.400 ;
        RECT 370.950 267.600 373.050 268.050 ;
        RECT 478.950 267.600 481.050 268.050 ;
        RECT 559.950 267.600 562.050 268.050 ;
        RECT 574.950 267.600 577.050 268.050 ;
        RECT 370.950 266.400 528.600 267.600 ;
        RECT 370.950 265.950 373.050 266.400 ;
        RECT 478.950 265.950 481.050 266.400 ;
        RECT 4.950 264.600 7.050 265.050 ;
        RECT 10.950 264.600 13.050 265.050 ;
        RECT 4.950 263.400 13.050 264.600 ;
        RECT 4.950 262.950 7.050 263.400 ;
        RECT 10.950 262.950 13.050 263.400 ;
        RECT 100.950 261.600 105.000 262.050 ;
        RECT 115.950 261.600 118.050 262.050 ;
        RECT 124.950 261.600 127.050 262.200 ;
        RECT 100.950 259.950 105.600 261.600 ;
        RECT 115.950 260.400 127.050 261.600 ;
        RECT 115.950 259.950 118.050 260.400 ;
        RECT 124.950 260.100 127.050 260.400 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 151.950 261.750 154.050 262.200 ;
        RECT 166.950 261.750 169.050 262.200 ;
        RECT 151.950 260.550 169.050 261.750 ;
        RECT 151.950 260.100 154.050 260.550 ;
        RECT 166.950 260.100 169.050 260.550 ;
        RECT 184.950 261.600 189.000 262.050 ;
        RECT 190.950 261.600 193.050 262.200 ;
        RECT 199.950 261.600 204.000 262.050 ;
        RECT 226.950 261.600 229.050 265.050 ;
        RECT 184.950 259.950 189.600 261.600 ;
        RECT 190.950 260.400 198.600 261.600 ;
        RECT 190.950 260.100 193.050 260.400 ;
        RECT 19.950 258.450 22.050 258.900 ;
        RECT 40.800 258.450 42.900 258.900 ;
        RECT 19.950 257.250 42.900 258.450 ;
        RECT 19.950 256.800 22.050 257.250 ;
        RECT 40.800 256.800 42.900 257.250 ;
        RECT 43.950 258.600 46.050 259.050 ;
        RECT 61.950 258.600 64.050 259.050 ;
        RECT 43.950 257.400 64.050 258.600 ;
        RECT 43.950 256.950 46.050 257.400 ;
        RECT 61.950 256.950 64.050 257.400 ;
        RECT 104.400 255.900 105.600 259.950 ;
        RECT 70.950 255.450 73.050 255.900 ;
        RECT 85.950 255.450 88.050 255.900 ;
        RECT 70.950 254.250 88.050 255.450 ;
        RECT 70.950 253.800 73.050 254.250 ;
        RECT 85.950 253.800 88.050 254.250 ;
        RECT 103.950 253.800 106.050 255.900 ;
        RECT 136.950 255.600 139.050 256.050 ;
        RECT 143.400 255.600 144.600 259.950 ;
        RECT 188.400 258.600 189.600 259.950 ;
        RECT 155.400 257.400 189.600 258.600 ;
        RECT 197.400 258.600 198.600 260.400 ;
        RECT 199.950 259.950 204.600 261.600 ;
        RECT 226.950 261.000 234.600 261.600 ;
        RECT 227.400 260.400 234.600 261.000 ;
        RECT 203.400 258.600 204.600 259.950 ;
        RECT 197.400 258.000 201.600 258.600 ;
        RECT 197.400 257.400 202.050 258.000 ;
        RECT 203.400 257.400 213.600 258.600 ;
        RECT 155.400 255.900 156.600 257.400 ;
        RECT 188.400 255.900 189.600 257.400 ;
        RECT 136.950 254.400 144.600 255.600 ;
        RECT 136.950 253.950 139.050 254.400 ;
        RECT 154.950 253.800 157.050 255.900 ;
        RECT 163.950 255.450 166.050 255.900 ;
        RECT 169.950 255.450 172.050 255.900 ;
        RECT 163.950 254.250 172.050 255.450 ;
        RECT 163.950 253.800 166.050 254.250 ;
        RECT 169.950 253.800 172.050 254.250 ;
        RECT 175.950 255.450 178.050 255.900 ;
        RECT 181.950 255.450 184.050 255.900 ;
        RECT 175.950 254.250 184.050 255.450 ;
        RECT 175.950 253.800 178.050 254.250 ;
        RECT 181.950 253.800 184.050 254.250 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 199.950 253.950 202.050 257.400 ;
        RECT 212.400 255.900 213.600 257.400 ;
        RECT 233.400 256.050 234.600 260.400 ;
        RECT 238.950 260.100 241.050 262.200 ;
        RECT 239.400 258.600 240.600 260.100 ;
        RECT 244.950 259.950 247.050 262.050 ;
        RECT 256.950 261.600 259.050 262.200 ;
        RECT 251.400 260.400 259.050 261.600 ;
        RECT 271.950 261.600 274.050 265.050 ;
        RECT 289.950 264.600 292.050 265.050 ;
        RECT 298.950 264.600 301.050 265.050 ;
        RECT 322.950 264.600 325.050 265.050 ;
        RECT 289.950 263.400 301.050 264.600 ;
        RECT 289.950 262.950 292.050 263.400 ;
        RECT 298.950 262.950 301.050 263.400 ;
        RECT 314.400 263.400 325.050 264.600 ;
        RECT 280.950 261.600 283.050 262.200 ;
        RECT 304.950 261.600 307.050 262.050 ;
        RECT 271.950 261.000 283.050 261.600 ;
        RECT 272.400 260.400 283.050 261.000 ;
        RECT 239.400 257.400 243.600 258.600 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 232.950 253.950 235.050 256.050 ;
        RECT 64.950 252.450 67.050 252.900 ;
        RECT 94.950 252.450 97.050 252.900 ;
        RECT 64.950 251.250 97.050 252.450 ;
        RECT 242.400 252.600 243.600 257.400 ;
        RECT 245.400 256.050 246.600 259.950 ;
        RECT 251.400 256.050 252.600 260.400 ;
        RECT 256.950 260.100 259.050 260.400 ;
        RECT 280.950 260.100 283.050 260.400 ;
        RECT 296.400 260.400 307.050 261.600 ;
        RECT 244.950 253.950 247.050 256.050 ;
        RECT 250.950 253.950 253.050 256.050 ;
        RECT 296.400 255.900 297.600 260.400 ;
        RECT 304.950 259.950 307.050 260.400 ;
        RECT 314.400 256.050 315.600 263.400 ;
        RECT 322.950 262.950 325.050 263.400 ;
        RECT 334.950 264.600 337.050 265.050 ;
        RECT 346.950 264.600 349.050 265.050 ;
        RECT 367.950 264.600 370.050 265.050 ;
        RECT 334.950 263.400 370.050 264.600 ;
        RECT 334.950 262.950 337.050 263.400 ;
        RECT 346.950 262.950 349.050 263.400 ;
        RECT 367.950 262.950 370.050 263.400 ;
        RECT 316.950 261.600 319.050 262.200 ;
        RECT 343.950 261.600 346.050 262.200 ;
        RECT 316.950 260.400 346.050 261.600 ;
        RECT 316.950 260.100 319.050 260.400 ;
        RECT 343.950 260.100 346.050 260.400 ;
        RECT 361.950 261.600 364.050 262.050 ;
        RECT 373.950 261.600 376.050 262.050 ;
        RECT 361.950 260.400 376.050 261.600 ;
        RECT 361.950 259.950 364.050 260.400 ;
        RECT 373.950 259.950 376.050 260.400 ;
        RECT 421.950 261.600 424.050 262.200 ;
        RECT 436.950 261.750 439.050 262.200 ;
        RECT 445.950 261.750 448.050 262.200 ;
        RECT 436.950 261.600 448.050 261.750 ;
        RECT 421.950 260.550 448.050 261.600 ;
        RECT 421.950 260.400 439.050 260.550 ;
        RECT 421.950 260.100 424.050 260.400 ;
        RECT 436.950 260.100 439.050 260.400 ;
        RECT 445.950 260.100 448.050 260.550 ;
        RECT 457.950 260.100 460.050 262.200 ;
        RECT 469.950 261.750 472.050 262.200 ;
        RECT 484.950 261.750 487.050 262.200 ;
        RECT 469.950 260.550 487.050 261.750 ;
        RECT 496.950 261.600 499.050 262.200 ;
        RECT 469.950 260.100 472.050 260.550 ;
        RECT 484.950 260.100 487.050 260.550 ;
        RECT 494.400 260.400 499.050 261.600 ;
        RECT 259.950 255.600 262.050 255.900 ;
        RECT 268.950 255.600 271.050 255.900 ;
        RECT 259.950 255.450 271.050 255.600 ;
        RECT 277.950 255.450 280.050 255.900 ;
        RECT 259.950 254.400 280.050 255.450 ;
        RECT 259.950 253.800 262.050 254.400 ;
        RECT 268.950 254.250 280.050 254.400 ;
        RECT 268.950 253.800 271.050 254.250 ;
        RECT 277.950 253.800 280.050 254.250 ;
        RECT 295.950 253.800 298.050 255.900 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 325.950 255.450 328.050 255.900 ;
        RECT 334.950 255.450 337.050 255.900 ;
        RECT 325.950 254.250 337.050 255.450 ;
        RECT 325.950 253.800 328.050 254.250 ;
        RECT 334.950 253.800 337.050 254.250 ;
        RECT 346.950 255.450 349.050 255.900 ;
        RECT 358.950 255.450 361.050 255.900 ;
        RECT 346.950 254.250 361.050 255.450 ;
        RECT 458.400 255.600 459.600 260.100 ;
        RECT 494.400 256.050 495.600 260.400 ;
        RECT 496.950 260.100 499.050 260.400 ;
        RECT 502.950 261.750 505.050 262.200 ;
        RECT 511.950 261.750 514.050 262.200 ;
        RECT 502.950 260.550 514.050 261.750 ;
        RECT 502.950 260.100 505.050 260.550 ;
        RECT 511.950 260.100 514.050 260.550 ;
        RECT 527.400 261.600 528.600 266.400 ;
        RECT 559.950 266.400 577.050 267.600 ;
        RECT 559.950 265.950 562.050 266.400 ;
        RECT 574.950 265.950 577.050 266.400 ;
        RECT 604.950 267.600 607.050 268.050 ;
        RECT 613.950 267.600 616.050 268.050 ;
        RECT 604.950 266.400 616.050 267.600 ;
        RECT 604.950 265.950 607.050 266.400 ;
        RECT 613.950 265.950 616.050 266.400 ;
        RECT 649.950 267.600 652.050 268.050 ;
        RECT 661.950 267.600 664.050 268.050 ;
        RECT 649.950 266.400 664.050 267.600 ;
        RECT 649.950 265.950 652.050 266.400 ;
        RECT 661.950 265.950 664.050 266.400 ;
        RECT 715.950 267.600 718.050 268.050 ;
        RECT 748.950 267.600 751.050 268.050 ;
        RECT 715.950 266.400 751.050 267.600 ;
        RECT 715.950 265.950 718.050 266.400 ;
        RECT 748.950 265.950 751.050 266.400 ;
        RECT 754.950 267.600 757.050 268.050 ;
        RECT 802.950 267.600 805.050 268.050 ;
        RECT 754.950 266.400 805.050 267.600 ;
        RECT 754.950 265.950 757.050 266.400 ;
        RECT 802.950 265.950 805.050 266.400 ;
        RECT 862.950 267.600 865.050 268.050 ;
        RECT 874.950 267.600 877.050 268.050 ;
        RECT 862.950 266.400 877.050 267.600 ;
        RECT 862.950 265.950 865.050 266.400 ;
        RECT 874.950 265.950 877.050 266.400 ;
        RECT 886.950 267.600 889.050 268.050 ;
        RECT 916.950 267.600 919.050 268.050 ;
        RECT 886.950 266.400 919.050 267.600 ;
        RECT 886.950 265.950 889.050 266.400 ;
        RECT 916.950 265.950 919.050 266.400 ;
        RECT 529.950 264.600 532.050 265.050 ;
        RECT 553.950 264.600 556.050 265.050 ;
        RECT 529.950 263.400 556.050 264.600 ;
        RECT 529.950 262.950 532.050 263.400 ;
        RECT 553.950 262.950 556.050 263.400 ;
        RECT 583.950 264.600 586.050 265.050 ;
        RECT 589.950 264.600 592.050 265.050 ;
        RECT 583.950 263.400 592.050 264.600 ;
        RECT 583.950 262.950 586.050 263.400 ;
        RECT 589.950 262.950 592.050 263.400 ;
        RECT 700.950 262.950 703.050 265.050 ;
        RECT 784.950 264.600 787.050 265.050 ;
        RECT 793.950 264.600 796.050 265.050 ;
        RECT 784.950 263.400 796.050 264.600 ;
        RECT 784.950 262.950 787.050 263.400 ;
        RECT 793.950 262.950 796.050 263.400 ;
        RECT 853.950 264.600 856.050 265.050 ;
        RECT 859.950 264.600 862.050 265.050 ;
        RECT 853.950 263.400 862.050 264.600 ;
        RECT 853.950 262.950 856.050 263.400 ;
        RECT 859.950 262.950 862.050 263.400 ;
        RECT 550.950 261.600 553.050 262.050 ;
        RECT 556.950 261.600 559.050 262.200 ;
        RECT 527.400 260.400 559.050 261.600 ;
        RECT 550.950 259.950 553.050 260.400 ;
        RECT 556.950 260.100 559.050 260.400 ;
        RECT 562.950 261.600 565.050 262.200 ;
        RECT 580.950 261.600 583.050 262.200 ;
        RECT 586.950 261.600 589.050 262.050 ;
        RECT 562.950 260.400 579.600 261.600 ;
        RECT 562.950 260.100 565.050 260.400 ;
        RECT 481.950 255.600 484.050 255.900 ;
        RECT 458.400 254.400 484.050 255.600 ;
        RECT 346.950 253.800 349.050 254.250 ;
        RECT 358.950 253.800 361.050 254.250 ;
        RECT 481.950 253.800 484.050 254.400 ;
        RECT 493.950 253.950 496.050 256.050 ;
        RECT 578.400 255.900 579.600 260.400 ;
        RECT 580.950 260.400 589.050 261.600 ;
        RECT 580.950 260.100 583.050 260.400 ;
        RECT 586.950 259.950 589.050 260.400 ;
        RECT 607.950 261.600 610.050 262.050 ;
        RECT 625.950 261.600 628.050 262.050 ;
        RECT 607.950 260.400 615.600 261.600 ;
        RECT 607.950 259.950 610.050 260.400 ;
        RECT 505.950 255.600 508.050 255.900 ;
        RECT 520.950 255.600 523.050 255.900 ;
        RECT 505.950 254.400 523.050 255.600 ;
        RECT 505.950 253.800 508.050 254.400 ;
        RECT 520.950 253.800 523.050 254.400 ;
        RECT 577.950 253.800 580.050 255.900 ;
        RECT 583.950 255.600 586.050 255.900 ;
        RECT 595.950 255.600 598.050 255.900 ;
        RECT 601.950 255.600 604.050 256.050 ;
        RECT 583.950 254.400 604.050 255.600 ;
        RECT 583.950 253.800 586.050 254.400 ;
        RECT 595.950 253.800 598.050 254.400 ;
        RECT 601.950 253.950 604.050 254.400 ;
        RECT 614.400 253.050 615.600 260.400 ;
        RECT 620.400 260.400 628.050 261.600 ;
        RECT 620.400 255.600 621.600 260.400 ;
        RECT 625.950 259.950 628.050 260.400 ;
        RECT 637.950 261.750 640.050 262.200 ;
        RECT 649.950 261.750 652.050 262.200 ;
        RECT 637.950 260.550 652.050 261.750 ;
        RECT 637.950 260.100 640.050 260.550 ;
        RECT 649.950 260.100 652.050 260.550 ;
        RECT 655.950 261.600 658.050 262.200 ;
        RECT 664.950 261.600 667.050 262.050 ;
        RECT 670.950 261.600 673.050 262.200 ;
        RECT 681.000 261.600 685.050 262.050 ;
        RECT 655.950 260.400 660.600 261.600 ;
        RECT 655.950 260.100 658.050 260.400 ;
        RECT 622.950 258.600 625.050 259.050 ;
        RECT 622.950 257.400 648.600 258.600 ;
        RECT 622.950 256.950 625.050 257.400 ;
        RECT 647.400 255.900 648.600 257.400 ;
        RECT 659.400 256.050 660.600 260.400 ;
        RECT 664.950 260.400 673.050 261.600 ;
        RECT 664.950 259.950 667.050 260.400 ;
        RECT 670.950 260.100 673.050 260.400 ;
        RECT 680.400 259.950 685.050 261.600 ;
        RECT 688.950 261.600 693.000 262.050 ;
        RECT 688.950 259.950 693.600 261.600 ;
        RECT 634.950 255.600 637.050 255.900 ;
        RECT 620.400 254.400 637.050 255.600 ;
        RECT 634.950 253.800 637.050 254.400 ;
        RECT 646.950 253.800 649.050 255.900 ;
        RECT 658.950 253.950 661.050 256.050 ;
        RECT 680.400 255.900 681.600 259.950 ;
        RECT 692.400 255.900 693.600 259.950 ;
        RECT 679.950 253.800 682.050 255.900 ;
        RECT 691.950 253.800 694.050 255.900 ;
        RECT 701.400 253.050 702.600 262.950 ;
        RECT 703.950 259.950 706.050 262.050 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 721.950 261.600 724.050 262.200 ;
        RECT 733.950 261.600 736.050 262.200 ;
        RECT 721.950 260.400 736.050 261.600 ;
        RECT 721.950 260.100 724.050 260.400 ;
        RECT 733.950 260.100 736.050 260.400 ;
        RECT 739.950 261.600 742.050 262.200 ;
        RECT 757.950 261.600 760.050 262.200 ;
        RECT 739.950 260.400 760.050 261.600 ;
        RECT 739.950 260.100 742.050 260.400 ;
        RECT 757.950 260.100 760.050 260.400 ;
        RECT 763.950 260.100 766.050 262.200 ;
        RECT 781.950 260.100 784.050 262.200 ;
        RECT 704.400 256.050 705.600 259.950 ;
        RECT 710.400 256.050 711.600 259.950 ;
        RECT 764.400 258.600 765.600 260.100 ;
        RECT 782.400 258.600 783.600 260.100 ;
        RECT 811.950 259.950 814.050 262.050 ;
        RECT 832.950 259.950 835.050 262.050 ;
        RECT 838.950 261.600 841.050 262.050 ;
        RECT 844.950 261.600 847.050 262.200 ;
        RECT 838.950 260.400 847.050 261.600 ;
        RECT 838.950 259.950 841.050 260.400 ;
        RECT 844.950 260.100 847.050 260.400 ;
        RECT 850.950 260.100 853.050 262.200 ;
        RECT 764.400 257.400 783.600 258.600 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 709.950 253.950 712.050 256.050 ;
        RECT 718.950 255.450 721.050 255.900 ;
        RECT 727.950 255.450 730.050 256.050 ;
        RECT 718.950 254.250 730.050 255.450 ;
        RECT 718.950 253.800 721.050 254.250 ;
        RECT 727.950 253.950 730.050 254.250 ;
        RECT 742.950 255.450 745.050 255.900 ;
        RECT 751.950 255.450 754.050 255.900 ;
        RECT 742.950 254.250 754.050 255.450 ;
        RECT 742.950 253.800 745.050 254.250 ;
        RECT 751.950 253.800 754.050 254.250 ;
        RECT 775.950 253.950 778.050 257.400 ;
        RECT 812.400 256.050 813.600 259.950 ;
        RECT 833.400 256.050 834.600 259.950 ;
        RECT 793.950 255.450 796.050 255.900 ;
        RECT 799.950 255.450 802.050 255.900 ;
        RECT 793.950 254.250 802.050 255.450 ;
        RECT 793.950 253.800 796.050 254.250 ;
        RECT 799.950 253.800 802.050 254.250 ;
        RECT 811.950 253.950 814.050 256.050 ;
        RECT 832.950 253.950 835.050 256.050 ;
        RECT 851.400 255.600 852.600 260.100 ;
        RECT 880.950 259.950 883.050 262.050 ;
        RECT 892.950 261.600 895.050 262.200 ;
        RECT 887.400 260.400 895.050 261.600 ;
        RECT 881.400 256.050 882.600 259.950 ;
        RECT 856.800 255.600 858.900 256.050 ;
        RECT 851.400 254.400 858.900 255.600 ;
        RECT 856.800 253.950 858.900 254.400 ;
        RECT 859.950 255.450 862.050 255.900 ;
        RECT 871.950 255.450 874.050 255.900 ;
        RECT 859.950 254.250 874.050 255.450 ;
        RECT 859.950 253.800 862.050 254.250 ;
        RECT 871.950 253.800 874.050 254.250 ;
        RECT 880.950 253.950 883.050 256.050 ;
        RECT 253.950 252.600 256.050 253.050 ;
        RECT 242.400 251.400 256.050 252.600 ;
        RECT 64.950 250.800 67.050 251.250 ;
        RECT 94.950 250.800 97.050 251.250 ;
        RECT 253.950 250.950 256.050 251.400 ;
        RECT 490.950 252.600 493.050 253.050 ;
        RECT 499.950 252.600 502.050 253.050 ;
        RECT 490.950 251.400 502.050 252.600 ;
        RECT 490.950 250.950 493.050 251.400 ;
        RECT 499.950 250.950 502.050 251.400 ;
        RECT 613.950 250.950 616.050 253.050 ;
        RECT 649.950 252.600 652.050 253.050 ;
        RECT 673.950 252.600 676.050 253.050 ;
        RECT 649.950 251.400 676.050 252.600 ;
        RECT 649.950 250.950 652.050 251.400 ;
        RECT 673.950 250.950 676.050 251.400 ;
        RECT 700.950 250.950 703.050 253.050 ;
        RECT 736.950 252.600 739.050 253.050 ;
        RECT 769.950 252.600 772.050 253.050 ;
        RECT 736.950 251.400 772.050 252.600 ;
        RECT 736.950 250.950 739.050 251.400 ;
        RECT 769.950 250.950 772.050 251.400 ;
        RECT 778.950 252.600 781.050 253.050 ;
        RECT 794.400 252.600 795.600 253.800 ;
        RECT 778.950 251.400 795.600 252.600 ;
        RECT 847.950 252.600 850.050 253.050 ;
        RECT 860.400 252.600 861.600 253.800 ;
        RECT 847.950 251.400 861.600 252.600 ;
        RECT 778.950 250.950 781.050 251.400 ;
        RECT 847.950 250.950 850.050 251.400 ;
        RECT 79.950 249.600 82.050 250.050 ;
        RECT 97.950 249.600 100.050 250.050 ;
        RECT 79.950 248.400 100.050 249.600 ;
        RECT 79.950 247.950 82.050 248.400 ;
        RECT 97.950 247.950 100.050 248.400 ;
        RECT 136.950 249.600 139.050 250.050 ;
        RECT 157.950 249.600 160.050 250.050 ;
        RECT 136.950 248.400 160.050 249.600 ;
        RECT 136.950 247.950 139.050 248.400 ;
        RECT 157.950 247.950 160.050 248.400 ;
        RECT 193.950 249.600 196.050 250.050 ;
        RECT 217.950 249.600 220.050 250.050 ;
        RECT 226.950 249.600 229.050 250.050 ;
        RECT 235.950 249.600 238.050 250.050 ;
        RECT 193.950 248.400 238.050 249.600 ;
        RECT 193.950 247.950 196.050 248.400 ;
        RECT 217.950 247.950 220.050 248.400 ;
        RECT 226.950 247.950 229.050 248.400 ;
        RECT 235.950 247.950 238.050 248.400 ;
        RECT 400.950 249.600 403.050 250.050 ;
        RECT 424.950 249.600 427.050 250.050 ;
        RECT 400.950 248.400 427.050 249.600 ;
        RECT 400.950 247.950 403.050 248.400 ;
        RECT 424.950 247.950 427.050 248.400 ;
        RECT 511.950 249.600 514.050 250.050 ;
        RECT 538.950 249.600 541.050 250.050 ;
        RECT 511.950 248.400 541.050 249.600 ;
        RECT 511.950 247.950 514.050 248.400 ;
        RECT 538.950 247.950 541.050 248.400 ;
        RECT 853.950 249.600 856.050 249.900 ;
        RECT 877.950 249.600 880.050 250.050 ;
        RECT 887.400 249.600 888.600 260.400 ;
        RECT 892.950 260.100 895.050 260.400 ;
        RECT 910.950 261.750 913.050 262.200 ;
        RECT 916.950 261.750 919.050 262.200 ;
        RECT 910.950 260.550 919.050 261.750 ;
        RECT 910.950 260.100 913.050 260.550 ;
        RECT 916.950 260.100 919.050 260.550 ;
        RECT 922.950 261.600 925.050 262.200 ;
        RECT 928.950 261.600 931.050 262.050 ;
        RECT 922.950 260.400 931.050 261.600 ;
        RECT 922.950 260.100 925.050 260.400 ;
        RECT 928.950 259.950 931.050 260.400 ;
        RECT 901.950 255.450 904.050 255.900 ;
        RECT 925.950 255.450 928.050 255.900 ;
        RECT 901.950 254.250 928.050 255.450 ;
        RECT 901.950 253.800 904.050 254.250 ;
        RECT 925.950 253.800 928.050 254.250 ;
        RECT 853.950 248.400 880.050 249.600 ;
        RECT 98.400 246.600 99.600 247.950 ;
        RECT 106.950 246.600 109.050 247.050 ;
        RECT 98.400 245.400 109.050 246.600 ;
        RECT 106.950 244.950 109.050 245.400 ;
        RECT 112.950 246.600 115.050 247.050 ;
        RECT 163.950 246.600 166.050 247.050 ;
        RECT 112.950 245.400 166.050 246.600 ;
        RECT 236.400 246.600 237.600 247.950 ;
        RECT 853.950 247.800 856.050 248.400 ;
        RECT 877.950 247.950 880.050 248.400 ;
        RECT 884.400 248.400 888.600 249.600 ;
        RECT 889.950 249.600 892.050 250.050 ;
        RECT 928.950 249.600 931.050 250.050 ;
        RECT 889.950 248.400 931.050 249.600 ;
        RECT 307.950 246.600 310.050 247.050 ;
        RECT 236.400 245.400 310.050 246.600 ;
        RECT 112.950 244.950 115.050 245.400 ;
        RECT 163.950 244.950 166.050 245.400 ;
        RECT 307.950 244.950 310.050 245.400 ;
        RECT 445.950 246.600 448.050 247.050 ;
        RECT 463.950 246.600 466.050 247.050 ;
        RECT 445.950 245.400 466.050 246.600 ;
        RECT 445.950 244.950 448.050 245.400 ;
        RECT 463.950 244.950 466.050 245.400 ;
        RECT 604.950 246.600 607.050 247.050 ;
        RECT 652.950 246.600 655.050 247.050 ;
        RECT 745.950 246.600 748.050 247.050 ;
        RECT 604.950 245.400 748.050 246.600 ;
        RECT 604.950 244.950 607.050 245.400 ;
        RECT 652.950 244.950 655.050 245.400 ;
        RECT 745.950 244.950 748.050 245.400 ;
        RECT 877.950 246.600 880.050 246.900 ;
        RECT 884.400 246.600 885.600 248.400 ;
        RECT 889.950 247.950 892.050 248.400 ;
        RECT 928.950 247.950 931.050 248.400 ;
        RECT 877.950 245.400 885.600 246.600 ;
        RECT 877.950 244.800 880.050 245.400 ;
        RECT 133.950 243.600 136.050 244.050 ;
        RECT 301.950 243.600 304.050 244.050 ;
        RECT 133.950 242.400 304.050 243.600 ;
        RECT 133.950 241.950 136.050 242.400 ;
        RECT 301.950 241.950 304.050 242.400 ;
        RECT 319.950 243.600 322.050 244.050 ;
        RECT 346.950 243.600 349.050 244.050 ;
        RECT 319.950 242.400 349.050 243.600 ;
        RECT 319.950 241.950 322.050 242.400 ;
        RECT 346.950 241.950 349.050 242.400 ;
        RECT 418.950 243.600 421.050 244.050 ;
        RECT 442.950 243.600 445.050 244.050 ;
        RECT 496.950 243.600 499.050 244.050 ;
        RECT 418.950 242.400 499.050 243.600 ;
        RECT 418.950 241.950 421.050 242.400 ;
        RECT 442.950 241.950 445.050 242.400 ;
        RECT 496.950 241.950 499.050 242.400 ;
        RECT 592.950 243.600 595.050 244.050 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 592.950 242.400 652.050 243.600 ;
        RECT 592.950 241.950 595.050 242.400 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 775.950 243.600 778.050 244.050 ;
        RECT 838.950 243.600 841.050 244.050 ;
        RECT 775.950 242.400 841.050 243.600 ;
        RECT 775.950 241.950 778.050 242.400 ;
        RECT 838.950 241.950 841.050 242.400 ;
        RECT 895.950 243.600 898.050 244.050 ;
        RECT 934.950 243.600 937.050 244.050 ;
        RECT 895.950 242.400 937.050 243.600 ;
        RECT 895.950 241.950 898.050 242.400 ;
        RECT 934.950 241.950 937.050 242.400 ;
        RECT 76.950 240.600 79.050 241.050 ;
        RECT 97.950 240.600 100.050 241.050 ;
        RECT 76.950 239.400 100.050 240.600 ;
        RECT 76.950 238.950 79.050 239.400 ;
        RECT 97.950 238.950 100.050 239.400 ;
        RECT 448.950 240.600 451.050 241.050 ;
        RECT 562.950 240.600 565.050 241.050 ;
        RECT 448.950 239.400 565.050 240.600 ;
        RECT 448.950 238.950 451.050 239.400 ;
        RECT 562.950 238.950 565.050 239.400 ;
        RECT 589.950 240.600 592.050 241.050 ;
        RECT 610.950 240.600 613.050 241.050 ;
        RECT 589.950 239.400 613.050 240.600 ;
        RECT 589.950 238.950 592.050 239.400 ;
        RECT 610.950 238.950 613.050 239.400 ;
        RECT 805.950 240.600 808.050 241.050 ;
        RECT 826.950 240.600 829.050 241.050 ;
        RECT 850.950 240.600 853.050 241.050 ;
        RECT 805.950 239.400 853.050 240.600 ;
        RECT 805.950 238.950 808.050 239.400 ;
        RECT 826.950 238.950 829.050 239.400 ;
        RECT 850.950 238.950 853.050 239.400 ;
        RECT 160.950 237.600 163.050 238.050 ;
        RECT 277.950 237.600 280.050 238.050 ;
        RECT 160.950 236.400 280.050 237.600 ;
        RECT 160.950 235.950 163.050 236.400 ;
        RECT 277.950 235.950 280.050 236.400 ;
        RECT 283.950 237.600 286.050 238.050 ;
        RECT 319.950 237.600 322.050 238.050 ;
        RECT 283.950 236.400 322.050 237.600 ;
        RECT 283.950 235.950 286.050 236.400 ;
        RECT 319.950 235.950 322.050 236.400 ;
        RECT 559.950 237.600 562.050 238.050 ;
        RECT 616.950 237.600 619.050 238.050 ;
        RECT 628.950 237.600 631.050 238.050 ;
        RECT 559.950 236.400 631.050 237.600 ;
        RECT 559.950 235.950 562.050 236.400 ;
        RECT 616.950 235.950 619.050 236.400 ;
        RECT 628.950 235.950 631.050 236.400 ;
        RECT 643.950 237.600 646.050 238.050 ;
        RECT 733.950 237.600 736.050 238.050 ;
        RECT 643.950 236.400 736.050 237.600 ;
        RECT 643.950 235.950 646.050 236.400 ;
        RECT 733.950 235.950 736.050 236.400 ;
        RECT 784.950 237.600 787.050 238.050 ;
        RECT 799.950 237.600 802.050 238.050 ;
        RECT 889.950 237.600 892.050 238.050 ;
        RECT 784.950 236.400 892.050 237.600 ;
        RECT 784.950 235.950 787.050 236.400 ;
        RECT 799.950 235.950 802.050 236.400 ;
        RECT 889.950 235.950 892.050 236.400 ;
        RECT 88.950 234.600 91.050 235.050 ;
        RECT 115.950 234.600 118.050 235.050 ;
        RECT 88.950 233.400 118.050 234.600 ;
        RECT 88.950 232.950 91.050 233.400 ;
        RECT 115.950 232.950 118.050 233.400 ;
        RECT 421.950 234.600 424.050 235.050 ;
        RECT 520.950 234.600 523.050 235.050 ;
        RECT 421.950 233.400 523.050 234.600 ;
        RECT 421.950 232.950 424.050 233.400 ;
        RECT 520.950 232.950 523.050 233.400 ;
        RECT 562.950 234.600 565.050 235.050 ;
        RECT 619.950 234.600 622.050 235.050 ;
        RECT 562.950 233.400 622.050 234.600 ;
        RECT 562.950 232.950 565.050 233.400 ;
        RECT 619.950 232.950 622.050 233.400 ;
        RECT 679.950 234.600 682.050 235.050 ;
        RECT 739.950 234.600 742.050 235.050 ;
        RECT 679.950 233.400 742.050 234.600 ;
        RECT 679.950 232.950 682.050 233.400 ;
        RECT 739.950 232.950 742.050 233.400 ;
        RECT 814.950 234.600 817.050 235.050 ;
        RECT 841.950 234.600 844.050 235.050 ;
        RECT 814.950 233.400 844.050 234.600 ;
        RECT 814.950 232.950 817.050 233.400 ;
        RECT 841.950 232.950 844.050 233.400 ;
        RECT 859.950 234.600 862.050 235.050 ;
        RECT 898.950 234.600 901.050 235.050 ;
        RECT 859.950 233.400 901.050 234.600 ;
        RECT 859.950 232.950 862.050 233.400 ;
        RECT 898.950 232.950 901.050 233.400 ;
        RECT 82.950 231.600 85.050 232.050 ;
        RECT 121.950 231.600 124.050 232.050 ;
        RECT 82.950 230.400 124.050 231.600 ;
        RECT 82.950 229.950 85.050 230.400 ;
        RECT 121.950 229.950 124.050 230.400 ;
        RECT 148.950 231.600 151.050 232.050 ;
        RECT 208.950 231.600 211.050 232.050 ;
        RECT 148.950 230.400 211.050 231.600 ;
        RECT 148.950 229.950 151.050 230.400 ;
        RECT 208.950 229.950 211.050 230.400 ;
        RECT 256.950 231.600 259.050 232.050 ;
        RECT 289.950 231.600 292.050 232.050 ;
        RECT 256.950 230.400 292.050 231.600 ;
        RECT 256.950 229.950 259.050 230.400 ;
        RECT 289.950 229.950 292.050 230.400 ;
        RECT 340.950 231.600 343.050 232.050 ;
        RECT 379.950 231.600 382.050 232.050 ;
        RECT 418.950 231.600 421.050 232.050 ;
        RECT 748.950 231.600 751.050 232.050 ;
        RECT 340.950 230.400 751.050 231.600 ;
        RECT 340.950 229.950 343.050 230.400 ;
        RECT 379.950 229.950 382.050 230.400 ;
        RECT 418.950 229.950 421.050 230.400 ;
        RECT 748.950 229.950 751.050 230.400 ;
        RECT 907.950 231.600 910.050 232.050 ;
        RECT 928.950 231.600 931.050 232.050 ;
        RECT 907.950 230.400 931.050 231.600 ;
        RECT 907.950 229.950 910.050 230.400 ;
        RECT 928.950 229.950 931.050 230.400 ;
        RECT 424.950 228.600 427.050 229.050 ;
        RECT 469.950 228.600 472.050 229.050 ;
        RECT 424.950 227.400 472.050 228.600 ;
        RECT 424.950 226.950 427.050 227.400 ;
        RECT 469.950 226.950 472.050 227.400 ;
        RECT 547.950 228.600 550.050 229.050 ;
        RECT 568.950 228.600 571.050 229.050 ;
        RECT 547.950 227.400 571.050 228.600 ;
        RECT 547.950 226.950 550.050 227.400 ;
        RECT 568.950 226.950 571.050 227.400 ;
        RECT 640.950 228.600 643.050 229.050 ;
        RECT 646.950 228.600 649.050 229.050 ;
        RECT 640.950 227.400 649.050 228.600 ;
        RECT 640.950 226.950 643.050 227.400 ;
        RECT 646.950 226.950 649.050 227.400 ;
        RECT 862.950 228.600 865.050 229.050 ;
        RECT 892.950 228.600 895.050 229.050 ;
        RECT 862.950 227.400 895.050 228.600 ;
        RECT 862.950 226.950 865.050 227.400 ;
        RECT 892.950 226.950 895.050 227.400 ;
        RECT 913.950 228.600 916.050 229.050 ;
        RECT 922.950 228.600 925.050 229.050 ;
        RECT 913.950 227.400 925.050 228.600 ;
        RECT 913.950 226.950 916.050 227.400 ;
        RECT 922.950 226.950 925.050 227.400 ;
        RECT 202.950 225.600 205.050 226.050 ;
        RECT 214.950 225.600 217.050 226.050 ;
        RECT 202.950 224.400 217.050 225.600 ;
        RECT 202.950 223.950 205.050 224.400 ;
        RECT 214.950 223.950 217.050 224.400 ;
        RECT 229.950 225.600 232.050 226.050 ;
        RECT 241.950 225.600 244.050 226.050 ;
        RECT 229.950 224.400 244.050 225.600 ;
        RECT 229.950 223.950 232.050 224.400 ;
        RECT 241.950 223.950 244.050 224.400 ;
        RECT 439.950 225.600 442.050 226.050 ;
        RECT 454.950 225.600 457.050 226.050 ;
        RECT 439.950 224.400 457.050 225.600 ;
        RECT 439.950 223.950 442.050 224.400 ;
        RECT 454.950 223.950 457.050 224.400 ;
        RECT 481.950 225.600 484.050 226.050 ;
        RECT 490.950 225.600 493.050 226.050 ;
        RECT 481.950 224.400 493.050 225.600 ;
        RECT 481.950 223.950 484.050 224.400 ;
        RECT 490.950 223.950 493.050 224.400 ;
        RECT 604.950 225.600 607.050 226.050 ;
        RECT 667.950 225.600 670.050 226.050 ;
        RECT 604.950 224.400 670.050 225.600 ;
        RECT 604.950 223.950 607.050 224.400 ;
        RECT 667.950 223.950 670.050 224.400 ;
        RECT 679.950 225.600 682.050 226.050 ;
        RECT 685.950 225.600 688.050 226.050 ;
        RECT 679.950 224.400 688.050 225.600 ;
        RECT 679.950 223.950 682.050 224.400 ;
        RECT 685.950 223.950 688.050 224.400 ;
        RECT 766.950 225.600 769.050 226.050 ;
        RECT 823.950 225.600 826.050 226.050 ;
        RECT 847.950 225.600 850.050 226.050 ;
        RECT 766.950 224.400 850.050 225.600 ;
        RECT 766.950 223.950 769.050 224.400 ;
        RECT 823.950 223.950 826.050 224.400 ;
        RECT 847.950 223.950 850.050 224.400 ;
        RECT 94.950 222.600 97.050 223.050 ;
        RECT 151.950 222.600 154.050 223.050 ;
        RECT 94.950 221.400 154.050 222.600 ;
        RECT 94.950 220.950 97.050 221.400 ;
        RECT 151.950 220.950 154.050 221.400 ;
        RECT 184.950 222.600 187.050 223.050 ;
        RECT 199.950 222.600 202.050 223.050 ;
        RECT 184.950 221.400 202.050 222.600 ;
        RECT 184.950 220.950 187.050 221.400 ;
        RECT 199.950 220.950 202.050 221.400 ;
        RECT 247.950 222.600 250.050 223.050 ;
        RECT 265.950 222.600 268.050 223.050 ;
        RECT 247.950 221.400 268.050 222.600 ;
        RECT 247.950 220.950 250.050 221.400 ;
        RECT 265.950 220.950 268.050 221.400 ;
        RECT 271.950 222.600 274.050 223.050 ;
        RECT 280.950 222.600 283.050 223.050 ;
        RECT 271.950 221.400 283.050 222.600 ;
        RECT 271.950 220.950 274.050 221.400 ;
        RECT 280.950 220.950 283.050 221.400 ;
        RECT 298.950 222.600 301.050 223.050 ;
        RECT 313.950 222.600 316.050 223.050 ;
        RECT 298.950 221.400 316.050 222.600 ;
        RECT 298.950 220.950 301.050 221.400 ;
        RECT 313.950 220.950 316.050 221.400 ;
        RECT 334.950 222.600 337.050 223.050 ;
        RECT 421.950 222.600 424.050 223.050 ;
        RECT 334.950 221.400 424.050 222.600 ;
        RECT 334.950 220.950 337.050 221.400 ;
        RECT 421.950 220.950 424.050 221.400 ;
        RECT 430.950 222.600 433.050 223.050 ;
        RECT 478.950 222.600 481.050 223.050 ;
        RECT 502.950 222.600 505.050 223.050 ;
        RECT 430.950 221.400 505.050 222.600 ;
        RECT 430.950 220.950 433.050 221.400 ;
        RECT 478.950 220.950 481.050 221.400 ;
        RECT 502.950 220.950 505.050 221.400 ;
        RECT 571.950 222.600 574.050 223.050 ;
        RECT 577.950 222.600 580.050 223.050 ;
        RECT 592.950 222.600 595.050 223.050 ;
        RECT 571.950 221.400 595.050 222.600 ;
        RECT 668.400 222.600 669.600 223.950 ;
        RECT 676.950 222.600 679.050 223.050 ;
        RECT 668.400 221.400 679.050 222.600 ;
        RECT 571.950 220.950 574.050 221.400 ;
        RECT 577.950 220.950 580.050 221.400 ;
        RECT 592.950 220.950 595.050 221.400 ;
        RECT 676.950 220.950 679.050 221.400 ;
        RECT 703.950 222.600 706.050 223.050 ;
        RECT 787.950 222.600 790.050 223.050 ;
        RECT 703.950 221.400 790.050 222.600 ;
        RECT 703.950 220.950 706.050 221.400 ;
        RECT 787.950 220.950 790.050 221.400 ;
        RECT 856.950 222.600 859.050 223.050 ;
        RECT 886.950 222.600 889.050 223.050 ;
        RECT 856.950 221.400 889.050 222.600 ;
        RECT 856.950 220.950 859.050 221.400 ;
        RECT 886.950 220.950 889.050 221.400 ;
        RECT 19.950 219.600 22.050 220.050 ;
        RECT 40.950 219.600 43.050 220.050 ;
        RECT 97.950 219.600 100.050 220.050 ;
        RECT 19.950 218.400 43.050 219.600 ;
        RECT 19.950 217.950 22.050 218.400 ;
        RECT 40.950 217.950 43.050 218.400 ;
        RECT 44.400 218.400 100.050 219.600 ;
        RECT 44.400 216.600 45.600 218.400 ;
        RECT 97.950 217.950 100.050 218.400 ;
        RECT 286.950 219.600 289.050 220.050 ;
        RECT 292.950 219.600 295.050 220.050 ;
        RECT 286.950 218.400 295.050 219.600 ;
        RECT 286.950 217.950 289.050 218.400 ;
        RECT 292.950 217.950 295.050 218.400 ;
        RECT 304.950 219.600 307.050 220.050 ;
        RECT 316.950 219.600 319.050 220.050 ;
        RECT 304.950 218.400 319.050 219.600 ;
        RECT 304.950 217.950 307.050 218.400 ;
        RECT 316.950 217.950 319.050 218.400 ;
        RECT 550.950 219.600 553.050 220.050 ;
        RECT 604.950 219.600 607.050 220.050 ;
        RECT 550.950 218.400 607.050 219.600 ;
        RECT 550.950 217.950 553.050 218.400 ;
        RECT 17.400 215.400 45.600 216.600 ;
        RECT 88.950 216.600 91.050 217.050 ;
        RECT 232.950 216.750 235.050 217.200 ;
        RECT 241.950 216.750 244.050 217.200 ;
        RECT 88.950 216.000 96.600 216.600 ;
        RECT 88.950 215.400 97.050 216.000 ;
        RECT 13.950 213.600 16.050 213.900 ;
        RECT 17.400 213.600 18.600 215.400 ;
        RECT 88.950 214.950 91.050 215.400 ;
        RECT 13.950 212.400 18.600 213.600 ;
        RECT 43.950 213.600 46.050 214.050 ;
        RECT 43.950 212.400 54.600 213.600 ;
        RECT 13.950 211.800 16.050 212.400 ;
        RECT 43.950 211.950 46.050 212.400 ;
        RECT 53.400 210.600 54.600 212.400 ;
        RECT 94.950 211.950 97.050 215.400 ;
        RECT 232.950 215.550 244.050 216.750 ;
        RECT 232.950 215.100 235.050 215.550 ;
        RECT 241.950 215.100 244.050 215.550 ;
        RECT 277.950 216.600 280.050 217.050 ;
        RECT 346.950 216.600 349.050 217.050 ;
        RECT 277.950 215.400 349.050 216.600 ;
        RECT 242.400 211.050 243.600 215.100 ;
        RECT 277.950 214.950 280.050 215.400 ;
        RECT 346.950 214.950 349.050 215.400 ;
        RECT 361.950 216.600 364.050 217.200 ;
        RECT 379.950 216.600 382.050 217.200 ;
        RECT 361.950 215.400 382.050 216.600 ;
        RECT 361.950 215.100 364.050 215.400 ;
        RECT 379.950 215.100 382.050 215.400 ;
        RECT 397.950 215.100 400.050 217.200 ;
        RECT 403.950 216.750 406.050 217.200 ;
        RECT 409.950 216.750 412.050 217.200 ;
        RECT 403.950 215.550 412.050 216.750 ;
        RECT 403.950 215.100 406.050 215.550 ;
        RECT 409.950 215.100 412.050 215.550 ;
        RECT 445.950 216.750 448.050 217.200 ;
        RECT 451.950 216.750 454.050 217.200 ;
        RECT 445.950 215.550 454.050 216.750 ;
        RECT 445.950 215.100 448.050 215.550 ;
        RECT 451.950 215.100 454.050 215.550 ;
        RECT 61.950 210.600 64.050 211.050 ;
        RECT 73.950 210.600 76.050 211.050 ;
        RECT 53.400 209.400 57.600 210.600 ;
        RECT 56.400 208.050 57.600 209.400 ;
        RECT 61.950 209.400 76.050 210.600 ;
        RECT 61.950 208.950 64.050 209.400 ;
        RECT 73.950 208.950 76.050 209.400 ;
        RECT 85.950 210.600 88.050 210.900 ;
        RECT 91.950 210.600 94.050 211.050 ;
        RECT 85.950 209.400 94.050 210.600 ;
        RECT 85.950 208.800 88.050 209.400 ;
        RECT 91.950 208.950 94.050 209.400 ;
        RECT 241.950 208.950 244.050 211.050 ;
        RECT 280.950 210.450 283.050 210.900 ;
        RECT 289.950 210.450 292.050 210.900 ;
        RECT 280.950 209.250 292.050 210.450 ;
        RECT 280.950 208.800 283.050 209.250 ;
        RECT 289.950 208.800 292.050 209.250 ;
        RECT 301.950 210.600 304.050 211.050 ;
        RECT 313.950 210.600 316.050 210.900 ;
        RECT 301.950 209.400 316.050 210.600 ;
        RECT 301.950 208.950 304.050 209.400 ;
        RECT 313.950 208.800 316.050 209.400 ;
        RECT 325.950 210.450 328.050 210.900 ;
        RECT 337.950 210.450 340.050 210.900 ;
        RECT 325.950 209.250 340.050 210.450 ;
        RECT 325.950 208.800 328.050 209.250 ;
        RECT 337.950 208.800 340.050 209.250 ;
        RECT 346.950 210.600 349.050 211.050 ;
        RECT 358.950 210.600 361.050 210.900 ;
        RECT 346.950 209.400 361.050 210.600 ;
        RECT 346.950 208.950 349.050 209.400 ;
        RECT 358.950 208.800 361.050 209.400 ;
        RECT 391.950 210.600 394.050 211.050 ;
        RECT 398.400 210.600 399.600 215.100 ;
        RECT 463.950 213.600 466.050 217.050 ;
        RECT 472.950 216.750 475.050 217.200 ;
        RECT 484.950 216.750 487.050 217.200 ;
        RECT 472.950 215.550 487.050 216.750 ;
        RECT 472.950 215.100 475.050 215.550 ;
        RECT 484.950 215.100 487.050 215.550 ;
        RECT 496.950 216.600 499.050 217.050 ;
        RECT 541.950 216.750 544.050 217.200 ;
        RECT 550.950 216.750 553.050 216.900 ;
        RECT 496.950 215.400 507.600 216.600 ;
        RECT 496.950 214.950 499.050 215.400 ;
        RECT 506.400 213.600 507.600 215.400 ;
        RECT 541.950 215.550 553.050 216.750 ;
        RECT 541.950 215.100 544.050 215.550 ;
        RECT 550.950 214.800 553.050 215.550 ;
        RECT 556.950 216.750 559.050 217.200 ;
        RECT 565.950 216.750 568.050 217.200 ;
        RECT 556.950 215.550 568.050 216.750 ;
        RECT 556.950 215.100 559.050 215.550 ;
        RECT 565.950 215.100 568.050 215.550 ;
        RECT 583.950 216.600 586.050 217.200 ;
        RECT 583.950 215.400 591.600 216.600 ;
        RECT 583.950 215.100 586.050 215.400 ;
        RECT 463.950 213.000 504.600 213.600 ;
        RECT 464.400 212.400 504.600 213.000 ;
        RECT 506.400 212.400 522.600 213.600 ;
        RECT 391.950 209.400 399.600 210.600 ;
        RECT 409.950 210.600 412.050 211.050 ;
        RECT 415.950 210.600 418.050 210.900 ;
        RECT 409.950 209.400 418.050 210.600 ;
        RECT 391.950 208.950 394.050 209.400 ;
        RECT 409.950 208.950 412.050 209.400 ;
        RECT 415.950 208.800 418.050 209.400 ;
        RECT 430.950 210.450 433.050 210.900 ;
        RECT 436.950 210.450 439.050 210.900 ;
        RECT 430.950 209.250 439.050 210.450 ;
        RECT 430.950 208.800 433.050 209.250 ;
        RECT 436.950 208.800 439.050 209.250 ;
        RECT 451.950 210.450 454.050 210.900 ;
        RECT 460.950 210.600 463.050 210.900 ;
        RECT 475.950 210.600 478.050 210.900 ;
        RECT 460.950 210.450 478.050 210.600 ;
        RECT 451.950 209.400 478.050 210.450 ;
        RECT 451.950 209.250 463.050 209.400 ;
        RECT 451.950 208.800 454.050 209.250 ;
        RECT 460.950 208.800 463.050 209.250 ;
        RECT 475.950 208.800 478.050 209.400 ;
        RECT 490.950 210.450 493.050 210.900 ;
        RECT 499.950 210.450 502.050 210.900 ;
        RECT 490.950 209.250 502.050 210.450 ;
        RECT 503.400 210.600 504.600 212.400 ;
        RECT 517.950 210.600 520.050 210.900 ;
        RECT 503.400 209.400 520.050 210.600 ;
        RECT 521.400 210.600 522.600 212.400 ;
        RECT 538.950 210.600 541.050 210.900 ;
        RECT 521.400 209.400 541.050 210.600 ;
        RECT 490.950 208.800 493.050 209.250 ;
        RECT 499.950 208.800 502.050 209.250 ;
        RECT 517.950 208.800 520.050 209.400 ;
        RECT 538.950 208.800 541.050 209.400 ;
        RECT 56.400 206.400 61.050 208.050 ;
        RECT 57.000 205.950 61.050 206.400 ;
        RECT 142.950 207.600 145.050 208.050 ;
        RECT 169.950 207.600 172.050 208.050 ;
        RECT 142.950 206.400 172.050 207.600 ;
        RECT 142.950 205.950 145.050 206.400 ;
        RECT 169.950 205.950 172.050 206.400 ;
        RECT 235.950 207.600 238.050 208.050 ;
        RECT 274.950 207.600 277.050 208.050 ;
        RECT 235.950 206.400 277.050 207.600 ;
        RECT 235.950 205.950 238.050 206.400 ;
        RECT 274.950 205.950 277.050 206.400 ;
        RECT 364.950 207.600 367.050 208.050 ;
        RECT 394.950 207.600 397.050 208.050 ;
        RECT 364.950 206.400 397.050 207.600 ;
        RECT 364.950 205.950 367.050 206.400 ;
        RECT 394.950 205.950 397.050 206.400 ;
        RECT 421.950 207.600 424.050 208.050 ;
        RECT 439.950 207.600 442.050 208.050 ;
        RECT 421.950 206.400 442.050 207.600 ;
        RECT 421.950 205.950 424.050 206.400 ;
        RECT 439.950 205.950 442.050 206.400 ;
        RECT 526.950 207.600 529.050 208.050 ;
        RECT 559.950 207.600 562.050 208.050 ;
        RECT 526.950 206.400 562.050 207.600 ;
        RECT 590.400 207.600 591.600 215.400 ;
        RECT 593.400 210.600 594.600 218.400 ;
        RECT 604.950 217.950 607.050 218.400 ;
        RECT 652.950 219.600 655.050 220.050 ;
        RECT 661.950 219.600 664.050 220.050 ;
        RECT 652.950 218.400 664.050 219.600 ;
        RECT 652.950 217.950 655.050 218.400 ;
        RECT 661.950 217.950 664.050 218.400 ;
        RECT 838.950 219.600 841.050 220.050 ;
        RECT 838.950 218.400 846.600 219.600 ;
        RECT 838.950 217.950 841.050 218.400 ;
        RECT 646.950 216.600 649.050 217.200 ;
        RECT 697.950 216.600 700.050 217.200 ;
        RECT 724.950 216.600 727.050 217.200 ;
        RECT 646.950 215.400 727.050 216.600 ;
        RECT 646.950 215.100 649.050 215.400 ;
        RECT 697.950 215.100 700.050 215.400 ;
        RECT 724.950 215.100 727.050 215.400 ;
        RECT 745.950 216.600 748.050 217.200 ;
        RECT 760.950 216.600 763.050 217.200 ;
        RECT 745.950 215.400 763.050 216.600 ;
        RECT 745.950 215.100 748.050 215.400 ;
        RECT 760.950 215.100 763.050 215.400 ;
        RECT 766.950 216.600 769.050 217.200 ;
        RECT 775.950 216.750 778.050 217.200 ;
        RECT 781.950 216.750 784.050 217.200 ;
        RECT 775.950 216.600 784.050 216.750 ;
        RECT 766.950 215.550 784.050 216.600 ;
        RECT 766.950 215.400 778.050 215.550 ;
        RECT 766.950 215.100 769.050 215.400 ;
        RECT 775.950 215.100 778.050 215.400 ;
        RECT 781.950 215.100 784.050 215.550 ;
        RECT 845.400 210.900 846.600 218.400 ;
        RECT 883.950 217.950 886.050 220.050 ;
        RECT 889.950 217.950 892.050 220.050 ;
        RECT 850.950 214.950 853.050 217.050 ;
        RECT 859.950 216.600 862.050 217.050 ;
        RECT 880.950 216.600 883.050 217.050 ;
        RECT 859.950 215.400 870.600 216.600 ;
        RECT 859.950 214.950 862.050 215.400 ;
        RECT 598.950 210.600 601.050 210.900 ;
        RECT 593.400 209.400 601.050 210.600 ;
        RECT 598.950 208.800 601.050 209.400 ;
        RECT 604.950 210.450 607.050 210.900 ;
        RECT 613.950 210.450 616.050 210.900 ;
        RECT 604.950 209.250 616.050 210.450 ;
        RECT 604.950 208.800 607.050 209.250 ;
        RECT 613.950 208.800 616.050 209.250 ;
        RECT 643.950 210.450 646.050 210.900 ;
        RECT 652.950 210.600 655.050 210.900 ;
        RECT 682.950 210.600 685.050 210.900 ;
        RECT 709.950 210.600 712.050 210.900 ;
        RECT 652.950 210.450 712.050 210.600 ;
        RECT 643.950 209.400 712.050 210.450 ;
        RECT 643.950 209.250 655.050 209.400 ;
        RECT 643.950 208.800 646.050 209.250 ;
        RECT 652.950 208.800 655.050 209.250 ;
        RECT 682.950 208.800 685.050 209.400 ;
        RECT 709.950 208.800 712.050 209.400 ;
        RECT 733.950 210.450 736.050 210.900 ;
        RECT 742.950 210.450 745.050 210.900 ;
        RECT 733.950 209.250 745.050 210.450 ;
        RECT 733.950 208.800 736.050 209.250 ;
        RECT 742.950 208.800 745.050 209.250 ;
        RECT 844.950 208.800 847.050 210.900 ;
        RECT 851.400 210.600 852.600 214.950 ;
        RECT 869.400 210.900 870.600 215.400 ;
        RECT 875.400 215.400 883.050 216.600 ;
        RECT 875.400 211.050 876.600 215.400 ;
        RECT 880.950 214.950 883.050 215.400 ;
        RECT 884.400 213.600 885.600 217.950 ;
        RECT 881.400 213.000 885.600 213.600 ;
        RECT 880.950 212.400 885.600 213.000 ;
        RECT 862.950 210.600 865.050 210.900 ;
        RECT 851.400 209.400 865.050 210.600 ;
        RECT 862.950 208.800 865.050 209.400 ;
        RECT 868.950 208.800 871.050 210.900 ;
        RECT 874.950 208.950 877.050 211.050 ;
        RECT 880.950 208.950 883.050 212.400 ;
        RECT 595.950 207.600 598.050 208.050 ;
        RECT 590.400 206.400 598.050 207.600 ;
        RECT 526.950 205.950 529.050 206.400 ;
        RECT 559.950 205.950 562.050 206.400 ;
        RECT 595.950 205.950 598.050 206.400 ;
        RECT 763.950 207.600 766.050 208.050 ;
        RECT 778.950 207.600 781.050 208.050 ;
        RECT 763.950 206.400 781.050 207.600 ;
        RECT 763.950 205.950 766.050 206.400 ;
        RECT 778.950 205.950 781.050 206.400 ;
        RECT 793.950 207.600 796.050 208.050 ;
        RECT 808.950 207.600 811.050 208.050 ;
        RECT 820.950 207.600 823.050 208.050 ;
        RECT 793.950 206.400 823.050 207.600 ;
        RECT 793.950 205.950 796.050 206.400 ;
        RECT 808.950 205.950 811.050 206.400 ;
        RECT 820.950 205.950 823.050 206.400 ;
        RECT 883.950 207.600 886.050 208.050 ;
        RECT 890.400 207.600 891.600 217.950 ;
        RECT 892.950 216.600 895.050 217.050 ;
        RECT 898.950 216.600 901.050 217.050 ;
        RECT 892.950 215.400 901.050 216.600 ;
        RECT 892.950 214.950 895.050 215.400 ;
        RECT 898.950 214.950 901.050 215.400 ;
        RECT 904.950 215.100 907.050 217.200 ;
        RECT 910.950 216.750 913.050 217.200 ;
        RECT 919.950 216.750 922.050 217.200 ;
        RECT 910.950 215.550 922.050 216.750 ;
        RECT 910.950 215.100 913.050 215.550 ;
        RECT 919.950 215.100 922.050 215.550 ;
        RECT 895.950 210.600 898.050 211.050 ;
        RECT 905.400 210.600 906.600 215.100 ;
        RECT 895.950 209.400 906.600 210.600 ;
        RECT 907.950 210.450 910.050 210.900 ;
        RECT 928.950 210.450 931.050 210.900 ;
        RECT 895.950 208.950 898.050 209.400 ;
        RECT 907.950 209.250 931.050 210.450 ;
        RECT 907.950 208.800 910.050 209.250 ;
        RECT 928.950 208.800 931.050 209.250 ;
        RECT 883.950 206.400 891.600 207.600 ;
        RECT 910.950 207.600 913.050 208.050 ;
        RECT 922.950 207.600 925.050 208.050 ;
        RECT 910.950 206.400 925.050 207.600 ;
        RECT 883.950 205.950 886.050 206.400 ;
        RECT 910.950 205.950 913.050 206.400 ;
        RECT 922.950 205.950 925.050 206.400 ;
        RECT 10.950 204.600 13.050 205.050 ;
        RECT 16.950 204.600 19.050 205.050 ;
        RECT 10.950 203.400 19.050 204.600 ;
        RECT 10.950 202.950 13.050 203.400 ;
        RECT 16.950 202.950 19.050 203.400 ;
        RECT 304.950 204.600 307.050 205.050 ;
        RECT 313.950 204.600 316.050 205.050 ;
        RECT 304.950 203.400 316.050 204.600 ;
        RECT 304.950 202.950 307.050 203.400 ;
        RECT 313.950 202.950 316.050 203.400 ;
        RECT 466.950 204.600 469.050 205.050 ;
        RECT 481.950 204.600 484.050 205.050 ;
        RECT 505.950 204.600 508.050 205.050 ;
        RECT 466.950 203.400 508.050 204.600 ;
        RECT 466.950 202.950 469.050 203.400 ;
        RECT 481.950 202.950 484.050 203.400 ;
        RECT 505.950 202.950 508.050 203.400 ;
        RECT 523.950 204.600 526.050 205.050 ;
        RECT 544.950 204.600 547.050 205.050 ;
        RECT 580.950 204.600 583.050 205.050 ;
        RECT 658.950 204.600 661.050 205.050 ;
        RECT 523.950 203.400 583.050 204.600 ;
        RECT 523.950 202.950 526.050 203.400 ;
        RECT 544.950 202.950 547.050 203.400 ;
        RECT 580.950 202.950 583.050 203.400 ;
        RECT 584.400 203.400 661.050 204.600 ;
        RECT 4.950 201.600 7.050 202.050 ;
        RECT 10.950 201.600 13.050 201.900 ;
        RECT 4.950 200.400 13.050 201.600 ;
        RECT 4.950 199.950 7.050 200.400 ;
        RECT 10.950 199.800 13.050 200.400 ;
        RECT 208.950 201.600 211.050 202.050 ;
        RECT 217.950 201.600 220.050 202.050 ;
        RECT 208.950 200.400 220.050 201.600 ;
        RECT 208.950 199.950 211.050 200.400 ;
        RECT 217.950 199.950 220.050 200.400 ;
        RECT 247.950 201.600 250.050 202.050 ;
        RECT 283.950 201.600 286.050 202.050 ;
        RECT 247.950 200.400 286.050 201.600 ;
        RECT 247.950 199.950 250.050 200.400 ;
        RECT 283.950 199.950 286.050 200.400 ;
        RECT 337.950 201.600 340.050 202.050 ;
        RECT 364.950 201.600 367.050 202.050 ;
        RECT 337.950 200.400 367.050 201.600 ;
        RECT 337.950 199.950 340.050 200.400 ;
        RECT 364.950 199.950 367.050 200.400 ;
        RECT 376.950 201.600 379.050 202.050 ;
        RECT 406.950 201.600 409.050 202.050 ;
        RECT 376.950 200.400 409.050 201.600 ;
        RECT 376.950 199.950 379.050 200.400 ;
        RECT 406.950 199.950 409.050 200.400 ;
        RECT 505.950 201.600 508.050 201.900 ;
        RECT 517.950 201.600 520.050 202.050 ;
        RECT 505.950 200.400 520.050 201.600 ;
        RECT 505.950 199.800 508.050 200.400 ;
        RECT 517.950 199.950 520.050 200.400 ;
        RECT 550.950 201.600 553.050 202.050 ;
        RECT 584.400 201.600 585.600 203.400 ;
        RECT 658.950 202.950 661.050 203.400 ;
        RECT 748.950 204.600 751.050 205.050 ;
        RECT 760.950 204.600 763.050 205.050 ;
        RECT 748.950 203.400 763.050 204.600 ;
        RECT 748.950 202.950 751.050 203.400 ;
        RECT 760.950 202.950 763.050 203.400 ;
        RECT 766.950 204.600 769.050 205.050 ;
        RECT 775.950 204.600 778.050 205.050 ;
        RECT 766.950 203.400 778.050 204.600 ;
        RECT 766.950 202.950 769.050 203.400 ;
        RECT 775.950 202.950 778.050 203.400 ;
        RECT 898.950 204.600 901.050 205.050 ;
        RECT 913.950 204.600 916.050 205.050 ;
        RECT 898.950 203.400 916.050 204.600 ;
        RECT 898.950 202.950 901.050 203.400 ;
        RECT 913.950 202.950 916.050 203.400 ;
        RECT 550.950 200.400 585.600 201.600 ;
        RECT 592.950 201.600 595.050 202.050 ;
        RECT 646.950 201.600 649.050 202.050 ;
        RECT 592.950 200.400 649.050 201.600 ;
        RECT 550.950 199.950 553.050 200.400 ;
        RECT 592.950 199.950 595.050 200.400 ;
        RECT 646.950 199.950 649.050 200.400 ;
        RECT 661.950 201.600 664.050 202.050 ;
        RECT 769.950 201.600 772.050 202.050 ;
        RECT 661.950 200.400 772.050 201.600 ;
        RECT 661.950 199.950 664.050 200.400 ;
        RECT 769.950 199.950 772.050 200.400 ;
        RECT 781.950 201.600 784.050 202.050 ;
        RECT 829.950 201.600 832.050 201.900 ;
        RECT 781.950 200.400 832.050 201.600 ;
        RECT 781.950 199.950 784.050 200.400 ;
        RECT 829.950 199.800 832.050 200.400 ;
        RECT 862.950 201.600 865.050 202.050 ;
        RECT 889.950 201.600 892.050 202.050 ;
        RECT 862.950 200.400 892.050 201.600 ;
        RECT 862.950 199.950 865.050 200.400 ;
        RECT 889.950 199.950 892.050 200.400 ;
        RECT 49.950 198.600 52.050 199.050 ;
        RECT 94.950 198.600 97.050 199.050 ;
        RECT 133.950 198.600 136.050 199.050 ;
        RECT 49.950 197.400 97.050 198.600 ;
        RECT 49.950 196.950 52.050 197.400 ;
        RECT 94.950 196.950 97.050 197.400 ;
        RECT 98.400 197.400 136.050 198.600 ;
        RECT 70.950 195.600 73.050 196.050 ;
        RECT 98.400 195.600 99.600 197.400 ;
        RECT 133.950 196.950 136.050 197.400 ;
        RECT 181.950 198.600 184.050 199.050 ;
        RECT 187.950 198.600 190.050 199.050 ;
        RECT 223.950 198.600 226.050 199.050 ;
        RECT 181.950 197.400 226.050 198.600 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 187.950 196.950 190.050 197.400 ;
        RECT 223.950 196.950 226.050 197.400 ;
        RECT 454.950 198.600 457.050 199.050 ;
        RECT 463.950 198.600 466.050 199.050 ;
        RECT 454.950 197.400 466.050 198.600 ;
        RECT 454.950 196.950 457.050 197.400 ;
        RECT 463.950 196.950 466.050 197.400 ;
        RECT 493.950 198.600 496.050 199.050 ;
        RECT 613.950 198.600 616.050 199.050 ;
        RECT 652.950 198.600 655.050 199.050 ;
        RECT 493.950 197.400 655.050 198.600 ;
        RECT 493.950 196.950 496.050 197.400 ;
        RECT 613.950 196.950 616.050 197.400 ;
        RECT 652.950 196.950 655.050 197.400 ;
        RECT 658.950 198.600 661.050 199.050 ;
        RECT 772.950 198.600 775.050 199.050 ;
        RECT 658.950 197.400 775.050 198.600 ;
        RECT 658.950 196.950 661.050 197.400 ;
        RECT 772.950 196.950 775.050 197.400 ;
        RECT 841.950 198.600 844.050 199.050 ;
        RECT 856.950 198.600 859.050 199.050 ;
        RECT 841.950 197.400 859.050 198.600 ;
        RECT 841.950 196.950 844.050 197.400 ;
        RECT 856.950 196.950 859.050 197.400 ;
        RECT 871.950 198.600 874.050 199.050 ;
        RECT 886.950 198.600 889.050 199.050 ;
        RECT 871.950 197.400 889.050 198.600 ;
        RECT 871.950 196.950 874.050 197.400 ;
        RECT 886.950 196.950 889.050 197.400 ;
        RECT 70.950 194.400 99.600 195.600 ;
        RECT 127.950 195.600 130.050 196.050 ;
        RECT 157.950 195.600 160.050 196.050 ;
        RECT 127.950 194.400 160.050 195.600 ;
        RECT 70.950 193.950 73.050 194.400 ;
        RECT 127.950 193.950 130.050 194.400 ;
        RECT 157.950 193.950 160.050 194.400 ;
        RECT 355.950 195.600 358.050 196.050 ;
        RECT 412.950 195.600 415.050 196.050 ;
        RECT 487.950 195.600 490.050 196.050 ;
        RECT 355.950 194.400 490.050 195.600 ;
        RECT 355.950 193.950 358.050 194.400 ;
        RECT 412.950 193.950 415.050 194.400 ;
        RECT 487.950 193.950 490.050 194.400 ;
        RECT 496.950 195.600 499.050 196.050 ;
        RECT 550.800 195.600 552.900 196.050 ;
        RECT 496.950 194.400 552.900 195.600 ;
        RECT 496.950 193.950 499.050 194.400 ;
        RECT 550.800 193.950 552.900 194.400 ;
        RECT 553.950 195.600 556.050 196.050 ;
        RECT 565.950 195.600 568.050 196.050 ;
        RECT 553.950 194.400 568.050 195.600 ;
        RECT 553.950 193.950 556.050 194.400 ;
        RECT 565.950 193.950 568.050 194.400 ;
        RECT 595.950 195.600 598.050 196.050 ;
        RECT 619.950 195.600 622.050 196.050 ;
        RECT 595.950 194.400 622.050 195.600 ;
        RECT 595.950 193.950 598.050 194.400 ;
        RECT 619.950 193.950 622.050 194.400 ;
        RECT 784.950 195.600 787.050 196.050 ;
        RECT 859.950 195.600 862.050 196.050 ;
        RECT 784.950 194.400 862.050 195.600 ;
        RECT 784.950 193.950 787.050 194.400 ;
        RECT 859.950 193.950 862.050 194.400 ;
        RECT 865.950 195.600 868.050 196.050 ;
        RECT 877.950 195.600 880.050 196.050 ;
        RECT 886.950 195.600 889.050 195.900 ;
        RECT 865.950 194.400 889.050 195.600 ;
        RECT 865.950 193.950 868.050 194.400 ;
        RECT 877.950 193.950 880.050 194.400 ;
        RECT 886.950 193.800 889.050 194.400 ;
        RECT 82.950 192.600 85.050 193.050 ;
        RECT 103.950 192.600 106.050 193.050 ;
        RECT 82.950 191.400 106.050 192.600 ;
        RECT 82.950 190.950 85.050 191.400 ;
        RECT 103.950 190.950 106.050 191.400 ;
        RECT 115.950 192.600 118.050 193.050 ;
        RECT 154.950 192.600 157.050 193.050 ;
        RECT 115.950 191.400 157.050 192.600 ;
        RECT 115.950 190.950 118.050 191.400 ;
        RECT 154.950 190.950 157.050 191.400 ;
        RECT 169.950 192.600 172.050 193.050 ;
        RECT 196.950 192.600 199.050 193.050 ;
        RECT 169.950 191.400 199.050 192.600 ;
        RECT 169.950 190.950 172.050 191.400 ;
        RECT 196.950 190.950 199.050 191.400 ;
        RECT 301.950 192.600 304.050 193.050 ;
        RECT 364.950 192.600 367.050 193.050 ;
        RECT 301.950 191.400 367.050 192.600 ;
        RECT 301.950 190.950 304.050 191.400 ;
        RECT 364.950 190.950 367.050 191.400 ;
        RECT 370.950 192.600 373.050 193.050 ;
        RECT 397.950 192.600 400.050 193.050 ;
        RECT 370.950 191.400 400.050 192.600 ;
        RECT 370.950 190.950 373.050 191.400 ;
        RECT 397.950 190.950 400.050 191.400 ;
        RECT 421.950 192.600 424.050 193.050 ;
        RECT 442.950 192.600 445.050 193.050 ;
        RECT 421.950 191.400 445.050 192.600 ;
        RECT 421.950 190.950 424.050 191.400 ;
        RECT 442.950 190.950 445.050 191.400 ;
        RECT 466.950 192.600 469.050 193.050 ;
        RECT 478.950 192.600 481.050 193.050 ;
        RECT 466.950 191.400 481.050 192.600 ;
        RECT 466.950 190.950 469.050 191.400 ;
        RECT 478.950 190.950 481.050 191.400 ;
        RECT 514.950 192.600 517.050 193.050 ;
        RECT 532.950 192.600 535.050 193.050 ;
        RECT 547.950 192.600 550.050 193.050 ;
        RECT 514.950 191.400 550.050 192.600 ;
        RECT 514.950 190.950 517.050 191.400 ;
        RECT 532.950 190.950 535.050 191.400 ;
        RECT 547.950 190.950 550.050 191.400 ;
        RECT 568.950 192.600 571.050 193.050 ;
        RECT 574.950 192.600 577.050 193.050 ;
        RECT 568.950 191.400 577.050 192.600 ;
        RECT 568.950 190.950 571.050 191.400 ;
        RECT 574.950 190.950 577.050 191.400 ;
        RECT 664.950 192.600 667.050 193.050 ;
        RECT 844.950 192.600 847.050 193.050 ;
        RECT 895.950 192.600 898.050 193.050 ;
        RECT 664.950 191.400 898.050 192.600 ;
        RECT 664.950 190.950 667.050 191.400 ;
        RECT 844.950 190.950 847.050 191.400 ;
        RECT 895.950 190.950 898.050 191.400 ;
        RECT 31.950 189.600 34.050 190.050 ;
        RECT 37.950 189.600 40.050 190.050 ;
        RECT 31.950 188.400 40.050 189.600 ;
        RECT 31.950 187.950 34.050 188.400 ;
        RECT 37.950 187.950 40.050 188.400 ;
        RECT 46.950 189.600 49.050 190.050 ;
        RECT 55.950 189.600 58.050 190.050 ;
        RECT 46.950 188.400 58.050 189.600 ;
        RECT 46.950 187.950 49.050 188.400 ;
        RECT 55.950 187.950 58.050 188.400 ;
        RECT 64.950 189.600 67.050 190.050 ;
        RECT 109.950 189.600 112.050 190.050 ;
        RECT 64.950 188.400 112.050 189.600 ;
        RECT 64.950 187.950 67.050 188.400 ;
        RECT 109.950 187.950 112.050 188.400 ;
        RECT 205.950 189.600 208.050 190.050 ;
        RECT 214.950 189.600 217.050 190.050 ;
        RECT 205.950 188.400 217.050 189.600 ;
        RECT 205.950 187.950 208.050 188.400 ;
        RECT 214.950 187.950 217.050 188.400 ;
        RECT 223.950 189.600 226.050 190.050 ;
        RECT 241.950 189.600 244.050 190.050 ;
        RECT 223.950 188.400 244.050 189.600 ;
        RECT 223.950 187.950 226.050 188.400 ;
        RECT 241.950 187.950 244.050 188.400 ;
        RECT 250.950 189.600 253.050 190.050 ;
        RECT 256.950 189.600 259.050 190.050 ;
        RECT 250.950 188.400 259.050 189.600 ;
        RECT 250.950 187.950 253.050 188.400 ;
        RECT 256.950 187.950 259.050 188.400 ;
        RECT 262.950 189.600 265.050 190.050 ;
        RECT 286.950 189.600 289.050 190.050 ;
        RECT 298.950 189.600 301.050 190.050 ;
        RECT 262.950 188.400 301.050 189.600 ;
        RECT 262.950 187.950 265.050 188.400 ;
        RECT 286.950 187.950 289.050 188.400 ;
        RECT 298.950 187.950 301.050 188.400 ;
        RECT 418.950 189.600 421.050 190.050 ;
        RECT 448.950 189.600 451.050 190.050 ;
        RECT 418.950 188.400 451.050 189.600 ;
        RECT 418.950 187.950 421.050 188.400 ;
        RECT 448.950 187.950 451.050 188.400 ;
        RECT 457.950 189.600 460.050 190.050 ;
        RECT 472.950 189.600 475.050 190.050 ;
        RECT 496.950 189.600 499.050 190.050 ;
        RECT 457.950 188.400 499.050 189.600 ;
        RECT 457.950 187.950 460.050 188.400 ;
        RECT 472.950 187.950 475.050 188.400 ;
        RECT 496.950 187.950 499.050 188.400 ;
        RECT 553.950 189.600 556.050 190.050 ;
        RECT 565.950 189.600 568.050 190.050 ;
        RECT 553.950 188.400 568.050 189.600 ;
        RECT 553.950 187.950 556.050 188.400 ;
        RECT 565.950 187.950 568.050 188.400 ;
        RECT 625.950 189.600 628.050 190.050 ;
        RECT 634.950 189.600 637.050 190.050 ;
        RECT 625.950 188.400 637.050 189.600 ;
        RECT 625.950 187.950 628.050 188.400 ;
        RECT 634.950 187.950 637.050 188.400 ;
        RECT 691.950 189.600 694.050 190.050 ;
        RECT 700.950 189.600 703.050 190.050 ;
        RECT 691.950 188.400 703.050 189.600 ;
        RECT 691.950 187.950 694.050 188.400 ;
        RECT 700.950 187.950 703.050 188.400 ;
        RECT 715.950 189.600 718.050 190.050 ;
        RECT 754.950 189.600 757.050 190.050 ;
        RECT 715.950 188.400 757.050 189.600 ;
        RECT 715.950 187.950 718.050 188.400 ;
        RECT 754.950 187.950 757.050 188.400 ;
        RECT 856.950 189.600 859.050 190.050 ;
        RECT 865.950 189.600 868.050 190.050 ;
        RECT 856.950 188.400 868.050 189.600 ;
        RECT 856.950 187.950 859.050 188.400 ;
        RECT 865.950 187.950 868.050 188.400 ;
        RECT 70.950 186.600 73.050 187.050 ;
        RECT 44.400 185.400 73.050 186.600 ;
        RECT 16.950 183.600 19.050 184.050 ;
        RECT 37.950 183.600 40.050 184.050 ;
        RECT 16.950 182.400 40.050 183.600 ;
        RECT 16.950 181.950 19.050 182.400 ;
        RECT 37.950 181.950 40.050 182.400 ;
        RECT 44.400 180.600 45.600 185.400 ;
        RECT 70.950 184.950 73.050 185.400 ;
        RECT 118.950 186.600 121.050 187.050 ;
        RECT 148.950 186.600 151.050 187.050 ;
        RECT 169.800 186.600 171.900 187.050 ;
        RECT 118.950 185.400 171.900 186.600 ;
        RECT 118.950 184.950 121.050 185.400 ;
        RECT 148.950 184.950 151.050 185.400 ;
        RECT 169.800 184.950 171.900 185.400 ;
        RECT 55.950 182.100 58.050 184.200 ;
        RECT 76.950 182.100 79.050 184.200 ;
        RECT 41.400 179.400 45.600 180.600 ;
        RECT 41.400 177.900 42.600 179.400 ;
        RECT 13.950 177.600 16.050 177.900 ;
        RECT 28.950 177.600 31.050 177.900 ;
        RECT 13.950 176.400 31.050 177.600 ;
        RECT 13.950 175.800 16.050 176.400 ;
        RECT 28.950 175.800 31.050 176.400 ;
        RECT 40.950 175.800 43.050 177.900 ;
        RECT 49.950 177.600 52.050 178.050 ;
        RECT 56.400 177.600 57.600 182.100 ;
        RECT 49.950 176.400 57.600 177.600 ;
        RECT 61.950 177.600 64.050 181.050 ;
        RECT 77.400 180.600 78.600 182.100 ;
        RECT 82.950 180.600 85.050 184.050 ;
        RECT 91.950 182.100 94.050 184.200 ;
        RECT 109.950 183.750 112.050 184.200 ;
        RECT 139.950 183.750 142.050 184.200 ;
        RECT 109.950 183.600 142.050 183.750 ;
        RECT 160.950 183.600 163.050 184.200 ;
        RECT 109.950 182.550 163.050 183.600 ;
        RECT 109.950 182.100 112.050 182.550 ;
        RECT 139.950 182.400 163.050 182.550 ;
        RECT 139.950 182.100 142.050 182.400 ;
        RECT 160.950 182.100 163.050 182.400 ;
        RECT 196.950 183.600 199.050 184.200 ;
        RECT 208.950 183.600 211.050 184.050 ;
        RECT 196.950 182.400 211.050 183.600 ;
        RECT 196.950 182.100 199.050 182.400 ;
        RECT 77.400 180.000 85.050 180.600 ;
        RECT 77.400 179.400 84.600 180.000 ;
        RECT 92.400 178.050 93.600 182.100 ;
        RECT 208.950 181.950 211.050 182.400 ;
        RECT 229.950 183.600 232.050 184.050 ;
        RECT 244.950 183.600 247.050 184.050 ;
        RECT 229.950 182.400 247.050 183.600 ;
        RECT 229.950 181.950 232.050 182.400 ;
        RECT 244.950 181.950 247.050 182.400 ;
        RECT 256.950 182.100 259.050 184.200 ;
        RECT 277.950 183.600 280.050 184.200 ;
        RECT 272.400 182.400 280.050 183.600 ;
        RECT 257.400 180.600 258.600 182.100 ;
        RECT 268.950 180.600 271.050 180.900 ;
        RECT 257.400 179.400 271.050 180.600 ;
        RECT 61.950 177.000 66.600 177.600 ;
        RECT 73.950 177.450 76.050 177.900 ;
        RECT 82.950 177.450 85.050 177.900 ;
        RECT 62.400 176.400 67.050 177.000 ;
        RECT 49.950 175.950 52.050 176.400 ;
        RECT 52.950 174.600 55.050 175.050 ;
        RECT 61.800 174.600 63.900 175.050 ;
        RECT 52.950 173.400 63.900 174.600 ;
        RECT 52.950 172.950 55.050 173.400 ;
        RECT 61.800 172.950 63.900 173.400 ;
        RECT 64.950 172.950 67.050 176.400 ;
        RECT 73.950 176.250 85.050 177.450 ;
        RECT 73.950 175.800 76.050 176.250 ;
        RECT 82.950 175.800 85.050 176.250 ;
        RECT 88.950 176.400 93.600 178.050 ;
        RECT 112.950 177.600 115.050 178.050 ;
        RECT 127.950 177.600 130.050 178.050 ;
        RECT 112.950 176.400 130.050 177.600 ;
        RECT 88.950 175.950 93.000 176.400 ;
        RECT 112.950 175.950 115.050 176.400 ;
        RECT 127.950 175.950 130.050 176.400 ;
        RECT 142.950 177.600 145.050 177.900 ;
        RECT 157.950 177.600 160.050 177.900 ;
        RECT 142.950 176.400 160.050 177.600 ;
        RECT 142.950 175.800 145.050 176.400 ;
        RECT 157.950 175.800 160.050 176.400 ;
        RECT 208.950 177.450 211.050 177.900 ;
        RECT 214.950 177.450 217.050 177.900 ;
        RECT 208.950 176.250 217.050 177.450 ;
        RECT 208.950 175.800 211.050 176.250 ;
        RECT 214.950 175.800 217.050 176.250 ;
        RECT 238.950 177.600 241.050 177.900 ;
        RECT 257.400 177.600 258.600 179.400 ;
        RECT 268.950 178.800 271.050 179.400 ;
        RECT 238.950 176.400 258.600 177.600 ;
        RECT 238.950 175.800 241.050 176.400 ;
        RECT 272.400 175.050 273.600 182.400 ;
        RECT 277.950 182.100 280.050 182.400 ;
        RECT 292.950 182.100 295.050 184.200 ;
        RECT 319.950 183.600 322.050 184.050 ;
        RECT 346.950 183.750 349.050 184.200 ;
        RECT 352.950 183.750 355.050 184.200 ;
        RECT 319.950 182.400 327.600 183.600 ;
        RECT 293.400 180.600 294.600 182.100 ;
        RECT 319.950 181.950 322.050 182.400 ;
        RECT 322.950 180.600 325.050 181.050 ;
        RECT 293.400 179.400 325.050 180.600 ;
        RECT 322.950 178.950 325.050 179.400 ;
        RECT 280.950 177.450 283.050 177.900 ;
        RECT 286.950 177.450 289.050 177.900 ;
        RECT 280.950 176.250 289.050 177.450 ;
        RECT 280.950 175.800 283.050 176.250 ;
        RECT 286.950 175.800 289.050 176.250 ;
        RECT 301.950 177.450 304.050 177.900 ;
        RECT 310.950 177.450 313.050 177.900 ;
        RECT 301.950 176.250 313.050 177.450 ;
        RECT 326.400 177.600 327.600 182.400 ;
        RECT 346.950 182.550 355.050 183.750 ;
        RECT 346.950 182.100 349.050 182.550 ;
        RECT 352.950 182.100 355.050 182.550 ;
        RECT 370.950 183.750 373.050 184.200 ;
        RECT 382.950 183.750 385.050 184.200 ;
        RECT 370.950 182.550 385.050 183.750 ;
        RECT 370.950 182.100 373.050 182.550 ;
        RECT 382.950 182.100 385.050 182.550 ;
        RECT 391.950 182.100 394.050 184.200 ;
        RECT 392.400 180.600 393.600 182.100 ;
        RECT 400.950 181.950 403.050 184.050 ;
        RECT 430.950 183.600 433.050 184.200 ;
        RECT 410.400 182.400 433.050 183.600 ;
        RECT 338.400 179.400 393.600 180.600 ;
        RECT 331.950 177.600 334.050 177.900 ;
        RECT 326.400 176.400 334.050 177.600 ;
        RECT 301.950 175.800 304.050 176.250 ;
        RECT 310.950 175.800 313.050 176.250 ;
        RECT 331.950 175.800 334.050 176.400 ;
        RECT 338.400 175.050 339.600 179.400 ;
        RECT 373.950 177.450 376.050 177.900 ;
        RECT 379.950 177.450 382.050 177.900 ;
        RECT 373.950 176.250 382.050 177.450 ;
        RECT 401.400 177.600 402.600 181.950 ;
        RECT 410.400 177.900 411.600 182.400 ;
        RECT 430.950 182.100 433.050 182.400 ;
        RECT 442.950 183.600 445.050 184.050 ;
        RECT 469.950 183.600 472.050 187.050 ;
        RECT 475.950 186.600 478.050 187.050 ;
        RECT 490.950 186.600 493.050 187.050 ;
        RECT 580.950 186.600 583.050 187.050 ;
        RECT 589.950 186.600 592.050 187.050 ;
        RECT 475.950 185.400 493.050 186.600 ;
        RECT 475.950 184.950 478.050 185.400 ;
        RECT 490.950 184.950 493.050 185.400 ;
        RECT 572.400 185.400 592.050 186.600 ;
        RECT 572.400 184.200 573.600 185.400 ;
        RECT 580.950 184.950 583.050 185.400 ;
        RECT 589.950 184.950 592.050 185.400 ;
        RECT 604.950 186.600 607.050 187.050 ;
        RECT 610.950 186.600 613.050 187.050 ;
        RECT 604.950 185.400 613.050 186.600 ;
        RECT 604.950 184.950 607.050 185.400 ;
        RECT 610.950 184.950 613.050 185.400 ;
        RECT 706.950 186.600 709.050 187.050 ;
        RECT 712.950 186.600 715.050 187.050 ;
        RECT 706.950 185.400 715.050 186.600 ;
        RECT 706.950 184.950 709.050 185.400 ;
        RECT 712.950 184.950 715.050 185.400 ;
        RECT 778.950 186.600 781.050 187.050 ;
        RECT 805.950 186.600 808.050 187.050 ;
        RECT 778.950 185.400 808.050 186.600 ;
        RECT 778.950 184.950 781.050 185.400 ;
        RECT 805.950 184.950 808.050 185.400 ;
        RECT 817.950 186.600 820.050 187.050 ;
        RECT 832.950 186.600 835.050 187.050 ;
        RECT 817.950 185.400 835.050 186.600 ;
        RECT 817.950 184.950 820.050 185.400 ;
        RECT 832.950 184.950 835.050 185.400 ;
        RECT 865.950 186.600 868.050 186.900 ;
        RECT 874.950 186.600 877.050 187.050 ;
        RECT 909.000 186.600 913.050 187.050 ;
        RECT 865.950 185.400 877.050 186.600 ;
        RECT 865.950 184.800 868.050 185.400 ;
        RECT 874.950 184.950 877.050 185.400 ;
        RECT 908.400 184.950 913.050 186.600 ;
        RECT 919.950 184.950 922.050 187.050 ;
        RECT 484.950 183.600 487.050 184.050 ;
        RECT 538.950 183.600 541.050 184.200 ;
        RECT 442.950 182.400 487.050 183.600 ;
        RECT 442.950 181.950 445.050 182.400 ;
        RECT 484.950 181.950 487.050 182.400 ;
        RECT 527.400 182.400 541.050 183.600 ;
        RECT 527.400 181.050 528.600 182.400 ;
        RECT 538.950 182.100 541.050 182.400 ;
        RECT 571.950 182.100 574.050 184.200 ;
        RECT 586.950 183.600 589.050 184.200 ;
        RECT 584.400 182.400 589.050 183.600 ;
        RECT 523.950 179.400 528.600 181.050 ;
        RECT 577.950 180.600 580.050 181.050 ;
        RECT 584.400 180.600 585.600 182.400 ;
        RECT 586.950 182.100 589.050 182.400 ;
        RECT 592.950 183.750 595.050 184.200 ;
        RECT 601.950 183.750 604.050 184.200 ;
        RECT 592.950 182.550 604.050 183.750 ;
        RECT 634.950 183.600 637.050 184.200 ;
        RECT 652.950 183.600 655.050 184.200 ;
        RECT 592.950 182.100 595.050 182.550 ;
        RECT 601.950 182.100 604.050 182.550 ;
        RECT 629.400 182.400 637.050 183.600 ;
        RECT 577.950 179.400 585.600 180.600 ;
        RECT 523.950 178.950 528.000 179.400 ;
        RECT 577.950 178.950 580.050 179.400 ;
        RECT 629.400 178.050 630.600 182.400 ;
        RECT 634.950 182.100 637.050 182.400 ;
        RECT 638.400 182.400 655.050 183.600 ;
        RECT 403.950 177.600 406.050 177.900 ;
        RECT 401.400 176.400 406.050 177.600 ;
        RECT 373.950 175.800 376.050 176.250 ;
        RECT 379.950 175.800 382.050 176.250 ;
        RECT 403.950 175.800 406.050 176.400 ;
        RECT 409.950 175.800 412.050 177.900 ;
        RECT 457.950 177.450 460.050 177.900 ;
        RECT 463.950 177.450 466.050 177.900 ;
        RECT 457.950 176.250 466.050 177.450 ;
        RECT 457.950 175.800 460.050 176.250 ;
        RECT 463.950 175.800 466.050 176.250 ;
        RECT 487.950 177.450 490.050 177.900 ;
        RECT 493.950 177.450 496.050 177.900 ;
        RECT 487.950 176.250 496.050 177.450 ;
        RECT 487.950 175.800 490.050 176.250 ;
        RECT 493.950 175.800 496.050 176.250 ;
        RECT 520.950 177.450 523.050 177.900 ;
        RECT 550.950 177.450 553.050 177.900 ;
        RECT 520.950 176.250 553.050 177.450 ;
        RECT 520.950 175.800 523.050 176.250 ;
        RECT 550.950 175.800 553.050 176.250 ;
        RECT 556.950 175.800 559.050 177.900 ;
        RECT 628.950 175.950 631.050 178.050 ;
        RECT 638.400 177.900 639.600 182.400 ;
        RECT 652.950 182.100 655.050 182.400 ;
        RECT 670.950 183.600 673.050 184.050 ;
        RECT 700.950 183.600 703.050 184.200 ;
        RECT 670.950 182.400 703.050 183.600 ;
        RECT 670.950 181.950 673.050 182.400 ;
        RECT 700.950 182.100 703.050 182.400 ;
        RECT 709.950 181.950 712.050 184.050 ;
        RECT 733.950 183.600 736.050 184.050 ;
        RECT 742.950 183.600 745.050 184.200 ;
        RECT 733.950 182.400 745.050 183.600 ;
        RECT 733.950 181.950 736.050 182.400 ;
        RECT 742.950 182.100 745.050 182.400 ;
        RECT 751.950 183.600 754.050 184.050 ;
        RECT 763.950 183.600 766.050 184.200 ;
        RECT 781.950 183.600 784.050 184.200 ;
        RECT 751.950 182.400 766.050 183.600 ;
        RECT 751.950 181.950 754.050 182.400 ;
        RECT 763.950 182.100 766.050 182.400 ;
        RECT 776.400 182.400 784.050 183.600 ;
        RECT 710.400 178.050 711.600 181.950 ;
        RECT 776.400 181.050 777.600 182.400 ;
        RECT 781.950 182.100 784.050 182.400 ;
        RECT 787.950 183.750 790.050 184.200 ;
        RECT 796.950 183.750 799.050 184.200 ;
        RECT 787.950 182.550 799.050 183.750 ;
        RECT 787.950 182.100 790.050 182.550 ;
        RECT 796.950 182.100 799.050 182.550 ;
        RECT 823.950 182.100 826.050 184.200 ;
        RECT 844.950 183.600 849.000 184.050 ;
        RECT 859.950 183.600 862.050 184.050 ;
        RECT 908.400 183.600 909.600 184.950 ;
        RECT 916.950 183.600 919.050 184.200 ;
        RECT 716.400 180.000 723.600 180.600 ;
        RECT 715.950 179.400 723.600 180.000 ;
        RECT 637.950 175.800 640.050 177.900 ;
        RECT 709.950 175.950 712.050 178.050 ;
        RECT 715.950 175.950 718.050 179.400 ;
        RECT 722.400 177.900 723.600 179.400 ;
        RECT 772.950 179.400 777.600 181.050 ;
        RECT 799.950 180.600 802.050 181.050 ;
        RECT 824.400 180.600 825.600 182.100 ;
        RECT 844.950 181.950 849.600 183.600 ;
        RECT 859.950 182.400 870.600 183.600 ;
        RECT 859.950 181.950 862.050 182.400 ;
        RECT 799.950 179.400 825.600 180.600 ;
        RECT 772.950 178.950 777.000 179.400 ;
        RECT 799.950 178.950 802.050 179.400 ;
        RECT 848.400 177.900 849.600 181.950 ;
        RECT 869.400 180.600 870.600 182.400 ;
        RECT 896.400 182.400 909.600 183.600 ;
        RECT 911.400 182.400 919.050 183.600 ;
        RECT 896.400 180.600 897.600 182.400 ;
        RECT 911.400 180.600 912.600 182.400 ;
        RECT 916.950 182.100 919.050 182.400 ;
        RECT 869.400 179.400 897.600 180.600 ;
        RECT 908.400 180.000 912.600 180.600 ;
        RECT 907.950 179.400 912.600 180.000 ;
        RECT 869.400 177.900 870.600 179.400 ;
        RECT 721.950 175.800 724.050 177.900 ;
        RECT 745.950 177.600 748.050 177.900 ;
        RECT 754.950 177.600 757.050 177.900 ;
        RECT 745.950 177.450 757.050 177.600 ;
        RECT 760.950 177.450 763.050 177.900 ;
        RECT 745.950 176.400 763.050 177.450 ;
        RECT 745.950 175.800 748.050 176.400 ;
        RECT 754.950 176.250 763.050 176.400 ;
        RECT 754.950 175.800 757.050 176.250 ;
        RECT 760.950 175.800 763.050 176.250 ;
        RECT 790.950 175.800 793.050 177.900 ;
        RECT 832.950 177.450 835.050 177.900 ;
        RECT 838.950 177.450 841.050 177.900 ;
        RECT 832.950 176.250 841.050 177.450 ;
        RECT 832.950 175.800 835.050 176.250 ;
        RECT 838.950 175.800 841.050 176.250 ;
        RECT 847.950 175.800 850.050 177.900 ;
        RECT 868.950 175.800 871.050 177.900 ;
        RECT 898.950 177.450 901.050 177.900 ;
        RECT 904.800 177.450 906.900 177.900 ;
        RECT 898.950 176.250 906.900 177.450 ;
        RECT 898.950 175.800 901.050 176.250 ;
        RECT 904.800 175.800 906.900 176.250 ;
        RECT 907.950 175.950 910.050 179.400 ;
        RECT 920.400 177.900 921.600 184.950 ;
        RECT 919.950 175.800 922.050 177.900 ;
        RECT 79.950 174.600 82.050 175.050 ;
        RECT 97.950 174.600 100.050 175.050 ;
        RECT 106.950 174.600 109.050 175.050 ;
        RECT 79.950 173.400 109.050 174.600 ;
        RECT 79.950 172.950 82.050 173.400 ;
        RECT 97.950 172.950 100.050 173.400 ;
        RECT 106.950 172.950 109.050 173.400 ;
        RECT 178.950 174.600 181.050 175.050 ;
        RECT 193.950 174.600 196.050 175.050 ;
        RECT 178.950 173.400 196.050 174.600 ;
        RECT 178.950 172.950 181.050 173.400 ;
        RECT 193.950 172.950 196.050 173.400 ;
        RECT 205.950 174.600 208.050 175.050 ;
        RECT 220.950 174.600 223.050 175.050 ;
        RECT 205.950 173.400 223.050 174.600 ;
        RECT 205.950 172.950 208.050 173.400 ;
        RECT 220.950 172.950 223.050 173.400 ;
        RECT 268.950 173.400 273.600 175.050 ;
        RECT 334.950 173.400 339.600 175.050 ;
        RECT 352.950 174.600 355.050 175.050 ;
        RECT 367.950 174.600 370.050 175.050 ;
        RECT 352.950 173.400 370.050 174.600 ;
        RECT 268.950 172.950 273.000 173.400 ;
        RECT 334.950 172.950 339.000 173.400 ;
        RECT 352.950 172.950 355.050 173.400 ;
        RECT 367.950 172.950 370.050 173.400 ;
        RECT 382.950 174.600 385.050 175.050 ;
        RECT 388.950 174.600 391.050 175.050 ;
        RECT 382.950 173.400 391.050 174.600 ;
        RECT 382.950 172.950 385.050 173.400 ;
        RECT 388.950 172.950 391.050 173.400 ;
        RECT 529.950 174.600 532.050 175.050 ;
        RECT 535.950 174.600 538.050 175.050 ;
        RECT 557.400 174.600 558.600 175.800 ;
        RECT 529.950 173.400 558.600 174.600 ;
        RECT 607.950 174.600 610.050 175.050 ;
        RECT 631.950 174.600 634.050 175.050 ;
        RECT 649.950 174.600 652.050 175.050 ;
        RECT 607.950 173.400 652.050 174.600 ;
        RECT 529.950 172.950 532.050 173.400 ;
        RECT 535.950 172.950 538.050 173.400 ;
        RECT 607.950 172.950 610.050 173.400 ;
        RECT 631.950 172.950 634.050 173.400 ;
        RECT 649.950 172.950 652.050 173.400 ;
        RECT 679.950 174.600 682.050 175.050 ;
        RECT 718.950 174.600 721.050 175.050 ;
        RECT 679.950 173.400 721.050 174.600 ;
        RECT 679.950 172.950 682.050 173.400 ;
        RECT 718.950 172.950 721.050 173.400 ;
        RECT 730.950 174.600 733.050 175.050 ;
        RECT 739.950 174.600 742.050 175.050 ;
        RECT 730.950 173.400 742.050 174.600 ;
        RECT 791.400 174.600 792.600 175.800 ;
        RECT 802.950 174.600 805.050 175.050 ;
        RECT 791.400 173.400 805.050 174.600 ;
        RECT 730.950 172.950 733.050 173.400 ;
        RECT 739.950 172.950 742.050 173.400 ;
        RECT 802.950 172.950 805.050 173.400 ;
        RECT 853.950 174.600 856.050 175.050 ;
        RECT 874.950 174.600 877.050 175.050 ;
        RECT 853.950 173.400 877.050 174.600 ;
        RECT 853.950 172.950 856.050 173.400 ;
        RECT 874.950 172.950 877.050 173.400 ;
        RECT 100.950 171.600 103.050 172.050 ;
        RECT 115.950 171.600 118.050 172.050 ;
        RECT 100.950 170.400 118.050 171.600 ;
        RECT 100.950 169.950 103.050 170.400 ;
        RECT 115.950 169.950 118.050 170.400 ;
        RECT 322.950 171.600 325.050 172.050 ;
        RECT 331.950 171.600 334.050 172.050 ;
        RECT 340.950 171.600 343.050 172.050 ;
        RECT 322.950 170.400 343.050 171.600 ;
        RECT 322.950 169.950 325.050 170.400 ;
        RECT 331.950 169.950 334.050 170.400 ;
        RECT 340.950 169.950 343.050 170.400 ;
        RECT 364.950 171.600 367.050 172.050 ;
        RECT 403.950 171.600 406.050 172.050 ;
        RECT 364.950 170.400 406.050 171.600 ;
        RECT 364.950 169.950 367.050 170.400 ;
        RECT 403.950 169.950 406.050 170.400 ;
        RECT 427.950 171.600 430.050 172.050 ;
        RECT 436.950 171.600 439.050 172.050 ;
        RECT 427.950 170.400 439.050 171.600 ;
        RECT 427.950 169.950 430.050 170.400 ;
        RECT 436.950 169.950 439.050 170.400 ;
        RECT 481.950 171.600 484.050 172.050 ;
        RECT 499.950 171.600 502.050 172.050 ;
        RECT 481.950 170.400 502.050 171.600 ;
        RECT 481.950 169.950 484.050 170.400 ;
        RECT 499.950 169.950 502.050 170.400 ;
        RECT 574.950 171.600 577.050 172.050 ;
        RECT 595.950 171.600 598.050 172.050 ;
        RECT 574.950 170.400 598.050 171.600 ;
        RECT 574.950 169.950 577.050 170.400 ;
        RECT 595.950 169.950 598.050 170.400 ;
        RECT 661.950 171.600 664.050 172.050 ;
        RECT 682.950 171.600 685.050 172.050 ;
        RECT 661.950 170.400 685.050 171.600 ;
        RECT 661.950 169.950 664.050 170.400 ;
        RECT 682.950 169.950 685.050 170.400 ;
        RECT 886.950 171.600 889.050 172.050 ;
        RECT 913.950 171.600 916.050 172.050 ;
        RECT 886.950 170.400 916.050 171.600 ;
        RECT 886.950 169.950 889.050 170.400 ;
        RECT 913.950 169.950 916.050 170.400 ;
        RECT 19.950 168.600 22.050 169.050 ;
        RECT 34.950 168.600 37.050 169.050 ;
        RECT 19.950 167.400 37.050 168.600 ;
        RECT 19.950 166.950 22.050 167.400 ;
        RECT 34.950 166.950 37.050 167.400 ;
        RECT 49.950 168.600 52.050 169.050 ;
        RECT 88.950 168.600 91.050 169.050 ;
        RECT 49.950 167.400 91.050 168.600 ;
        RECT 49.950 166.950 52.050 167.400 ;
        RECT 88.950 166.950 91.050 167.400 ;
        RECT 94.950 168.600 97.050 169.050 ;
        RECT 109.950 168.600 112.050 169.050 ;
        RECT 94.950 167.400 112.050 168.600 ;
        RECT 94.950 166.950 97.050 167.400 ;
        RECT 109.950 166.950 112.050 167.400 ;
        RECT 163.950 168.600 166.050 169.050 ;
        RECT 199.950 168.600 202.050 169.050 ;
        RECT 265.950 168.600 268.050 169.050 ;
        RECT 163.950 167.400 268.050 168.600 ;
        RECT 163.950 166.950 166.050 167.400 ;
        RECT 199.950 166.950 202.050 167.400 ;
        RECT 265.950 166.950 268.050 167.400 ;
        RECT 622.950 168.600 625.050 169.050 ;
        RECT 700.950 168.600 703.050 169.050 ;
        RECT 622.950 167.400 703.050 168.600 ;
        RECT 622.950 166.950 625.050 167.400 ;
        RECT 700.950 166.950 703.050 167.400 ;
        RECT 706.950 168.600 709.050 169.050 ;
        RECT 766.950 168.600 769.050 169.050 ;
        RECT 706.950 167.400 769.050 168.600 ;
        RECT 706.950 166.950 709.050 167.400 ;
        RECT 766.950 166.950 769.050 167.400 ;
        RECT 787.950 168.600 790.050 169.050 ;
        RECT 796.950 168.600 799.050 169.050 ;
        RECT 787.950 167.400 799.050 168.600 ;
        RECT 787.950 166.950 790.050 167.400 ;
        RECT 796.950 166.950 799.050 167.400 ;
        RECT 874.950 168.600 877.050 169.050 ;
        RECT 892.950 168.600 895.050 169.050 ;
        RECT 874.950 167.400 895.050 168.600 ;
        RECT 874.950 166.950 877.050 167.400 ;
        RECT 892.950 166.950 895.050 167.400 ;
        RECT 346.950 165.600 349.050 166.050 ;
        RECT 409.950 165.600 412.050 166.050 ;
        RECT 346.950 164.400 412.050 165.600 ;
        RECT 346.950 163.950 349.050 164.400 ;
        RECT 409.950 163.950 412.050 164.400 ;
        RECT 475.950 165.600 478.050 166.050 ;
        RECT 547.950 165.600 550.050 166.050 ;
        RECT 619.950 165.600 622.050 166.050 ;
        RECT 772.950 165.600 775.050 166.050 ;
        RECT 475.950 164.400 775.050 165.600 ;
        RECT 475.950 163.950 478.050 164.400 ;
        RECT 547.950 163.950 550.050 164.400 ;
        RECT 619.950 163.950 622.050 164.400 ;
        RECT 772.950 163.950 775.050 164.400 ;
        RECT 31.950 162.600 34.050 163.050 ;
        RECT 49.950 162.600 52.050 163.050 ;
        RECT 31.950 161.400 52.050 162.600 ;
        RECT 31.950 160.950 34.050 161.400 ;
        RECT 49.950 160.950 52.050 161.400 ;
        RECT 484.950 162.600 487.050 163.050 ;
        RECT 511.950 162.600 514.050 163.050 ;
        RECT 484.950 161.400 514.050 162.600 ;
        RECT 484.950 160.950 487.050 161.400 ;
        RECT 511.950 160.950 514.050 161.400 ;
        RECT 541.950 162.600 544.050 163.050 ;
        RECT 580.950 162.600 583.050 163.050 ;
        RECT 541.950 161.400 583.050 162.600 ;
        RECT 541.950 160.950 544.050 161.400 ;
        RECT 580.950 160.950 583.050 161.400 ;
        RECT 589.950 162.600 592.050 163.050 ;
        RECT 670.950 162.600 673.050 163.050 ;
        RECT 589.950 161.400 673.050 162.600 ;
        RECT 589.950 160.950 592.050 161.400 ;
        RECT 670.950 160.950 673.050 161.400 ;
        RECT 691.950 162.600 694.050 163.050 ;
        RECT 706.950 162.600 709.050 163.050 ;
        RECT 691.950 161.400 709.050 162.600 ;
        RECT 691.950 160.950 694.050 161.400 ;
        RECT 706.950 160.950 709.050 161.400 ;
        RECT 802.950 162.600 805.050 163.050 ;
        RECT 853.950 162.600 856.050 163.050 ;
        RECT 802.950 161.400 856.050 162.600 ;
        RECT 802.950 160.950 805.050 161.400 ;
        RECT 853.950 160.950 856.050 161.400 ;
        RECT 595.950 159.600 598.050 160.050 ;
        RECT 625.950 159.600 628.050 160.050 ;
        RECT 595.950 158.400 628.050 159.600 ;
        RECT 595.950 157.950 598.050 158.400 ;
        RECT 625.950 157.950 628.050 158.400 ;
        RECT 637.950 159.600 640.050 160.050 ;
        RECT 661.950 159.600 664.050 160.050 ;
        RECT 637.950 158.400 664.050 159.600 ;
        RECT 637.950 157.950 640.050 158.400 ;
        RECT 661.950 157.950 664.050 158.400 ;
        RECT 883.950 159.600 886.050 160.050 ;
        RECT 913.950 159.600 916.050 160.050 ;
        RECT 883.950 158.400 916.050 159.600 ;
        RECT 883.950 157.950 886.050 158.400 ;
        RECT 913.950 157.950 916.050 158.400 ;
        RECT 136.950 156.600 139.050 157.050 ;
        RECT 229.950 156.600 232.050 157.050 ;
        RECT 136.950 155.400 232.050 156.600 ;
        RECT 136.950 154.950 139.050 155.400 ;
        RECT 229.950 154.950 232.050 155.400 ;
        RECT 397.950 156.600 400.050 157.050 ;
        RECT 412.950 156.600 415.050 157.050 ;
        RECT 397.950 155.400 415.050 156.600 ;
        RECT 397.950 154.950 400.050 155.400 ;
        RECT 412.950 154.950 415.050 155.400 ;
        RECT 505.950 156.600 508.050 157.050 ;
        RECT 532.950 156.600 535.050 157.050 ;
        RECT 505.950 155.400 535.050 156.600 ;
        RECT 505.950 154.950 508.050 155.400 ;
        RECT 532.950 154.950 535.050 155.400 ;
        RECT 565.950 156.600 568.050 157.050 ;
        RECT 589.950 156.600 592.050 157.050 ;
        RECT 565.950 155.400 592.050 156.600 ;
        RECT 565.950 154.950 568.050 155.400 ;
        RECT 589.950 154.950 592.050 155.400 ;
        RECT 655.950 156.600 658.050 157.050 ;
        RECT 667.950 156.600 670.050 157.050 ;
        RECT 697.950 156.600 700.050 157.050 ;
        RECT 733.950 156.600 736.050 157.050 ;
        RECT 655.950 155.400 736.050 156.600 ;
        RECT 655.950 154.950 658.050 155.400 ;
        RECT 667.950 154.950 670.050 155.400 ;
        RECT 697.950 154.950 700.050 155.400 ;
        RECT 733.950 154.950 736.050 155.400 ;
        RECT 862.950 156.600 865.050 157.050 ;
        RECT 883.950 156.600 886.050 156.900 ;
        RECT 862.950 155.400 886.050 156.600 ;
        RECT 862.950 154.950 865.050 155.400 ;
        RECT 883.950 154.800 886.050 155.400 ;
        RECT 928.950 153.600 931.050 154.050 ;
        RECT 872.400 152.400 931.050 153.600 ;
        RECT 43.950 150.600 46.050 151.050 ;
        RECT 58.950 150.600 61.050 151.050 ;
        RECT 43.950 149.400 61.050 150.600 ;
        RECT 43.950 148.950 46.050 149.400 ;
        RECT 58.950 148.950 61.050 149.400 ;
        RECT 160.950 150.600 163.050 151.050 ;
        RECT 328.950 150.600 331.050 151.050 ;
        RECT 160.950 149.400 331.050 150.600 ;
        RECT 160.950 148.950 163.050 149.400 ;
        RECT 328.950 148.950 331.050 149.400 ;
        RECT 400.950 150.600 403.050 151.050 ;
        RECT 421.950 150.600 424.050 151.050 ;
        RECT 400.950 149.400 424.050 150.600 ;
        RECT 400.950 148.950 403.050 149.400 ;
        RECT 421.950 148.950 424.050 149.400 ;
        RECT 481.950 150.600 484.050 151.050 ;
        RECT 508.950 150.600 511.050 151.050 ;
        RECT 577.950 150.600 580.050 151.050 ;
        RECT 583.950 150.600 586.050 151.050 ;
        RECT 601.950 150.600 604.050 151.050 ;
        RECT 481.950 149.400 604.050 150.600 ;
        RECT 481.950 148.950 484.050 149.400 ;
        RECT 508.950 148.950 511.050 149.400 ;
        RECT 577.950 148.950 580.050 149.400 ;
        RECT 583.950 148.950 586.050 149.400 ;
        RECT 601.950 148.950 604.050 149.400 ;
        RECT 628.950 150.600 631.050 151.050 ;
        RECT 709.950 150.600 712.050 151.050 ;
        RECT 730.950 150.600 733.050 151.050 ;
        RECT 742.950 150.600 745.050 151.050 ;
        RECT 872.400 150.600 873.600 152.400 ;
        RECT 928.950 151.950 931.050 152.400 ;
        RECT 628.950 149.400 745.050 150.600 ;
        RECT 628.950 148.950 631.050 149.400 ;
        RECT 709.950 148.950 712.050 149.400 ;
        RECT 730.950 148.950 733.050 149.400 ;
        RECT 742.950 148.950 745.050 149.400 ;
        RECT 869.400 149.400 873.600 150.600 ;
        RECT 869.400 148.050 870.600 149.400 ;
        RECT 199.950 147.600 202.050 148.050 ;
        RECT 208.950 147.600 211.050 148.050 ;
        RECT 259.950 147.600 262.050 148.050 ;
        RECT 199.950 146.400 262.050 147.600 ;
        RECT 199.950 145.950 202.050 146.400 ;
        RECT 208.950 145.950 211.050 146.400 ;
        RECT 259.950 145.950 262.050 146.400 ;
        RECT 283.950 147.600 286.050 148.050 ;
        RECT 322.950 147.600 325.050 148.050 ;
        RECT 283.950 146.400 325.050 147.600 ;
        RECT 283.950 145.950 286.050 146.400 ;
        RECT 322.950 145.950 325.050 146.400 ;
        RECT 370.950 147.600 373.050 148.050 ;
        RECT 376.950 147.600 379.050 148.050 ;
        RECT 397.950 147.600 400.050 148.050 ;
        RECT 370.950 146.400 400.050 147.600 ;
        RECT 370.950 145.950 373.050 146.400 ;
        RECT 376.950 145.950 379.050 146.400 ;
        RECT 397.950 145.950 400.050 146.400 ;
        RECT 556.950 147.600 559.050 148.050 ;
        RECT 574.950 147.600 577.050 148.050 ;
        RECT 556.950 146.400 577.050 147.600 ;
        RECT 556.950 145.950 559.050 146.400 ;
        RECT 574.950 145.950 577.050 146.400 ;
        RECT 688.950 147.600 691.050 148.050 ;
        RECT 694.950 147.600 697.050 148.050 ;
        RECT 706.950 147.600 709.050 148.050 ;
        RECT 868.950 147.600 871.050 148.050 ;
        RECT 688.950 146.400 709.050 147.600 ;
        RECT 688.950 145.950 691.050 146.400 ;
        RECT 694.950 145.950 697.050 146.400 ;
        RECT 706.950 145.950 709.050 146.400 ;
        RECT 839.400 146.400 871.050 147.600 ;
        RECT 839.400 145.050 840.600 146.400 ;
        RECT 868.950 145.950 871.050 146.400 ;
        RECT 874.950 147.600 877.050 148.050 ;
        RECT 889.950 147.600 892.050 148.050 ;
        RECT 910.950 147.600 913.050 148.050 ;
        RECT 874.950 146.400 913.050 147.600 ;
        RECT 874.950 145.950 877.050 146.400 ;
        RECT 889.950 145.950 892.050 146.400 ;
        RECT 910.950 145.950 913.050 146.400 ;
        RECT 193.950 144.600 196.050 145.050 ;
        RECT 268.950 144.600 271.050 145.050 ;
        RECT 193.950 143.400 271.050 144.600 ;
        RECT 193.950 142.950 196.050 143.400 ;
        RECT 268.950 142.950 271.050 143.400 ;
        RECT 634.950 144.600 637.050 145.050 ;
        RECT 778.950 144.600 781.050 145.050 ;
        RECT 796.950 144.600 799.050 145.050 ;
        RECT 634.950 143.400 666.600 144.600 ;
        RECT 634.950 142.950 637.050 143.400 ;
        RECT 665.400 142.050 666.600 143.400 ;
        RECT 778.950 143.400 799.050 144.600 ;
        RECT 778.950 142.950 781.050 143.400 ;
        RECT 796.950 142.950 799.050 143.400 ;
        RECT 808.950 144.600 811.050 145.050 ;
        RECT 838.950 144.600 841.050 145.050 ;
        RECT 808.950 143.400 841.050 144.600 ;
        RECT 808.950 142.950 811.050 143.400 ;
        RECT 838.950 142.950 841.050 143.400 ;
        RECT 844.950 144.600 847.050 145.050 ;
        RECT 856.950 144.600 859.050 145.050 ;
        RECT 871.950 144.600 874.050 145.050 ;
        RECT 844.950 143.400 874.050 144.600 ;
        RECT 844.950 142.950 847.050 143.400 ;
        RECT 856.950 142.950 859.050 143.400 ;
        RECT 871.950 142.950 874.050 143.400 ;
        RECT 130.950 141.600 133.050 142.050 ;
        RECT 313.950 141.600 316.050 142.050 ;
        RECT 340.950 141.600 343.050 142.050 ;
        RECT 130.950 140.400 276.600 141.600 ;
        RECT 130.950 139.950 133.050 140.400 ;
        RECT 152.400 139.200 153.600 140.400 ;
        RECT 16.950 137.100 19.050 139.200 ;
        RECT 31.800 138.000 33.900 139.050 ;
        RECT 17.400 135.600 18.600 137.100 ;
        RECT 31.800 136.950 34.050 138.000 ;
        RECT 34.950 137.100 37.050 139.200 ;
        RECT 40.950 137.100 43.050 139.200 ;
        RECT 58.950 138.600 61.050 139.200 ;
        RECT 67.950 138.750 70.050 139.200 ;
        RECT 76.950 138.750 79.050 139.200 ;
        RECT 67.950 138.600 79.050 138.750 ;
        RECT 58.950 137.550 79.050 138.600 ;
        RECT 58.950 137.400 70.050 137.550 ;
        RECT 58.950 137.100 61.050 137.400 ;
        RECT 67.950 137.100 70.050 137.400 ;
        RECT 76.950 137.100 79.050 137.550 ;
        RECT 82.950 137.100 85.050 139.200 ;
        RECT 91.950 138.750 94.050 139.200 ;
        RECT 103.950 138.750 106.050 139.200 ;
        RECT 91.950 137.550 106.050 138.750 ;
        RECT 91.950 137.100 94.050 137.550 ;
        RECT 103.950 137.100 106.050 137.550 ;
        RECT 115.950 138.750 118.050 139.200 ;
        RECT 124.950 138.750 127.050 139.200 ;
        RECT 115.950 137.550 127.050 138.750 ;
        RECT 115.950 137.100 118.050 137.550 ;
        RECT 124.950 137.100 127.050 137.550 ;
        RECT 145.950 137.100 148.050 139.200 ;
        RECT 151.950 137.100 154.050 139.200 ;
        RECT 181.950 138.750 184.050 139.200 ;
        RECT 187.950 138.750 190.050 139.200 ;
        RECT 181.950 137.550 190.050 138.750 ;
        RECT 181.950 137.100 184.050 137.550 ;
        RECT 187.950 137.100 190.050 137.550 ;
        RECT 217.950 138.600 220.050 139.200 ;
        RECT 235.950 138.600 238.050 139.200 ;
        RECT 217.950 137.400 238.050 138.600 ;
        RECT 217.950 137.100 220.050 137.400 ;
        RECT 235.950 137.100 238.050 137.400 ;
        RECT 241.950 138.600 244.050 139.200 ;
        RECT 256.950 138.600 259.050 139.200 ;
        RECT 241.950 137.400 259.050 138.600 ;
        RECT 241.950 137.100 244.050 137.400 ;
        RECT 256.950 137.100 259.050 137.400 ;
        RECT 271.950 137.100 274.050 139.200 ;
        RECT 275.400 138.600 276.600 140.400 ;
        RECT 313.950 140.400 343.050 141.600 ;
        RECT 313.950 139.950 316.050 140.400 ;
        RECT 340.950 139.950 343.050 140.400 ;
        RECT 382.950 141.600 385.050 142.050 ;
        RECT 388.950 141.600 391.050 142.050 ;
        RECT 382.950 140.400 391.050 141.600 ;
        RECT 382.950 139.950 385.050 140.400 ;
        RECT 388.950 139.950 391.050 140.400 ;
        RECT 403.950 141.600 406.050 142.050 ;
        RECT 409.950 141.600 412.050 142.050 ;
        RECT 418.950 141.600 421.050 142.050 ;
        RECT 403.950 140.400 421.050 141.600 ;
        RECT 403.950 139.950 406.050 140.400 ;
        RECT 409.950 139.950 412.050 140.400 ;
        RECT 418.950 139.950 421.050 140.400 ;
        RECT 484.950 141.600 487.050 142.050 ;
        RECT 517.950 141.600 520.050 142.050 ;
        RECT 484.950 140.400 520.050 141.600 ;
        RECT 484.950 139.950 487.050 140.400 ;
        RECT 517.950 139.950 520.050 140.400 ;
        RECT 616.950 141.600 619.050 142.050 ;
        RECT 631.950 141.600 634.050 142.050 ;
        RECT 616.950 140.400 634.050 141.600 ;
        RECT 616.950 139.950 619.050 140.400 ;
        RECT 631.950 139.950 634.050 140.400 ;
        RECT 664.950 141.600 667.050 142.050 ;
        RECT 673.950 141.600 676.050 142.050 ;
        RECT 802.950 141.600 805.050 142.050 ;
        RECT 664.950 140.400 676.050 141.600 ;
        RECT 664.950 139.950 667.050 140.400 ;
        RECT 673.950 139.950 676.050 140.400 ;
        RECT 788.400 140.400 805.050 141.600 ;
        RECT 277.950 138.600 280.050 139.200 ;
        RECT 275.400 137.400 280.050 138.600 ;
        RECT 277.950 137.100 280.050 137.400 ;
        RECT 289.950 138.750 292.050 139.200 ;
        RECT 295.950 138.750 298.050 139.200 ;
        RECT 289.950 137.550 298.050 138.750 ;
        RECT 289.950 137.100 292.050 137.550 ;
        RECT 295.950 137.100 298.050 137.550 ;
        RECT 301.950 138.750 304.050 139.200 ;
        RECT 310.950 138.750 313.050 139.200 ;
        RECT 301.950 137.550 313.050 138.750 ;
        RECT 367.950 138.600 370.050 139.050 ;
        RECT 301.950 137.100 304.050 137.550 ;
        RECT 310.950 137.100 313.050 137.550 ;
        RECT 359.400 137.400 370.050 138.600 ;
        RECT 31.950 135.600 34.050 136.950 ;
        RECT 11.400 135.000 18.600 135.600 ;
        RECT 10.950 134.400 18.600 135.000 ;
        RECT 20.400 135.000 34.050 135.600 ;
        RECT 20.400 134.400 33.450 135.000 ;
        RECT 10.950 130.950 13.050 134.400 ;
        RECT 20.400 132.900 21.600 134.400 ;
        RECT 35.400 133.050 36.600 137.100 ;
        RECT 41.400 135.600 42.600 137.100 ;
        RECT 41.400 134.400 45.600 135.600 ;
        RECT 19.950 130.800 22.050 132.900 ;
        RECT 31.950 131.400 36.600 133.050 ;
        RECT 44.400 132.600 45.600 134.400 ;
        RECT 83.400 133.050 84.600 137.100 ;
        RECT 146.400 135.600 147.600 137.100 ;
        RECT 140.400 135.000 147.600 135.600 ;
        RECT 139.950 134.400 147.600 135.000 ;
        RECT 272.400 135.600 273.600 137.100 ;
        RECT 290.400 135.600 291.600 137.100 ;
        RECT 272.400 134.400 291.600 135.600 ;
        RECT 73.950 132.600 76.050 132.900 ;
        RECT 44.400 131.400 76.050 132.600 ;
        RECT 83.400 131.400 88.050 133.050 ;
        RECT 31.950 130.950 36.000 131.400 ;
        RECT 73.950 130.800 76.050 131.400 ;
        RECT 84.000 130.950 88.050 131.400 ;
        RECT 106.950 132.600 109.050 132.900 ;
        RECT 112.950 132.600 115.050 133.050 ;
        RECT 106.950 131.400 115.050 132.600 ;
        RECT 106.950 130.800 109.050 131.400 ;
        RECT 112.950 130.950 115.050 131.400 ;
        RECT 139.950 130.950 142.050 134.400 ;
        RECT 359.400 133.050 360.600 137.400 ;
        RECT 367.950 136.950 370.050 137.400 ;
        RECT 391.950 138.600 394.050 139.050 ;
        RECT 397.950 138.600 400.050 139.200 ;
        RECT 391.950 137.400 400.050 138.600 ;
        RECT 391.950 136.950 394.050 137.400 ;
        RECT 397.950 137.100 400.050 137.400 ;
        RECT 421.950 138.750 424.050 139.200 ;
        RECT 433.950 138.750 436.050 139.200 ;
        RECT 421.950 137.550 436.050 138.750 ;
        RECT 421.950 137.100 424.050 137.550 ;
        RECT 433.950 137.100 436.050 137.550 ;
        RECT 469.950 138.750 472.050 139.200 ;
        RECT 508.950 138.750 511.050 139.200 ;
        RECT 469.950 137.550 511.050 138.750 ;
        RECT 469.950 137.100 472.050 137.550 ;
        RECT 508.950 137.100 511.050 137.550 ;
        RECT 517.950 138.600 520.050 139.200 ;
        RECT 535.950 138.750 538.050 139.200 ;
        RECT 553.950 138.750 556.050 139.200 ;
        RECT 535.950 138.600 556.050 138.750 ;
        RECT 517.950 137.550 556.050 138.600 ;
        RECT 517.950 137.400 538.050 137.550 ;
        RECT 517.950 137.100 520.050 137.400 ;
        RECT 535.950 137.100 538.050 137.400 ;
        RECT 553.950 137.100 556.050 137.550 ;
        RECT 571.950 138.600 574.050 139.200 ;
        RECT 589.950 138.600 592.050 139.200 ;
        RECT 601.950 138.600 604.050 139.200 ;
        RECT 571.950 137.400 604.050 138.600 ;
        RECT 571.950 137.100 574.050 137.400 ;
        RECT 589.950 137.100 592.050 137.400 ;
        RECT 601.950 137.100 604.050 137.400 ;
        RECT 607.950 137.100 610.050 139.200 ;
        RECT 631.950 138.600 634.050 139.200 ;
        RECT 649.950 138.600 652.050 139.200 ;
        RECT 694.950 138.600 697.050 139.200 ;
        RECT 631.950 137.400 652.050 138.600 ;
        RECT 631.950 137.100 634.050 137.400 ;
        RECT 649.950 137.100 652.050 137.400 ;
        RECT 674.400 137.400 697.050 138.600 ;
        RECT 436.950 135.600 439.050 136.050 ;
        RECT 460.950 135.600 463.050 136.050 ;
        RECT 362.400 134.400 429.600 135.600 ;
        RECT 208.950 132.450 211.050 132.900 ;
        RECT 214.950 132.600 217.050 132.900 ;
        RECT 229.950 132.600 232.050 133.050 ;
        RECT 214.950 132.450 232.050 132.600 ;
        RECT 208.950 131.400 232.050 132.450 ;
        RECT 208.950 131.250 217.050 131.400 ;
        RECT 208.950 130.800 211.050 131.250 ;
        RECT 214.950 130.800 217.050 131.250 ;
        RECT 229.950 130.950 232.050 131.400 ;
        RECT 238.950 132.450 241.050 132.900 ;
        RECT 265.950 132.450 268.050 132.900 ;
        RECT 238.950 131.250 268.050 132.450 ;
        RECT 238.950 130.800 241.050 131.250 ;
        RECT 265.950 130.800 268.050 131.250 ;
        RECT 274.950 132.600 277.050 132.900 ;
        RECT 298.950 132.600 301.050 132.900 ;
        RECT 274.950 131.400 301.050 132.600 ;
        RECT 274.950 130.800 277.050 131.400 ;
        RECT 298.950 130.800 301.050 131.400 ;
        RECT 304.950 132.600 307.050 132.900 ;
        RECT 313.950 132.600 316.050 133.050 ;
        RECT 304.950 131.400 316.050 132.600 ;
        RECT 304.950 130.800 307.050 131.400 ;
        RECT 313.950 130.950 316.050 131.400 ;
        RECT 358.800 130.950 360.900 133.050 ;
        RECT 362.400 132.900 363.600 134.400 ;
        RECT 361.950 130.800 364.050 132.900 ;
        RECT 379.950 132.600 382.050 132.900 ;
        RECT 424.950 132.600 427.050 132.900 ;
        RECT 379.950 131.400 427.050 132.600 ;
        RECT 428.400 132.600 429.600 134.400 ;
        RECT 436.950 134.400 463.050 135.600 ;
        RECT 608.400 135.600 609.600 137.100 ;
        RECT 616.950 135.600 619.050 136.050 ;
        RECT 674.400 135.600 675.600 137.400 ;
        RECT 694.950 137.100 697.050 137.400 ;
        RECT 712.950 138.600 715.050 139.050 ;
        RECT 739.950 138.600 742.050 139.050 ;
        RECT 712.950 137.400 742.050 138.600 ;
        RECT 712.950 136.950 715.050 137.400 ;
        RECT 739.950 136.950 742.050 137.400 ;
        RECT 745.950 138.600 748.050 139.050 ;
        RECT 751.950 138.600 754.050 139.050 ;
        RECT 745.950 137.400 754.050 138.600 ;
        RECT 745.950 136.950 748.050 137.400 ;
        RECT 751.950 136.950 754.050 137.400 ;
        RECT 772.950 138.600 775.050 139.200 ;
        RECT 788.400 138.600 789.600 140.400 ;
        RECT 802.950 139.950 805.050 140.400 ;
        RECT 772.950 137.400 789.600 138.600 ;
        RECT 772.950 137.100 775.050 137.400 ;
        RECT 608.400 134.400 619.050 135.600 ;
        RECT 436.950 133.950 439.050 134.400 ;
        RECT 460.950 133.950 463.050 134.400 ;
        RECT 616.950 133.950 619.050 134.400 ;
        RECT 629.400 134.400 639.600 135.600 ;
        RECT 629.400 132.900 630.600 134.400 ;
        RECT 638.400 132.900 639.600 134.400 ;
        RECT 671.400 134.400 675.600 135.600 ;
        RECT 671.400 132.900 672.600 134.400 ;
        RECT 466.950 132.600 469.050 132.900 ;
        RECT 428.400 131.400 469.050 132.600 ;
        RECT 379.950 130.800 382.050 131.400 ;
        RECT 424.950 130.800 427.050 131.400 ;
        RECT 466.950 130.800 469.050 131.400 ;
        RECT 502.950 132.600 505.050 132.900 ;
        RECT 514.950 132.600 517.050 132.900 ;
        RECT 502.950 132.450 517.050 132.600 ;
        RECT 529.950 132.600 532.050 132.900 ;
        RECT 550.950 132.600 553.050 132.900 ;
        RECT 529.950 132.450 553.050 132.600 ;
        RECT 502.950 131.400 553.050 132.450 ;
        RECT 502.950 130.800 505.050 131.400 ;
        RECT 514.950 131.250 532.050 131.400 ;
        RECT 514.950 130.800 517.050 131.250 ;
        RECT 529.950 130.800 532.050 131.250 ;
        RECT 550.950 130.800 553.050 131.400 ;
        RECT 568.950 132.450 571.050 132.900 ;
        RECT 577.950 132.450 580.050 132.900 ;
        RECT 568.950 131.250 580.050 132.450 ;
        RECT 568.950 130.800 571.050 131.250 ;
        RECT 577.950 130.800 580.050 131.250 ;
        RECT 628.950 130.800 631.050 132.900 ;
        RECT 637.950 132.450 640.050 132.900 ;
        RECT 652.950 132.450 655.050 132.900 ;
        RECT 637.950 131.250 655.050 132.450 ;
        RECT 637.950 130.800 640.050 131.250 ;
        RECT 652.950 130.800 655.050 131.250 ;
        RECT 670.950 130.800 673.050 132.900 ;
        RECT 682.950 132.600 685.050 133.050 ;
        RECT 691.950 132.600 694.050 132.900 ;
        RECT 682.950 131.400 694.050 132.600 ;
        RECT 682.950 130.950 685.050 131.400 ;
        RECT 691.950 130.800 694.050 131.400 ;
        RECT 748.950 132.450 751.050 132.900 ;
        RECT 754.950 132.450 757.050 132.900 ;
        RECT 748.950 131.250 757.050 132.450 ;
        RECT 748.950 130.800 751.050 131.250 ;
        RECT 754.950 130.800 757.050 131.250 ;
        RECT 760.950 132.600 763.050 132.900 ;
        RECT 773.400 132.600 774.600 137.100 ;
        RECT 790.950 136.950 793.050 139.050 ;
        RECT 802.950 138.600 805.050 139.200 ;
        RECT 814.950 138.600 817.050 139.050 ;
        RECT 802.950 137.400 817.050 138.600 ;
        RECT 802.950 137.100 805.050 137.400 ;
        RECT 814.950 136.950 817.050 137.400 ;
        RECT 820.950 138.600 823.050 139.200 ;
        RECT 829.950 138.600 832.050 139.050 ;
        RECT 820.950 137.400 832.050 138.600 ;
        RECT 835.950 138.600 838.050 142.050 ;
        RECT 841.950 141.600 844.050 142.050 ;
        RECT 850.950 141.600 853.050 142.050 ;
        RECT 841.950 140.400 853.050 141.600 ;
        RECT 841.950 139.950 844.050 140.400 ;
        RECT 850.950 139.950 853.050 140.400 ;
        RECT 856.950 138.750 859.050 139.200 ;
        RECT 862.950 138.750 865.050 139.200 ;
        RECT 835.950 138.000 840.600 138.600 ;
        RECT 836.400 137.400 840.600 138.000 ;
        RECT 820.950 137.100 823.050 137.400 ;
        RECT 829.950 136.950 832.050 137.400 ;
        RECT 791.400 133.050 792.600 136.950 ;
        RECT 839.400 135.600 840.600 137.400 ;
        RECT 856.950 137.550 865.050 138.750 ;
        RECT 856.950 137.100 859.050 137.550 ;
        RECT 862.950 137.100 865.050 137.550 ;
        RECT 883.950 138.600 886.050 139.200 ;
        RECT 895.950 138.600 898.050 139.050 ;
        RECT 883.950 137.400 898.050 138.600 ;
        RECT 883.950 137.100 886.050 137.400 ;
        RECT 895.950 136.950 898.050 137.400 ;
        RECT 904.950 137.100 907.050 139.200 ;
        RECT 839.400 134.400 846.600 135.600 ;
        RECT 760.950 131.400 774.600 132.600 ;
        RECT 760.950 130.800 763.050 131.400 ;
        RECT 790.950 130.950 793.050 133.050 ;
        RECT 799.950 132.600 802.050 132.900 ;
        RECT 817.950 132.600 820.050 132.900 ;
        RECT 799.950 131.400 820.050 132.600 ;
        RECT 799.950 130.800 802.050 131.400 ;
        RECT 817.950 130.800 820.050 131.400 ;
        RECT 13.950 129.600 16.050 130.050 ;
        RECT 22.950 129.600 25.050 130.050 ;
        RECT 13.950 128.400 25.050 129.600 ;
        RECT 13.950 127.950 16.050 128.400 ;
        RECT 22.950 127.950 25.050 128.400 ;
        RECT 28.950 129.600 31.050 130.050 ;
        RECT 37.950 129.600 40.050 130.050 ;
        RECT 28.950 128.400 40.050 129.600 ;
        RECT 28.950 127.950 31.050 128.400 ;
        RECT 37.950 127.950 40.050 128.400 ;
        RECT 55.950 129.600 58.050 130.050 ;
        RECT 64.950 129.600 67.050 130.050 ;
        RECT 55.950 128.400 67.050 129.600 ;
        RECT 55.950 127.950 58.050 128.400 ;
        RECT 64.950 127.950 67.050 128.400 ;
        RECT 79.950 129.600 82.050 130.050 ;
        RECT 91.950 129.600 94.050 130.050 ;
        RECT 79.950 128.400 94.050 129.600 ;
        RECT 79.950 127.950 82.050 128.400 ;
        RECT 91.950 127.950 94.050 128.400 ;
        RECT 127.950 129.600 130.050 130.050 ;
        RECT 148.950 129.600 151.050 130.050 ;
        RECT 160.950 129.600 163.050 130.050 ;
        RECT 127.950 128.400 163.050 129.600 ;
        RECT 127.950 127.950 130.050 128.400 ;
        RECT 148.950 127.950 151.050 128.400 ;
        RECT 160.950 127.950 163.050 128.400 ;
        RECT 250.950 129.600 253.050 130.050 ;
        RECT 259.950 129.600 262.050 130.050 ;
        RECT 250.950 128.400 262.050 129.600 ;
        RECT 250.950 127.950 253.050 128.400 ;
        RECT 259.950 127.950 262.050 128.400 ;
        RECT 412.950 129.600 415.050 130.050 ;
        RECT 448.950 129.600 451.050 130.050 ;
        RECT 412.950 128.400 451.050 129.600 ;
        RECT 412.950 127.950 415.050 128.400 ;
        RECT 448.950 127.950 451.050 128.400 ;
        RECT 472.950 129.600 475.050 130.050 ;
        RECT 578.400 129.600 579.600 130.800 ;
        RECT 845.400 130.050 846.600 134.400 ;
        RECT 853.950 132.600 856.050 133.050 ;
        RECT 859.950 132.600 862.050 132.900 ;
        RECT 853.950 131.400 862.050 132.600 ;
        RECT 853.950 130.950 856.050 131.400 ;
        RECT 859.950 130.800 862.050 131.400 ;
        RECT 905.400 130.050 906.600 137.100 ;
        RECT 913.950 136.950 916.050 139.050 ;
        RECT 914.400 133.050 915.600 136.950 ;
        RECT 913.950 130.950 916.050 133.050 ;
        RECT 604.950 129.600 607.050 130.050 ;
        RECT 472.950 128.400 495.600 129.600 ;
        RECT 578.400 128.400 607.050 129.600 ;
        RECT 472.950 127.950 475.050 128.400 ;
        RECT 67.950 126.600 70.050 127.050 ;
        RECT 121.950 126.600 124.050 127.050 ;
        RECT 67.950 125.400 124.050 126.600 ;
        RECT 67.950 124.950 70.050 125.400 ;
        RECT 121.950 124.950 124.050 125.400 ;
        RECT 157.950 126.600 160.050 127.050 ;
        RECT 175.950 126.600 178.050 127.050 ;
        RECT 157.950 125.400 178.050 126.600 ;
        RECT 157.950 124.950 160.050 125.400 ;
        RECT 175.950 124.950 178.050 125.400 ;
        RECT 199.950 126.600 202.050 127.050 ;
        RECT 232.950 126.600 235.050 127.050 ;
        RECT 199.950 125.400 235.050 126.600 ;
        RECT 199.950 124.950 202.050 125.400 ;
        RECT 232.950 124.950 235.050 125.400 ;
        RECT 316.950 126.600 319.050 127.050 ;
        RECT 325.950 126.600 328.050 127.050 ;
        RECT 334.950 126.600 337.050 127.050 ;
        RECT 316.950 125.400 337.050 126.600 ;
        RECT 316.950 124.950 319.050 125.400 ;
        RECT 325.950 124.950 328.050 125.400 ;
        RECT 334.950 124.950 337.050 125.400 ;
        RECT 394.950 126.600 397.050 127.050 ;
        RECT 400.950 126.600 403.050 127.050 ;
        RECT 433.950 126.600 436.050 127.050 ;
        RECT 394.950 125.400 436.050 126.600 ;
        RECT 394.950 124.950 397.050 125.400 ;
        RECT 400.950 124.950 403.050 125.400 ;
        RECT 433.950 124.950 436.050 125.400 ;
        RECT 454.950 126.600 457.050 127.050 ;
        RECT 490.950 126.600 493.050 127.050 ;
        RECT 454.950 125.400 493.050 126.600 ;
        RECT 494.400 126.600 495.600 128.400 ;
        RECT 604.950 127.950 607.050 128.400 ;
        RECT 709.950 129.600 712.050 130.050 ;
        RECT 733.950 129.600 736.050 130.050 ;
        RECT 745.950 129.600 748.050 130.050 ;
        RECT 778.950 129.600 781.050 130.050 ;
        RECT 709.950 128.400 748.050 129.600 ;
        RECT 709.950 127.950 712.050 128.400 ;
        RECT 733.950 127.950 736.050 128.400 ;
        RECT 745.950 127.950 748.050 128.400 ;
        RECT 767.400 128.400 781.050 129.600 ;
        RECT 520.950 126.600 523.050 127.050 ;
        RECT 494.400 125.400 523.050 126.600 ;
        RECT 454.950 124.950 457.050 125.400 ;
        RECT 490.950 124.950 493.050 125.400 ;
        RECT 520.950 124.950 523.050 125.400 ;
        RECT 661.950 126.600 664.050 127.050 ;
        RECT 767.400 126.600 768.600 128.400 ;
        RECT 778.950 127.950 781.050 128.400 ;
        RECT 844.950 127.950 847.050 130.050 ;
        RECT 862.950 129.600 865.050 130.050 ;
        RECT 874.950 129.600 877.050 130.050 ;
        RECT 862.950 128.400 877.050 129.600 ;
        RECT 862.950 127.950 865.050 128.400 ;
        RECT 874.950 127.950 877.050 128.400 ;
        RECT 880.950 129.600 883.050 130.050 ;
        RECT 898.950 129.600 901.050 130.050 ;
        RECT 880.950 128.400 901.050 129.600 ;
        RECT 880.950 127.950 883.050 128.400 ;
        RECT 898.950 127.950 901.050 128.400 ;
        RECT 904.950 127.950 907.050 130.050 ;
        RECT 661.950 125.400 768.600 126.600 ;
        RECT 841.950 126.600 844.050 127.050 ;
        RECT 865.950 126.600 868.050 127.050 ;
        RECT 841.950 125.400 868.050 126.600 ;
        RECT 661.950 124.950 664.050 125.400 ;
        RECT 841.950 124.950 844.050 125.400 ;
        RECT 865.950 124.950 868.050 125.400 ;
        RECT 61.950 123.600 64.050 124.050 ;
        RECT 109.950 123.600 112.050 124.050 ;
        RECT 61.950 122.400 112.050 123.600 ;
        RECT 61.950 121.950 64.050 122.400 ;
        RECT 109.950 121.950 112.050 122.400 ;
        RECT 139.950 123.600 142.050 124.050 ;
        RECT 148.950 123.600 151.050 124.050 ;
        RECT 139.950 122.400 151.050 123.600 ;
        RECT 139.950 121.950 142.050 122.400 ;
        RECT 148.950 121.950 151.050 122.400 ;
        RECT 202.950 123.600 205.050 124.050 ;
        RECT 250.950 123.600 253.050 124.050 ;
        RECT 202.950 122.400 253.050 123.600 ;
        RECT 202.950 121.950 205.050 122.400 ;
        RECT 250.950 121.950 253.050 122.400 ;
        RECT 280.950 123.600 283.050 124.050 ;
        RECT 310.950 123.600 313.050 124.050 ;
        RECT 361.950 123.600 364.050 124.050 ;
        RECT 280.950 122.400 364.050 123.600 ;
        RECT 280.950 121.950 283.050 122.400 ;
        RECT 310.950 121.950 313.050 122.400 ;
        RECT 361.950 121.950 364.050 122.400 ;
        RECT 397.950 123.600 400.050 124.050 ;
        RECT 436.950 123.600 439.050 124.050 ;
        RECT 397.950 122.400 439.050 123.600 ;
        RECT 397.950 121.950 400.050 122.400 ;
        RECT 436.950 121.950 439.050 122.400 ;
        RECT 514.950 123.600 517.050 124.050 ;
        RECT 589.950 123.600 592.050 124.050 ;
        RECT 514.950 122.400 592.050 123.600 ;
        RECT 514.950 121.950 517.050 122.400 ;
        RECT 589.950 121.950 592.050 122.400 ;
        RECT 646.950 123.600 649.050 124.050 ;
        RECT 775.950 123.600 778.050 124.050 ;
        RECT 799.950 123.600 802.050 124.050 ;
        RECT 646.950 122.400 802.050 123.600 ;
        RECT 646.950 121.950 649.050 122.400 ;
        RECT 775.950 121.950 778.050 122.400 ;
        RECT 799.950 121.950 802.050 122.400 ;
        RECT 886.950 123.600 889.050 124.050 ;
        RECT 907.950 123.600 910.050 124.050 ;
        RECT 886.950 122.400 910.050 123.600 ;
        RECT 886.950 121.950 889.050 122.400 ;
        RECT 907.950 121.950 910.050 122.400 ;
        RECT 10.950 120.600 13.050 121.050 ;
        RECT 52.950 120.600 55.050 121.050 ;
        RECT 172.950 120.600 175.050 121.050 ;
        RECT 10.950 119.400 175.050 120.600 ;
        RECT 10.950 118.950 13.050 119.400 ;
        RECT 52.950 118.950 55.050 119.400 ;
        RECT 172.950 118.950 175.050 119.400 ;
        RECT 319.950 120.600 322.050 121.050 ;
        RECT 328.950 120.600 331.050 121.050 ;
        RECT 319.950 119.400 331.050 120.600 ;
        RECT 319.950 118.950 322.050 119.400 ;
        RECT 328.950 118.950 331.050 119.400 ;
        RECT 388.950 120.600 391.050 121.050 ;
        RECT 451.950 120.600 454.050 121.050 ;
        RECT 388.950 119.400 454.050 120.600 ;
        RECT 388.950 118.950 391.050 119.400 ;
        RECT 451.950 118.950 454.050 119.400 ;
        RECT 457.950 120.600 460.050 121.050 ;
        RECT 484.950 120.600 487.050 121.050 ;
        RECT 595.950 120.600 598.050 121.050 ;
        RECT 457.950 119.400 598.050 120.600 ;
        RECT 457.950 118.950 460.050 119.400 ;
        RECT 484.950 118.950 487.050 119.400 ;
        RECT 595.950 118.950 598.050 119.400 ;
        RECT 610.950 120.600 613.050 121.050 ;
        RECT 625.950 120.600 628.050 121.050 ;
        RECT 610.950 119.400 628.050 120.600 ;
        RECT 610.950 118.950 613.050 119.400 ;
        RECT 625.950 118.950 628.050 119.400 ;
        RECT 712.950 120.600 715.050 121.050 ;
        RECT 778.950 120.600 781.050 121.050 ;
        RECT 712.950 119.400 750.600 120.600 ;
        RECT 712.950 118.950 715.050 119.400 ;
        RECT 118.950 117.600 121.050 118.050 ;
        RECT 142.950 117.600 145.050 118.050 ;
        RECT 118.950 116.400 145.050 117.600 ;
        RECT 118.950 115.950 121.050 116.400 ;
        RECT 142.950 115.950 145.050 116.400 ;
        RECT 178.950 117.600 181.050 118.050 ;
        RECT 217.950 117.600 220.050 118.050 ;
        RECT 343.950 117.600 346.050 118.050 ;
        RECT 178.950 116.400 346.050 117.600 ;
        RECT 178.950 115.950 181.050 116.400 ;
        RECT 217.950 115.950 220.050 116.400 ;
        RECT 343.950 115.950 346.050 116.400 ;
        RECT 418.950 117.600 421.050 118.050 ;
        RECT 436.950 117.600 439.050 118.050 ;
        RECT 418.950 116.400 439.050 117.600 ;
        RECT 418.950 115.950 421.050 116.400 ;
        RECT 436.950 115.950 439.050 116.400 ;
        RECT 541.950 117.600 544.050 118.050 ;
        RECT 628.950 117.600 631.050 118.050 ;
        RECT 541.950 116.400 631.050 117.600 ;
        RECT 749.400 117.600 750.600 119.400 ;
        RECT 778.950 119.400 798.600 120.600 ;
        RECT 778.950 118.950 781.050 119.400 ;
        RECT 775.950 117.600 778.050 118.050 ;
        RECT 787.950 117.600 790.050 118.050 ;
        RECT 749.400 116.400 790.050 117.600 ;
        RECT 797.400 117.600 798.600 119.400 ;
        RECT 805.950 117.600 808.050 118.050 ;
        RECT 797.400 116.400 808.050 117.600 ;
        RECT 541.950 115.950 544.050 116.400 ;
        RECT 628.950 115.950 631.050 116.400 ;
        RECT 775.950 115.950 778.050 116.400 ;
        RECT 787.950 115.950 790.050 116.400 ;
        RECT 805.950 115.950 808.050 116.400 ;
        RECT 814.950 117.600 817.050 118.050 ;
        RECT 832.950 117.600 835.050 118.050 ;
        RECT 856.950 117.600 859.050 118.050 ;
        RECT 814.950 116.400 859.050 117.600 ;
        RECT 814.950 115.950 817.050 116.400 ;
        RECT 832.950 115.950 835.050 116.400 ;
        RECT 856.950 115.950 859.050 116.400 ;
        RECT 877.950 117.600 880.050 118.050 ;
        RECT 892.950 117.600 895.050 118.050 ;
        RECT 877.950 116.400 895.050 117.600 ;
        RECT 877.950 115.950 880.050 116.400 ;
        RECT 892.950 115.950 895.050 116.400 ;
        RECT 898.950 117.600 901.050 118.050 ;
        RECT 907.950 117.600 910.050 118.050 ;
        RECT 898.950 116.400 910.050 117.600 ;
        RECT 898.950 115.950 901.050 116.400 ;
        RECT 907.950 115.950 910.050 116.400 ;
        RECT 235.950 114.600 238.050 115.050 ;
        RECT 250.950 114.600 253.050 115.050 ;
        RECT 235.950 113.400 253.050 114.600 ;
        RECT 235.950 112.950 238.050 113.400 ;
        RECT 250.950 112.950 253.050 113.400 ;
        RECT 352.950 114.600 355.050 115.050 ;
        RECT 397.950 114.600 400.050 115.050 ;
        RECT 352.950 113.400 400.050 114.600 ;
        RECT 352.950 112.950 355.050 113.400 ;
        RECT 397.950 112.950 400.050 113.400 ;
        RECT 439.950 114.600 442.050 115.050 ;
        RECT 487.950 114.600 490.050 115.050 ;
        RECT 439.950 113.400 490.050 114.600 ;
        RECT 439.950 112.950 442.050 113.400 ;
        RECT 487.950 112.950 490.050 113.400 ;
        RECT 556.950 114.600 559.050 115.050 ;
        RECT 565.950 114.600 568.050 115.050 ;
        RECT 556.950 113.400 568.050 114.600 ;
        RECT 556.950 112.950 559.050 113.400 ;
        RECT 565.950 112.950 568.050 113.400 ;
        RECT 610.950 114.600 613.050 115.050 ;
        RECT 616.950 114.600 619.050 115.050 ;
        RECT 622.950 114.600 625.050 115.050 ;
        RECT 610.950 113.400 625.050 114.600 ;
        RECT 610.950 112.950 613.050 113.400 ;
        RECT 616.950 112.950 619.050 113.400 ;
        RECT 622.950 112.950 625.050 113.400 ;
        RECT 640.950 114.600 643.050 115.050 ;
        RECT 652.950 114.600 655.050 115.050 ;
        RECT 640.950 113.400 655.050 114.600 ;
        RECT 640.950 112.950 643.050 113.400 ;
        RECT 652.950 112.950 655.050 113.400 ;
        RECT 676.950 114.600 679.050 115.050 ;
        RECT 745.950 114.600 748.050 115.050 ;
        RECT 676.950 113.400 748.050 114.600 ;
        RECT 676.950 112.950 679.050 113.400 ;
        RECT 745.950 112.950 748.050 113.400 ;
        RECT 790.950 114.600 793.050 115.050 ;
        RECT 883.950 114.600 886.050 115.050 ;
        RECT 790.950 113.400 886.050 114.600 ;
        RECT 790.950 112.950 793.050 113.400 ;
        RECT 883.950 112.950 886.050 113.400 ;
        RECT 31.950 111.600 34.050 112.050 ;
        RECT 37.950 111.600 40.050 112.050 ;
        RECT 79.950 111.600 82.050 112.050 ;
        RECT 85.950 111.600 88.050 112.050 ;
        RECT 142.950 111.600 145.050 112.050 ;
        RECT 31.950 110.400 145.050 111.600 ;
        RECT 31.950 109.950 34.050 110.400 ;
        RECT 37.950 109.950 40.050 110.400 ;
        RECT 79.950 109.950 82.050 110.400 ;
        RECT 85.950 109.950 88.050 110.400 ;
        RECT 142.950 109.950 145.050 110.400 ;
        RECT 148.950 111.600 151.050 112.050 ;
        RECT 184.950 111.600 187.050 112.050 ;
        RECT 148.950 110.400 187.050 111.600 ;
        RECT 148.950 109.950 151.050 110.400 ;
        RECT 184.950 109.950 187.050 110.400 ;
        RECT 193.950 111.600 196.050 112.050 ;
        RECT 208.950 111.600 211.050 112.050 ;
        RECT 193.950 110.400 211.050 111.600 ;
        RECT 193.950 109.950 196.050 110.400 ;
        RECT 208.950 109.950 211.050 110.400 ;
        RECT 229.950 111.600 232.050 112.050 ;
        RECT 244.950 111.600 247.050 112.050 ;
        RECT 229.950 110.400 247.050 111.600 ;
        RECT 229.950 109.950 232.050 110.400 ;
        RECT 244.950 109.950 247.050 110.400 ;
        RECT 400.950 111.600 403.050 112.050 ;
        RECT 427.950 111.600 430.050 112.050 ;
        RECT 400.950 110.400 430.050 111.600 ;
        RECT 400.950 109.950 403.050 110.400 ;
        RECT 427.950 109.950 430.050 110.400 ;
        RECT 586.950 111.600 589.050 112.050 ;
        RECT 622.950 111.600 625.050 111.900 ;
        RECT 655.950 111.600 658.050 112.050 ;
        RECT 586.950 110.400 658.050 111.600 ;
        RECT 586.950 109.950 589.050 110.400 ;
        RECT 622.950 109.800 625.050 110.400 ;
        RECT 655.950 109.950 658.050 110.400 ;
        RECT 700.950 111.600 703.050 112.050 ;
        RECT 739.950 111.600 742.050 112.050 ;
        RECT 700.950 110.400 742.050 111.600 ;
        RECT 700.950 109.950 703.050 110.400 ;
        RECT 739.950 109.950 742.050 110.400 ;
        RECT 865.950 111.600 868.050 112.050 ;
        RECT 880.950 111.600 883.050 112.050 ;
        RECT 865.950 110.400 883.050 111.600 ;
        RECT 865.950 109.950 868.050 110.400 ;
        RECT 880.950 109.950 883.050 110.400 ;
        RECT 889.950 111.600 892.050 112.050 ;
        RECT 895.950 111.600 898.050 112.050 ;
        RECT 889.950 110.400 898.050 111.600 ;
        RECT 889.950 109.950 892.050 110.400 ;
        RECT 895.950 109.950 898.050 110.400 ;
        RECT 247.950 108.600 250.050 109.050 ;
        RECT 259.950 108.600 262.050 109.050 ;
        RECT 247.950 107.400 262.050 108.600 ;
        RECT 247.950 106.950 250.050 107.400 ;
        RECT 259.950 106.950 262.050 107.400 ;
        RECT 283.950 108.600 286.050 109.050 ;
        RECT 292.950 108.600 295.050 109.050 ;
        RECT 283.950 107.400 295.050 108.600 ;
        RECT 283.950 106.950 286.050 107.400 ;
        RECT 292.950 106.950 295.050 107.400 ;
        RECT 388.950 108.600 391.050 109.050 ;
        RECT 448.950 108.600 451.050 109.050 ;
        RECT 472.950 108.600 475.050 109.050 ;
        RECT 481.950 108.600 484.050 109.050 ;
        RECT 388.950 107.400 405.600 108.600 ;
        RECT 388.950 106.950 391.050 107.400 ;
        RECT 1.950 105.750 4.050 106.200 ;
        RECT 10.950 105.750 13.050 106.200 ;
        RECT 1.950 104.550 13.050 105.750 ;
        RECT 1.950 104.100 4.050 104.550 ;
        RECT 10.950 104.100 13.050 104.550 ;
        RECT 43.950 105.750 46.050 106.200 ;
        RECT 52.950 105.750 55.050 106.200 ;
        RECT 43.950 104.550 55.050 105.750 ;
        RECT 43.950 104.100 46.050 104.550 ;
        RECT 52.950 104.100 55.050 104.550 ;
        RECT 61.950 105.600 64.050 106.200 ;
        RECT 67.950 105.750 70.050 106.200 ;
        RECT 73.950 105.750 76.050 106.200 ;
        RECT 61.950 104.400 66.600 105.600 ;
        RECT 61.950 104.100 64.050 104.400 ;
        RECT 22.950 99.450 25.050 99.900 ;
        RECT 28.950 99.450 31.050 99.900 ;
        RECT 22.950 98.250 31.050 99.450 ;
        RECT 22.950 97.800 25.050 98.250 ;
        RECT 28.950 97.800 31.050 98.250 ;
        RECT 65.400 96.600 66.600 104.400 ;
        RECT 67.950 104.550 76.050 105.750 ;
        RECT 67.950 104.100 70.050 104.550 ;
        RECT 73.950 104.100 76.050 104.550 ;
        RECT 103.950 105.600 106.050 106.200 ;
        RECT 115.950 105.600 118.050 106.050 ;
        RECT 121.950 105.600 124.050 106.200 ;
        RECT 103.950 104.400 124.050 105.600 ;
        RECT 103.950 104.100 106.050 104.400 ;
        RECT 115.950 103.950 118.050 104.400 ;
        RECT 121.950 104.100 124.050 104.400 ;
        RECT 130.950 105.600 133.050 106.050 ;
        RECT 136.950 105.600 139.050 106.050 ;
        RECT 130.950 104.400 139.050 105.600 ;
        RECT 130.950 103.950 133.050 104.400 ;
        RECT 136.950 103.950 139.050 104.400 ;
        RECT 154.950 105.750 157.050 106.200 ;
        RECT 163.950 105.750 166.050 106.200 ;
        RECT 154.950 104.550 166.050 105.750 ;
        RECT 154.950 104.100 157.050 104.550 ;
        RECT 163.950 104.100 166.050 104.550 ;
        RECT 169.950 104.100 172.050 106.200 ;
        RECT 175.950 105.600 178.050 106.050 ;
        RECT 202.950 105.600 205.050 106.200 ;
        RECT 175.950 104.400 205.050 105.600 ;
        RECT 170.400 102.600 171.600 104.100 ;
        RECT 175.950 103.950 178.050 104.400 ;
        RECT 202.950 104.100 205.050 104.400 ;
        RECT 226.950 105.600 229.050 106.200 ;
        RECT 238.950 105.600 241.050 106.050 ;
        RECT 255.000 105.600 259.050 106.050 ;
        RECT 226.950 104.400 241.050 105.600 ;
        RECT 226.950 104.100 229.050 104.400 ;
        RECT 238.950 103.950 241.050 104.400 ;
        RECT 254.400 103.950 259.050 105.600 ;
        RECT 274.950 105.600 277.050 106.050 ;
        RECT 304.950 105.600 307.050 106.200 ;
        RECT 274.950 104.400 307.050 105.600 ;
        RECT 274.950 103.950 277.050 104.400 ;
        RECT 304.950 104.100 307.050 104.400 ;
        RECT 310.950 105.750 313.050 106.200 ;
        RECT 316.950 105.750 319.050 106.200 ;
        RECT 310.950 104.550 319.050 105.750 ;
        RECT 310.950 104.100 313.050 104.550 ;
        RECT 316.950 104.100 319.050 104.550 ;
        RECT 337.950 105.750 340.050 106.200 ;
        RECT 343.950 105.750 346.050 106.200 ;
        RECT 337.950 104.550 346.050 105.750 ;
        RECT 337.950 104.100 340.050 104.550 ;
        RECT 343.950 104.100 346.050 104.550 ;
        RECT 370.950 105.600 373.050 105.900 ;
        RECT 379.950 105.600 382.050 106.200 ;
        RECT 384.000 105.600 388.050 106.050 ;
        RECT 370.950 104.400 382.050 105.600 ;
        RECT 170.400 101.400 198.600 102.600 ;
        RECT 76.950 99.600 79.050 99.900 ;
        RECT 94.950 99.600 97.050 99.900 ;
        RECT 76.950 98.400 97.050 99.600 ;
        RECT 76.950 97.800 79.050 98.400 ;
        RECT 94.950 97.800 97.050 98.400 ;
        RECT 172.950 99.450 175.050 99.900 ;
        RECT 178.950 99.450 181.050 99.900 ;
        RECT 172.950 98.250 181.050 99.450 ;
        RECT 172.950 97.800 175.050 98.250 ;
        RECT 178.950 97.800 181.050 98.250 ;
        RECT 187.950 99.600 190.050 99.900 ;
        RECT 193.950 99.600 196.050 100.050 ;
        RECT 187.950 98.400 196.050 99.600 ;
        RECT 197.400 99.600 198.600 101.400 ;
        RECT 254.400 99.900 255.600 103.950 ;
        RECT 370.950 103.800 373.050 104.400 ;
        RECT 379.950 104.100 382.050 104.400 ;
        RECT 383.400 103.950 388.050 105.600 ;
        RECT 391.950 105.750 394.050 106.200 ;
        RECT 400.950 105.750 403.050 106.200 ;
        RECT 391.950 104.550 403.050 105.750 ;
        RECT 391.950 104.100 394.050 104.550 ;
        RECT 400.950 104.100 403.050 104.550 ;
        RECT 404.400 105.600 405.600 107.400 ;
        RECT 448.950 107.400 484.050 108.600 ;
        RECT 448.950 106.950 451.050 107.400 ;
        RECT 472.950 106.950 475.050 107.400 ;
        RECT 481.950 106.950 484.050 107.400 ;
        RECT 487.950 108.600 492.000 109.050 ;
        RECT 544.950 108.600 547.050 109.050 ;
        RECT 559.950 108.600 562.050 109.050 ;
        RECT 631.950 108.600 634.050 109.050 ;
        RECT 487.950 106.950 492.600 108.600 ;
        RECT 544.950 107.400 634.050 108.600 ;
        RECT 544.950 106.950 547.050 107.400 ;
        RECT 559.950 106.950 562.050 107.400 ;
        RECT 421.950 105.600 424.050 106.200 ;
        RECT 442.950 105.600 445.050 106.200 ;
        RECT 404.400 104.400 445.050 105.600 ;
        RECT 421.950 104.100 424.050 104.400 ;
        RECT 442.950 104.100 445.050 104.400 ;
        RECT 460.950 105.600 463.050 106.050 ;
        RECT 466.950 105.600 469.050 106.200 ;
        RECT 460.950 104.400 469.050 105.600 ;
        RECT 460.950 103.950 463.050 104.400 ;
        RECT 466.950 104.100 469.050 104.400 ;
        RECT 484.950 105.600 489.000 106.050 ;
        RECT 484.950 103.950 489.600 105.600 ;
        RECT 211.950 99.600 214.050 99.900 ;
        RECT 197.400 98.400 214.050 99.600 ;
        RECT 187.950 97.800 190.050 98.400 ;
        RECT 193.950 97.950 196.050 98.400 ;
        RECT 211.950 97.800 214.050 98.400 ;
        RECT 217.950 99.450 220.050 99.900 ;
        RECT 223.950 99.450 226.050 99.900 ;
        RECT 217.950 98.250 226.050 99.450 ;
        RECT 217.950 97.800 220.050 98.250 ;
        RECT 223.950 97.800 226.050 98.250 ;
        RECT 253.950 97.800 256.050 99.900 ;
        RECT 307.950 99.450 310.050 99.900 ;
        RECT 319.950 99.450 322.050 99.900 ;
        RECT 307.950 98.250 322.050 99.450 ;
        RECT 307.950 97.800 310.050 98.250 ;
        RECT 319.950 97.800 322.050 98.250 ;
        RECT 346.950 99.600 349.050 99.900 ;
        RECT 355.950 99.600 358.050 100.050 ;
        RECT 383.400 99.900 384.600 103.950 ;
        RECT 409.950 102.600 412.050 103.050 ;
        RECT 409.950 101.400 432.600 102.600 ;
        RECT 409.950 100.950 412.050 101.400 ;
        RECT 431.400 99.900 432.600 101.400 ;
        RECT 488.400 99.900 489.600 103.950 ;
        RECT 491.400 102.600 492.600 106.950 ;
        RECT 502.950 105.750 505.050 106.200 ;
        RECT 508.950 105.750 511.050 106.200 ;
        RECT 502.950 104.550 511.050 105.750 ;
        RECT 502.950 104.100 505.050 104.550 ;
        RECT 508.950 104.100 511.050 104.550 ;
        RECT 517.950 103.950 520.050 106.050 ;
        RECT 544.950 105.600 547.050 105.900 ;
        RECT 553.950 105.600 556.050 106.200 ;
        RECT 544.950 104.400 556.050 105.600 ;
        RECT 491.400 101.400 498.600 102.600 ;
        RECT 346.950 98.400 358.050 99.600 ;
        RECT 346.950 97.800 349.050 98.400 ;
        RECT 355.950 97.950 358.050 98.400 ;
        RECT 361.950 99.600 364.050 99.900 ;
        RECT 376.950 99.600 379.050 99.900 ;
        RECT 361.950 98.400 379.050 99.600 ;
        RECT 361.950 97.800 364.050 98.400 ;
        RECT 376.950 97.800 379.050 98.400 ;
        RECT 382.950 97.800 385.050 99.900 ;
        RECT 430.950 97.800 433.050 99.900 ;
        RECT 451.950 99.450 454.050 99.900 ;
        RECT 457.950 99.450 460.050 99.900 ;
        RECT 451.950 98.250 460.050 99.450 ;
        RECT 451.950 97.800 454.050 98.250 ;
        RECT 457.950 97.800 460.050 98.250 ;
        RECT 475.950 99.600 478.050 99.900 ;
        RECT 487.950 99.600 490.050 99.900 ;
        RECT 475.950 98.400 490.050 99.600 ;
        RECT 497.400 99.600 498.600 101.400 ;
        RECT 518.400 100.050 519.600 103.950 ;
        RECT 544.950 103.800 547.050 104.400 ;
        RECT 553.950 104.100 556.050 104.400 ;
        RECT 562.950 105.750 565.050 106.200 ;
        RECT 568.950 105.750 571.050 106.050 ;
        RECT 574.950 105.750 577.050 106.200 ;
        RECT 562.950 104.550 577.050 105.750 ;
        RECT 562.950 104.100 565.050 104.550 ;
        RECT 568.950 103.950 571.050 104.550 ;
        RECT 574.950 104.100 577.050 104.550 ;
        RECT 580.950 104.100 583.050 106.200 ;
        RECT 511.950 99.600 514.050 99.900 ;
        RECT 497.400 98.400 514.050 99.600 ;
        RECT 475.950 97.800 478.050 98.400 ;
        RECT 487.950 97.800 490.050 98.400 ;
        RECT 511.950 97.800 514.050 98.400 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 535.950 99.450 538.050 99.900 ;
        RECT 541.950 99.450 544.050 99.900 ;
        RECT 535.950 98.250 544.050 99.450 ;
        RECT 535.950 97.800 538.050 98.250 ;
        RECT 541.950 97.800 544.050 98.250 ;
        RECT 88.950 96.600 91.050 97.050 ;
        RECT 118.950 96.600 121.050 97.050 ;
        RECT 139.950 96.600 142.050 97.050 ;
        RECT 154.950 96.600 157.050 97.050 ;
        RECT 65.400 95.400 157.050 96.600 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 118.950 94.950 121.050 95.400 ;
        RECT 139.950 94.950 142.050 95.400 ;
        RECT 154.950 94.950 157.050 95.400 ;
        RECT 247.950 96.600 250.050 97.050 ;
        RECT 265.950 96.600 268.050 97.050 ;
        RECT 247.950 95.400 268.050 96.600 ;
        RECT 247.950 94.950 250.050 95.400 ;
        RECT 265.950 94.950 268.050 95.400 ;
        RECT 280.950 96.600 283.050 97.050 ;
        RECT 295.950 96.600 298.050 97.050 ;
        RECT 325.950 96.600 328.050 97.050 ;
        RECT 280.950 95.400 328.050 96.600 ;
        RECT 280.950 94.950 283.050 95.400 ;
        RECT 295.950 94.950 298.050 95.400 ;
        RECT 325.950 94.950 328.050 95.400 ;
        RECT 412.950 96.600 415.050 97.050 ;
        RECT 445.950 96.600 448.050 97.050 ;
        RECT 469.950 96.600 472.050 97.050 ;
        RECT 412.950 95.400 472.050 96.600 ;
        RECT 412.950 94.950 415.050 95.400 ;
        RECT 445.950 94.950 448.050 95.400 ;
        RECT 469.950 94.950 472.050 95.400 ;
        RECT 550.950 96.600 553.050 97.050 ;
        RECT 565.950 96.600 568.050 97.050 ;
        RECT 550.950 95.400 568.050 96.600 ;
        RECT 550.950 94.950 553.050 95.400 ;
        RECT 565.950 94.950 568.050 95.400 ;
        RECT 58.950 93.600 61.050 94.050 ;
        RECT 67.950 93.600 70.050 94.050 ;
        RECT 58.950 92.400 70.050 93.600 ;
        RECT 58.950 91.950 61.050 92.400 ;
        RECT 67.950 91.950 70.050 92.400 ;
        RECT 109.950 93.600 112.050 94.050 ;
        RECT 166.950 93.600 169.050 94.050 ;
        RECT 109.950 92.400 169.050 93.600 ;
        RECT 109.950 91.950 112.050 92.400 ;
        RECT 166.950 91.950 169.050 92.400 ;
        RECT 319.950 93.600 322.050 94.050 ;
        RECT 331.950 93.600 334.050 94.050 ;
        RECT 319.950 92.400 334.050 93.600 ;
        RECT 319.950 91.950 322.050 92.400 ;
        RECT 331.950 91.950 334.050 92.400 ;
        RECT 370.950 93.600 373.050 94.050 ;
        RECT 418.950 93.600 421.050 94.050 ;
        RECT 370.950 92.400 421.050 93.600 ;
        RECT 370.950 91.950 373.050 92.400 ;
        RECT 418.950 91.950 421.050 92.400 ;
        RECT 520.950 93.600 523.050 94.050 ;
        RECT 529.950 93.600 532.050 94.050 ;
        RECT 541.950 93.600 544.050 94.050 ;
        RECT 520.950 92.400 544.050 93.600 ;
        RECT 581.400 93.600 582.600 104.100 ;
        RECT 584.400 99.900 585.600 107.400 ;
        RECT 631.950 106.950 634.050 107.400 ;
        RECT 646.950 108.600 649.050 109.050 ;
        RECT 652.950 108.600 655.050 109.050 ;
        RECT 646.950 107.400 655.050 108.600 ;
        RECT 646.950 106.950 649.050 107.400 ;
        RECT 652.950 106.950 655.050 107.400 ;
        RECT 760.950 108.600 763.050 109.050 ;
        RECT 766.950 108.600 769.050 109.050 ;
        RECT 760.950 107.400 769.050 108.600 ;
        RECT 760.950 106.950 763.050 107.400 ;
        RECT 766.950 106.950 769.050 107.400 ;
        RECT 808.950 108.600 811.050 109.050 ;
        RECT 823.950 108.600 826.050 109.050 ;
        RECT 829.950 108.600 832.050 109.050 ;
        RECT 808.950 107.400 819.600 108.600 ;
        RECT 808.950 106.950 811.050 107.400 ;
        RECT 586.950 105.600 589.050 106.050 ;
        RECT 598.950 105.600 601.050 106.200 ;
        RECT 607.950 105.600 610.050 106.050 ;
        RECT 586.950 104.400 597.600 105.600 ;
        RECT 586.950 103.950 589.050 104.400 ;
        RECT 596.400 99.900 597.600 104.400 ;
        RECT 598.950 104.400 610.050 105.600 ;
        RECT 598.950 104.100 601.050 104.400 ;
        RECT 607.950 103.950 610.050 104.400 ;
        RECT 655.950 105.600 660.000 106.050 ;
        RECT 673.950 105.600 676.050 106.050 ;
        RECT 682.950 105.600 685.050 106.200 ;
        RECT 655.950 103.950 660.600 105.600 ;
        RECT 673.950 104.400 685.050 105.600 ;
        RECT 673.950 103.950 676.050 104.400 ;
        RECT 682.950 104.100 685.050 104.400 ;
        RECT 688.950 105.750 691.050 106.200 ;
        RECT 697.950 105.750 700.050 106.200 ;
        RECT 688.950 104.550 700.050 105.750 ;
        RECT 688.950 104.100 691.050 104.550 ;
        RECT 697.950 104.100 700.050 104.550 ;
        RECT 706.950 104.100 709.050 106.200 ;
        RECT 659.400 99.900 660.600 103.950 ;
        RECT 707.400 102.600 708.600 104.100 ;
        RECT 718.950 103.950 721.050 106.050 ;
        RECT 730.950 104.100 733.050 106.200 ;
        RECT 751.950 105.600 754.050 106.200 ;
        RECT 769.950 105.600 772.050 106.200 ;
        RECT 790.950 105.600 793.050 106.200 ;
        RECT 751.950 104.400 793.050 105.600 ;
        RECT 751.950 104.100 754.050 104.400 ;
        RECT 769.950 104.100 772.050 104.400 ;
        RECT 790.950 104.100 793.050 104.400 ;
        RECT 695.400 101.400 708.600 102.600 ;
        RECT 583.950 97.800 586.050 99.900 ;
        RECT 595.950 97.800 598.050 99.900 ;
        RECT 601.950 99.450 604.050 99.900 ;
        RECT 610.950 99.450 613.050 99.900 ;
        RECT 601.950 98.250 613.050 99.450 ;
        RECT 601.950 97.800 604.050 98.250 ;
        RECT 610.950 97.800 613.050 98.250 ;
        RECT 631.950 99.450 634.050 99.900 ;
        RECT 643.950 99.450 646.050 99.900 ;
        RECT 631.950 98.250 646.050 99.450 ;
        RECT 631.950 97.800 634.050 98.250 ;
        RECT 643.950 97.800 646.050 98.250 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 676.950 99.450 679.050 99.900 ;
        RECT 685.950 99.450 688.050 99.900 ;
        RECT 676.950 98.250 688.050 99.450 ;
        RECT 676.950 97.800 679.050 98.250 ;
        RECT 685.950 97.800 688.050 98.250 ;
        RECT 691.950 99.600 694.050 99.900 ;
        RECT 695.400 99.600 696.600 101.400 ;
        RECT 719.400 100.050 720.600 103.950 ;
        RECT 691.950 98.400 696.600 99.600 ;
        RECT 691.950 97.800 694.050 98.400 ;
        RECT 718.950 97.950 721.050 100.050 ;
        RECT 715.950 96.600 718.050 97.050 ;
        RECT 731.400 96.600 732.600 104.100 ;
        RECT 799.950 103.950 802.050 106.050 ;
        RECT 800.400 100.050 801.600 103.950 ;
        RECT 733.950 99.600 736.050 99.900 ;
        RECT 748.950 99.600 751.050 99.900 ;
        RECT 733.950 98.400 751.050 99.600 ;
        RECT 733.950 97.800 736.050 98.400 ;
        RECT 748.950 97.800 751.050 98.400 ;
        RECT 754.950 99.600 757.050 99.900 ;
        RECT 760.950 99.600 763.050 99.900 ;
        RECT 754.950 99.450 763.050 99.600 ;
        RECT 766.950 99.600 769.050 99.900 ;
        RECT 793.950 99.600 796.050 99.900 ;
        RECT 766.950 99.450 796.050 99.600 ;
        RECT 754.950 98.400 796.050 99.450 ;
        RECT 754.950 97.800 757.050 98.400 ;
        RECT 760.950 98.250 769.050 98.400 ;
        RECT 760.950 97.800 763.050 98.250 ;
        RECT 766.950 97.800 769.050 98.250 ;
        RECT 793.950 97.800 796.050 98.400 ;
        RECT 799.950 97.950 802.050 100.050 ;
        RECT 818.400 99.900 819.600 107.400 ;
        RECT 823.950 107.400 832.050 108.600 ;
        RECT 823.950 106.950 826.050 107.400 ;
        RECT 829.950 106.950 832.050 107.400 ;
        RECT 826.950 102.600 829.050 106.050 ;
        RECT 838.950 105.600 841.050 106.200 ;
        RECT 868.950 105.600 871.050 106.050 ;
        RECT 888.000 105.600 891.900 106.050 ;
        RECT 838.950 104.400 871.050 105.600 ;
        RECT 838.950 104.100 841.050 104.400 ;
        RECT 868.950 103.950 871.050 104.400 ;
        RECT 887.400 103.950 891.900 105.600 ;
        RECT 892.950 105.750 895.050 106.200 ;
        RECT 901.950 105.750 904.050 106.200 ;
        RECT 892.950 104.550 904.050 105.750 ;
        RECT 904.950 105.600 907.050 109.050 ;
        RECT 904.950 105.000 912.600 105.600 ;
        RECT 892.950 104.100 895.050 104.550 ;
        RECT 901.950 104.100 904.050 104.550 ;
        RECT 905.400 104.400 912.600 105.000 ;
        RECT 826.950 102.000 831.600 102.600 ;
        RECT 827.400 101.400 831.600 102.000 ;
        RECT 830.400 99.900 831.600 101.400 ;
        RECT 887.400 99.900 888.600 103.950 ;
        RECT 911.400 99.900 912.600 104.400 ;
        RECT 817.950 97.800 820.050 99.900 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 835.950 99.600 838.050 99.900 ;
        RECT 853.950 99.600 856.050 99.900 ;
        RECT 835.950 98.400 856.050 99.600 ;
        RECT 835.950 97.800 838.050 98.400 ;
        RECT 853.950 97.800 856.050 98.400 ;
        RECT 868.950 99.450 871.050 99.900 ;
        RECT 880.950 99.450 883.050 99.900 ;
        RECT 868.950 98.250 883.050 99.450 ;
        RECT 868.950 97.800 871.050 98.250 ;
        RECT 880.950 97.800 883.050 98.250 ;
        RECT 886.950 97.800 889.050 99.900 ;
        RECT 910.950 97.800 913.050 99.900 ;
        RECT 772.950 96.600 775.050 97.050 ;
        RECT 787.950 96.600 790.050 97.050 ;
        RECT 895.950 96.600 898.050 96.900 ;
        RECT 715.950 95.400 898.050 96.600 ;
        RECT 715.950 94.950 718.050 95.400 ;
        RECT 772.950 94.950 775.050 95.400 ;
        RECT 787.950 94.950 790.050 95.400 ;
        RECT 895.950 94.800 898.050 95.400 ;
        RECT 901.950 96.600 904.050 97.050 ;
        RECT 910.950 96.600 913.050 97.050 ;
        RECT 901.950 95.400 913.050 96.600 ;
        RECT 901.950 94.950 904.050 95.400 ;
        RECT 910.950 94.950 913.050 95.400 ;
        RECT 601.950 93.600 604.050 94.050 ;
        RECT 581.400 92.400 604.050 93.600 ;
        RECT 520.950 91.950 523.050 92.400 ;
        RECT 529.950 91.950 532.050 92.400 ;
        RECT 541.950 91.950 544.050 92.400 ;
        RECT 601.950 91.950 604.050 92.400 ;
        RECT 628.950 93.600 631.050 94.050 ;
        RECT 673.950 93.600 676.050 94.050 ;
        RECT 628.950 92.400 676.050 93.600 ;
        RECT 628.950 91.950 631.050 92.400 ;
        RECT 673.950 91.950 676.050 92.400 ;
        RECT 679.950 93.600 682.050 94.050 ;
        RECT 709.950 93.600 712.050 94.050 ;
        RECT 679.950 92.400 712.050 93.600 ;
        RECT 679.950 91.950 682.050 92.400 ;
        RECT 709.950 91.950 712.050 92.400 ;
        RECT 844.950 93.600 847.050 94.050 ;
        RECT 874.950 93.600 877.050 94.050 ;
        RECT 844.950 92.400 877.050 93.600 ;
        RECT 844.950 91.950 847.050 92.400 ;
        RECT 874.950 91.950 877.050 92.400 ;
        RECT 880.950 93.600 883.050 94.050 ;
        RECT 892.950 93.600 895.050 94.050 ;
        RECT 880.950 92.400 895.050 93.600 ;
        RECT 880.950 91.950 883.050 92.400 ;
        RECT 892.950 91.950 895.050 92.400 ;
        RECT 145.950 90.600 148.050 91.050 ;
        RECT 151.950 90.600 154.050 91.050 ;
        RECT 160.950 90.600 163.050 91.050 ;
        RECT 145.950 89.400 163.050 90.600 ;
        RECT 145.950 88.950 148.050 89.400 ;
        RECT 151.950 88.950 154.050 89.400 ;
        RECT 160.950 88.950 163.050 89.400 ;
        RECT 271.950 90.600 274.050 91.050 ;
        RECT 352.950 90.600 355.050 91.050 ;
        RECT 271.950 89.400 355.050 90.600 ;
        RECT 271.950 88.950 274.050 89.400 ;
        RECT 352.950 88.950 355.050 89.400 ;
        RECT 481.950 90.600 484.050 91.050 ;
        RECT 493.950 90.600 496.050 91.050 ;
        RECT 481.950 89.400 496.050 90.600 ;
        RECT 481.950 88.950 484.050 89.400 ;
        RECT 493.950 88.950 496.050 89.400 ;
        RECT 664.950 90.600 667.050 91.050 ;
        RECT 724.950 90.600 727.050 91.050 ;
        RECT 808.950 90.600 811.050 91.050 ;
        RECT 811.950 90.600 814.050 91.050 ;
        RECT 838.950 90.600 841.050 91.050 ;
        RECT 664.950 89.400 841.050 90.600 ;
        RECT 664.950 88.950 667.050 89.400 ;
        RECT 724.950 88.950 727.050 89.400 ;
        RECT 808.950 88.950 811.050 89.400 ;
        RECT 811.950 88.950 814.050 89.400 ;
        RECT 838.950 88.950 841.050 89.400 ;
        RECT 100.950 87.600 103.050 88.050 ;
        RECT 238.950 87.600 241.050 88.050 ;
        RECT 100.950 86.400 241.050 87.600 ;
        RECT 100.950 85.950 103.050 86.400 ;
        RECT 238.950 85.950 241.050 86.400 ;
        RECT 346.950 87.600 349.050 88.050 ;
        RECT 388.950 87.600 391.050 88.050 ;
        RECT 346.950 86.400 391.050 87.600 ;
        RECT 346.950 85.950 349.050 86.400 ;
        RECT 388.950 85.950 391.050 86.400 ;
        RECT 526.950 87.600 529.050 88.050 ;
        RECT 577.950 87.600 580.050 88.050 ;
        RECT 619.950 87.600 622.050 88.050 ;
        RECT 526.950 86.400 622.050 87.600 ;
        RECT 526.950 85.950 529.050 86.400 ;
        RECT 577.950 85.950 580.050 86.400 ;
        RECT 619.950 85.950 622.050 86.400 ;
        RECT 673.950 87.600 676.050 88.050 ;
        RECT 691.950 87.600 694.050 88.050 ;
        RECT 673.950 86.400 694.050 87.600 ;
        RECT 673.950 85.950 676.050 86.400 ;
        RECT 691.950 85.950 694.050 86.400 ;
        RECT 829.950 87.600 832.050 88.050 ;
        RECT 859.950 87.600 862.050 88.050 ;
        RECT 829.950 86.400 862.050 87.600 ;
        RECT 829.950 85.950 832.050 86.400 ;
        RECT 859.950 85.950 862.050 86.400 ;
        RECT 868.950 87.600 871.050 88.050 ;
        RECT 904.950 87.600 907.050 88.050 ;
        RECT 868.950 86.400 907.050 87.600 ;
        RECT 868.950 85.950 871.050 86.400 ;
        RECT 904.950 85.950 907.050 86.400 ;
        RECT 331.950 84.600 334.050 85.050 ;
        RECT 415.950 84.600 418.050 85.050 ;
        RECT 460.950 84.600 463.050 85.050 ;
        RECT 331.950 83.400 463.050 84.600 ;
        RECT 331.950 82.950 334.050 83.400 ;
        RECT 415.950 82.950 418.050 83.400 ;
        RECT 460.950 82.950 463.050 83.400 ;
        RECT 697.950 84.600 700.050 85.050 ;
        RECT 703.950 84.600 706.050 85.050 ;
        RECT 697.950 83.400 706.050 84.600 ;
        RECT 697.950 82.950 700.050 83.400 ;
        RECT 703.950 82.950 706.050 83.400 ;
        RECT 589.950 81.600 592.050 82.050 ;
        RECT 679.950 81.600 682.050 82.050 ;
        RECT 589.950 80.400 682.050 81.600 ;
        RECT 589.950 79.950 592.050 80.400 ;
        RECT 679.950 79.950 682.050 80.400 ;
        RECT 847.950 81.600 850.050 82.050 ;
        RECT 856.950 81.600 859.050 82.050 ;
        RECT 847.950 80.400 859.050 81.600 ;
        RECT 847.950 79.950 850.050 80.400 ;
        RECT 856.950 79.950 859.050 80.400 ;
        RECT 211.950 78.600 214.050 79.050 ;
        RECT 229.950 78.600 232.050 79.050 ;
        RECT 274.950 78.600 277.050 79.050 ;
        RECT 211.950 77.400 277.050 78.600 ;
        RECT 211.950 76.950 214.050 77.400 ;
        RECT 229.950 76.950 232.050 77.400 ;
        RECT 274.950 76.950 277.050 77.400 ;
        RECT 376.950 78.600 379.050 79.050 ;
        RECT 400.950 78.600 403.050 79.050 ;
        RECT 439.950 78.600 442.050 79.050 ;
        RECT 544.950 78.600 547.050 79.050 ;
        RECT 376.950 77.400 547.050 78.600 ;
        RECT 376.950 76.950 379.050 77.400 ;
        RECT 400.950 76.950 403.050 77.400 ;
        RECT 439.950 76.950 442.050 77.400 ;
        RECT 544.950 76.950 547.050 77.400 ;
        RECT 688.950 78.600 691.050 79.050 ;
        RECT 796.950 78.600 799.050 79.050 ;
        RECT 688.950 77.400 799.050 78.600 ;
        RECT 688.950 76.950 691.050 77.400 ;
        RECT 796.950 76.950 799.050 77.400 ;
        RECT 1.950 75.600 4.050 76.050 ;
        RECT 37.950 75.600 40.050 76.050 ;
        RECT 148.950 75.600 151.050 76.050 ;
        RECT 196.950 75.600 199.050 76.050 ;
        RECT 1.950 74.400 199.050 75.600 ;
        RECT 1.950 73.950 4.050 74.400 ;
        RECT 37.950 73.950 40.050 74.400 ;
        RECT 148.950 73.950 151.050 74.400 ;
        RECT 196.950 73.950 199.050 74.400 ;
        RECT 586.950 75.600 589.050 76.050 ;
        RECT 607.950 75.600 610.050 76.050 ;
        RECT 586.950 74.400 610.050 75.600 ;
        RECT 586.950 73.950 589.050 74.400 ;
        RECT 607.950 73.950 610.050 74.400 ;
        RECT 640.950 75.600 643.050 76.050 ;
        RECT 655.950 75.600 658.050 76.050 ;
        RECT 853.950 75.600 856.050 76.050 ;
        RECT 640.950 74.400 856.050 75.600 ;
        RECT 640.950 73.950 643.050 74.400 ;
        RECT 655.950 73.950 658.050 74.400 ;
        RECT 853.950 73.950 856.050 74.400 ;
        RECT 871.950 75.600 874.050 76.050 ;
        RECT 877.950 75.600 880.050 76.050 ;
        RECT 871.950 74.400 880.050 75.600 ;
        RECT 871.950 73.950 874.050 74.400 ;
        RECT 877.950 73.950 880.050 74.400 ;
        RECT 340.950 72.600 343.050 73.050 ;
        RECT 355.950 72.600 358.050 73.050 ;
        RECT 397.950 72.600 400.050 73.050 ;
        RECT 340.950 71.400 400.050 72.600 ;
        RECT 340.950 70.950 343.050 71.400 ;
        RECT 355.950 70.950 358.050 71.400 ;
        RECT 397.950 70.950 400.050 71.400 ;
        RECT 739.950 72.600 742.050 73.050 ;
        RECT 751.950 72.600 754.050 73.050 ;
        RECT 757.950 72.600 760.050 73.050 ;
        RECT 739.950 71.400 760.050 72.600 ;
        RECT 739.950 70.950 742.050 71.400 ;
        RECT 751.950 70.950 754.050 71.400 ;
        RECT 757.950 70.950 760.050 71.400 ;
        RECT 775.950 72.600 778.050 73.050 ;
        RECT 835.950 72.600 838.050 73.050 ;
        RECT 775.950 71.400 838.050 72.600 ;
        RECT 775.950 70.950 778.050 71.400 ;
        RECT 835.950 70.950 838.050 71.400 ;
        RECT 847.950 72.600 850.050 73.050 ;
        RECT 874.950 72.600 877.050 72.900 ;
        RECT 847.950 71.400 877.050 72.600 ;
        RECT 847.950 70.950 850.050 71.400 ;
        RECT 874.950 70.800 877.050 71.400 ;
        RECT 100.950 69.600 103.050 70.050 ;
        RECT 127.950 69.600 130.050 70.050 ;
        RECT 100.950 68.400 130.050 69.600 ;
        RECT 100.950 67.950 103.050 68.400 ;
        RECT 127.950 67.950 130.050 68.400 ;
        RECT 202.950 69.600 205.050 70.050 ;
        RECT 286.950 69.600 289.050 70.050 ;
        RECT 307.950 69.600 310.050 70.050 ;
        RECT 337.950 69.600 340.050 70.050 ;
        RECT 388.950 69.600 391.050 70.050 ;
        RECT 202.950 68.400 225.600 69.600 ;
        RECT 202.950 67.950 205.050 68.400 ;
        RECT 224.400 67.050 225.600 68.400 ;
        RECT 286.950 68.400 391.050 69.600 ;
        RECT 286.950 67.950 289.050 68.400 ;
        RECT 307.950 67.950 310.050 68.400 ;
        RECT 337.950 67.950 340.050 68.400 ;
        RECT 388.950 67.950 391.050 68.400 ;
        RECT 427.950 69.600 430.050 70.050 ;
        RECT 469.950 69.600 472.050 70.050 ;
        RECT 427.950 68.400 472.050 69.600 ;
        RECT 427.950 67.950 430.050 68.400 ;
        RECT 469.950 67.950 472.050 68.400 ;
        RECT 499.950 69.600 502.050 70.050 ;
        RECT 532.950 69.600 535.050 70.050 ;
        RECT 553.950 69.600 556.050 70.050 ;
        RECT 571.950 69.600 574.050 70.050 ;
        RECT 499.950 68.400 574.050 69.600 ;
        RECT 499.950 67.950 502.050 68.400 ;
        RECT 532.950 67.950 535.050 68.400 ;
        RECT 553.950 67.950 556.050 68.400 ;
        RECT 571.950 67.950 574.050 68.400 ;
        RECT 601.950 69.600 604.050 70.050 ;
        RECT 607.950 69.600 610.050 70.050 ;
        RECT 634.950 69.600 637.050 70.050 ;
        RECT 694.950 69.600 697.050 70.050 ;
        RECT 601.950 68.400 637.050 69.600 ;
        RECT 601.950 67.950 604.050 68.400 ;
        RECT 607.950 67.950 610.050 68.400 ;
        RECT 634.950 67.950 637.050 68.400 ;
        RECT 641.400 68.400 697.050 69.600 ;
        RECT 85.950 66.600 88.050 66.900 ;
        RECT 130.950 66.600 133.050 67.050 ;
        RECT 85.950 65.400 133.050 66.600 ;
        RECT 85.950 64.800 88.050 65.400 ;
        RECT 130.950 64.950 133.050 65.400 ;
        RECT 223.950 66.600 226.050 67.050 ;
        RECT 259.950 66.600 262.050 67.050 ;
        RECT 223.950 65.400 262.050 66.600 ;
        RECT 223.950 64.950 226.050 65.400 ;
        RECT 259.950 64.950 262.050 65.400 ;
        RECT 394.950 66.600 397.050 67.050 ;
        RECT 412.950 66.600 415.050 67.050 ;
        RECT 394.950 65.400 415.050 66.600 ;
        RECT 394.950 64.950 397.050 65.400 ;
        RECT 412.950 64.950 415.050 65.400 ;
        RECT 424.950 66.600 427.050 67.050 ;
        RECT 433.950 66.600 436.050 67.050 ;
        RECT 424.950 65.400 436.050 66.600 ;
        RECT 424.950 64.950 427.050 65.400 ;
        RECT 433.950 64.950 436.050 65.400 ;
        RECT 628.950 66.600 631.050 67.050 ;
        RECT 641.400 66.600 642.600 68.400 ;
        RECT 694.950 67.950 697.050 68.400 ;
        RECT 883.950 69.600 886.050 70.050 ;
        RECT 898.950 69.600 901.050 70.050 ;
        RECT 883.950 68.400 901.050 69.600 ;
        RECT 883.950 67.950 886.050 68.400 ;
        RECT 898.950 67.950 901.050 68.400 ;
        RECT 907.950 69.600 910.050 70.050 ;
        RECT 916.950 69.600 919.050 70.050 ;
        RECT 907.950 68.400 919.050 69.600 ;
        RECT 907.950 67.950 910.050 68.400 ;
        RECT 916.950 67.950 919.050 68.400 ;
        RECT 736.950 66.600 739.050 67.050 ;
        RECT 628.950 65.400 642.600 66.600 ;
        RECT 719.400 65.400 739.050 66.600 ;
        RECT 628.950 64.950 631.050 65.400 ;
        RECT 13.950 63.600 16.050 64.050 ;
        RECT 28.950 63.600 31.050 64.200 ;
        RECT 13.950 62.400 31.050 63.600 ;
        RECT 13.950 61.950 16.050 62.400 ;
        RECT 28.950 62.100 31.050 62.400 ;
        RECT 46.950 63.600 49.050 64.050 ;
        RECT 64.950 63.600 67.050 64.050 ;
        RECT 46.950 62.400 67.050 63.600 ;
        RECT 46.950 61.950 49.050 62.400 ;
        RECT 64.950 61.950 67.050 62.400 ;
        RECT 211.950 63.600 214.050 64.050 ;
        RECT 235.950 63.600 238.050 64.050 ;
        RECT 211.950 62.400 238.050 63.600 ;
        RECT 211.950 61.950 214.050 62.400 ;
        RECT 235.950 61.950 238.050 62.400 ;
        RECT 346.950 63.600 349.050 64.050 ;
        RECT 478.950 63.600 481.050 64.050 ;
        RECT 487.950 63.600 490.050 64.050 ;
        RECT 346.950 62.400 426.600 63.600 ;
        RECT 346.950 61.950 349.050 62.400 ;
        RECT 31.950 60.600 34.050 61.050 ;
        RECT 67.950 60.600 70.050 61.050 ;
        RECT 76.950 60.600 79.050 61.200 ;
        RECT 31.950 59.400 79.050 60.600 ;
        RECT 31.950 58.950 34.050 59.400 ;
        RECT 67.950 58.950 70.050 59.400 ;
        RECT 76.950 59.100 79.050 59.400 ;
        RECT 88.950 58.950 91.050 61.050 ;
        RECT 94.950 60.600 97.050 61.200 ;
        RECT 109.950 60.600 112.050 61.050 ;
        RECT 115.950 60.600 118.050 61.050 ;
        RECT 94.950 59.400 118.050 60.600 ;
        RECT 94.950 59.100 97.050 59.400 ;
        RECT 109.950 58.950 112.050 59.400 ;
        RECT 115.950 58.950 118.050 59.400 ;
        RECT 136.950 59.100 139.050 61.200 ;
        RECT 142.950 59.100 145.050 61.200 ;
        RECT 157.950 59.100 160.050 61.200 ;
        RECT 163.950 59.100 166.050 61.200 ;
        RECT 175.950 60.600 178.050 61.200 ;
        RECT 184.950 60.600 187.050 61.050 ;
        RECT 241.950 60.600 244.050 61.200 ;
        RECT 175.950 59.400 187.050 60.600 ;
        RECT 175.950 59.100 178.050 59.400 ;
        RECT 1.950 54.450 4.050 54.900 ;
        RECT 16.950 54.450 19.050 54.900 ;
        RECT 1.950 53.250 19.050 54.450 ;
        RECT 1.950 52.800 4.050 53.250 ;
        RECT 16.950 52.800 19.050 53.250 ;
        RECT 22.950 54.600 25.050 55.050 ;
        RECT 28.950 54.600 31.050 54.900 ;
        RECT 22.950 53.400 31.050 54.600 ;
        RECT 22.950 52.950 25.050 53.400 ;
        RECT 28.950 52.800 31.050 53.400 ;
        RECT 58.950 54.450 61.050 54.900 ;
        RECT 67.950 54.450 70.050 54.900 ;
        RECT 58.950 53.250 70.050 54.450 ;
        RECT 58.950 52.800 61.050 53.250 ;
        RECT 67.950 52.800 70.050 53.250 ;
        RECT 73.950 54.450 76.050 54.900 ;
        RECT 85.950 54.450 88.050 54.900 ;
        RECT 73.950 53.250 88.050 54.450 ;
        RECT 89.400 54.600 90.600 58.950 ;
        RECT 137.400 57.600 138.600 59.100 ;
        RECT 131.400 56.400 138.600 57.600 ;
        RECT 143.400 57.600 144.600 59.100 ;
        RECT 158.400 57.600 159.600 59.100 ;
        RECT 143.400 56.400 159.600 57.600 ;
        RECT 91.950 54.600 94.050 54.900 ;
        RECT 89.400 53.400 94.050 54.600 ;
        RECT 73.950 52.800 76.050 53.250 ;
        RECT 85.950 52.800 88.050 53.250 ;
        RECT 91.950 52.800 94.050 53.400 ;
        RECT 118.950 54.600 121.050 54.900 ;
        RECT 131.400 54.600 132.600 56.400 ;
        RECT 158.400 55.050 159.600 56.400 ;
        RECT 118.950 53.400 132.600 54.600 ;
        RECT 154.950 53.400 159.600 55.050 ;
        RECT 164.400 55.050 165.600 59.100 ;
        RECT 184.950 58.950 187.050 59.400 ;
        RECT 236.400 59.400 244.050 60.600 ;
        RECT 236.400 58.050 237.600 59.400 ;
        RECT 241.950 59.100 244.050 59.400 ;
        RECT 256.950 60.750 259.050 61.200 ;
        RECT 265.950 60.750 268.050 61.200 ;
        RECT 256.950 59.550 268.050 60.750 ;
        RECT 256.950 59.100 259.050 59.550 ;
        RECT 265.950 59.100 268.050 59.550 ;
        RECT 271.950 60.600 274.050 61.200 ;
        RECT 277.950 60.600 280.050 61.050 ;
        RECT 271.950 59.400 280.050 60.600 ;
        RECT 271.950 59.100 274.050 59.400 ;
        RECT 277.950 58.950 280.050 59.400 ;
        RECT 292.950 60.750 295.050 61.200 ;
        RECT 301.950 60.750 304.050 61.200 ;
        RECT 292.950 59.550 304.050 60.750 ;
        RECT 292.950 59.100 295.050 59.550 ;
        RECT 301.950 59.100 304.050 59.550 ;
        RECT 313.950 60.750 316.050 61.200 ;
        RECT 322.950 60.750 325.050 61.200 ;
        RECT 313.950 59.550 325.050 60.750 ;
        RECT 313.950 59.100 316.050 59.550 ;
        RECT 322.950 59.100 325.050 59.550 ;
        RECT 382.950 59.100 385.050 61.200 ;
        RECT 391.950 60.750 394.050 61.200 ;
        RECT 406.950 60.750 409.050 61.200 ;
        RECT 391.950 60.600 409.050 60.750 ;
        RECT 391.950 59.550 417.600 60.600 ;
        RECT 391.950 59.100 394.050 59.550 ;
        RECT 406.950 59.400 417.600 59.550 ;
        RECT 406.950 59.100 409.050 59.400 ;
        RECT 232.950 56.400 237.600 58.050 ;
        RECT 335.400 56.400 348.600 57.600 ;
        RECT 232.950 55.950 237.000 56.400 ;
        RECT 164.400 53.400 169.050 55.050 ;
        RECT 118.950 52.800 121.050 53.400 ;
        RECT 154.950 52.950 159.000 53.400 ;
        RECT 165.000 52.950 169.050 53.400 ;
        RECT 178.950 54.600 181.050 54.900 ;
        RECT 193.950 54.600 196.050 54.900 ;
        RECT 178.950 53.400 196.050 54.600 ;
        RECT 178.950 52.800 181.050 53.400 ;
        RECT 193.950 52.800 196.050 53.400 ;
        RECT 199.950 54.600 202.050 54.900 ;
        RECT 211.950 54.600 214.050 54.900 ;
        RECT 199.950 54.450 214.050 54.600 ;
        RECT 220.950 54.450 223.050 54.900 ;
        RECT 199.950 53.400 223.050 54.450 ;
        RECT 199.950 52.800 202.050 53.400 ;
        RECT 211.950 53.250 223.050 53.400 ;
        RECT 211.950 52.800 214.050 53.250 ;
        RECT 220.950 52.800 223.050 53.250 ;
        RECT 226.950 54.600 229.050 54.900 ;
        RECT 238.950 54.600 241.050 54.900 ;
        RECT 226.950 53.400 241.050 54.600 ;
        RECT 226.950 52.800 229.050 53.400 ;
        RECT 238.950 52.800 241.050 53.400 ;
        RECT 253.950 54.600 256.050 55.050 ;
        RECT 283.950 54.600 286.050 55.050 ;
        RECT 253.950 53.400 286.050 54.600 ;
        RECT 253.950 52.950 256.050 53.400 ;
        RECT 283.950 52.950 286.050 53.400 ;
        RECT 289.950 54.600 292.050 54.900 ;
        RECT 298.800 54.600 300.900 55.050 ;
        RECT 289.950 53.400 300.900 54.600 ;
        RECT 289.950 52.800 292.050 53.400 ;
        RECT 298.800 52.950 300.900 53.400 ;
        RECT 301.950 54.600 304.050 55.050 ;
        RECT 316.950 54.600 319.050 55.050 ;
        RECT 335.400 54.900 336.600 56.400 ;
        RECT 347.400 54.900 348.600 56.400 ;
        RECT 301.950 53.400 319.050 54.600 ;
        RECT 301.950 52.950 304.050 53.400 ;
        RECT 316.950 52.950 319.050 53.400 ;
        RECT 334.950 52.800 337.050 54.900 ;
        RECT 346.950 54.450 349.050 54.900 ;
        RECT 358.950 54.450 361.050 54.900 ;
        RECT 346.950 53.250 361.050 54.450 ;
        RECT 383.400 54.600 384.600 59.100 ;
        RECT 416.400 55.050 417.600 59.400 ;
        RECT 418.950 59.100 421.050 61.200 ;
        RECT 403.950 54.600 406.050 54.900 ;
        RECT 383.400 53.400 406.050 54.600 ;
        RECT 346.950 52.800 349.050 53.250 ;
        RECT 358.950 52.800 361.050 53.250 ;
        RECT 403.950 52.800 406.050 53.400 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 133.950 51.600 136.050 52.050 ;
        RECT 151.950 51.600 154.050 52.050 ;
        RECT 133.950 50.400 154.050 51.600 ;
        RECT 133.950 49.950 136.050 50.400 ;
        RECT 151.950 49.950 154.050 50.400 ;
        RECT 244.950 51.600 247.050 52.050 ;
        RECT 256.950 51.600 259.050 52.050 ;
        RECT 244.950 50.400 259.050 51.600 ;
        RECT 244.950 49.950 247.050 50.400 ;
        RECT 256.950 49.950 259.050 50.400 ;
        RECT 310.950 51.600 313.050 52.050 ;
        RECT 406.950 51.600 409.050 52.050 ;
        RECT 419.400 51.600 420.600 59.100 ;
        RECT 425.400 54.600 426.600 62.400 ;
        RECT 478.950 62.400 490.050 63.600 ;
        RECT 478.950 61.950 481.050 62.400 ;
        RECT 487.950 61.950 490.050 62.400 ;
        RECT 499.950 63.600 502.050 64.050 ;
        RECT 508.950 63.600 511.050 64.050 ;
        RECT 499.950 62.400 511.050 63.600 ;
        RECT 499.950 61.950 502.050 62.400 ;
        RECT 508.950 61.950 511.050 62.400 ;
        RECT 595.950 63.600 598.050 64.050 ;
        RECT 619.950 63.600 622.050 64.050 ;
        RECT 688.950 63.600 691.050 64.050 ;
        RECT 595.950 62.400 691.050 63.600 ;
        RECT 595.950 61.950 598.050 62.400 ;
        RECT 619.950 61.950 622.050 62.400 ;
        RECT 688.950 61.950 691.050 62.400 ;
        RECT 706.950 63.600 709.050 64.050 ;
        RECT 719.400 63.600 720.600 65.400 ;
        RECT 736.950 64.950 739.050 65.400 ;
        RECT 868.950 66.600 871.050 67.050 ;
        RECT 904.950 66.600 907.050 67.050 ;
        RECT 868.950 65.400 907.050 66.600 ;
        RECT 868.950 64.950 871.050 65.400 ;
        RECT 904.950 64.950 907.050 65.400 ;
        RECT 706.950 62.400 720.600 63.600 ;
        RECT 790.950 63.600 793.050 64.050 ;
        RECT 799.950 63.600 802.050 64.050 ;
        RECT 826.950 63.600 829.050 64.050 ;
        RECT 790.950 62.400 829.050 63.600 ;
        RECT 706.950 61.950 709.050 62.400 ;
        RECT 790.950 61.950 793.050 62.400 ;
        RECT 799.950 61.950 802.050 62.400 ;
        RECT 826.950 61.950 829.050 62.400 ;
        RECT 913.950 63.600 916.050 64.050 ;
        RECT 925.950 63.600 928.050 64.050 ;
        RECT 913.950 62.400 928.050 63.600 ;
        RECT 913.950 61.950 916.050 62.400 ;
        RECT 925.950 61.950 928.050 62.400 ;
        RECT 436.950 60.750 439.050 61.200 ;
        RECT 445.950 60.750 448.050 61.200 ;
        RECT 436.950 59.550 448.050 60.750 ;
        RECT 436.950 59.100 439.050 59.550 ;
        RECT 445.950 59.100 448.050 59.550 ;
        RECT 469.950 60.750 472.050 61.200 ;
        RECT 475.950 60.750 478.050 61.200 ;
        RECT 469.950 59.550 478.050 60.750 ;
        RECT 469.950 59.100 472.050 59.550 ;
        RECT 475.950 59.100 478.050 59.550 ;
        RECT 493.950 60.750 496.050 61.200 ;
        RECT 517.950 60.750 520.050 61.200 ;
        RECT 493.950 59.550 520.050 60.750 ;
        RECT 493.950 59.100 496.050 59.550 ;
        RECT 517.950 59.100 520.050 59.550 ;
        RECT 547.950 60.600 550.050 61.200 ;
        RECT 577.950 60.600 580.050 61.200 ;
        RECT 613.950 60.600 616.050 61.200 ;
        RECT 547.950 59.400 580.050 60.600 ;
        RECT 547.950 59.100 550.050 59.400 ;
        RECT 577.950 59.100 580.050 59.400 ;
        RECT 611.400 59.400 616.050 60.600 ;
        RECT 611.400 57.600 612.600 59.400 ;
        RECT 613.950 59.100 616.050 59.400 ;
        RECT 652.950 60.750 655.050 61.200 ;
        RECT 661.950 60.750 664.050 61.200 ;
        RECT 652.950 60.600 664.050 60.750 ;
        RECT 682.950 60.600 685.050 61.200 ;
        RECT 652.950 59.550 685.050 60.600 ;
        RECT 652.950 59.100 655.050 59.550 ;
        RECT 661.950 59.400 685.050 59.550 ;
        RECT 661.950 59.100 664.050 59.400 ;
        RECT 682.950 59.100 685.050 59.400 ;
        RECT 715.950 60.600 718.050 61.050 ;
        RECT 721.950 60.600 724.050 61.200 ;
        RECT 715.950 59.400 724.050 60.600 ;
        RECT 715.950 58.950 718.050 59.400 ;
        RECT 721.950 59.100 724.050 59.400 ;
        RECT 730.950 60.600 733.050 61.200 ;
        RECT 745.950 60.600 748.050 61.200 ;
        RECT 730.950 59.400 748.050 60.600 ;
        RECT 730.950 59.100 733.050 59.400 ;
        RECT 745.950 59.100 748.050 59.400 ;
        RECT 850.950 60.750 853.050 61.200 ;
        RECT 862.950 60.750 865.050 61.200 ;
        RECT 850.950 59.550 865.050 60.750 ;
        RECT 850.950 59.100 853.050 59.550 ;
        RECT 862.950 59.100 865.050 59.550 ;
        RECT 868.950 60.600 871.050 61.050 ;
        RECT 874.950 60.600 877.050 61.050 ;
        RECT 868.950 59.400 877.050 60.600 ;
        RECT 868.950 58.950 871.050 59.400 ;
        RECT 874.950 58.950 877.050 59.400 ;
        RECT 895.950 59.100 898.050 61.200 ;
        RECT 896.400 57.600 897.600 59.100 ;
        RECT 904.950 58.950 907.050 61.050 ;
        RECT 919.950 58.950 922.050 61.050 ;
        RECT 569.400 56.400 588.600 57.600 ;
        RECT 430.950 54.600 433.050 55.050 ;
        RECT 425.400 53.400 433.050 54.600 ;
        RECT 430.950 52.950 433.050 53.400 ;
        RECT 466.950 54.600 469.050 54.900 ;
        RECT 478.950 54.600 481.050 55.050 ;
        RECT 466.950 53.400 481.050 54.600 ;
        RECT 466.950 52.800 469.050 53.400 ;
        RECT 478.950 52.950 481.050 53.400 ;
        RECT 550.950 54.600 553.050 54.900 ;
        RECT 569.400 54.600 570.600 56.400 ;
        RECT 587.400 55.050 588.600 56.400 ;
        RECT 605.400 56.400 612.600 57.600 ;
        RECT 890.400 56.400 897.600 57.600 ;
        RECT 586.950 54.600 589.050 55.050 ;
        RECT 550.950 53.400 570.600 54.600 ;
        RECT 578.400 53.400 589.050 54.600 ;
        RECT 550.950 52.800 553.050 53.400 ;
        RECT 578.400 52.050 579.600 53.400 ;
        RECT 586.950 52.950 589.050 53.400 ;
        RECT 598.950 54.600 601.050 54.900 ;
        RECT 605.400 54.600 606.600 56.400 ;
        RECT 598.950 53.400 606.600 54.600 ;
        RECT 607.950 54.450 610.050 54.900 ;
        RECT 616.950 54.450 619.050 54.900 ;
        RECT 598.950 52.800 601.050 53.400 ;
        RECT 607.950 53.250 619.050 54.450 ;
        RECT 607.950 52.800 610.050 53.250 ;
        RECT 616.950 52.800 619.050 53.250 ;
        RECT 718.950 54.450 721.050 54.900 ;
        RECT 727.950 54.450 730.050 54.900 ;
        RECT 718.950 53.250 730.050 54.450 ;
        RECT 718.950 52.800 721.050 53.250 ;
        RECT 727.950 52.800 730.050 53.250 ;
        RECT 736.950 54.450 739.050 54.900 ;
        RECT 742.950 54.450 745.050 54.900 ;
        RECT 736.950 53.250 745.050 54.450 ;
        RECT 736.950 52.800 739.050 53.250 ;
        RECT 742.950 52.800 745.050 53.250 ;
        RECT 757.950 54.450 760.050 54.900 ;
        RECT 763.950 54.450 766.050 54.900 ;
        RECT 757.950 53.250 766.050 54.450 ;
        RECT 757.950 52.800 760.050 53.250 ;
        RECT 763.950 52.800 766.050 53.250 ;
        RECT 787.950 54.600 790.050 54.900 ;
        RECT 796.950 54.600 799.050 55.050 ;
        RECT 787.950 53.400 799.050 54.600 ;
        RECT 787.950 52.800 790.050 53.400 ;
        RECT 796.950 52.950 799.050 53.400 ;
        RECT 853.950 54.600 856.050 55.050 ;
        RECT 859.950 54.600 862.050 55.050 ;
        RECT 853.950 53.400 862.050 54.600 ;
        RECT 853.950 52.950 856.050 53.400 ;
        RECT 859.950 52.950 862.050 53.400 ;
        RECT 310.950 51.000 321.600 51.600 ;
        RECT 310.950 50.400 322.050 51.000 ;
        RECT 310.950 49.950 313.050 50.400 ;
        RECT 52.950 48.600 55.050 49.050 ;
        RECT 109.950 48.600 112.050 49.050 ;
        RECT 52.950 47.400 112.050 48.600 ;
        RECT 52.950 46.950 55.050 47.400 ;
        RECT 109.950 46.950 112.050 47.400 ;
        RECT 154.950 48.600 157.050 49.050 ;
        RECT 181.950 48.600 184.050 49.050 ;
        RECT 268.950 48.600 271.050 49.050 ;
        RECT 154.950 47.400 271.050 48.600 ;
        RECT 154.950 46.950 157.050 47.400 ;
        RECT 181.950 46.950 184.050 47.400 ;
        RECT 268.950 46.950 271.050 47.400 ;
        RECT 319.950 46.950 322.050 50.400 ;
        RECT 406.950 50.400 420.600 51.600 ;
        RECT 433.950 51.600 436.050 52.050 ;
        RECT 448.950 51.600 451.050 52.050 ;
        RECT 460.950 51.600 463.050 52.050 ;
        RECT 433.950 50.400 463.050 51.600 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 433.950 49.950 436.050 50.400 ;
        RECT 448.950 49.950 451.050 50.400 ;
        RECT 460.950 49.950 463.050 50.400 ;
        RECT 574.950 50.400 579.600 52.050 ;
        RECT 580.950 51.600 583.050 52.050 ;
        RECT 598.950 51.600 601.050 52.050 ;
        RECT 580.950 50.400 601.050 51.600 ;
        RECT 574.950 49.950 579.000 50.400 ;
        RECT 580.950 49.950 583.050 50.400 ;
        RECT 598.950 49.950 601.050 50.400 ;
        RECT 619.950 51.600 622.050 52.050 ;
        RECT 664.950 51.600 667.050 52.050 ;
        RECT 679.950 51.600 682.050 52.050 ;
        RECT 619.950 50.400 682.050 51.600 ;
        RECT 619.950 49.950 622.050 50.400 ;
        RECT 664.950 49.950 667.050 50.400 ;
        RECT 679.950 49.950 682.050 50.400 ;
        RECT 703.950 51.600 706.050 52.050 ;
        RECT 719.400 51.600 720.600 52.800 ;
        RECT 890.400 52.050 891.600 56.400 ;
        RECT 892.950 54.600 895.050 54.900 ;
        RECT 905.400 54.600 906.600 58.950 ;
        RECT 892.950 53.400 906.600 54.600 ;
        RECT 916.950 54.600 919.050 54.900 ;
        RECT 920.400 54.600 921.600 58.950 ;
        RECT 916.950 53.400 921.600 54.600 ;
        RECT 892.950 52.800 895.050 53.400 ;
        RECT 916.950 52.800 919.050 53.400 ;
        RECT 703.950 50.400 720.600 51.600 ;
        RECT 799.950 51.600 802.050 52.050 ;
        RECT 805.950 51.600 808.050 52.050 ;
        RECT 817.950 51.600 820.050 52.050 ;
        RECT 799.950 50.400 820.050 51.600 ;
        RECT 703.950 49.950 706.050 50.400 ;
        RECT 799.950 49.950 802.050 50.400 ;
        RECT 805.950 49.950 808.050 50.400 ;
        RECT 817.950 49.950 820.050 50.400 ;
        RECT 823.950 51.600 826.050 52.050 ;
        RECT 841.950 51.600 844.050 52.050 ;
        RECT 823.950 50.400 844.050 51.600 ;
        RECT 823.950 49.950 826.050 50.400 ;
        RECT 841.950 49.950 844.050 50.400 ;
        RECT 871.950 51.600 874.050 52.050 ;
        RECT 880.950 51.600 883.050 52.050 ;
        RECT 871.950 50.400 883.050 51.600 ;
        RECT 871.950 49.950 874.050 50.400 ;
        RECT 880.950 49.950 883.050 50.400 ;
        RECT 889.950 49.950 892.050 52.050 ;
        RECT 352.950 48.600 355.050 49.050 ;
        RECT 379.950 48.600 382.050 49.050 ;
        RECT 391.800 48.600 393.900 49.050 ;
        RECT 352.950 47.400 393.900 48.600 ;
        RECT 352.950 46.950 355.050 47.400 ;
        RECT 379.950 46.950 382.050 47.400 ;
        RECT 391.800 46.950 393.900 47.400 ;
        RECT 394.950 48.600 397.050 49.050 ;
        RECT 400.950 48.600 403.050 49.050 ;
        RECT 394.950 47.400 403.050 48.600 ;
        RECT 394.950 46.950 397.050 47.400 ;
        RECT 400.950 46.950 403.050 47.400 ;
        RECT 415.950 48.600 418.050 49.050 ;
        RECT 421.950 48.600 424.050 49.050 ;
        RECT 415.950 47.400 424.050 48.600 ;
        RECT 415.950 46.950 418.050 47.400 ;
        RECT 421.950 46.950 424.050 47.400 ;
        RECT 475.950 48.600 478.050 49.050 ;
        RECT 523.950 48.600 526.050 49.050 ;
        RECT 475.950 47.400 526.050 48.600 ;
        RECT 475.950 46.950 478.050 47.400 ;
        RECT 523.950 46.950 526.050 47.400 ;
        RECT 556.950 48.600 559.050 49.050 ;
        RECT 571.950 48.600 574.050 49.050 ;
        RECT 556.950 47.400 574.050 48.600 ;
        RECT 556.950 46.950 559.050 47.400 ;
        RECT 571.950 46.950 574.050 47.400 ;
        RECT 577.950 48.600 580.050 49.050 ;
        RECT 595.800 48.600 597.900 49.050 ;
        RECT 577.950 47.400 597.900 48.600 ;
        RECT 599.400 48.600 600.600 49.950 ;
        RECT 637.950 48.600 640.050 49.050 ;
        RECT 599.400 47.400 640.050 48.600 ;
        RECT 577.950 46.950 580.050 47.400 ;
        RECT 595.800 46.950 597.900 47.400 ;
        RECT 637.950 46.950 640.050 47.400 ;
        RECT 688.950 48.600 691.050 49.050 ;
        RECT 697.950 48.600 700.050 49.050 ;
        RECT 688.950 47.400 700.050 48.600 ;
        RECT 688.950 46.950 691.050 47.400 ;
        RECT 697.950 46.950 700.050 47.400 ;
        RECT 706.950 48.600 709.050 49.050 ;
        RECT 757.950 48.600 760.050 49.050 ;
        RECT 706.950 47.400 760.050 48.600 ;
        RECT 706.950 46.950 709.050 47.400 ;
        RECT 757.950 46.950 760.050 47.400 ;
        RECT 856.950 48.600 859.050 49.050 ;
        RECT 895.950 48.600 898.050 49.050 ;
        RECT 856.950 47.400 898.050 48.600 ;
        RECT 856.950 46.950 859.050 47.400 ;
        RECT 895.950 46.950 898.050 47.400 ;
        RECT 910.950 48.600 913.050 49.050 ;
        RECT 934.950 48.600 937.050 49.050 ;
        RECT 910.950 47.400 937.050 48.600 ;
        RECT 910.950 46.950 913.050 47.400 ;
        RECT 934.950 46.950 937.050 47.400 ;
        RECT 184.950 45.600 187.050 46.050 ;
        RECT 208.950 45.600 211.050 46.050 ;
        RECT 184.950 44.400 211.050 45.600 ;
        RECT 184.950 43.950 187.050 44.400 ;
        RECT 208.950 43.950 211.050 44.400 ;
        RECT 214.950 45.600 217.050 46.050 ;
        RECT 253.950 45.600 256.050 46.050 ;
        RECT 214.950 44.400 256.050 45.600 ;
        RECT 214.950 43.950 217.050 44.400 ;
        RECT 253.950 43.950 256.050 44.400 ;
        RECT 388.950 45.600 391.050 46.050 ;
        RECT 460.950 45.600 463.050 46.050 ;
        RECT 388.950 44.400 463.050 45.600 ;
        RECT 388.950 43.950 391.050 44.400 ;
        RECT 460.950 43.950 463.050 44.400 ;
        RECT 541.950 45.600 544.050 46.050 ;
        RECT 547.950 45.600 550.050 46.050 ;
        RECT 541.950 44.400 550.050 45.600 ;
        RECT 541.950 43.950 544.050 44.400 ;
        RECT 547.950 43.950 550.050 44.400 ;
        RECT 592.950 45.600 595.050 46.050 ;
        RECT 610.950 45.600 613.050 46.050 ;
        RECT 592.950 44.400 613.050 45.600 ;
        RECT 592.950 43.950 595.050 44.400 ;
        RECT 610.950 43.950 613.050 44.400 ;
        RECT 646.950 45.600 649.050 46.050 ;
        RECT 685.950 45.600 688.050 46.050 ;
        RECT 646.950 44.400 688.050 45.600 ;
        RECT 646.950 43.950 649.050 44.400 ;
        RECT 685.950 43.950 688.050 44.400 ;
        RECT 694.950 45.600 697.050 46.050 ;
        RECT 853.950 45.600 856.050 46.050 ;
        RECT 694.950 44.400 856.050 45.600 ;
        RECT 694.950 43.950 697.050 44.400 ;
        RECT 853.950 43.950 856.050 44.400 ;
        RECT 859.950 45.600 862.050 46.050 ;
        RECT 874.950 45.600 877.050 46.050 ;
        RECT 859.950 44.400 877.050 45.600 ;
        RECT 859.950 43.950 862.050 44.400 ;
        RECT 874.950 43.950 877.050 44.400 ;
        RECT 139.950 42.600 142.050 43.050 ;
        RECT 166.950 42.600 169.050 43.050 ;
        RECT 337.950 42.600 340.050 43.050 ;
        RECT 466.950 42.600 469.050 43.050 ;
        RECT 139.950 41.400 264.600 42.600 ;
        RECT 139.950 40.950 142.050 41.400 ;
        RECT 166.950 40.950 169.050 41.400 ;
        RECT 263.400 40.050 264.600 41.400 ;
        RECT 337.950 41.400 469.050 42.600 ;
        RECT 337.950 40.950 340.050 41.400 ;
        RECT 466.950 40.950 469.050 41.400 ;
        RECT 502.950 42.600 505.050 43.050 ;
        RECT 526.950 42.600 529.050 43.050 ;
        RECT 502.950 41.400 529.050 42.600 ;
        RECT 502.950 40.950 505.050 41.400 ;
        RECT 526.950 40.950 529.050 41.400 ;
        RECT 565.950 42.600 568.050 43.050 ;
        RECT 628.950 42.600 631.050 43.050 ;
        RECT 565.950 41.400 631.050 42.600 ;
        RECT 565.950 40.950 568.050 41.400 ;
        RECT 628.950 40.950 631.050 41.400 ;
        RECT 643.950 42.600 646.050 43.050 ;
        RECT 691.950 42.600 694.050 43.050 ;
        RECT 643.950 41.400 694.050 42.600 ;
        RECT 643.950 40.950 646.050 41.400 ;
        RECT 691.950 40.950 694.050 41.400 ;
        RECT 775.950 42.600 778.050 43.050 ;
        RECT 781.950 42.600 784.050 43.050 ;
        RECT 793.950 42.600 796.050 43.050 ;
        RECT 775.950 41.400 796.050 42.600 ;
        RECT 775.950 40.950 778.050 41.400 ;
        RECT 781.950 40.950 784.050 41.400 ;
        RECT 793.950 40.950 796.050 41.400 ;
        RECT 127.950 39.600 130.050 40.050 ;
        RECT 160.950 39.600 163.050 40.050 ;
        RECT 127.950 38.400 163.050 39.600 ;
        RECT 127.950 37.950 130.050 38.400 ;
        RECT 160.950 37.950 163.050 38.400 ;
        RECT 196.950 39.600 199.050 40.050 ;
        RECT 226.950 39.600 229.050 40.050 ;
        RECT 196.950 38.400 229.050 39.600 ;
        RECT 196.950 37.950 199.050 38.400 ;
        RECT 226.950 37.950 229.050 38.400 ;
        RECT 262.950 39.600 265.050 40.050 ;
        RECT 286.950 39.600 289.050 40.050 ;
        RECT 310.950 39.600 313.050 40.050 ;
        RECT 397.950 39.600 400.050 40.050 ;
        RECT 490.950 39.600 493.050 40.050 ;
        RECT 262.950 38.400 313.050 39.600 ;
        RECT 262.950 37.950 265.050 38.400 ;
        RECT 286.950 37.950 289.050 38.400 ;
        RECT 310.950 37.950 313.050 38.400 ;
        RECT 392.400 38.400 493.050 39.600 ;
        RECT 352.950 36.600 355.050 37.050 ;
        RECT 392.400 36.600 393.600 38.400 ;
        RECT 397.950 37.950 400.050 38.400 ;
        RECT 490.950 37.950 493.050 38.400 ;
        RECT 592.950 39.600 595.050 40.050 ;
        RECT 644.400 39.600 645.600 40.950 ;
        RECT 592.950 38.400 645.600 39.600 ;
        RECT 712.950 39.600 715.050 40.050 ;
        RECT 727.950 39.600 730.050 40.050 ;
        RECT 769.950 39.600 772.050 40.050 ;
        RECT 712.950 38.400 772.050 39.600 ;
        RECT 592.950 37.950 595.050 38.400 ;
        RECT 712.950 37.950 715.050 38.400 ;
        RECT 727.950 37.950 730.050 38.400 ;
        RECT 769.950 37.950 772.050 38.400 ;
        RECT 811.950 39.600 814.050 40.050 ;
        RECT 841.950 39.600 844.050 40.050 ;
        RECT 811.950 38.400 844.050 39.600 ;
        RECT 811.950 37.950 814.050 38.400 ;
        RECT 841.950 37.950 844.050 38.400 ;
        RECT 856.950 39.600 859.050 40.050 ;
        RECT 868.950 39.600 871.050 40.050 ;
        RECT 856.950 38.400 871.050 39.600 ;
        RECT 856.950 37.950 859.050 38.400 ;
        RECT 868.950 37.950 871.050 38.400 ;
        RECT 352.950 35.400 393.600 36.600 ;
        RECT 400.950 36.600 403.050 37.050 ;
        RECT 454.950 36.600 457.050 37.050 ;
        RECT 499.950 36.600 502.050 37.050 ;
        RECT 400.950 35.400 502.050 36.600 ;
        RECT 352.950 34.950 355.050 35.400 ;
        RECT 400.950 34.950 403.050 35.400 ;
        RECT 454.950 34.950 457.050 35.400 ;
        RECT 499.950 34.950 502.050 35.400 ;
        RECT 568.950 36.600 571.050 37.050 ;
        RECT 586.950 36.600 589.050 37.050 ;
        RECT 568.950 35.400 589.050 36.600 ;
        RECT 568.950 34.950 571.050 35.400 ;
        RECT 586.950 34.950 589.050 35.400 ;
        RECT 601.950 36.600 604.050 37.050 ;
        RECT 646.950 36.600 649.050 37.050 ;
        RECT 601.950 35.400 649.050 36.600 ;
        RECT 601.950 34.950 604.050 35.400 ;
        RECT 646.950 34.950 649.050 35.400 ;
        RECT 658.950 36.600 661.050 37.050 ;
        RECT 670.950 36.600 673.050 37.050 ;
        RECT 658.950 35.400 673.050 36.600 ;
        RECT 658.950 34.950 661.050 35.400 ;
        RECT 670.950 34.950 673.050 35.400 ;
        RECT 700.950 36.600 703.050 37.050 ;
        RECT 706.950 36.600 709.050 37.050 ;
        RECT 700.950 35.400 709.050 36.600 ;
        RECT 842.400 36.600 843.600 37.950 ;
        RECT 850.950 36.600 853.050 37.050 ;
        RECT 865.950 36.600 868.050 37.050 ;
        RECT 842.400 35.400 868.050 36.600 ;
        RECT 700.950 34.950 703.050 35.400 ;
        RECT 706.950 34.950 709.050 35.400 ;
        RECT 850.950 34.950 853.050 35.400 ;
        RECT 865.950 34.950 868.050 35.400 ;
        RECT 874.950 36.600 877.050 37.050 ;
        RECT 883.950 36.600 886.050 37.050 ;
        RECT 922.950 36.600 925.050 37.050 ;
        RECT 874.950 35.400 925.050 36.600 ;
        RECT 874.950 34.950 877.050 35.400 ;
        RECT 883.950 34.950 886.050 35.400 ;
        RECT 922.950 34.950 925.050 35.400 ;
        RECT 34.950 33.600 37.050 34.050 ;
        RECT 73.950 33.600 76.050 34.050 ;
        RECT 34.950 32.400 76.050 33.600 ;
        RECT 34.950 31.950 37.050 32.400 ;
        RECT 73.950 31.950 76.050 32.400 ;
        RECT 97.950 33.600 100.050 34.050 ;
        RECT 106.950 33.600 109.050 34.050 ;
        RECT 118.950 33.600 121.050 34.050 ;
        RECT 154.950 33.600 157.050 34.050 ;
        RECT 163.950 33.600 166.050 34.050 ;
        RECT 193.950 33.600 196.050 34.050 ;
        RECT 211.950 33.600 214.050 34.050 ;
        RECT 97.950 32.400 114.600 33.600 ;
        RECT 97.950 31.950 100.050 32.400 ;
        RECT 106.950 31.950 109.050 32.400 ;
        RECT 113.400 30.600 114.600 32.400 ;
        RECT 118.950 32.400 214.050 33.600 ;
        RECT 118.950 31.950 121.050 32.400 ;
        RECT 154.950 31.950 157.050 32.400 ;
        RECT 163.950 31.950 166.050 32.400 ;
        RECT 193.950 31.950 196.050 32.400 ;
        RECT 211.950 31.950 214.050 32.400 ;
        RECT 226.950 33.600 229.050 34.050 ;
        RECT 232.950 33.600 235.050 34.050 ;
        RECT 226.950 32.400 235.050 33.600 ;
        RECT 226.950 31.950 229.050 32.400 ;
        RECT 232.950 31.950 235.050 32.400 ;
        RECT 283.950 33.600 286.050 34.050 ;
        RECT 325.950 33.600 328.050 34.050 ;
        RECT 283.950 32.400 328.050 33.600 ;
        RECT 283.950 31.950 286.050 32.400 ;
        RECT 325.950 31.950 328.050 32.400 ;
        RECT 331.950 33.600 334.050 34.050 ;
        RECT 364.950 33.600 367.050 34.050 ;
        RECT 385.950 33.600 388.050 34.050 ;
        RECT 331.950 32.400 348.600 33.600 ;
        RECT 331.950 31.950 334.050 32.400 ;
        RECT 124.950 30.600 127.050 31.050 ;
        RECT 113.400 29.400 127.050 30.600 ;
        RECT 124.950 28.950 127.050 29.400 ;
        RECT 214.950 28.950 217.050 31.050 ;
        RECT 235.950 28.950 238.050 31.050 ;
        RECT 280.950 30.600 283.050 31.050 ;
        RECT 331.950 30.600 334.050 30.900 ;
        RECT 280.950 29.400 334.050 30.600 ;
        RECT 347.400 30.600 348.600 32.400 ;
        RECT 364.950 32.400 388.050 33.600 ;
        RECT 364.950 31.950 367.050 32.400 ;
        RECT 385.950 31.950 388.050 32.400 ;
        RECT 400.950 33.600 403.050 33.900 ;
        RECT 409.950 33.600 412.050 34.050 ;
        RECT 400.950 32.400 412.050 33.600 ;
        RECT 400.950 31.800 403.050 32.400 ;
        RECT 409.950 31.950 412.050 32.400 ;
        RECT 466.950 33.600 469.050 34.050 ;
        RECT 484.950 33.600 487.050 34.050 ;
        RECT 496.950 33.600 499.050 34.050 ;
        RECT 466.950 32.400 499.050 33.600 ;
        RECT 466.950 31.950 469.050 32.400 ;
        RECT 484.950 31.950 487.050 32.400 ;
        RECT 496.950 31.950 499.050 32.400 ;
        RECT 508.950 33.600 511.050 34.050 ;
        RECT 562.950 33.600 565.050 34.050 ;
        RECT 616.950 33.600 619.050 34.050 ;
        RECT 508.950 32.400 619.050 33.600 ;
        RECT 508.950 31.950 511.050 32.400 ;
        RECT 562.950 31.950 565.050 32.400 ;
        RECT 616.950 31.950 619.050 32.400 ;
        RECT 664.950 33.600 667.050 34.050 ;
        RECT 673.950 33.600 676.050 34.050 ;
        RECT 664.950 32.400 676.050 33.600 ;
        RECT 664.950 31.950 667.050 32.400 ;
        RECT 673.950 31.950 676.050 32.400 ;
        RECT 679.950 33.600 682.050 34.050 ;
        RECT 685.950 33.600 688.050 34.050 ;
        RECT 679.950 32.400 688.050 33.600 ;
        RECT 679.950 31.950 682.050 32.400 ;
        RECT 685.950 31.950 688.050 32.400 ;
        RECT 748.950 33.600 751.050 34.050 ;
        RECT 802.950 33.600 805.050 34.050 ;
        RECT 814.950 33.600 817.050 34.050 ;
        RECT 835.950 33.600 838.050 34.050 ;
        RECT 748.950 32.400 838.050 33.600 ;
        RECT 748.950 31.950 751.050 32.400 ;
        RECT 802.950 31.950 805.050 32.400 ;
        RECT 814.950 31.950 817.050 32.400 ;
        RECT 835.950 31.950 838.050 32.400 ;
        RECT 358.950 30.600 361.050 31.050 ;
        RECT 370.950 30.600 373.050 31.050 ;
        RECT 347.400 29.400 361.050 30.600 ;
        RECT 280.950 28.950 283.050 29.400 ;
        RECT 4.950 27.750 7.050 28.200 ;
        RECT 13.950 27.750 16.050 28.200 ;
        RECT 4.950 26.550 16.050 27.750 ;
        RECT 4.950 26.100 7.050 26.550 ;
        RECT 13.950 26.100 16.050 26.550 ;
        RECT 37.950 27.750 40.050 28.200 ;
        RECT 43.950 27.750 46.050 28.200 ;
        RECT 37.950 26.550 46.050 27.750 ;
        RECT 37.950 26.100 40.050 26.550 ;
        RECT 43.950 26.100 46.050 26.550 ;
        RECT 55.950 27.750 58.050 28.200 ;
        RECT 64.950 27.750 67.050 28.200 ;
        RECT 55.950 26.550 67.050 27.750 ;
        RECT 55.950 26.100 58.050 26.550 ;
        RECT 64.950 26.100 67.050 26.550 ;
        RECT 73.950 27.600 76.050 28.200 ;
        RECT 109.950 27.600 112.050 28.200 ;
        RECT 73.950 26.400 112.050 27.600 ;
        RECT 73.950 26.100 76.050 26.400 ;
        RECT 109.950 26.100 112.050 26.400 ;
        RECT 130.950 26.100 133.050 28.200 ;
        RECT 175.950 27.750 178.050 28.200 ;
        RECT 187.950 27.750 190.050 28.200 ;
        RECT 175.950 26.550 190.050 27.750 ;
        RECT 175.950 26.100 178.050 26.550 ;
        RECT 187.950 26.100 190.050 26.550 ;
        RECT 110.400 24.600 111.600 26.100 ;
        RECT 131.400 24.600 132.600 26.100 ;
        RECT 110.400 23.400 132.600 24.600 ;
        RECT 61.950 21.600 64.050 22.050 ;
        RECT 70.950 21.600 73.050 21.900 ;
        RECT 61.950 20.400 73.050 21.600 ;
        RECT 61.950 19.950 64.050 20.400 ;
        RECT 70.950 19.800 73.050 20.400 ;
        RECT 79.950 21.600 82.050 22.050 ;
        RECT 106.950 21.600 109.050 21.900 ;
        RECT 79.950 21.450 109.050 21.600 ;
        RECT 118.950 21.450 121.050 21.900 ;
        RECT 79.950 20.400 121.050 21.450 ;
        RECT 79.950 19.950 82.050 20.400 ;
        RECT 106.950 20.250 121.050 20.400 ;
        RECT 106.950 19.800 109.050 20.250 ;
        RECT 118.950 19.800 121.050 20.250 ;
        RECT 163.950 21.450 166.050 21.900 ;
        RECT 172.950 21.450 175.050 21.900 ;
        RECT 163.950 20.250 175.050 21.450 ;
        RECT 163.950 19.800 166.050 20.250 ;
        RECT 172.950 19.800 175.050 20.250 ;
        RECT 187.950 21.600 190.050 22.050 ;
        RECT 215.400 21.900 216.600 28.950 ;
        RECT 217.950 27.600 220.050 28.200 ;
        RECT 223.950 27.600 226.050 28.050 ;
        RECT 217.950 26.400 226.050 27.600 ;
        RECT 217.950 26.100 220.050 26.400 ;
        RECT 223.950 25.950 226.050 26.400 ;
        RECT 236.400 21.900 237.600 28.950 ;
        RECT 331.950 28.800 334.050 29.400 ;
        RECT 358.950 28.950 361.050 29.400 ;
        RECT 362.400 29.400 373.050 30.600 ;
        RECT 238.950 27.600 241.050 28.200 ;
        RECT 256.950 27.600 259.050 28.200 ;
        RECT 238.950 26.400 259.050 27.600 ;
        RECT 238.950 26.100 241.050 26.400 ;
        RECT 256.950 26.100 259.050 26.400 ;
        RECT 262.950 27.600 265.050 28.200 ;
        RECT 286.950 27.600 291.000 28.050 ;
        RECT 292.950 27.600 295.050 28.200 ;
        RECT 325.950 27.600 328.050 28.050 ;
        RECT 262.950 26.400 282.600 27.600 ;
        RECT 262.950 26.100 265.050 26.400 ;
        RECT 281.400 25.050 282.600 26.400 ;
        RECT 286.950 25.950 291.600 27.600 ;
        RECT 292.950 26.400 328.050 27.600 ;
        RECT 292.950 26.100 295.050 26.400 ;
        RECT 325.950 25.950 328.050 26.400 ;
        RECT 281.400 23.400 286.050 25.050 ;
        RECT 282.000 22.950 286.050 23.400 ;
        RECT 290.400 21.900 291.600 25.950 ;
        RECT 362.400 21.900 363.600 29.400 ;
        RECT 370.950 28.950 373.050 29.400 ;
        RECT 388.950 30.600 391.050 31.050 ;
        RECT 412.950 30.600 415.050 31.050 ;
        RECT 388.950 29.400 415.050 30.600 ;
        RECT 388.950 28.950 391.050 29.400 ;
        RECT 412.950 28.950 415.050 29.400 ;
        RECT 517.950 30.600 520.050 31.050 ;
        RECT 622.950 30.600 625.050 31.050 ;
        RECT 658.950 30.600 661.050 31.050 ;
        RECT 517.950 29.400 661.050 30.600 ;
        RECT 517.950 28.950 520.050 29.400 ;
        RECT 373.950 27.600 376.050 28.050 ;
        RECT 382.950 27.600 385.050 28.200 ;
        RECT 373.950 26.400 385.050 27.600 ;
        RECT 373.950 25.950 376.050 26.400 ;
        RECT 382.950 26.100 385.050 26.400 ;
        RECT 448.950 27.600 451.050 28.200 ;
        RECT 475.950 27.600 478.050 28.050 ;
        RECT 484.950 27.600 487.050 28.200 ;
        RECT 448.950 26.400 465.600 27.600 ;
        RECT 448.950 26.100 451.050 26.400 ;
        RECT 464.400 24.600 465.600 26.400 ;
        RECT 475.950 26.400 487.050 27.600 ;
        RECT 475.950 25.950 478.050 26.400 ;
        RECT 484.950 26.100 487.050 26.400 ;
        RECT 493.950 27.600 496.050 28.050 ;
        RECT 502.950 27.600 505.050 28.200 ;
        RECT 493.950 26.400 505.050 27.600 ;
        RECT 493.950 25.950 496.050 26.400 ;
        RECT 502.950 26.100 505.050 26.400 ;
        RECT 532.950 27.600 535.050 28.200 ;
        RECT 553.950 27.750 556.050 28.200 ;
        RECT 568.950 27.750 571.050 28.200 ;
        RECT 553.950 27.600 571.050 27.750 ;
        RECT 532.950 26.550 571.050 27.600 ;
        RECT 532.950 26.400 556.050 26.550 ;
        RECT 532.950 26.100 535.050 26.400 ;
        RECT 553.950 26.100 556.050 26.400 ;
        RECT 568.950 26.100 571.050 26.550 ;
        RECT 464.400 23.400 468.600 24.600 ;
        RECT 193.950 21.600 196.050 21.900 ;
        RECT 208.950 21.600 211.050 21.900 ;
        RECT 187.950 20.400 211.050 21.600 ;
        RECT 187.950 19.950 190.050 20.400 ;
        RECT 193.950 19.800 196.050 20.400 ;
        RECT 208.950 19.800 211.050 20.400 ;
        RECT 214.950 19.800 217.050 21.900 ;
        RECT 226.950 21.450 229.050 21.900 ;
        RECT 235.950 21.450 238.050 21.900 ;
        RECT 226.950 20.250 238.050 21.450 ;
        RECT 226.950 19.800 229.050 20.250 ;
        RECT 235.950 19.800 238.050 20.250 ;
        RECT 253.950 21.600 256.050 21.900 ;
        RECT 274.950 21.600 277.050 21.900 ;
        RECT 253.950 20.400 277.050 21.600 ;
        RECT 253.950 19.800 256.050 20.400 ;
        RECT 274.950 19.800 277.050 20.400 ;
        RECT 289.950 19.800 292.050 21.900 ;
        RECT 295.950 21.600 298.050 21.900 ;
        RECT 307.950 21.600 310.050 21.900 ;
        RECT 295.950 20.400 310.050 21.600 ;
        RECT 295.950 19.800 298.050 20.400 ;
        RECT 307.950 19.800 310.050 20.400 ;
        RECT 313.950 21.450 316.050 21.900 ;
        RECT 319.950 21.450 322.050 21.900 ;
        RECT 313.950 20.250 322.050 21.450 ;
        RECT 313.950 19.800 316.050 20.250 ;
        RECT 319.950 19.800 322.050 20.250 ;
        RECT 325.950 21.450 328.050 21.900 ;
        RECT 334.950 21.450 337.050 21.900 ;
        RECT 325.950 20.250 337.050 21.450 ;
        RECT 325.950 19.800 328.050 20.250 ;
        RECT 334.950 19.800 337.050 20.250 ;
        RECT 349.950 21.450 352.050 21.900 ;
        RECT 355.950 21.450 358.050 21.900 ;
        RECT 349.950 20.250 358.050 21.450 ;
        RECT 349.950 19.800 352.050 20.250 ;
        RECT 355.950 19.800 358.050 20.250 ;
        RECT 361.950 19.800 364.050 21.900 ;
        RECT 370.950 21.450 373.050 21.900 ;
        RECT 379.950 21.450 382.050 21.900 ;
        RECT 370.950 20.250 382.050 21.450 ;
        RECT 370.950 19.800 373.050 20.250 ;
        RECT 379.950 19.800 382.050 20.250 ;
        RECT 391.950 21.600 394.050 22.050 ;
        RECT 430.950 21.600 433.050 22.050 ;
        RECT 391.950 20.400 433.050 21.600 ;
        RECT 391.950 19.950 394.050 20.400 ;
        RECT 430.950 19.950 433.050 20.400 ;
        RECT 439.950 21.450 442.050 21.900 ;
        RECT 454.950 21.450 457.050 21.900 ;
        RECT 439.950 20.250 457.050 21.450 ;
        RECT 467.400 21.600 468.600 23.400 ;
        RECT 572.400 21.900 573.600 29.400 ;
        RECT 622.950 28.950 625.050 29.400 ;
        RECT 658.950 28.950 661.050 29.400 ;
        RECT 718.950 30.600 721.050 31.050 ;
        RECT 745.950 30.600 748.050 31.050 ;
        RECT 718.950 29.400 748.050 30.600 ;
        RECT 718.950 28.950 721.050 29.400 ;
        RECT 745.950 28.950 748.050 29.400 ;
        RECT 760.950 30.600 763.050 31.050 ;
        RECT 772.950 30.600 775.050 31.050 ;
        RECT 760.950 29.400 775.050 30.600 ;
        RECT 760.950 28.950 763.050 29.400 ;
        RECT 772.950 28.950 775.050 29.400 ;
        RECT 820.950 30.600 823.050 31.050 ;
        RECT 847.950 30.600 850.050 31.050 ;
        RECT 856.950 30.600 859.050 31.050 ;
        RECT 820.950 29.400 859.050 30.600 ;
        RECT 820.950 28.950 823.050 29.400 ;
        RECT 847.950 28.950 850.050 29.400 ;
        RECT 856.950 28.950 859.050 29.400 ;
        RECT 865.950 30.600 868.050 31.050 ;
        RECT 874.950 30.600 877.050 31.050 ;
        RECT 865.950 29.400 877.050 30.600 ;
        RECT 865.950 28.950 868.050 29.400 ;
        RECT 874.950 28.950 877.050 29.400 ;
        RECT 886.950 30.600 889.050 31.050 ;
        RECT 928.950 30.600 931.050 31.050 ;
        RECT 886.950 29.400 931.050 30.600 ;
        RECT 886.950 28.950 889.050 29.400 ;
        RECT 928.950 28.950 931.050 29.400 ;
        RECT 574.950 27.600 577.050 28.200 ;
        RECT 574.950 26.400 579.600 27.600 ;
        RECT 574.950 26.100 577.050 26.400 ;
        RECT 469.950 21.600 472.050 21.900 ;
        RECT 481.950 21.600 484.050 21.900 ;
        RECT 467.400 20.400 484.050 21.600 ;
        RECT 439.950 19.800 442.050 20.250 ;
        RECT 454.950 19.800 457.050 20.250 ;
        RECT 469.950 19.800 472.050 20.400 ;
        RECT 481.950 19.800 484.050 20.400 ;
        RECT 535.950 21.600 538.050 21.900 ;
        RECT 556.950 21.600 559.050 21.900 ;
        RECT 535.950 21.450 559.050 21.600 ;
        RECT 562.950 21.450 565.050 21.900 ;
        RECT 535.950 20.400 565.050 21.450 ;
        RECT 535.950 19.800 538.050 20.400 ;
        RECT 556.950 20.250 565.050 20.400 ;
        RECT 556.950 19.800 559.050 20.250 ;
        RECT 562.950 19.800 565.050 20.250 ;
        RECT 571.950 19.800 574.050 21.900 ;
        RECT 578.400 19.050 579.600 26.400 ;
        RECT 580.950 26.100 583.050 28.200 ;
        RECT 592.950 27.600 595.050 28.050 ;
        RECT 592.950 26.400 600.600 27.600 ;
        RECT 581.400 24.600 582.600 26.100 ;
        RECT 592.950 25.950 595.050 26.400 ;
        RECT 589.950 24.600 592.050 25.050 ;
        RECT 581.400 23.400 592.050 24.600 ;
        RECT 589.950 22.950 592.050 23.400 ;
        RECT 599.400 21.900 600.600 26.400 ;
        RECT 607.950 25.950 610.050 28.050 ;
        RECT 637.950 26.100 640.050 28.200 ;
        RECT 706.950 27.600 709.050 28.200 ;
        RECT 677.400 26.400 709.050 27.600 ;
        RECT 608.400 22.050 609.600 25.950 ;
        RECT 638.400 24.600 639.600 26.100 ;
        RECT 677.400 24.600 678.600 26.400 ;
        RECT 706.950 26.100 709.050 26.400 ;
        RECT 712.950 24.600 715.050 28.050 ;
        RECT 775.950 27.600 778.050 28.200 ;
        RECT 784.950 27.600 787.050 28.050 ;
        RECT 775.950 26.400 787.050 27.600 ;
        RECT 775.950 26.100 778.050 26.400 ;
        RECT 784.950 25.950 787.050 26.400 ;
        RECT 859.950 26.100 862.050 28.200 ;
        RECT 626.400 23.400 678.600 24.600 ;
        RECT 598.950 19.800 601.050 21.900 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 626.400 21.900 627.600 23.400 ;
        RECT 677.400 21.900 678.600 23.400 ;
        RECT 710.400 24.000 715.050 24.600 ;
        RECT 826.950 24.600 829.050 25.050 ;
        RECT 860.400 24.600 861.600 26.100 ;
        RECT 868.950 24.600 871.050 28.050 ;
        RECT 710.400 23.400 714.600 24.000 ;
        RECT 826.950 23.400 861.600 24.600 ;
        RECT 863.400 24.000 871.050 24.600 ;
        RECT 863.400 23.400 870.600 24.000 ;
        RECT 710.400 21.900 711.600 23.400 ;
        RECT 826.950 22.950 829.050 23.400 ;
        RECT 845.400 21.900 846.600 23.400 ;
        RECT 863.400 21.900 864.600 23.400 ;
        RECT 625.950 19.800 628.050 21.900 ;
        RECT 640.950 21.600 643.050 21.900 ;
        RECT 655.950 21.600 658.050 21.900 ;
        RECT 640.950 20.400 658.050 21.600 ;
        RECT 640.950 19.800 643.050 20.400 ;
        RECT 655.950 19.800 658.050 20.400 ;
        RECT 661.950 21.450 664.050 21.900 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 661.950 20.250 673.050 21.450 ;
        RECT 661.950 19.800 664.050 20.250 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 676.950 19.800 679.050 21.900 ;
        RECT 682.950 21.450 685.050 21.900 ;
        RECT 691.950 21.450 694.050 21.900 ;
        RECT 682.950 20.250 694.050 21.450 ;
        RECT 682.950 19.800 685.050 20.250 ;
        RECT 691.950 19.800 694.050 20.250 ;
        RECT 709.950 19.800 712.050 21.900 ;
        RECT 718.950 21.450 721.050 21.900 ;
        RECT 724.950 21.450 727.050 21.900 ;
        RECT 718.950 20.250 727.050 21.450 ;
        RECT 718.950 19.800 721.050 20.250 ;
        RECT 724.950 19.800 727.050 20.250 ;
        RECT 760.950 21.450 763.050 21.900 ;
        RECT 766.950 21.450 769.050 21.900 ;
        RECT 760.950 20.250 769.050 21.450 ;
        RECT 760.950 19.800 763.050 20.250 ;
        RECT 766.950 19.800 769.050 20.250 ;
        RECT 784.950 21.450 787.050 21.900 ;
        RECT 790.950 21.450 793.050 21.900 ;
        RECT 784.950 20.250 793.050 21.450 ;
        RECT 784.950 19.800 787.050 20.250 ;
        RECT 790.950 19.800 793.050 20.250 ;
        RECT 796.950 21.450 799.050 21.900 ;
        RECT 802.950 21.450 805.050 21.900 ;
        RECT 796.950 20.250 805.050 21.450 ;
        RECT 796.950 19.800 799.050 20.250 ;
        RECT 802.950 19.800 805.050 20.250 ;
        RECT 844.950 19.800 847.050 21.900 ;
        RECT 850.950 21.450 853.050 21.900 ;
        RECT 856.950 21.450 859.050 21.900 ;
        RECT 850.950 20.250 859.050 21.450 ;
        RECT 850.950 19.800 853.050 20.250 ;
        RECT 856.950 19.800 859.050 20.250 ;
        RECT 862.950 19.800 865.050 21.900 ;
        RECT 874.950 21.450 877.050 21.900 ;
        RECT 880.950 21.450 883.050 21.900 ;
        RECT 874.950 20.250 883.050 21.450 ;
        RECT 874.950 19.800 877.050 20.250 ;
        RECT 880.950 19.800 883.050 20.250 ;
        RECT 886.950 21.450 889.050 21.900 ;
        RECT 898.950 21.450 901.050 21.900 ;
        RECT 886.950 20.250 901.050 21.450 ;
        RECT 886.950 19.800 889.050 20.250 ;
        RECT 898.950 19.800 901.050 20.250 ;
        RECT 385.950 18.600 388.050 19.050 ;
        RECT 541.950 18.600 544.050 19.050 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 385.950 17.400 405.600 18.600 ;
        RECT 385.950 16.950 388.050 17.400 ;
        RECT 404.400 16.050 405.600 17.400 ;
        RECT 541.950 17.400 553.050 18.600 ;
        RECT 541.950 16.950 544.050 17.400 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 574.950 17.400 579.600 19.050 ;
        RECT 589.950 18.600 592.050 19.050 ;
        RECT 790.950 18.600 793.050 19.050 ;
        RECT 808.950 18.600 811.050 19.050 ;
        RECT 832.950 18.600 835.050 19.050 ;
        RECT 589.950 17.400 606.600 18.600 ;
        RECT 574.950 16.950 579.000 17.400 ;
        RECT 589.950 16.950 592.050 17.400 ;
        RECT 605.400 16.050 606.600 17.400 ;
        RECT 790.950 17.400 835.050 18.600 ;
        RECT 790.950 16.950 793.050 17.400 ;
        RECT 808.950 16.950 811.050 17.400 ;
        RECT 832.950 16.950 835.050 17.400 ;
        RECT 85.950 15.600 88.050 16.050 ;
        RECT 112.950 15.600 115.050 16.050 ;
        RECT 85.950 14.400 115.050 15.600 ;
        RECT 85.950 13.950 88.050 14.400 ;
        RECT 112.950 13.950 115.050 14.400 ;
        RECT 127.950 15.600 130.050 16.050 ;
        RECT 148.950 15.600 151.050 16.050 ;
        RECT 127.950 14.400 151.050 15.600 ;
        RECT 127.950 13.950 130.050 14.400 ;
        RECT 148.950 13.950 151.050 14.400 ;
        RECT 178.950 15.600 181.050 16.050 ;
        RECT 241.950 15.600 244.050 16.050 ;
        RECT 373.950 15.600 376.050 16.050 ;
        RECT 178.950 14.400 376.050 15.600 ;
        RECT 178.950 13.950 181.050 14.400 ;
        RECT 241.950 13.950 244.050 14.400 ;
        RECT 373.950 13.950 376.050 14.400 ;
        RECT 403.950 15.600 406.050 16.050 ;
        RECT 424.950 15.600 427.050 16.050 ;
        RECT 403.950 14.400 427.050 15.600 ;
        RECT 403.950 13.950 406.050 14.400 ;
        RECT 424.950 13.950 427.050 14.400 ;
        RECT 463.950 15.600 466.050 16.050 ;
        RECT 592.950 15.600 595.050 16.050 ;
        RECT 598.950 15.600 601.050 16.050 ;
        RECT 463.950 14.400 501.600 15.600 ;
        RECT 463.950 13.950 466.050 14.400 ;
        RECT 223.950 12.600 226.050 13.050 ;
        RECT 238.950 12.600 241.050 13.050 ;
        RECT 223.950 11.400 241.050 12.600 ;
        RECT 223.950 10.950 226.050 11.400 ;
        RECT 238.950 10.950 241.050 11.400 ;
        RECT 322.950 12.600 325.050 13.050 ;
        RECT 391.950 12.600 394.050 13.050 ;
        RECT 322.950 11.400 394.050 12.600 ;
        RECT 322.950 10.950 325.050 11.400 ;
        RECT 391.950 10.950 394.050 11.400 ;
        RECT 430.950 12.600 433.050 13.050 ;
        RECT 493.950 12.600 496.050 13.050 ;
        RECT 430.950 11.400 496.050 12.600 ;
        RECT 500.400 12.600 501.600 14.400 ;
        RECT 592.950 14.400 601.050 15.600 ;
        RECT 592.950 13.950 595.050 14.400 ;
        RECT 598.950 13.950 601.050 14.400 ;
        RECT 604.950 15.600 607.050 16.050 ;
        RECT 640.950 15.600 643.050 16.050 ;
        RECT 604.950 14.400 643.050 15.600 ;
        RECT 604.950 13.950 607.050 14.400 ;
        RECT 640.950 13.950 643.050 14.400 ;
        RECT 715.950 15.600 718.050 16.050 ;
        RECT 730.950 15.600 733.050 16.050 ;
        RECT 742.950 15.600 745.050 16.050 ;
        RECT 715.950 14.400 745.050 15.600 ;
        RECT 715.950 13.950 718.050 14.400 ;
        RECT 730.950 13.950 733.050 14.400 ;
        RECT 742.950 13.950 745.050 14.400 ;
        RECT 838.950 15.600 841.050 16.050 ;
        RECT 871.950 15.600 874.050 16.050 ;
        RECT 838.950 14.400 874.050 15.600 ;
        RECT 838.950 13.950 841.050 14.400 ;
        RECT 871.950 13.950 874.050 14.400 ;
        RECT 901.950 15.600 904.050 16.050 ;
        RECT 931.950 15.600 934.050 16.050 ;
        RECT 901.950 14.400 934.050 15.600 ;
        RECT 901.950 13.950 904.050 14.400 ;
        RECT 931.950 13.950 934.050 14.400 ;
        RECT 574.950 12.600 577.050 13.050 ;
        RECT 500.400 11.400 577.050 12.600 ;
        RECT 430.950 10.950 433.050 11.400 ;
        RECT 493.950 10.950 496.050 11.400 ;
        RECT 574.950 10.950 577.050 11.400 ;
        RECT 619.950 12.600 622.050 13.050 ;
        RECT 670.950 12.600 673.050 13.050 ;
        RECT 619.950 11.400 673.050 12.600 ;
        RECT 619.950 10.950 622.050 11.400 ;
        RECT 670.950 10.950 673.050 11.400 ;
        RECT 577.950 9.600 580.050 10.050 ;
        RECT 610.950 9.600 613.050 10.050 ;
        RECT 577.950 8.400 613.050 9.600 ;
        RECT 577.950 7.950 580.050 8.400 ;
        RECT 610.950 7.950 613.050 8.400 ;
        RECT 703.950 9.600 706.050 10.050 ;
        RECT 736.950 9.600 739.050 10.050 ;
        RECT 703.950 8.400 739.050 9.600 ;
        RECT 703.950 7.950 706.050 8.400 ;
        RECT 736.950 7.950 739.050 8.400 ;
        RECT 895.950 9.600 898.050 10.050 ;
        RECT 910.950 9.600 913.050 10.050 ;
        RECT 895.950 8.400 913.050 9.600 ;
        RECT 895.950 7.950 898.050 8.400 ;
        RECT 910.950 7.950 913.050 8.400 ;
        RECT 112.950 6.600 115.050 7.050 ;
        RECT 157.950 6.600 160.050 7.050 ;
        RECT 112.950 5.400 160.050 6.600 ;
        RECT 112.950 4.950 115.050 5.400 ;
        RECT 157.950 4.950 160.050 5.400 ;
        RECT 475.950 6.600 478.050 7.050 ;
        RECT 505.950 6.600 508.050 7.050 ;
        RECT 475.950 5.400 508.050 6.600 ;
        RECT 475.950 4.950 478.050 5.400 ;
        RECT 505.950 4.950 508.050 5.400 ;
  END
END ALU_wrapper
END LIBRARY

