/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module ALU_wrapper(
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    output Done_o,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input clk,
    input reset
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire BI_0_bF$buf0 ;
wire BI_0_bF$buf1 ;
wire BI_0_bF$buf2 ;
wire BI_0_bF$buf3 ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire \u_ALU.AI7  ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire ABCmd_i_2_bF$buf0 ;
wire ABCmd_i_2_bF$buf1 ;
wire ABCmd_i_2_bF$buf2 ;
wire ABCmd_i_2_bF$buf3 ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _705__bF$buf0 ;
wire _705__bF$buf1 ;
wire _705__bF$buf2 ;
wire _705__bF$buf3 ;
wire _878_ ;
wire _458_ ;
wire _32__bF$buf0 ;
wire _32__bF$buf1 ;
wire _32__bF$buf2 ;
wire _32__bF$buf3 ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire Done_o ;
wire _740_ ;
wire _320_ ;
wire AI_5_bF$buf0 ;
wire AI_5_bF$buf1 ;
wire AI_5_bF$buf2 ;
wire AI_5_bF$buf3 ;
wire _56_ ;
wire _605_ ;
wire BI_4_bF$buf0 ;
wire BI_4_bF$buf1 ;
wire BI_4_bF$buf2 ;
wire BI_4_bF$buf3 ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire [7:0] _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _713_ ;
wire [7:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire BI_1_bF$buf0 ;
wire BI_1_bF$buf1 ;
wire BI_1_bF$buf2 ;
wire BI_1_bF$buf3 ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [2:0] state ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire BI_3_bF$buf0 ;
wire BI_3_bF$buf1 ;
wire BI_3_bF$buf2 ;
wire BI_3_bF$buf3 ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire [2:0] _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _0__bF$buf0 ;
wire _0__bF$buf1 ;
wire _0__bF$buf2 ;
wire _0__bF$buf3 ;
wire _0__bF$buf4 ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert41 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf0)
);

BUFX2 BUFX2_insert40 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf1)
);

BUFX2 BUFX2_insert39 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf2)
);

BUFX2 BUFX2_insert38 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf3)
);

BUFX2 BUFX2_insert37 (
    .A(BI[1]),
    .Y(BI_1_bF$buf0)
);

BUFX2 BUFX2_insert36 (
    .A(BI[1]),
    .Y(BI_1_bF$buf1)
);

BUFX2 BUFX2_insert35 (
    .A(BI[1]),
    .Y(BI_1_bF$buf2)
);

BUFX2 BUFX2_insert34 (
    .A(BI[1]),
    .Y(BI_1_bF$buf3)
);

BUFX2 BUFX2_insert33 (
    .A(BI[4]),
    .Y(BI_4_bF$buf0)
);

BUFX2 BUFX2_insert32 (
    .A(BI[4]),
    .Y(BI_4_bF$buf1)
);

BUFX2 BUFX2_insert31 (
    .A(BI[4]),
    .Y(BI_4_bF$buf2)
);

BUFX2 BUFX2_insert30 (
    .A(BI[4]),
    .Y(BI_4_bF$buf3)
);

BUFX2 BUFX2_insert29 (
    .A(_32_),
    .Y(_32__bF$buf0)
);

BUFX2 BUFX2_insert28 (
    .A(_32_),
    .Y(_32__bF$buf1)
);

BUFX2 BUFX2_insert27 (
    .A(_32_),
    .Y(_32__bF$buf2)
);

BUFX2 BUFX2_insert26 (
    .A(_32_),
    .Y(_32__bF$buf3)
);

BUFX2 BUFX2_insert25 (
    .A(AI[5]),
    .Y(AI_5_bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .A(AI[5]),
    .Y(AI_5_bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .A(AI[5]),
    .Y(AI_5_bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .A(AI[5]),
    .Y(AI_5_bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .A(_0_),
    .Y(_0__bF$buf0)
);

BUFX2 BUFX2_insert20 (
    .A(_0_),
    .Y(_0__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .A(_0_),
    .Y(_0__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .A(_0_),
    .Y(_0__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .A(_0_),
    .Y(_0__bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .A(_705_),
    .Y(_705__bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .A(_705_),
    .Y(_705__bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .A(_705_),
    .Y(_705__bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .A(_705_),
    .Y(_705__bF$buf3)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .A(BI[0]),
    .Y(BI_0_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .A(BI[0]),
    .Y(BI_0_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .A(BI[0]),
    .Y(BI_0_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .A(BI[0]),
    .Y(BI_0_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .A(BI[3]),
    .Y(BI_3_bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .A(BI[3]),
    .Y(BI_3_bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .A(BI[3]),
    .Y(BI_3_bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .A(BI[3]),
    .Y(BI_3_bF$buf3)
);

INVX1 _1000_ (
    .A(_105_),
    .Y(_106_)
);

AND2X2 _1001_ (
    .A(BI_3_bF$buf3),
    .B(AI[2]),
    .Y(_107_)
);

NAND2X1 _1002_ (
    .A(_60_),
    .B(_107_),
    .Y(_108_)
);

INVX1 _1003_ (
    .A(AI[2]),
    .Y(_109_)
);

OAI21X1 _1004_ (
    .A(_58_),
    .B(_109_),
    .C(_82_),
    .Y(_110_)
);

NAND3X1 _1005_ (
    .A(_110_),
    .B(_106_),
    .C(_108_),
    .Y(_111_)
);

OAI21X1 _1006_ (
    .A(_58_),
    .B(_109_),
    .C(_60_),
    .Y(_112_)
);

INVX1 _1007_ (
    .A(AI[1]),
    .Y(_113_)
);

OAI21X1 _1008_ (
    .A(_83_),
    .B(_113_),
    .C(_107_),
    .Y(_114_)
);

NAND3X1 _1009_ (
    .A(_105_),
    .B(_112_),
    .C(_114_),
    .Y(_115_)
);

AND2X2 _1010_ (
    .A(_115_),
    .B(_111_),
    .Y(_116_)
);

NAND3X1 _1011_ (
    .A(_100_),
    .B(_104_),
    .C(_116_),
    .Y(_117_)
);

AOI21X1 _1012_ (
    .A(_102_),
    .B(_103_),
    .C(_101_),
    .Y(_118_)
);

AOI21X1 _1013_ (
    .A(_99_),
    .B(_96_),
    .C(_89_),
    .Y(_119_)
);

NAND2X1 _1014_ (
    .A(_111_),
    .B(_115_),
    .Y(_120_)
);

OAI21X1 _1015_ (
    .A(_118_),
    .B(_119_),
    .C(_120_),
    .Y(_121_)
);

NAND3X1 _1016_ (
    .A(_117_),
    .B(_121_),
    .C(_88_),
    .Y(_122_)
);

AOI21X1 _1017_ (
    .A(_121_),
    .B(_117_),
    .C(_88_),
    .Y(_123_)
);

OAI21X1 _1018_ (
    .A(_61_),
    .B(_123_),
    .C(_122_),
    .Y(_124_)
);

AOI21X1 _1019_ (
    .A(_104_),
    .B(_116_),
    .C(_118_),
    .Y(_125_)
);

OAI21X1 _1020_ (
    .A(_92_),
    .B(_94_),
    .C(_91_),
    .Y(_126_)
);

AND2X2 _1021_ (
    .A(BI_1_bF$buf3),
    .B(AI[6]),
    .Y(_127_)
);

NAND2X1 _1022_ (
    .A(_90_),
    .B(_127_),
    .Y(_128_)
);

INVX1 _1023_ (
    .A(BI_1_bF$buf2),
    .Y(_129_)
);

INVX2 _1024_ (
    .A(AI_5_bF$buf3),
    .Y(_130_)
);

NAND2X1 _1025_ (
    .A(BI_0_bF$buf3),
    .B(AI[6]),
    .Y(_131_)
);

OAI21X1 _1026_ (
    .A(_129_),
    .B(_130_),
    .C(_131_),
    .Y(_132_)
);

NAND2X1 _1027_ (
    .A(BI[2]),
    .B(AI[4]),
    .Y(_133_)
);

INVX1 _1028_ (
    .A(_133_),
    .Y(_134_)
);

NAND3X1 _1029_ (
    .A(_132_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

NOR2X1 _1030_ (
    .A(_97_),
    .B(_131_),
    .Y(_136_)
);

AOI22X1 _1031_ (
    .A(BI_0_bF$buf2),
    .B(AI[6]),
    .C(BI_1_bF$buf1),
    .D(AI_5_bF$buf2),
    .Y(_137_)
);

OAI21X1 _1032_ (
    .A(_137_),
    .B(_136_),
    .C(_133_),
    .Y(_138_)
);

AOI21X1 _1033_ (
    .A(_138_),
    .B(_135_),
    .C(_126_),
    .Y(_139_)
);

AOI21X1 _1034_ (
    .A(_93_),
    .B(_95_),
    .C(_98_),
    .Y(_140_)
);

OAI21X1 _1035_ (
    .A(_137_),
    .B(_136_),
    .C(_134_),
    .Y(_141_)
);

NAND3X1 _1036_ (
    .A(_132_),
    .B(_133_),
    .C(_128_),
    .Y(_142_)
);

AOI21X1 _1037_ (
    .A(_141_),
    .B(_142_),
    .C(_140_),
    .Y(_143_)
);

NAND2X1 _1038_ (
    .A(BI[5]),
    .B(AI[1]),
    .Y(_144_)
);

INVX1 _1039_ (
    .A(_144_),
    .Y(_145_)
);

AND2X2 _1040_ (
    .A(BI_4_bF$buf3),
    .B(AI[2]),
    .Y(_146_)
);

AND2X2 _1041_ (
    .A(BI_3_bF$buf2),
    .B(AI[3]),
    .Y(_147_)
);

NAND2X1 _1042_ (
    .A(_146_),
    .B(_147_),
    .Y(_148_)
);

INVX2 _1043_ (
    .A(AI[3]),
    .Y(_149_)
);

NAND2X1 _1044_ (
    .A(BI_4_bF$buf2),
    .B(AI[2]),
    .Y(_150_)
);

OAI21X1 _1045_ (
    .A(_58_),
    .B(_149_),
    .C(_150_),
    .Y(_151_)
);

NAND3X1 _1046_ (
    .A(_151_),
    .B(_145_),
    .C(_148_),
    .Y(_152_)
);

OAI21X1 _1047_ (
    .A(_58_),
    .B(_149_),
    .C(_146_),
    .Y(_153_)
);

OAI21X1 _1048_ (
    .A(_83_),
    .B(_109_),
    .C(_147_),
    .Y(_154_)
);

NAND3X1 _1049_ (
    .A(_144_),
    .B(_153_),
    .C(_154_),
    .Y(_155_)
);

AND2X2 _1050_ (
    .A(_155_),
    .B(_152_),
    .Y(_156_)
);

OAI21X1 _1051_ (
    .A(_139_),
    .B(_143_),
    .C(_156_),
    .Y(_157_)
);

NAND3X1 _1052_ (
    .A(_142_),
    .B(_141_),
    .C(_140_),
    .Y(_158_)
);

NAND3X1 _1053_ (
    .A(_126_),
    .B(_135_),
    .C(_138_),
    .Y(_159_)
);

NAND2X1 _1054_ (
    .A(_152_),
    .B(_155_),
    .Y(_160_)
);

NAND3X1 _1055_ (
    .A(_160_),
    .B(_159_),
    .C(_158_),
    .Y(_161_)
);

NAND3X1 _1056_ (
    .A(_161_),
    .B(_125_),
    .C(_157_),
    .Y(_162_)
);

OAI21X1 _1057_ (
    .A(_120_),
    .B(_119_),
    .C(_100_),
    .Y(_163_)
);

NAND3X1 _1058_ (
    .A(_159_),
    .B(_158_),
    .C(_156_),
    .Y(_164_)
);

OAI21X1 _1059_ (
    .A(_139_),
    .B(_143_),
    .C(_160_),
    .Y(_165_)
);

NAND3X1 _1060_ (
    .A(_164_),
    .B(_165_),
    .C(_163_),
    .Y(_166_)
);

INVX4 _1061_ (
    .A(BI[6]),
    .Y(_167_)
);

NOR2X1 _1062_ (
    .A(_57_),
    .B(_167_),
    .Y(_168_)
);

OAI21X1 _1063_ (
    .A(_84_),
    .B(_150_),
    .C(_111_),
    .Y(_169_)
);

XNOR2X1 _1064_ (
    .A(_169_),
    .B(_168_),
    .Y(_170_)
);

INVX1 _1065_ (
    .A(_170_),
    .Y(_171_)
);

NAND3X1 _1066_ (
    .A(_162_),
    .B(_166_),
    .C(_171_),
    .Y(_172_)
);

AOI21X1 _1067_ (
    .A(_165_),
    .B(_164_),
    .C(_163_),
    .Y(_173_)
);

AOI21X1 _1068_ (
    .A(_157_),
    .B(_161_),
    .C(_125_),
    .Y(_174_)
);

OAI21X1 _1069_ (
    .A(_174_),
    .B(_173_),
    .C(_170_),
    .Y(_175_)
);

NAND3X1 _1070_ (
    .A(_172_),
    .B(_175_),
    .C(_124_),
    .Y(_176_)
);

NAND2X1 _1071_ (
    .A(_168_),
    .B(_169_),
    .Y(_177_)
);

INVX1 _1072_ (
    .A(_177_),
    .Y(_178_)
);

OAI21X1 _1073_ (
    .A(_170_),
    .B(_173_),
    .C(_166_),
    .Y(_179_)
);

AOI21X1 _1074_ (
    .A(_158_),
    .B(_156_),
    .C(_143_),
    .Y(_180_)
);

OAI21X1 _1075_ (
    .A(_137_),
    .B(_133_),
    .C(_128_),
    .Y(_181_)
);

NAND3X1 _1076_ (
    .A(BI_0_bF$buf1),
    .B(\u_ALU.AI7 ),
    .C(_127_),
    .Y(_182_)
);

AOI22X1 _1077_ (
    .A(BI_0_bF$buf0),
    .B(\u_ALU.AI7 ),
    .C(BI_1_bF$buf0),
    .D(AI[6]),
    .Y(_183_)
);

INVX1 _1078_ (
    .A(_183_),
    .Y(_184_)
);

NAND2X1 _1079_ (
    .A(BI[2]),
    .B(AI_5_bF$buf1),
    .Y(_185_)
);

INVX1 _1080_ (
    .A(_185_),
    .Y(_186_)
);

NAND3X1 _1081_ (
    .A(_184_),
    .B(_186_),
    .C(_182_),
    .Y(_187_)
);

NAND2X1 _1082_ (
    .A(BI_1_bF$buf3),
    .B(\u_ALU.AI7 ),
    .Y(_188_)
);

NOR2X1 _1083_ (
    .A(_131_),
    .B(_188_),
    .Y(_189_)
);

OAI21X1 _1084_ (
    .A(_183_),
    .B(_189_),
    .C(_185_),
    .Y(_190_)
);

AOI21X1 _1085_ (
    .A(_190_),
    .B(_187_),
    .C(_181_),
    .Y(_191_)
);

OAI21X1 _1086_ (
    .A(_183_),
    .B(_189_),
    .C(_186_),
    .Y(_192_)
);

NAND3X1 _1087_ (
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_193_)
);

AOI22X1 _1088_ (
    .A(_128_),
    .B(_135_),
    .C(_192_),
    .D(_193_),
    .Y(_194_)
);

NAND2X1 _1089_ (
    .A(BI[5]),
    .B(AI[2]),
    .Y(_195_)
);

INVX1 _1090_ (
    .A(_195_),
    .Y(_196_)
);

AND2X2 _1091_ (
    .A(BI_4_bF$buf1),
    .B(AI[3]),
    .Y(_197_)
);

AND2X2 _1092_ (
    .A(BI_3_bF$buf1),
    .B(AI[4]),
    .Y(_198_)
);

NAND2X1 _1093_ (
    .A(_197_),
    .B(_198_),
    .Y(_199_)
);

AOI22X1 _1094_ (
    .A(BI_3_bF$buf0),
    .B(AI[4]),
    .C(BI_4_bF$buf0),
    .D(AI[3]),
    .Y(_200_)
);

INVX1 _1095_ (
    .A(_200_),
    .Y(_201_)
);

NAND3X1 _1096_ (
    .A(_196_),
    .B(_201_),
    .C(_199_),
    .Y(_202_)
);

OAI21X1 _1097_ (
    .A(_58_),
    .B(_74_),
    .C(_197_),
    .Y(_203_)
);

OAI21X1 _1098_ (
    .A(_83_),
    .B(_149_),
    .C(_198_),
    .Y(_204_)
);

NAND3X1 _1099_ (
    .A(_195_),
    .B(_203_),
    .C(_204_),
    .Y(_205_)
);

AND2X2 _1100_ (
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

OAI21X1 _1101_ (
    .A(_194_),
    .B(_191_),
    .C(_206_),
    .Y(_207_)
);

AOI21X1 _1102_ (
    .A(_132_),
    .B(_134_),
    .C(_136_),
    .Y(_208_)
);

NAND3X1 _1103_ (
    .A(_193_),
    .B(_192_),
    .C(_208_),
    .Y(_209_)
);

NAND3X1 _1104_ (
    .A(_181_),
    .B(_187_),
    .C(_190_),
    .Y(_210_)
);

NAND2X1 _1105_ (
    .A(_202_),
    .B(_205_),
    .Y(_211_)
);

NAND3X1 _1106_ (
    .A(_211_),
    .B(_210_),
    .C(_209_),
    .Y(_212_)
);

NAND3X1 _1107_ (
    .A(_212_),
    .B(_207_),
    .C(_180_),
    .Y(_213_)
);

OAI21X1 _1108_ (
    .A(_160_),
    .B(_139_),
    .C(_159_),
    .Y(_214_)
);

NAND3X1 _1109_ (
    .A(_210_),
    .B(_209_),
    .C(_206_),
    .Y(_215_)
);

OAI21X1 _1110_ (
    .A(_194_),
    .B(_191_),
    .C(_211_),
    .Y(_216_)
);

NAND3X1 _1111_ (
    .A(_215_),
    .B(_214_),
    .C(_216_),
    .Y(_217_)
);

NAND2X1 _1112_ (
    .A(AI[0]),
    .B(BI[7]),
    .Y(_218_)
);

INVX1 _1113_ (
    .A(_218_),
    .Y(_219_)
);

AOI22X1 _1114_ (
    .A(_107_),
    .B(_197_),
    .C(_151_),
    .D(_145_),
    .Y(_220_)
);

INVX1 _1115_ (
    .A(_220_),
    .Y(_221_)
);

OAI21X1 _1116_ (
    .A(_167_),
    .B(_113_),
    .C(_221_),
    .Y(_222_)
);

NOR2X1 _1117_ (
    .A(_167_),
    .B(_113_),
    .Y(_223_)
);

NAND2X1 _1118_ (
    .A(_223_),
    .B(_220_),
    .Y(_224_)
);

NAND3X1 _1119_ (
    .A(_219_),
    .B(_224_),
    .C(_222_),
    .Y(_225_)
);

NAND2X1 _1120_ (
    .A(_223_),
    .B(_221_),
    .Y(_226_)
);

OAI21X1 _1121_ (
    .A(_167_),
    .B(_113_),
    .C(_220_),
    .Y(_227_)
);

NAND3X1 _1122_ (
    .A(_218_),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

NAND2X1 _1123_ (
    .A(_228_),
    .B(_225_),
    .Y(_229_)
);

NAND3X1 _1124_ (
    .A(_229_),
    .B(_213_),
    .C(_217_),
    .Y(_230_)
);

AOI21X1 _1125_ (
    .A(_216_),
    .B(_215_),
    .C(_214_),
    .Y(_231_)
);

AOI21X1 _1126_ (
    .A(_207_),
    .B(_212_),
    .C(_180_),
    .Y(_232_)
);

NAND3X1 _1127_ (
    .A(_219_),
    .B(_227_),
    .C(_226_),
    .Y(_233_)
);

NAND3X1 _1128_ (
    .A(_218_),
    .B(_224_),
    .C(_222_),
    .Y(_234_)
);

NAND2X1 _1129_ (
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

OAI21X1 _1130_ (
    .A(_231_),
    .B(_232_),
    .C(_235_),
    .Y(_236_)
);

AOI21X1 _1131_ (
    .A(_236_),
    .B(_230_),
    .C(_179_),
    .Y(_237_)
);

AOI21X1 _1132_ (
    .A(_162_),
    .B(_171_),
    .C(_174_),
    .Y(_238_)
);

OAI21X1 _1133_ (
    .A(_231_),
    .B(_232_),
    .C(_229_),
    .Y(_239_)
);

NAND3X1 _1134_ (
    .A(_235_),
    .B(_213_),
    .C(_217_),
    .Y(_240_)
);

AOI21X1 _1135_ (
    .A(_239_),
    .B(_240_),
    .C(_238_),
    .Y(_241_)
);

OAI21X1 _1136_ (
    .A(_241_),
    .B(_237_),
    .C(_178_),
    .Y(_242_)
);

NAND3X1 _1137_ (
    .A(_240_),
    .B(_239_),
    .C(_238_),
    .Y(_243_)
);

NAND3X1 _1138_ (
    .A(_230_),
    .B(_236_),
    .C(_179_),
    .Y(_244_)
);

NAND3X1 _1139_ (
    .A(_177_),
    .B(_243_),
    .C(_244_),
    .Y(_245_)
);

AOI21X1 _1140_ (
    .A(_242_),
    .B(_245_),
    .C(_176_),
    .Y(_246_)
);

INVX1 _1141_ (
    .A(_246_),
    .Y(_247_)
);

INVX1 _1142_ (
    .A(_61_),
    .Y(_248_)
);

NOR2X1 _1143_ (
    .A(_62_),
    .B(_63_),
    .Y(_249_)
);

INVX1 _1144_ (
    .A(_65_),
    .Y(_250_)
);

OAI21X1 _1145_ (
    .A(_73_),
    .B(_149_),
    .C(_62_),
    .Y(_251_)
);

AOI21X1 _1146_ (
    .A(_250_),
    .B(_251_),
    .C(_249_),
    .Y(_252_)
);

OAI21X1 _1147_ (
    .A(_77_),
    .B(_78_),
    .C(_69_),
    .Y(_253_)
);

NAND3X1 _1148_ (
    .A(_68_),
    .B(_75_),
    .C(_72_),
    .Y(_254_)
);

AOI21X1 _1149_ (
    .A(_254_),
    .B(_253_),
    .C(_252_),
    .Y(_255_)
);

AND2X2 _1150_ (
    .A(_61_),
    .B(_85_),
    .Y(_256_)
);

NAND3X1 _1151_ (
    .A(_252_),
    .B(_253_),
    .C(_254_),
    .Y(_257_)
);

AOI21X1 _1152_ (
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

OAI21X1 _1153_ (
    .A(_118_),
    .B(_119_),
    .C(_116_),
    .Y(_259_)
);

NAND3X1 _1154_ (
    .A(_120_),
    .B(_100_),
    .C(_104_),
    .Y(_260_)
);

NAND3X1 _1155_ (
    .A(_260_),
    .B(_259_),
    .C(_258_),
    .Y(_261_)
);

NAND3X1 _1156_ (
    .A(_248_),
    .B(_122_),
    .C(_261_),
    .Y(_262_)
);

OAI21X1 _1157_ (
    .A(_174_),
    .B(_173_),
    .C(_171_),
    .Y(_263_)
);

NAND3X1 _1158_ (
    .A(_170_),
    .B(_162_),
    .C(_166_),
    .Y(_264_)
);

AOI22X1 _1159_ (
    .A(_122_),
    .B(_262_),
    .C(_263_),
    .D(_264_),
    .Y(_265_)
);

NAND3X1 _1160_ (
    .A(_178_),
    .B(_243_),
    .C(_244_),
    .Y(_266_)
);

OAI21X1 _1161_ (
    .A(_241_),
    .B(_237_),
    .C(_177_),
    .Y(_267_)
);

AOI21X1 _1162_ (
    .A(_267_),
    .B(_266_),
    .C(_265_),
    .Y(_268_)
);

NAND3X1 _1163_ (
    .A(_256_),
    .B(_257_),
    .C(_80_),
    .Y(_269_)
);

NAND3X1 _1164_ (
    .A(_251_),
    .B(_250_),
    .C(_64_),
    .Y(_270_)
);

NAND2X1 _1165_ (
    .A(BI_0_bF$buf3),
    .B(AI[1]),
    .Y(_271_)
);

OR2X2 _1166_ (
    .A(_62_),
    .B(_271_),
    .Y(_272_)
);

NAND2X1 _1167_ (
    .A(AI[0]),
    .B(BI[2]),
    .Y(_273_)
);

AOI22X1 _1168_ (
    .A(BI_0_bF$buf2),
    .B(AI[2]),
    .C(BI_1_bF$buf2),
    .D(AI[1]),
    .Y(_274_)
);

OAI21X1 _1169_ (
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(_275_)
);

OAI21X1 _1170_ (
    .A(_249_),
    .B(_66_),
    .C(_65_),
    .Y(_276_)
);

NAND3X1 _1171_ (
    .A(_276_),
    .B(_275_),
    .C(_270_),
    .Y(_277_)
);

AOI21X1 _1172_ (
    .A(_270_),
    .B(_276_),
    .C(_275_),
    .Y(_278_)
);

OAI21X1 _1173_ (
    .A(_81_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

OAI21X1 _1174_ (
    .A(_255_),
    .B(_87_),
    .C(_86_),
    .Y(_280_)
);

NAND3X1 _1175_ (
    .A(_269_),
    .B(_279_),
    .C(_280_),
    .Y(_281_)
);

INVX1 _1176_ (
    .A(_281_),
    .Y(_282_)
);

AOI22X1 _1177_ (
    .A(_80_),
    .B(_269_),
    .C(_259_),
    .D(_260_),
    .Y(_283_)
);

OAI21X1 _1178_ (
    .A(_283_),
    .B(_123_),
    .C(_61_),
    .Y(_284_)
);

NAND3X1 _1179_ (
    .A(_262_),
    .B(_282_),
    .C(_284_),
    .Y(_285_)
);

AOI21X1 _1180_ (
    .A(_175_),
    .B(_172_),
    .C(_124_),
    .Y(_286_)
);

NOR3X1 _1181_ (
    .A(_285_),
    .B(_265_),
    .C(_286_),
    .Y(_287_)
);

INVX1 _1182_ (
    .A(_278_),
    .Y(_288_)
);

NAND3X1 _1183_ (
    .A(_59_),
    .B(_277_),
    .C(_288_),
    .Y(_289_)
);

INVX1 _1184_ (
    .A(_274_),
    .Y(_290_)
);

OAI21X1 _1185_ (
    .A(_62_),
    .B(_271_),
    .C(_290_),
    .Y(_291_)
);

OR2X2 _1186_ (
    .A(_291_),
    .B(_273_),
    .Y(_292_)
);

NAND2X1 _1187_ (
    .A(AI[0]),
    .B(BI_1_bF$buf1),
    .Y(_293_)
);

NOR2X1 _1188_ (
    .A(_271_),
    .B(_293_),
    .Y(_294_)
);

INVX1 _1189_ (
    .A(BI[2]),
    .Y(_295_)
);

OAI21X1 _1190_ (
    .A(_57_),
    .B(_295_),
    .C(_291_),
    .Y(_296_)
);

NAND3X1 _1191_ (
    .A(_294_),
    .B(_296_),
    .C(_292_),
    .Y(_297_)
);

INVX1 _1192_ (
    .A(_297_),
    .Y(_298_)
);

INVX1 _1193_ (
    .A(_277_),
    .Y(_299_)
);

OAI21X1 _1194_ (
    .A(_278_),
    .B(_299_),
    .C(_81_),
    .Y(_300_)
);

NAND3X1 _1195_ (
    .A(_298_),
    .B(_289_),
    .C(_300_),
    .Y(_301_)
);

AOI21X1 _1196_ (
    .A(_280_),
    .B(_269_),
    .C(_279_),
    .Y(_302_)
);

NOR3X1 _1197_ (
    .A(_302_),
    .B(_301_),
    .C(_282_),
    .Y(_303_)
);

OAI21X1 _1198_ (
    .A(_283_),
    .B(_123_),
    .C(_248_),
    .Y(_304_)
);

NAND3X1 _1199_ (
    .A(_61_),
    .B(_122_),
    .C(_261_),
    .Y(_305_)
);

NAND3X1 _1200_ (
    .A(_281_),
    .B(_305_),
    .C(_304_),
    .Y(_306_)
);

NAND3X1 _1201_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_307_)
);

INVX1 _1202_ (
    .A(_307_),
    .Y(_308_)
);

OAI21X1 _1203_ (
    .A(_265_),
    .B(_286_),
    .C(_285_),
    .Y(_309_)
);

AOI21X1 _1204_ (
    .A(_308_),
    .B(_309_),
    .C(_287_),
    .Y(_310_)
);

OAI21X1 _1205_ (
    .A(_268_),
    .B(_310_),
    .C(_247_),
    .Y(_311_)
);

AOI21X1 _1206_ (
    .A(_178_),
    .B(_243_),
    .C(_241_),
    .Y(_312_)
);

NAND2X1 _1207_ (
    .A(_226_),
    .B(_233_),
    .Y(_313_)
);

OAI21X1 _1208_ (
    .A(_235_),
    .B(_231_),
    .C(_217_),
    .Y(_314_)
);

NAND2X1 _1209_ (
    .A(BI[7]),
    .B(AI[1]),
    .Y(_315_)
);

INVX1 _1210_ (
    .A(_315_),
    .Y(_316_)
);

NOR2X1 _1211_ (
    .A(_109_),
    .B(_167_),
    .Y(_317_)
);

OAI21X1 _1212_ (
    .A(_195_),
    .B(_200_),
    .C(_199_),
    .Y(_318_)
);

NAND2X1 _1213_ (
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

OR2X2 _1214_ (
    .A(_318_),
    .B(_317_),
    .Y(_320_)
);

NAND3X1 _1215_ (
    .A(_316_),
    .B(_319_),
    .C(_320_),
    .Y(_321_)
);

AND2X2 _1216_ (
    .A(_318_),
    .B(_317_),
    .Y(_322_)
);

NOR2X1 _1217_ (
    .A(_317_),
    .B(_318_),
    .Y(_323_)
);

OAI21X1 _1218_ (
    .A(_323_),
    .B(_322_),
    .C(_315_),
    .Y(_324_)
);

NAND2X1 _1219_ (
    .A(_324_),
    .B(_321_),
    .Y(_325_)
);

AOI21X1 _1220_ (
    .A(_206_),
    .B(_209_),
    .C(_194_),
    .Y(_326_)
);

NAND2X1 _1221_ (
    .A(BI[5]),
    .B(AI[3]),
    .Y(_327_)
);

AND2X2 _1222_ (
    .A(BI_4_bF$buf3),
    .B(AI[4]),
    .Y(_328_)
);

OAI21X1 _1223_ (
    .A(_130_),
    .B(_58_),
    .C(_328_),
    .Y(_329_)
);

AND2X2 _1224_ (
    .A(AI_5_bF$buf0),
    .B(BI_3_bF$buf3),
    .Y(_330_)
);

OAI21X1 _1225_ (
    .A(_83_),
    .B(_74_),
    .C(_330_),
    .Y(_331_)
);

NAND3X1 _1226_ (
    .A(_327_),
    .B(_329_),
    .C(_331_),
    .Y(_332_)
);

INVX1 _1227_ (
    .A(_327_),
    .Y(_333_)
);

NAND2X1 _1228_ (
    .A(_328_),
    .B(_330_),
    .Y(_334_)
);

AOI22X1 _1229_ (
    .A(AI_5_bF$buf3),
    .B(BI_3_bF$buf2),
    .C(BI_4_bF$buf2),
    .D(AI[4]),
    .Y(_335_)
);

INVX1 _1230_ (
    .A(_335_),
    .Y(_336_)
);

NAND3X1 _1231_ (
    .A(_333_),
    .B(_336_),
    .C(_334_),
    .Y(_337_)
);

NAND2X1 _1232_ (
    .A(_337_),
    .B(_332_),
    .Y(_338_)
);

AOI21X1 _1233_ (
    .A(_184_),
    .B(_186_),
    .C(_189_),
    .Y(_339_)
);

NAND2X1 _1234_ (
    .A(BI[2]),
    .B(AI[6]),
    .Y(_340_)
);

XOR2X1 _1235_ (
    .A(_188_),
    .B(_340_),
    .Y(_341_)
);

NAND2X1 _1236_ (
    .A(_341_),
    .B(_339_),
    .Y(_342_)
);

OAI21X1 _1237_ (
    .A(_183_),
    .B(_185_),
    .C(_182_),
    .Y(_343_)
);

XNOR2X1 _1238_ (
    .A(_188_),
    .B(_340_),
    .Y(_344_)
);

NAND2X1 _1239_ (
    .A(_343_),
    .B(_344_),
    .Y(_345_)
);

NAND3X1 _1240_ (
    .A(_345_),
    .B(_338_),
    .C(_342_),
    .Y(_346_)
);

AND2X2 _1241_ (
    .A(_332_),
    .B(_337_),
    .Y(_347_)
);

NAND2X1 _1242_ (
    .A(_343_),
    .B(_341_),
    .Y(_348_)
);

NAND2X1 _1243_ (
    .A(_344_),
    .B(_339_),
    .Y(_349_)
);

NAND3X1 _1244_ (
    .A(_348_),
    .B(_349_),
    .C(_347_),
    .Y(_350_)
);

NAND3X1 _1245_ (
    .A(_346_),
    .B(_350_),
    .C(_326_),
    .Y(_351_)
);

OAI21X1 _1246_ (
    .A(_211_),
    .B(_191_),
    .C(_210_),
    .Y(_352_)
);

AOI22X1 _1247_ (
    .A(_332_),
    .B(_337_),
    .C(_349_),
    .D(_348_),
    .Y(_353_)
);

AOI21X1 _1248_ (
    .A(_342_),
    .B(_345_),
    .C(_338_),
    .Y(_354_)
);

OAI21X1 _1249_ (
    .A(_353_),
    .B(_354_),
    .C(_352_),
    .Y(_355_)
);

NAND3X1 _1250_ (
    .A(_325_),
    .B(_355_),
    .C(_351_),
    .Y(_356_)
);

AND2X2 _1251_ (
    .A(_321_),
    .B(_324_),
    .Y(_357_)
);

NAND3X1 _1252_ (
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_358_)
);

OAI21X1 _1253_ (
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_359_)
);

NAND3X1 _1254_ (
    .A(_359_),
    .B(_358_),
    .C(_357_),
    .Y(_360_)
);

NAND3X1 _1255_ (
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_361_)
);

AOI21X1 _1256_ (
    .A(_213_),
    .B(_229_),
    .C(_232_),
    .Y(_362_)
);

AOI22X1 _1257_ (
    .A(_321_),
    .B(_324_),
    .C(_358_),
    .D(_359_),
    .Y(_363_)
);

AOI21X1 _1258_ (
    .A(_351_),
    .B(_355_),
    .C(_325_),
    .Y(_364_)
);

OAI21X1 _1259_ (
    .A(_363_),
    .B(_364_),
    .C(_362_),
    .Y(_365_)
);

AOI21X1 _1260_ (
    .A(_361_),
    .B(_365_),
    .C(_313_),
    .Y(_366_)
);

INVX1 _1261_ (
    .A(_313_),
    .Y(_367_)
);

NAND3X1 _1262_ (
    .A(_356_),
    .B(_360_),
    .C(_362_),
    .Y(_368_)
);

OAI21X1 _1263_ (
    .A(_363_),
    .B(_364_),
    .C(_314_),
    .Y(_369_)
);

AOI21X1 _1264_ (
    .A(_368_),
    .B(_369_),
    .C(_367_),
    .Y(_370_)
);

OAI21X1 _1265_ (
    .A(_366_),
    .B(_370_),
    .C(_312_),
    .Y(_371_)
);

OAI21X1 _1266_ (
    .A(_177_),
    .B(_237_),
    .C(_244_),
    .Y(_372_)
);

NAND3X1 _1267_ (
    .A(_367_),
    .B(_369_),
    .C(_368_),
    .Y(_373_)
);

NAND3X1 _1268_ (
    .A(_313_),
    .B(_365_),
    .C(_361_),
    .Y(_374_)
);

NAND3X1 _1269_ (
    .A(_373_),
    .B(_374_),
    .C(_372_),
    .Y(_375_)
);

AND2X2 _1270_ (
    .A(_371_),
    .B(_375_),
    .Y(_376_)
);

XOR2X1 _1271_ (
    .A(_311_),
    .B(_376_),
    .Y(_377_)
);

NOR2X1 _1272_ (
    .A(ABCmd_i[7]),
    .B(HC),
    .Y(_378_)
);

NOR2X1 _1273_ (
    .A(_378_),
    .B(_715_),
    .Y(_379_)
);

OAI21X1 _1274_ (
    .A(_54_),
    .B(_377_),
    .C(_379_),
    .Y(_380_)
);

AOI21X1 _1275_ (
    .A(BI_0_bF$buf1),
    .B(AI[0]),
    .C(_54_),
    .Y(_381_)
);

OAI21X1 _1276_ (
    .A(ACC[0]),
    .B(ABCmd_i[7]),
    .C(_715_),
    .Y(_382_)
);

OAI21X1 _1277_ (
    .A(_381_),
    .B(_382_),
    .C(_380_),
    .Y(_383_)
);

NAND2X1 _1278_ (
    .A(_700_),
    .B(_383_),
    .Y(_384_)
);

OAI21X1 _1279_ (
    .A(_56_),
    .B(_700_),
    .C(_384_),
    .Y(_9_)
);

INVX1 _1280_ (
    .A(_886_[1]),
    .Y(_385_)
);

INVX1 _1281_ (
    .A(AN),
    .Y(_386_)
);

OAI21X1 _1282_ (
    .A(state[1]),
    .B(_712_),
    .C(ABCmd_i[7]),
    .Y(_387_)
);

OAI21X1 _1283_ (
    .A(_386_),
    .B(_715_),
    .C(_387_),
    .Y(_388_)
);

NAND3X1 _1284_ (
    .A(_176_),
    .B(_245_),
    .C(_242_),
    .Y(_389_)
);

INVX1 _1285_ (
    .A(_285_),
    .Y(_390_)
);

NAND2X1 _1286_ (
    .A(_172_),
    .B(_175_),
    .Y(_391_)
);

NAND3X1 _1287_ (
    .A(_122_),
    .B(_262_),
    .C(_391_),
    .Y(_392_)
);

NAND3X1 _1288_ (
    .A(_176_),
    .B(_390_),
    .C(_392_),
    .Y(_393_)
);

AOI21X1 _1289_ (
    .A(_392_),
    .B(_176_),
    .C(_390_),
    .Y(_394_)
);

OAI21X1 _1290_ (
    .A(_307_),
    .B(_394_),
    .C(_393_),
    .Y(_395_)
);

AOI21X1 _1291_ (
    .A(_395_),
    .B(_389_),
    .C(_246_),
    .Y(_396_)
);

NAND2X1 _1292_ (
    .A(_375_),
    .B(_371_),
    .Y(_397_)
);

OAI21X1 _1293_ (
    .A(_397_),
    .B(_396_),
    .C(_375_),
    .Y(_398_)
);

INVX1 _1294_ (
    .A(_361_),
    .Y(_399_)
);

AOI21X1 _1295_ (
    .A(_313_),
    .B(_365_),
    .C(_399_),
    .Y(_400_)
);

OAI21X1 _1296_ (
    .A(_315_),
    .B(_323_),
    .C(_319_),
    .Y(_401_)
);

INVX1 _1297_ (
    .A(_401_),
    .Y(_402_)
);

AOI21X1 _1298_ (
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_403_)
);

OAI21X1 _1299_ (
    .A(_325_),
    .B(_403_),
    .C(_358_),
    .Y(_404_)
);

NAND2X1 _1300_ (
    .A(AI[2]),
    .B(BI[7]),
    .Y(_405_)
);

NOR2X1 _1301_ (
    .A(_149_),
    .B(_167_),
    .Y(_406_)
);

NAND2X1 _1302_ (
    .A(BI_3_bF$buf1),
    .B(AI[4]),
    .Y(_407_)
);

NAND2X1 _1303_ (
    .A(AI_5_bF$buf2),
    .B(BI_4_bF$buf1),
    .Y(_408_)
);

OAI22X1 _1304_ (
    .A(_407_),
    .B(_408_),
    .C(_327_),
    .D(_335_),
    .Y(_409_)
);

XNOR2X1 _1305_ (
    .A(_409_),
    .B(_406_),
    .Y(_410_)
);

XNOR2X1 _1306_ (
    .A(_410_),
    .B(_405_),
    .Y(_411_)
);

NOR2X1 _1307_ (
    .A(_344_),
    .B(_339_),
    .Y(_412_)
);

AOI21X1 _1308_ (
    .A(_347_),
    .B(_349_),
    .C(_412_),
    .Y(_413_)
);

NAND2X1 _1309_ (
    .A(\u_ALU.AI7 ),
    .B(BI[2]),
    .Y(_414_)
);

NAND2X1 _1310_ (
    .A(AI[4]),
    .B(BI[5]),
    .Y(_415_)
);

INVX1 _1311_ (
    .A(_415_),
    .Y(_416_)
);

AND2X2 _1312_ (
    .A(AI_5_bF$buf1),
    .B(BI_4_bF$buf0),
    .Y(_417_)
);

AND2X2 _1313_ (
    .A(AI[6]),
    .B(BI_3_bF$buf0),
    .Y(_418_)
);

NAND2X1 _1314_ (
    .A(_417_),
    .B(_418_),
    .Y(_419_)
);

AOI22X1 _1315_ (
    .A(AI[6]),
    .B(BI_3_bF$buf3),
    .C(AI_5_bF$buf0),
    .D(BI_4_bF$buf3),
    .Y(_420_)
);

INVX1 _1316_ (
    .A(_420_),
    .Y(_421_)
);

AOI21X1 _1317_ (
    .A(_419_),
    .B(_421_),
    .C(_416_),
    .Y(_422_)
);

INVX2 _1318_ (
    .A(AI[6]),
    .Y(_423_)
);

OAI21X1 _1319_ (
    .A(_423_),
    .B(_58_),
    .C(_417_),
    .Y(_424_)
);

OAI21X1 _1320_ (
    .A(_130_),
    .B(_83_),
    .C(_418_),
    .Y(_425_)
);

AOI21X1 _1321_ (
    .A(_424_),
    .B(_425_),
    .C(_415_),
    .Y(_426_)
);

OAI22X1 _1322_ (
    .A(_127_),
    .B(_414_),
    .C(_422_),
    .D(_426_),
    .Y(_427_)
);

NAND3X1 _1323_ (
    .A(_415_),
    .B(_424_),
    .C(_425_),
    .Y(_428_)
);

NAND3X1 _1324_ (
    .A(_416_),
    .B(_421_),
    .C(_419_),
    .Y(_429_)
);

NOR2X1 _1325_ (
    .A(_414_),
    .B(_127_),
    .Y(_430_)
);

NAND3X1 _1326_ (
    .A(_430_),
    .B(_429_),
    .C(_428_),
    .Y(_431_)
);

NAND2X1 _1327_ (
    .A(_431_),
    .B(_427_),
    .Y(_432_)
);

NOR2X1 _1328_ (
    .A(_432_),
    .B(_413_),
    .Y(_433_)
);

NOR2X1 _1329_ (
    .A(_343_),
    .B(_341_),
    .Y(_434_)
);

OAI21X1 _1330_ (
    .A(_338_),
    .B(_434_),
    .C(_348_),
    .Y(_435_)
);

AOI21X1 _1331_ (
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_436_)
);

OAI21X1 _1332_ (
    .A(_436_),
    .B(_433_),
    .C(_411_),
    .Y(_437_)
);

XOR2X1 _1333_ (
    .A(_410_),
    .B(_405_),
    .Y(_438_)
);

NAND3X1 _1334_ (
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_439_)
);

NAND2X1 _1335_ (
    .A(_432_),
    .B(_413_),
    .Y(_440_)
);

NAND3X1 _1336_ (
    .A(_438_),
    .B(_440_),
    .C(_439_),
    .Y(_441_)
);

NAND3X1 _1337_ (
    .A(_441_),
    .B(_437_),
    .C(_404_),
    .Y(_442_)
);

NOR3X1 _1338_ (
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_443_)
);

AOI21X1 _1339_ (
    .A(_357_),
    .B(_359_),
    .C(_443_),
    .Y(_444_)
);

AOI21X1 _1340_ (
    .A(_439_),
    .B(_440_),
    .C(_438_),
    .Y(_445_)
);

NAND3X1 _1341_ (
    .A(_427_),
    .B(_431_),
    .C(_413_),
    .Y(_446_)
);

OAI21X1 _1342_ (
    .A(_412_),
    .B(_354_),
    .C(_432_),
    .Y(_447_)
);

AOI21X1 _1343_ (
    .A(_446_),
    .B(_447_),
    .C(_411_),
    .Y(_448_)
);

OAI21X1 _1344_ (
    .A(_445_),
    .B(_448_),
    .C(_444_),
    .Y(_449_)
);

NAND3X1 _1345_ (
    .A(_402_),
    .B(_442_),
    .C(_449_),
    .Y(_450_)
);

NAND3X1 _1346_ (
    .A(_437_),
    .B(_441_),
    .C(_444_),
    .Y(_451_)
);

OAI21X1 _1347_ (
    .A(_445_),
    .B(_448_),
    .C(_404_),
    .Y(_452_)
);

NAND3X1 _1348_ (
    .A(_401_),
    .B(_452_),
    .C(_451_),
    .Y(_453_)
);

NAND3X1 _1349_ (
    .A(_450_),
    .B(_453_),
    .C(_400_),
    .Y(_454_)
);

AOI21X1 _1350_ (
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_455_)
);

OAI21X1 _1351_ (
    .A(_367_),
    .B(_455_),
    .C(_361_),
    .Y(_456_)
);

NAND3X1 _1352_ (
    .A(_401_),
    .B(_442_),
    .C(_449_),
    .Y(_457_)
);

NAND3X1 _1353_ (
    .A(_402_),
    .B(_452_),
    .C(_451_),
    .Y(_458_)
);

NAND3X1 _1354_ (
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_459_)
);

NAND2X1 _1355_ (
    .A(_459_),
    .B(_454_),
    .Y(_460_)
);

AND2X2 _1356_ (
    .A(_398_),
    .B(_460_),
    .Y(_461_)
);

OAI21X1 _1357_ (
    .A(_460_),
    .B(_398_),
    .C(ABCmd_i[7]),
    .Y(_462_)
);

OAI21X1 _1358_ (
    .A(_462_),
    .B(_461_),
    .C(_388_),
    .Y(_463_)
);

AND2X2 _1359_ (
    .A(_271_),
    .B(_293_),
    .Y(_464_)
);

NAND2X1 _1360_ (
    .A(ACC[1]),
    .B(_54_),
    .Y(_465_)
);

OAI21X1 _1361_ (
    .A(_271_),
    .B(_293_),
    .C(ABCmd_i[7]),
    .Y(_466_)
);

OAI21X1 _1362_ (
    .A(_466_),
    .B(_464_),
    .C(_465_),
    .Y(_467_)
);

AOI21X1 _1363_ (
    .A(_467_),
    .B(_703_),
    .C(_712_),
    .Y(_468_)
);

AOI22X1 _1364_ (
    .A(_385_),
    .B(_712_),
    .C(_463_),
    .D(_468_),
    .Y(_10_)
);

OAI21X1 _1365_ (
    .A(state[0]),
    .B(_699_),
    .C(_886_[2]),
    .Y(_469_)
);

AOI21X1 _1366_ (
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_470_)
);

AOI22X1 _1367_ (
    .A(_361_),
    .B(_374_),
    .C(_453_),
    .D(_450_),
    .Y(_471_)
);

NOR2X1 _1368_ (
    .A(_471_),
    .B(_470_),
    .Y(_472_)
);

NAND3X1 _1369_ (
    .A(_376_),
    .B(_472_),
    .C(_311_),
    .Y(_473_)
);

AOI21X1 _1370_ (
    .A(_375_),
    .B(_459_),
    .C(_470_),
    .Y(_474_)
);

INVX1 _1371_ (
    .A(_474_),
    .Y(_475_)
);

NAND2X1 _1372_ (
    .A(_406_),
    .B(_409_),
    .Y(_476_)
);

OAI21X1 _1373_ (
    .A(_405_),
    .B(_410_),
    .C(_476_),
    .Y(_477_)
);

INVX1 _1374_ (
    .A(_477_),
    .Y(_478_)
);

AOI21X1 _1375_ (
    .A(_438_),
    .B(_440_),
    .C(_433_),
    .Y(_479_)
);

NAND2X1 _1376_ (
    .A(AI[3]),
    .B(BI[7]),
    .Y(_480_)
);

INVX1 _1377_ (
    .A(_480_),
    .Y(_481_)
);

NOR2X1 _1378_ (
    .A(_74_),
    .B(_167_),
    .Y(_482_)
);

OAI21X1 _1379_ (
    .A(_415_),
    .B(_420_),
    .C(_419_),
    .Y(_483_)
);

NAND2X1 _1380_ (
    .A(_482_),
    .B(_483_),
    .Y(_484_)
);

OR2X2 _1381_ (
    .A(_483_),
    .B(_482_),
    .Y(_485_)
);

NAND3X1 _1382_ (
    .A(_481_),
    .B(_484_),
    .C(_485_),
    .Y(_486_)
);

AND2X2 _1383_ (
    .A(_483_),
    .B(_482_),
    .Y(_487_)
);

NOR2X1 _1384_ (
    .A(_482_),
    .B(_483_),
    .Y(_488_)
);

OAI21X1 _1385_ (
    .A(_488_),
    .B(_487_),
    .C(_480_),
    .Y(_489_)
);

NAND2X1 _1386_ (
    .A(_489_),
    .B(_486_),
    .Y(_490_)
);

OR2X2 _1387_ (
    .A(_188_),
    .B(_340_),
    .Y(_491_)
);

NAND2X1 _1388_ (
    .A(AI_5_bF$buf3),
    .B(BI[5]),
    .Y(_492_)
);

NAND2X1 _1389_ (
    .A(AI[6]),
    .B(BI_3_bF$buf2),
    .Y(_493_)
);

NAND2X1 _1390_ (
    .A(\u_ALU.AI7 ),
    .B(BI_4_bF$buf2),
    .Y(_494_)
);

AOI22X1 _1391_ (
    .A(\u_ALU.AI7 ),
    .B(BI_3_bF$buf1),
    .C(AI[6]),
    .D(BI_4_bF$buf1),
    .Y(_495_)
);

INVX1 _1392_ (
    .A(_495_),
    .Y(_496_)
);

OAI21X1 _1393_ (
    .A(_493_),
    .B(_494_),
    .C(_496_),
    .Y(_497_)
);

XNOR2X1 _1394_ (
    .A(_497_),
    .B(_492_),
    .Y(_498_)
);

AOI21X1 _1395_ (
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_499_)
);

NAND3X1 _1396_ (
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_500_)
);

INVX1 _1397_ (
    .A(_500_),
    .Y(_501_)
);

OAI21X1 _1398_ (
    .A(_499_),
    .B(_501_),
    .C(_490_),
    .Y(_502_)
);

AND2X2 _1399_ (
    .A(_486_),
    .B(_489_),
    .Y(_503_)
);

NAND2X1 _1400_ (
    .A(_491_),
    .B(_431_),
    .Y(_504_)
);

INVX1 _1401_ (
    .A(_498_),
    .Y(_505_)
);

NAND2X1 _1402_ (
    .A(_504_),
    .B(_505_),
    .Y(_506_)
);

NAND3X1 _1403_ (
    .A(_506_),
    .B(_500_),
    .C(_503_),
    .Y(_507_)
);

NAND3X1 _1404_ (
    .A(_502_),
    .B(_507_),
    .C(_479_),
    .Y(_508_)
);

OAI21X1 _1405_ (
    .A(_411_),
    .B(_436_),
    .C(_439_),
    .Y(_509_)
);

AOI22X1 _1406_ (
    .A(_486_),
    .B(_489_),
    .C(_506_),
    .D(_500_),
    .Y(_510_)
);

OR2X2 _1407_ (
    .A(_504_),
    .B(_498_),
    .Y(_511_)
);

NAND2X1 _1408_ (
    .A(_498_),
    .B(_504_),
    .Y(_512_)
);

AOI21X1 _1409_ (
    .A(_511_),
    .B(_512_),
    .C(_490_),
    .Y(_513_)
);

OAI21X1 _1410_ (
    .A(_510_),
    .B(_513_),
    .C(_509_),
    .Y(_514_)
);

NAND3X1 _1411_ (
    .A(_478_),
    .B(_514_),
    .C(_508_),
    .Y(_515_)
);

NAND3X1 _1412_ (
    .A(_507_),
    .B(_502_),
    .C(_509_),
    .Y(_516_)
);

OAI21X1 _1413_ (
    .A(_510_),
    .B(_513_),
    .C(_479_),
    .Y(_517_)
);

NAND3X1 _1414_ (
    .A(_477_),
    .B(_516_),
    .C(_517_),
    .Y(_518_)
);

NAND2X1 _1415_ (
    .A(_518_),
    .B(_515_),
    .Y(_519_)
);

NAND3X1 _1416_ (
    .A(_442_),
    .B(_457_),
    .C(_519_),
    .Y(_520_)
);

AOI21X1 _1417_ (
    .A(_437_),
    .B(_441_),
    .C(_404_),
    .Y(_521_)
);

OAI21X1 _1418_ (
    .A(_402_),
    .B(_521_),
    .C(_442_),
    .Y(_522_)
);

NAND3X1 _1419_ (
    .A(_515_),
    .B(_518_),
    .C(_522_),
    .Y(_523_)
);

NAND2X1 _1420_ (
    .A(_523_),
    .B(_520_),
    .Y(_524_)
);

AOI21X1 _1421_ (
    .A(_473_),
    .B(_475_),
    .C(_524_),
    .Y(_525_)
);

NAND2X1 _1422_ (
    .A(_376_),
    .B(_472_),
    .Y(_526_)
);

OAI21X1 _1423_ (
    .A(_396_),
    .B(_526_),
    .C(_475_),
    .Y(_527_)
);

INVX1 _1424_ (
    .A(_524_),
    .Y(_528_)
);

NOR2X1 _1425_ (
    .A(_528_),
    .B(_527_),
    .Y(_529_)
);

OAI21X1 _1426_ (
    .A(_525_),
    .B(_529_),
    .C(ABCmd_i[7]),
    .Y(_530_)
);

NOR2X1 _1427_ (
    .A(ABCmd_i[7]),
    .B(AZ),
    .Y(_531_)
);

NOR2X1 _1428_ (
    .A(_531_),
    .B(_715_),
    .Y(_532_)
);

AOI21X1 _1429_ (
    .A(_292_),
    .B(_296_),
    .C(_294_),
    .Y(_533_)
);

OAI21X1 _1430_ (
    .A(_533_),
    .B(_298_),
    .C(ABCmd_i[7]),
    .Y(_534_)
);

NOR2X1 _1431_ (
    .A(ABCmd_i[7]),
    .B(ACC[2]),
    .Y(_535_)
);

NOR2X1 _1432_ (
    .A(_535_),
    .B(_25_),
    .Y(_536_)
);

AOI22X1 _1433_ (
    .A(_534_),
    .B(_536_),
    .C(_530_),
    .D(_532_),
    .Y(_537_)
);

OAI21X1 _1434_ (
    .A(_712_),
    .B(_537_),
    .C(_469_),
    .Y(_11_)
);

INVX1 _1435_ (
    .A(_886_[3]),
    .Y(_538_)
);

INVX1 _1436_ (
    .A(AV),
    .Y(_539_)
);

OAI21X1 _1437_ (
    .A(_539_),
    .B(_715_),
    .C(_387_),
    .Y(_540_)
);

INVX1 _1438_ (
    .A(_523_),
    .Y(_541_)
);

OAI21X1 _1439_ (
    .A(_480_),
    .B(_488_),
    .C(_484_),
    .Y(_542_)
);

INVX1 _1440_ (
    .A(_542_),
    .Y(_543_)
);

AOI21X1 _1441_ (
    .A(_503_),
    .B(_500_),
    .C(_499_),
    .Y(_544_)
);

NAND2X1 _1442_ (
    .A(AI[4]),
    .B(BI[7]),
    .Y(_545_)
);

INVX1 _1443_ (
    .A(_545_),
    .Y(_546_)
);

NOR2X1 _1444_ (
    .A(_130_),
    .B(_167_),
    .Y(_547_)
);

OAI22X1 _1445_ (
    .A(_493_),
    .B(_494_),
    .C(_492_),
    .D(_495_),
    .Y(_548_)
);

NAND2X1 _1446_ (
    .A(_547_),
    .B(_548_),
    .Y(_549_)
);

NOR2X1 _1447_ (
    .A(_547_),
    .B(_548_),
    .Y(_550_)
);

INVX1 _1448_ (
    .A(_550_),
    .Y(_551_)
);

NAND3X1 _1449_ (
    .A(_546_),
    .B(_549_),
    .C(_551_),
    .Y(_552_)
);

INVX1 _1450_ (
    .A(_549_),
    .Y(_553_)
);

OAI21X1 _1451_ (
    .A(_550_),
    .B(_553_),
    .C(_545_),
    .Y(_554_)
);

NAND2X1 _1452_ (
    .A(AI[6]),
    .B(BI_4_bF$buf0),
    .Y(_555_)
);

NAND2X1 _1453_ (
    .A(\u_ALU.AI7 ),
    .B(BI[5]),
    .Y(_556_)
);

OR2X2 _1454_ (
    .A(_555_),
    .B(_556_),
    .Y(_557_)
);

INVX1 _1455_ (
    .A(BI[5]),
    .Y(_558_)
);

OAI21X1 _1456_ (
    .A(_423_),
    .B(_558_),
    .C(_494_),
    .Y(_559_)
);

AND2X2 _1457_ (
    .A(_557_),
    .B(_559_),
    .Y(_560_)
);

AOI21X1 _1458_ (
    .A(_552_),
    .B(_554_),
    .C(_560_),
    .Y(_561_)
);

INVX1 _1459_ (
    .A(_561_),
    .Y(_562_)
);

NAND3X1 _1460_ (
    .A(_560_),
    .B(_554_),
    .C(_552_),
    .Y(_563_)
);

NAND3X1 _1461_ (
    .A(_562_),
    .B(_563_),
    .C(_544_),
    .Y(_564_)
);

OAI21X1 _1462_ (
    .A(_490_),
    .B(_501_),
    .C(_506_),
    .Y(_565_)
);

INVX1 _1463_ (
    .A(_563_),
    .Y(_566_)
);

OAI21X1 _1464_ (
    .A(_561_),
    .B(_566_),
    .C(_565_),
    .Y(_567_)
);

NAND3X1 _1465_ (
    .A(_543_),
    .B(_567_),
    .C(_564_),
    .Y(_568_)
);

NAND3X1 _1466_ (
    .A(_563_),
    .B(_562_),
    .C(_565_),
    .Y(_569_)
);

OAI21X1 _1467_ (
    .A(_561_),
    .B(_566_),
    .C(_544_),
    .Y(_570_)
);

NAND3X1 _1468_ (
    .A(_542_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

NAND2X1 _1469_ (
    .A(_571_),
    .B(_568_),
    .Y(_572_)
);

NAND3X1 _1470_ (
    .A(_516_),
    .B(_518_),
    .C(_572_),
    .Y(_573_)
);

AOI21X1 _1471_ (
    .A(_502_),
    .B(_507_),
    .C(_509_),
    .Y(_574_)
);

OAI21X1 _1472_ (
    .A(_478_),
    .B(_574_),
    .C(_516_),
    .Y(_575_)
);

NAND3X1 _1473_ (
    .A(_568_),
    .B(_571_),
    .C(_575_),
    .Y(_576_)
);

NAND2X1 _1474_ (
    .A(_576_),
    .B(_573_),
    .Y(_577_)
);

NOR3X1 _1475_ (
    .A(_541_),
    .B(_577_),
    .C(_525_),
    .Y(_578_)
);

AOI21X1 _1476_ (
    .A(_527_),
    .B(_528_),
    .C(_541_),
    .Y(_579_)
);

INVX1 _1477_ (
    .A(_577_),
    .Y(_580_)
);

OAI21X1 _1478_ (
    .A(_580_),
    .B(_579_),
    .C(ABCmd_i[7]),
    .Y(_581_)
);

OAI21X1 _1479_ (
    .A(_578_),
    .B(_581_),
    .C(_540_),
    .Y(_582_)
);

NAND2X1 _1480_ (
    .A(_289_),
    .B(_300_),
    .Y(_583_)
);

NAND2X1 _1481_ (
    .A(_297_),
    .B(_583_),
    .Y(_584_)
);

NAND2X1 _1482_ (
    .A(_301_),
    .B(_584_),
    .Y(_585_)
);

NAND2X1 _1483_ (
    .A(ACC[3]),
    .B(_54_),
    .Y(_586_)
);

OAI21X1 _1484_ (
    .A(_54_),
    .B(_585_),
    .C(_586_),
    .Y(_587_)
);

AOI21X1 _1485_ (
    .A(_587_),
    .B(_703_),
    .C(_712_),
    .Y(_588_)
);

AOI22X1 _1486_ (
    .A(_538_),
    .B(_712_),
    .C(_582_),
    .D(_588_),
    .Y(_12_)
);

INVX1 _1487_ (
    .A(_886_[4]),
    .Y(_589_)
);

OAI21X1 _1488_ (
    .A(_545_),
    .B(_550_),
    .C(_549_),
    .Y(_590_)
);

INVX1 _1489_ (
    .A(_590_),
    .Y(_591_)
);

INVX1 _1490_ (
    .A(\u_ALU.AI7 ),
    .Y(_592_)
);

NAND2X1 _1491_ (
    .A(AI_5_bF$buf2),
    .B(BI[7]),
    .Y(_593_)
);

OAI21X1 _1492_ (
    .A(_423_),
    .B(_167_),
    .C(_557_),
    .Y(_594_)
);

OAI21X1 _1493_ (
    .A(_167_),
    .B(_557_),
    .C(_594_),
    .Y(_595_)
);

OR2X2 _1494_ (
    .A(_595_),
    .B(_593_),
    .Y(_596_)
);

INVX1 _1495_ (
    .A(BI[7]),
    .Y(_597_)
);

OAI21X1 _1496_ (
    .A(_130_),
    .B(_597_),
    .C(_595_),
    .Y(_598_)
);

NAND2X1 _1497_ (
    .A(_598_),
    .B(_596_),
    .Y(_599_)
);

OAI21X1 _1498_ (
    .A(_592_),
    .B(_558_),
    .C(_599_),
    .Y(_600_)
);

INVX1 _1499_ (
    .A(_556_),
    .Y(_601_)
);

NAND3X1 _1500_ (
    .A(_601_),
    .B(_598_),
    .C(_596_),
    .Y(_602_)
);

NAND2X1 _1501_ (
    .A(_602_),
    .B(_600_),
    .Y(_603_)
);

NOR2X1 _1502_ (
    .A(_563_),
    .B(_603_),
    .Y(_604_)
);

NAND2X1 _1503_ (
    .A(_563_),
    .B(_603_),
    .Y(_605_)
);

INVX1 _1504_ (
    .A(_605_),
    .Y(_606_)
);

OAI21X1 _1505_ (
    .A(_604_),
    .B(_606_),
    .C(_591_),
    .Y(_607_)
);

OR2X2 _1506_ (
    .A(_603_),
    .B(_563_),
    .Y(_608_)
);

NAND3X1 _1507_ (
    .A(_590_),
    .B(_605_),
    .C(_608_),
    .Y(_609_)
);

NAND2X1 _1508_ (
    .A(_609_),
    .B(_607_),
    .Y(_610_)
);

NAND3X1 _1509_ (
    .A(_569_),
    .B(_571_),
    .C(_610_),
    .Y(_611_)
);

NAND2X1 _1510_ (
    .A(_569_),
    .B(_571_),
    .Y(_612_)
);

NAND3X1 _1511_ (
    .A(_612_),
    .B(_609_),
    .C(_607_),
    .Y(_613_)
);

NAND2X1 _1512_ (
    .A(_613_),
    .B(_611_),
    .Y(_614_)
);

NOR2X1 _1513_ (
    .A(_397_),
    .B(_460_),
    .Y(_615_)
);

NOR2X1 _1514_ (
    .A(_577_),
    .B(_524_),
    .Y(_616_)
);

NAND3X1 _1515_ (
    .A(_311_),
    .B(_616_),
    .C(_615_),
    .Y(_617_)
);

NAND2X1 _1516_ (
    .A(_576_),
    .B(_523_),
    .Y(_618_)
);

AOI22X1 _1517_ (
    .A(_573_),
    .B(_618_),
    .C(_616_),
    .D(_474_),
    .Y(_619_)
);

AOI21X1 _1518_ (
    .A(_619_),
    .B(_617_),
    .C(_614_),
    .Y(_620_)
);

NAND2X1 _1519_ (
    .A(_573_),
    .B(_618_),
    .Y(_621_)
);

OAI21X1 _1520_ (
    .A(_524_),
    .B(_577_),
    .C(_621_),
    .Y(_622_)
);

AOI21X1 _1521_ (
    .A(_573_),
    .B(_618_),
    .C(_474_),
    .Y(_623_)
);

OAI21X1 _1522_ (
    .A(_396_),
    .B(_526_),
    .C(_623_),
    .Y(_624_)
);

AOI22X1 _1523_ (
    .A(_611_),
    .B(_613_),
    .C(_624_),
    .D(_622_),
    .Y(_625_)
);

OAI21X1 _1524_ (
    .A(_625_),
    .B(_620_),
    .C(ABCmd_i[7]),
    .Y(_626_)
);

OR2X2 _1525_ (
    .A(ABCmd_i[7]),
    .B(CO),
    .Y(_627_)
);

NAND3X1 _1526_ (
    .A(_25_),
    .B(_627_),
    .C(_626_),
    .Y(_628_)
);

INVX1 _1527_ (
    .A(_303_),
    .Y(_629_)
);

OAI21X1 _1528_ (
    .A(_302_),
    .B(_282_),
    .C(_301_),
    .Y(_630_)
);

NAND2X1 _1529_ (
    .A(_630_),
    .B(_629_),
    .Y(_631_)
);

NAND2X1 _1530_ (
    .A(ACC[4]),
    .B(_54_),
    .Y(_632_)
);

OAI21X1 _1531_ (
    .A(_54_),
    .B(_631_),
    .C(_632_),
    .Y(_633_)
);

AOI21X1 _1532_ (
    .A(_633_),
    .B(_703_),
    .C(_712_),
    .Y(_634_)
);

AOI22X1 _1533_ (
    .A(_589_),
    .B(_712_),
    .C(_628_),
    .D(_634_),
    .Y(_13_)
);

INVX1 _1534_ (
    .A(_886_[5]),
    .Y(_635_)
);

INVX1 _1535_ (
    .A(_387_),
    .Y(_636_)
);

NAND2X1 _1536_ (
    .A(_622_),
    .B(_624_),
    .Y(_637_)
);

INVX1 _1537_ (
    .A(_613_),
    .Y(_638_)
);

AOI21X1 _1538_ (
    .A(_590_),
    .B(_605_),
    .C(_604_),
    .Y(_639_)
);

OAI21X1 _1539_ (
    .A(_167_),
    .B(_557_),
    .C(_596_),
    .Y(_640_)
);

NOR2X1 _1540_ (
    .A(_592_),
    .B(_597_),
    .Y(_641_)
);

NAND3X1 _1541_ (
    .A(AI[6]),
    .B(BI[6]),
    .C(_641_),
    .Y(_642_)
);

OAI22X1 _1542_ (
    .A(_592_),
    .B(_167_),
    .C(_423_),
    .D(_597_),
    .Y(_643_)
);

NAND2X1 _1543_ (
    .A(_643_),
    .B(_642_),
    .Y(_644_)
);

XNOR2X1 _1544_ (
    .A(_602_),
    .B(_644_),
    .Y(_645_)
);

XOR2X1 _1545_ (
    .A(_645_),
    .B(_640_),
    .Y(_646_)
);

XOR2X1 _1546_ (
    .A(_639_),
    .B(_646_),
    .Y(_647_)
);

NOR2X1 _1547_ (
    .A(_638_),
    .B(_647_),
    .Y(_648_)
);

OAI21X1 _1548_ (
    .A(_614_),
    .B(_637_),
    .C(_648_),
    .Y(_649_)
);

OAI21X1 _1549_ (
    .A(_638_),
    .B(_620_),
    .C(_647_),
    .Y(_650_)
);

NAND3X1 _1550_ (
    .A(_636_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

AOI21X1 _1551_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_652_)
);

OAI21X1 _1552_ (
    .A(_652_),
    .B(_308_),
    .C(ABCmd_i[7]),
    .Y(_653_)
);

INVX1 _1553_ (
    .A(ACC[5]),
    .Y(_654_)
);

AOI21X1 _1554_ (
    .A(_54_),
    .B(_654_),
    .C(state[1]),
    .Y(_655_)
);

AOI21X1 _1555_ (
    .A(_653_),
    .B(_655_),
    .C(_712_),
    .Y(_656_)
);

AOI22X1 _1556_ (
    .A(_635_),
    .B(_712_),
    .C(_651_),
    .D(_656_),
    .Y(_14_)
);

INVX1 _1557_ (
    .A(_886_[6]),
    .Y(_657_)
);

NAND3X1 _1558_ (
    .A(_613_),
    .B(_647_),
    .C(_611_),
    .Y(_658_)
);

INVX1 _1559_ (
    .A(_658_),
    .Y(_659_)
);

NAND3X1 _1560_ (
    .A(_622_),
    .B(_659_),
    .C(_624_),
    .Y(_660_)
);

NAND2X1 _1561_ (
    .A(_638_),
    .B(_647_),
    .Y(_661_)
);

OAI21X1 _1562_ (
    .A(_639_),
    .B(_646_),
    .C(_661_),
    .Y(_662_)
);

INVX1 _1563_ (
    .A(_662_),
    .Y(_663_)
);

INVX1 _1564_ (
    .A(_645_),
    .Y(_664_)
);

NAND2X1 _1565_ (
    .A(_640_),
    .B(_664_),
    .Y(_665_)
);

OAI21X1 _1566_ (
    .A(_602_),
    .B(_644_),
    .C(_665_),
    .Y(_666_)
);

OAI21X1 _1567_ (
    .A(_423_),
    .B(_167_),
    .C(_641_),
    .Y(_667_)
);

XOR2X1 _1568_ (
    .A(_666_),
    .B(_667_),
    .Y(_668_)
);

NAND3X1 _1569_ (
    .A(_668_),
    .B(_663_),
    .C(_660_),
    .Y(_669_)
);

AOI21X1 _1570_ (
    .A(_619_),
    .B(_617_),
    .C(_658_),
    .Y(_670_)
);

INVX1 _1571_ (
    .A(_668_),
    .Y(_671_)
);

OAI21X1 _1572_ (
    .A(_662_),
    .B(_670_),
    .C(_671_),
    .Y(_672_)
);

NAND3X1 _1573_ (
    .A(_636_),
    .B(_669_),
    .C(_672_),
    .Y(_673_)
);

NAND2X1 _1574_ (
    .A(_309_),
    .B(_393_),
    .Y(_674_)
);

NOR2X1 _1575_ (
    .A(_307_),
    .B(_674_),
    .Y(_675_)
);

AOI21X1 _1576_ (
    .A(_393_),
    .B(_309_),
    .C(_308_),
    .Y(_676_)
);

OAI21X1 _1577_ (
    .A(_676_),
    .B(_675_),
    .C(ABCmd_i[7]),
    .Y(_677_)
);

NOR2X1 _1578_ (
    .A(ABCmd_i[7]),
    .B(ACC[6]),
    .Y(_678_)
);

NOR2X1 _1579_ (
    .A(_678_),
    .B(_25_),
    .Y(_679_)
);

AOI21X1 _1580_ (
    .A(_677_),
    .B(_679_),
    .C(_712_),
    .Y(_680_)
);

AOI22X1 _1581_ (
    .A(_657_),
    .B(_712_),
    .C(_673_),
    .D(_680_),
    .Y(_15_)
);

INVX1 _1582_ (
    .A(_886_[7]),
    .Y(_681_)
);

AOI21X1 _1583_ (
    .A(_660_),
    .B(_663_),
    .C(_668_),
    .Y(_682_)
);

NAND3X1 _1584_ (
    .A(_641_),
    .B(_642_),
    .C(_666_),
    .Y(_683_)
);

NAND2X1 _1585_ (
    .A(_642_),
    .B(_683_),
    .Y(_684_)
);

OAI21X1 _1586_ (
    .A(_684_),
    .B(_682_),
    .C(_636_),
    .Y(_685_)
);

NAND2X1 _1587_ (
    .A(_389_),
    .B(_247_),
    .Y(_686_)
);

XNOR2X1 _1588_ (
    .A(_686_),
    .B(_310_),
    .Y(_687_)
);

NAND2X1 _1589_ (
    .A(AN),
    .B(_54_),
    .Y(_688_)
);

OAI21X1 _1590_ (
    .A(_54_),
    .B(_687_),
    .C(_688_),
    .Y(_689_)
);

AOI21X1 _1591_ (
    .A(_689_),
    .B(_703_),
    .C(_712_),
    .Y(_690_)
);

AOI22X1 _1592_ (
    .A(_681_),
    .B(_712_),
    .C(_685_),
    .D(_690_),
    .Y(_16_)
);

NAND2X1 _1593_ (
    .A(AI[0]),
    .B(_705__bF$buf3),
    .Y(_691_)
);

OAI21X1 _1594_ (
    .A(_40_),
    .B(_705__bF$buf2),
    .C(_691_),
    .Y(_17_)
);

NAND2X1 _1595_ (
    .A(AI[1]),
    .B(_705__bF$buf1),
    .Y(_692_)
);

OAI21X1 _1596_ (
    .A(_42_),
    .B(_705__bF$buf0),
    .C(_692_),
    .Y(_18_)
);

NAND2X1 _1597_ (
    .A(AI[2]),
    .B(_705__bF$buf3),
    .Y(_693_)
);

OAI21X1 _1598_ (
    .A(_44_),
    .B(_705__bF$buf2),
    .C(_693_),
    .Y(_19_)
);

NAND2X1 _1599_ (
    .A(AI[3]),
    .B(_705__bF$buf1),
    .Y(_694_)
);

OAI21X1 _1600_ (
    .A(_46_),
    .B(_705__bF$buf0),
    .C(_694_),
    .Y(_20_)
);

NAND2X1 _1601_ (
    .A(AI[4]),
    .B(_705__bF$buf3),
    .Y(_695_)
);

OAI21X1 _1602_ (
    .A(_48_),
    .B(_705__bF$buf2),
    .C(_695_),
    .Y(_21_)
);

NAND2X1 _1603_ (
    .A(AI_5_bF$buf1),
    .B(_705__bF$buf1),
    .Y(_696_)
);

OAI21X1 _1604_ (
    .A(_50_),
    .B(_705__bF$buf0),
    .C(_696_),
    .Y(_22_)
);

NAND2X1 _1605_ (
    .A(AI[6]),
    .B(_705__bF$buf3),
    .Y(_697_)
);

OAI21X1 _1606_ (
    .A(_52_),
    .B(_705__bF$buf2),
    .C(_697_),
    .Y(_23_)
);

NAND2X1 _1607_ (
    .A(\u_ALU.AI7 ),
    .B(_705__bF$buf1),
    .Y(_698_)
);

OAI21X1 _1608_ (
    .A(_54_),
    .B(_705__bF$buf0),
    .C(_698_),
    .Y(_24_)
);

DFFSR _1609_ (
    .CLK(clk_bF$buf4),
    .D(_1_),
    .Q(BI[0]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1610_ (
    .CLK(clk_bF$buf3),
    .D(_2_),
    .Q(BI[1]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1611_ (
    .CLK(clk_bF$buf2),
    .D(_3_),
    .Q(BI[2]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1612_ (
    .CLK(clk_bF$buf1),
    .D(_4_),
    .Q(BI[3]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1613_ (
    .CLK(clk_bF$buf0),
    .D(_5_),
    .Q(BI[4]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1614_ (
    .CLK(clk_bF$buf4),
    .D(_6_),
    .Q(BI[5]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1615_ (
    .CLK(clk_bF$buf3),
    .D(_7_),
    .Q(BI[6]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1616_ (
    .CLK(clk_bF$buf2),
    .D(_8_),
    .Q(BI[7]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1617_ (
    .CLK(clk_bF$buf1),
    .D(_9_),
    .Q(_886_[0]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1618_ (
    .CLK(clk_bF$buf0),
    .D(_10_),
    .Q(_886_[1]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1619_ (
    .CLK(clk_bF$buf4),
    .D(_11_),
    .Q(_886_[2]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1620_ (
    .CLK(clk_bF$buf3),
    .D(_12_),
    .Q(_886_[3]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1621_ (
    .CLK(clk_bF$buf2),
    .D(_13_),
    .Q(_886_[4]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1622_ (
    .CLK(clk_bF$buf1),
    .D(_14_),
    .Q(_886_[5]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1623_ (
    .CLK(clk_bF$buf0),
    .D(_15_),
    .Q(_886_[6]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1624_ (
    .CLK(clk_bF$buf4),
    .D(_16_),
    .Q(_886_[7]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1625_ (
    .CLK(clk_bF$buf3),
    .D(_17_),
    .Q(AI[0]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1626_ (
    .CLK(clk_bF$buf2),
    .D(_18_),
    .Q(AI[1]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1627_ (
    .CLK(clk_bF$buf1),
    .D(_19_),
    .Q(AI[2]),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1628_ (
    .CLK(clk_bF$buf0),
    .D(_20_),
    .Q(AI[3]),
    .R(_0__bF$buf0),
    .S(vdd)
);

DFFSR _1629_ (
    .CLK(clk_bF$buf4),
    .D(_21_),
    .Q(AI[4]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1630_ (
    .CLK(clk_bF$buf3),
    .D(_22_),
    .Q(AI[5]),
    .R(_0__bF$buf3),
    .S(vdd)
);

DFFSR _1631_ (
    .CLK(clk_bF$buf2),
    .D(_23_),
    .Q(AI[6]),
    .R(_0__bF$buf2),
    .S(vdd)
);

DFFSR _1632_ (
    .CLK(clk_bF$buf1),
    .D(_24_),
    .Q(\u_ALU.AI7 ),
    .R(_0__bF$buf1),
    .S(vdd)
);

DFFSR _1633_ (
    .CLK(clk_bF$buf0),
    .D(_888_[0]),
    .Q(state[0]),
    .R(vdd),
    .S(_0__bF$buf0)
);

DFFSR _1634_ (
    .CLK(clk_bF$buf4),
    .D(_888_[1]),
    .Q(state[1]),
    .R(_0__bF$buf4),
    .S(vdd)
);

DFFSR _1635_ (
    .CLK(clk_bF$buf3),
    .D(_888_[2]),
    .Q(state[2]),
    .R(_0__bF$buf3),
    .S(vdd)
);

INVX1 _1636_ (
    .A(ABCmd_i_2_bF$buf3),
    .Y(_824_)
);

INVX4 _1637_ (
    .A(ABCmd_i[3]),
    .Y(_825_)
);

OAI21X1 _1638_ (
    .A(_824_),
    .B(_825_),
    .C(ABCmd_i[4]),
    .Y(_826_)
);

NOR2X1 _1639_ (
    .A(ABCmd_i[5]),
    .B(_826_),
    .Y(_827_)
);

INVX1 _1640_ (
    .A(_827_),
    .Y(_828_)
);

INVX2 _1641_ (
    .A(ABCmd_i[1]),
    .Y(_829_)
);

NAND2X1 _1642_ (
    .A(ABCmd_i[0]),
    .B(_829_),
    .Y(_830_)
);

INVX2 _1643_ (
    .A(ABCmd_i[0]),
    .Y(_831_)
);

NAND2X1 _1644_ (
    .A(BI_0_bF$buf0),
    .B(_831_),
    .Y(_832_)
);

NAND2X1 _1645_ (
    .A(AI[0]),
    .B(ABCmd_i[1]),
    .Y(_833_)
);

AOI22X1 _1646_ (
    .A(BI_0_bF$buf3),
    .B(_833_),
    .C(_830_),
    .D(_832_),
    .Y(_834_)
);

INVX2 _1647_ (
    .A(ABCmd_i[5]),
    .Y(_835_)
);

INVX1 _1648_ (
    .A(BI_0_bF$buf2),
    .Y(_836_)
);

INVX1 _1649_ (
    .A(AI[0]),
    .Y(_837_)
);

OAI21X1 _1650_ (
    .A(ABCmd_i[0]),
    .B(_836_),
    .C(_837_),
    .Y(_838_)
);

NAND2X1 _1651_ (
    .A(_835_),
    .B(_838_),
    .Y(_839_)
);

NAND2X1 _1652_ (
    .A(AI[1]),
    .B(ABCmd_i[5]),
    .Y(_840_)
);

OAI21X1 _1653_ (
    .A(_834_),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

OAI21X1 _1654_ (
    .A(BI_0_bF$buf1),
    .B(ABCmd_i_2_bF$buf2),
    .C(_825_),
    .Y(_842_)
);

AOI21X1 _1655_ (
    .A(BI_0_bF$buf0),
    .B(ABCmd_i_2_bF$buf1),
    .C(_842_),
    .Y(_843_)
);

NOR2X1 _1656_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(_825_),
    .Y(_844_)
);

OAI21X1 _1657_ (
    .A(_844_),
    .B(_843_),
    .C(_841_),
    .Y(_845_)
);

OAI21X1 _1658_ (
    .A(_841_),
    .B(_843_),
    .C(_845_),
    .Y(_846_)
);

XOR2X1 _1659_ (
    .A(_846_),
    .B(_828_),
    .Y(ACC[0])
);

NOR2X1 _1660_ (
    .A(_843_),
    .B(_841_),
    .Y(_847_)
);

OAI21X1 _1661_ (
    .A(_828_),
    .B(_847_),
    .C(_845_),
    .Y(_848_)
);

NAND2X1 _1662_ (
    .A(ABCmd_i[5]),
    .B(AI[2]),
    .Y(_849_)
);

NAND3X1 _1663_ (
    .A(AI[1]),
    .B(BI_1_bF$buf0),
    .C(_831_),
    .Y(_850_)
);

AOI22X1 _1664_ (
    .A(_829_),
    .B(BI_1_bF$buf3),
    .C(_850_),
    .D(_830_),
    .Y(_851_)
);

INVX1 _1665_ (
    .A(BI_1_bF$buf2),
    .Y(_852_)
);

NOR2X1 _1666_ (
    .A(ABCmd_i[0]),
    .B(_852_),
    .Y(_853_)
);

OAI21X1 _1667_ (
    .A(AI[1]),
    .B(_853_),
    .C(_835_),
    .Y(_854_)
);

OAI21X1 _1668_ (
    .A(_851_),
    .B(_854_),
    .C(_849_),
    .Y(_855_)
);

OAI21X1 _1669_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_1_bF$buf1),
    .C(_825_),
    .Y(_856_)
);

AOI21X1 _1670_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_1_bF$buf0),
    .C(_856_),
    .Y(_857_)
);

INVX1 _1671_ (
    .A(_857_),
    .Y(_858_)
);

OAI21X1 _1672_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .C(_858_),
    .Y(_859_)
);

MUX2X1 _1673_ (
    .A(_859_),
    .B(_858_),
    .S(_855_),
    .Y(_860_)
);

NAND2X1 _1674_ (
    .A(_860_),
    .B(_848_),
    .Y(_861_)
);

INVX1 _1675_ (
    .A(_842_),
    .Y(_862_)
);

OAI21X1 _1676_ (
    .A(_836_),
    .B(_824_),
    .C(_862_),
    .Y(_863_)
);

OAI21X1 _1677_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(_825_),
    .C(_863_),
    .Y(_864_)
);

MUX2X1 _1678_ (
    .A(ABCmd_i[1]),
    .B(_836_),
    .S(ABCmd_i[0]),
    .Y(_865_)
);

NAND2X1 _1679_ (
    .A(BI_0_bF$buf3),
    .B(_833_),
    .Y(_866_)
);

NAND2X1 _1680_ (
    .A(_866_),
    .B(_865_),
    .Y(_867_)
);

AOI21X1 _1681_ (
    .A(_832_),
    .B(_837_),
    .C(ABCmd_i[5]),
    .Y(_868_)
);

NAND2X1 _1682_ (
    .A(_868_),
    .B(_867_),
    .Y(_869_)
);

NAND3X1 _1683_ (
    .A(_840_),
    .B(_863_),
    .C(_869_),
    .Y(_870_)
);

AOI22X1 _1684_ (
    .A(_841_),
    .B(_864_),
    .C(_870_),
    .D(_827_),
    .Y(_871_)
);

OAI21X1 _1685_ (
    .A(_844_),
    .B(_857_),
    .C(_855_),
    .Y(_872_)
);

OAI21X1 _1686_ (
    .A(_855_),
    .B(_857_),
    .C(_872_),
    .Y(_873_)
);

NAND2X1 _1687_ (
    .A(_871_),
    .B(_873_),
    .Y(_874_)
);

NAND2X1 _1688_ (
    .A(_874_),
    .B(_861_),
    .Y(_875_)
);

INVX1 _1689_ (
    .A(_875_),
    .Y(ACC[1])
);

NOR2X1 _1690_ (
    .A(_857_),
    .B(_855_),
    .Y(_876_)
);

OAI21X1 _1691_ (
    .A(_876_),
    .B(_871_),
    .C(_872_),
    .Y(_877_)
);

NAND2X1 _1692_ (
    .A(ABCmd_i[5]),
    .B(AI[3]),
    .Y(_878_)
);

NAND3X1 _1693_ (
    .A(AI[2]),
    .B(BI[2]),
    .C(_831_),
    .Y(_879_)
);

AOI22X1 _1694_ (
    .A(_829_),
    .B(BI[2]),
    .C(_879_),
    .D(_830_),
    .Y(_880_)
);

INVX1 _1695_ (
    .A(BI[2]),
    .Y(_881_)
);

NOR2X1 _1696_ (
    .A(ABCmd_i[0]),
    .B(_881_),
    .Y(_882_)
);

OAI21X1 _1697_ (
    .A(AI[2]),
    .B(_882_),
    .C(_835_),
    .Y(_883_)
);

OAI21X1 _1698_ (
    .A(_880_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

OAI21X1 _1699_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[2]),
    .C(_825_),
    .Y(_885_)
);

AOI21X1 _1700_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI[2]),
    .C(_885_),
    .Y(_716_)
);

OAI21X1 _1701_ (
    .A(_844_),
    .B(_716_),
    .C(_884_),
    .Y(_717_)
);

OAI21X1 _1702_ (
    .A(_884_),
    .B(_716_),
    .C(_717_),
    .Y(_718_)
);

XOR2X1 _1703_ (
    .A(_877_),
    .B(_718_),
    .Y(_719_)
);

INVX1 _1704_ (
    .A(_719_),
    .Y(ACC[2])
);

INVX1 _1705_ (
    .A(_716_),
    .Y(_720_)
);

OAI21X1 _1706_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .C(_720_),
    .Y(_721_)
);

INVX1 _1707_ (
    .A(_718_),
    .Y(_722_)
);

AOI22X1 _1708_ (
    .A(_884_),
    .B(_721_),
    .C(_877_),
    .D(_722_),
    .Y(_723_)
);

NAND2X1 _1709_ (
    .A(ABCmd_i[5]),
    .B(AI[4]),
    .Y(_724_)
);

AND2X2 _1710_ (
    .A(_831_),
    .B(BI_3_bF$buf0),
    .Y(_725_)
);

NAND2X1 _1711_ (
    .A(AI[3]),
    .B(_725_),
    .Y(_726_)
);

AOI22X1 _1712_ (
    .A(_829_),
    .B(BI_3_bF$buf3),
    .C(_726_),
    .D(_830_),
    .Y(_727_)
);

OAI21X1 _1713_ (
    .A(AI[3]),
    .B(_725_),
    .C(_835_),
    .Y(_728_)
);

OAI21X1 _1714_ (
    .A(_728_),
    .B(_727_),
    .C(_724_),
    .Y(_729_)
);

OAI21X1 _1715_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI_3_bF$buf2),
    .C(_825_),
    .Y(_730_)
);

AOI21X1 _1716_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI_3_bF$buf1),
    .C(_730_),
    .Y(_731_)
);

OAI21X1 _1717_ (
    .A(_844_),
    .B(_731_),
    .C(_729_),
    .Y(_732_)
);

OAI21X1 _1718_ (
    .A(_729_),
    .B(_731_),
    .C(_732_),
    .Y(_733_)
);

XOR2X1 _1719_ (
    .A(_723_),
    .B(_733_),
    .Y(ACC[3])
);

XNOR2X1 _1720_ (
    .A(_723_),
    .B(_733_),
    .Y(_734_)
);

NAND2X1 _1721_ (
    .A(_718_),
    .B(_877_),
    .Y(_735_)
);

NAND3X1 _1722_ (
    .A(_872_),
    .B(_722_),
    .C(_861_),
    .Y(_736_)
);

NAND3X1 _1723_ (
    .A(_735_),
    .B(_875_),
    .C(_736_),
    .Y(_737_)
);

NAND2X1 _1724_ (
    .A(ABCmd_i[6]),
    .B(_737_),
    .Y(_738_)
);

OAI21X1 _1725_ (
    .A(_733_),
    .B(_723_),
    .C(_732_),
    .Y(_739_)
);

INVX1 _1726_ (
    .A(_739_),
    .Y(_740_)
);

OAI21X1 _1727_ (
    .A(_738_),
    .B(_734_),
    .C(_740_),
    .Y(HC)
);

NAND2X1 _1728_ (
    .A(ABCmd_i[5]),
    .B(AI_5_bF$buf0),
    .Y(_741_)
);

AND2X2 _1729_ (
    .A(_831_),
    .B(BI_4_bF$buf3),
    .Y(_742_)
);

NAND2X1 _1730_ (
    .A(AI[4]),
    .B(_742_),
    .Y(_743_)
);

AOI22X1 _1731_ (
    .A(_829_),
    .B(BI_4_bF$buf2),
    .C(_743_),
    .D(_830_),
    .Y(_744_)
);

OAI21X1 _1732_ (
    .A(AI[4]),
    .B(_742_),
    .C(_835_),
    .Y(_745_)
);

OAI21X1 _1733_ (
    .A(_745_),
    .B(_744_),
    .C(_741_),
    .Y(_746_)
);

OAI21X1 _1734_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_4_bF$buf1),
    .C(_825_),
    .Y(_747_)
);

AOI21X1 _1735_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI_4_bF$buf0),
    .C(_747_),
    .Y(_748_)
);

OAI21X1 _1736_ (
    .A(_844_),
    .B(_748_),
    .C(_746_),
    .Y(_749_)
);

OAI21X1 _1737_ (
    .A(_746_),
    .B(_748_),
    .C(_749_),
    .Y(_750_)
);

INVX1 _1738_ (
    .A(_750_),
    .Y(_751_)
);

XOR2X1 _1739_ (
    .A(HC),
    .B(_751_),
    .Y(ACC[4])
);

INVX1 _1740_ (
    .A(_749_),
    .Y(_752_)
);

AOI21X1 _1741_ (
    .A(HC),
    .B(_751_),
    .C(_752_),
    .Y(_753_)
);

NAND2X1 _1742_ (
    .A(ABCmd_i[5]),
    .B(AI[6]),
    .Y(_754_)
);

AND2X2 _1743_ (
    .A(_831_),
    .B(BI[5]),
    .Y(_755_)
);

NAND2X1 _1744_ (
    .A(AI_5_bF$buf3),
    .B(_755_),
    .Y(_756_)
);

AOI22X1 _1745_ (
    .A(_829_),
    .B(BI[5]),
    .C(_756_),
    .D(_830_),
    .Y(_757_)
);

OAI21X1 _1746_ (
    .A(AI_5_bF$buf2),
    .B(_755_),
    .C(_835_),
    .Y(_758_)
);

OAI21X1 _1747_ (
    .A(_758_),
    .B(_757_),
    .C(_754_),
    .Y(_759_)
);

OAI21X1 _1748_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[5]),
    .C(_825_),
    .Y(_760_)
);

AOI21X1 _1749_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[5]),
    .C(_760_),
    .Y(_761_)
);

OAI21X1 _1750_ (
    .A(_844_),
    .B(_761_),
    .C(_759_),
    .Y(_762_)
);

OAI21X1 _1751_ (
    .A(_759_),
    .B(_761_),
    .C(_762_),
    .Y(_763_)
);

INVX1 _1752_ (
    .A(_763_),
    .Y(_764_)
);

XOR2X1 _1753_ (
    .A(_753_),
    .B(_764_),
    .Y(_765_)
);

INVX1 _1754_ (
    .A(_765_),
    .Y(ACC[5])
);

OAI21X1 _1755_ (
    .A(_763_),
    .B(_753_),
    .C(_762_),
    .Y(_766_)
);

INVX1 _1756_ (
    .A(\u_ALU.AI7 ),
    .Y(_767_)
);

AND2X2 _1757_ (
    .A(_831_),
    .B(BI[6]),
    .Y(_768_)
);

NAND2X1 _1758_ (
    .A(AI[6]),
    .B(_768_),
    .Y(_769_)
);

AOI22X1 _1759_ (
    .A(_829_),
    .B(BI[6]),
    .C(_769_),
    .D(_830_),
    .Y(_770_)
);

OAI21X1 _1760_ (
    .A(AI[6]),
    .B(_768_),
    .C(_835_),
    .Y(_771_)
);

OAI22X1 _1761_ (
    .A(_835_),
    .B(_767_),
    .C(_771_),
    .D(_770_),
    .Y(_772_)
);

OAI21X1 _1762_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI[6]),
    .C(_825_),
    .Y(_773_)
);

AOI21X1 _1763_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI[6]),
    .C(_773_),
    .Y(_774_)
);

OAI21X1 _1764_ (
    .A(_844_),
    .B(_774_),
    .C(_772_),
    .Y(_775_)
);

OAI21X1 _1765_ (
    .A(_772_),
    .B(_774_),
    .C(_775_),
    .Y(_776_)
);

NAND2X1 _1766_ (
    .A(_776_),
    .B(_766_),
    .Y(_777_)
);

INVX1 _1767_ (
    .A(ABCmd_i[6]),
    .Y(_778_)
);

AOI21X1 _1768_ (
    .A(_719_),
    .B(_875_),
    .C(_778_),
    .Y(_779_)
);

AOI21X1 _1769_ (
    .A(_779_),
    .B(ACC[3]),
    .C(_739_),
    .Y(_780_)
);

OAI21X1 _1770_ (
    .A(_750_),
    .B(_780_),
    .C(_749_),
    .Y(_781_)
);

OR2X2 _1771_ (
    .A(_761_),
    .B(_844_),
    .Y(_782_)
);

AOI22X1 _1772_ (
    .A(_759_),
    .B(_782_),
    .C(_781_),
    .D(_764_),
    .Y(_783_)
);

INVX1 _1773_ (
    .A(_776_),
    .Y(_784_)
);

NAND2X1 _1774_ (
    .A(_784_),
    .B(_783_),
    .Y(_785_)
);

NAND2X1 _1775_ (
    .A(_777_),
    .B(_785_),
    .Y(ACC[6])
);

OAI21X1 _1776_ (
    .A(_776_),
    .B(_783_),
    .C(_775_),
    .Y(_786_)
);

NAND2X1 _1777_ (
    .A(ABCmd_i[5]),
    .B(ABCmd_i[4]),
    .Y(_787_)
);

AND2X2 _1778_ (
    .A(_831_),
    .B(BI[7]),
    .Y(_788_)
);

NAND2X1 _1779_ (
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .Y(_789_)
);

AOI22X1 _1780_ (
    .A(_829_),
    .B(BI[7]),
    .C(_789_),
    .D(_830_),
    .Y(_790_)
);

OAI21X1 _1781_ (
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .C(_835_),
    .Y(_791_)
);

OAI21X1 _1782_ (
    .A(_791_),
    .B(_790_),
    .C(_787_),
    .Y(_792_)
);

OAI21X1 _1783_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[7]),
    .C(_825_),
    .Y(_793_)
);

AOI21X1 _1784_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[7]),
    .C(_793_),
    .Y(_794_)
);

OAI21X1 _1785_ (
    .A(_844_),
    .B(_794_),
    .C(_792_),
    .Y(_795_)
);

OAI21X1 _1786_ (
    .A(_792_),
    .B(_794_),
    .C(_795_),
    .Y(_796_)
);

NAND2X1 _1787_ (
    .A(_796_),
    .B(_786_),
    .Y(_797_)
);

NAND2X1 _1788_ (
    .A(_784_),
    .B(_766_),
    .Y(_798_)
);

INVX1 _1789_ (
    .A(_796_),
    .Y(_799_)
);

NAND3X1 _1790_ (
    .A(_775_),
    .B(_799_),
    .C(_798_),
    .Y(_800_)
);

NAND2X1 _1791_ (
    .A(_800_),
    .B(_797_),
    .Y(AN)
);

NOR2X1 _1792_ (
    .A(ACC[0]),
    .B(_737_),
    .Y(_801_)
);

NAND2X1 _1793_ (
    .A(_734_),
    .B(_801_),
    .Y(_802_)
);

NOR2X1 _1794_ (
    .A(_802_),
    .B(ACC[4]),
    .Y(_803_)
);

NAND3X1 _1795_ (
    .A(_765_),
    .B(_777_),
    .C(_785_),
    .Y(_804_)
);

NOR2X1 _1796_ (
    .A(_804_),
    .B(AN),
    .Y(_805_)
);

AND2X2 _1797_ (
    .A(_805_),
    .B(_803_),
    .Y(AZ)
);

NAND3X1 _1798_ (
    .A(_775_),
    .B(_796_),
    .C(_798_),
    .Y(_806_)
);

NAND2X1 _1799_ (
    .A(_799_),
    .B(_786_),
    .Y(_807_)
);

NAND2X1 _1800_ (
    .A(_806_),
    .B(_807_),
    .Y(_808_)
);

NAND2X1 _1801_ (
    .A(ABCmd_i[6]),
    .B(_804_),
    .Y(_809_)
);

NOR2X1 _1802_ (
    .A(_837_),
    .B(_835_),
    .Y(_810_)
);

OAI21X1 _1803_ (
    .A(_775_),
    .B(_796_),
    .C(_795_),
    .Y(_811_)
);

NOR2X1 _1804_ (
    .A(_796_),
    .B(_776_),
    .Y(_812_)
);

AOI21X1 _1805_ (
    .A(_766_),
    .B(_812_),
    .C(_811_),
    .Y(_813_)
);

XOR2X1 _1806_ (
    .A(_813_),
    .B(_810_),
    .Y(_814_)
);

OAI21X1 _1807_ (
    .A(_809_),
    .B(_808_),
    .C(_814_),
    .Y(CO)
);

NAND3X1 _1808_ (
    .A(ABCmd_i[6]),
    .B(_804_),
    .C(AN),
    .Y(_815_)
);

AOI21X1 _1809_ (
    .A(_792_),
    .B(_844_),
    .C(_794_),
    .Y(_816_)
);

XOR2X1 _1810_ (
    .A(_816_),
    .B(_767_),
    .Y(_817_)
);

NAND3X1 _1811_ (
    .A(_800_),
    .B(_817_),
    .C(_797_),
    .Y(_818_)
);

INVX1 _1812_ (
    .A(_817_),
    .Y(_819_)
);

NAND3X1 _1813_ (
    .A(_806_),
    .B(_819_),
    .C(_807_),
    .Y(_820_)
);

NAND2X1 _1814_ (
    .A(_818_),
    .B(_820_),
    .Y(_821_)
);

NAND3X1 _1815_ (
    .A(_814_),
    .B(_815_),
    .C(_821_),
    .Y(_822_)
);

NAND3X1 _1816_ (
    .A(_818_),
    .B(_820_),
    .C(CO),
    .Y(_823_)
);

NAND2X1 _1817_ (
    .A(_822_),
    .B(_823_),
    .Y(AV)
);

BUFX2 _1818_ (
    .A(_886_[0]),
    .Y(ACC_o[0])
);

BUFX2 _1819_ (
    .A(_886_[1]),
    .Y(ACC_o[1])
);

BUFX2 _1820_ (
    .A(_886_[2]),
    .Y(ACC_o[2])
);

BUFX2 _1821_ (
    .A(_886_[3]),
    .Y(ACC_o[3])
);

BUFX2 _1822_ (
    .A(_886_[4]),
    .Y(ACC_o[4])
);

BUFX2 _1823_ (
    .A(_886_[5]),
    .Y(ACC_o[5])
);

BUFX2 _1824_ (
    .A(_886_[6]),
    .Y(ACC_o[6])
);

BUFX2 _1825_ (
    .A(_886_[7]),
    .Y(ACC_o[7])
);

BUFX2 _1826_ (
    .A(_887_),
    .Y(Done_o)
);

INVX1 _889_ (
    .A(state[2]),
    .Y(_699_)
);

NOR2X1 _890_ (
    .A(state[0]),
    .B(_699_),
    .Y(_700_)
);

NAND2X1 _891_ (
    .A(state[1]),
    .B(_700_),
    .Y(_701_)
);

INVX1 _892_ (
    .A(_701_),
    .Y(_887_)
);

INVX1 _893_ (
    .A(state[0]),
    .Y(_702_)
);

INVX2 _894_ (
    .A(state[1]),
    .Y(_703_)
);

NOR2X1 _895_ (
    .A(state[2]),
    .B(_703_),
    .Y(_704_)
);

NAND2X1 _896_ (
    .A(_702_),
    .B(_704_),
    .Y(_705_)
);

INVX1 _897_ (
    .A(_705__bF$buf3),
    .Y(_706_)
);

NOR2X1 _898_ (
    .A(state[2]),
    .B(_702_),
    .Y(_707_)
);

AOI21X1 _899_ (
    .A(_703_),
    .B(_707_),
    .C(_887_),
    .Y(_708_)
);

NOR2X1 _900_ (
    .A(LoadCmd_i),
    .B(_708_),
    .Y(_709_)
);

OAI21X1 _901_ (
    .A(_706_),
    .B(_709_),
    .C(LoadB_i),
    .Y(_710_)
);

INVX1 _902_ (
    .A(LoadA_i),
    .Y(_711_)
);

INVX4 _903_ (
    .A(_700_),
    .Y(_712_)
);

OAI21X1 _904_ (
    .A(state[1]),
    .B(state[0]),
    .C(_699_),
    .Y(_713_)
);

INVX1 _905_ (
    .A(LoadB_i),
    .Y(_714_)
);

NOR2X1 _906_ (
    .A(state[1]),
    .B(_712_),
    .Y(_715_)
);

INVX1 _907_ (
    .A(_715_),
    .Y(_25_)
);

INVX1 _908_ (
    .A(LoadCmd_i),
    .Y(_26_)
);

OAI21X1 _909_ (
    .A(_707_),
    .B(_887_),
    .C(_26_),
    .Y(_27_)
);

OAI21X1 _910_ (
    .A(_714_),
    .B(_25_),
    .C(_27_),
    .Y(_28_)
);

AOI22X1 _911_ (
    .A(_712_),
    .B(_713_),
    .C(_28_),
    .D(_711_),
    .Y(_29_)
);

NAND2X1 _912_ (
    .A(_29_),
    .B(_710_),
    .Y(_888_[0])
);

OAI21X1 _913_ (
    .A(LoadA_i),
    .B(LoadB_i),
    .C(_26_),
    .Y(_30_)
);

OAI21X1 _914_ (
    .A(_30_),
    .B(_708_),
    .C(_25_),
    .Y(_31_)
);

NAND2X1 _915_ (
    .A(state[1]),
    .B(_707_),
    .Y(_32_)
);

NOR2X1 _916_ (
    .A(LoadA_i),
    .B(_26_),
    .Y(_33_)
);

NOR2X1 _917_ (
    .A(LoadB_i),
    .B(_26_),
    .Y(_34_)
);

OAI22X1 _918_ (
    .A(_33_),
    .B(_32__bF$buf3),
    .C(_705__bF$buf2),
    .D(_34_),
    .Y(_35_)
);

OR2X2 _919_ (
    .A(_31_),
    .B(_35_),
    .Y(_888_[1])
);

INVX1 _920_ (
    .A(_32__bF$buf2),
    .Y(_36_)
);

AOI22X1 _921_ (
    .A(_36_),
    .B(_33_),
    .C(_706_),
    .D(_34_),
    .Y(_37_)
);

NAND3X1 _922_ (
    .A(_711_),
    .B(_714_),
    .C(_715_),
    .Y(_38_)
);

AND2X2 _923_ (
    .A(_37_),
    .B(_38_),
    .Y(_39_)
);

OAI21X1 _924_ (
    .A(_26_),
    .B(_708_),
    .C(_39_),
    .Y(_888_[2])
);

INVX8 _925_ (
    .A(reset),
    .Y(_0_)
);

INVX1 _926_ (
    .A(ABCmd_i[0]),
    .Y(_40_)
);

NAND2X1 _927_ (
    .A(BI_0_bF$buf2),
    .B(_32__bF$buf1),
    .Y(_41_)
);

OAI21X1 _928_ (
    .A(_40_),
    .B(_32__bF$buf0),
    .C(_41_),
    .Y(_1_)
);

INVX1 _929_ (
    .A(ABCmd_i[1]),
    .Y(_42_)
);

NAND2X1 _930_ (
    .A(BI_1_bF$buf3),
    .B(_32__bF$buf3),
    .Y(_43_)
);

OAI21X1 _931_ (
    .A(_42_),
    .B(_32__bF$buf2),
    .C(_43_),
    .Y(_2_)
);

INVX1 _932_ (
    .A(ABCmd_i_2_bF$buf2),
    .Y(_44_)
);

NAND2X1 _933_ (
    .A(BI[2]),
    .B(_32__bF$buf1),
    .Y(_45_)
);

OAI21X1 _934_ (
    .A(_44_),
    .B(_32__bF$buf0),
    .C(_45_),
    .Y(_3_)
);

INVX1 _935_ (
    .A(ABCmd_i[3]),
    .Y(_46_)
);

NAND2X1 _936_ (
    .A(BI_3_bF$buf0),
    .B(_32__bF$buf3),
    .Y(_47_)
);

OAI21X1 _937_ (
    .A(_46_),
    .B(_32__bF$buf2),
    .C(_47_),
    .Y(_4_)
);

INVX1 _938_ (
    .A(ABCmd_i[4]),
    .Y(_48_)
);

NAND2X1 _939_ (
    .A(BI_4_bF$buf3),
    .B(_32__bF$buf1),
    .Y(_49_)
);

OAI21X1 _940_ (
    .A(_48_),
    .B(_32__bF$buf0),
    .C(_49_),
    .Y(_5_)
);

INVX1 _941_ (
    .A(ABCmd_i[5]),
    .Y(_50_)
);

NAND2X1 _942_ (
    .A(BI[5]),
    .B(_32__bF$buf3),
    .Y(_51_)
);

OAI21X1 _943_ (
    .A(_50_),
    .B(_32__bF$buf2),
    .C(_51_),
    .Y(_6_)
);

INVX1 _944_ (
    .A(ABCmd_i[6]),
    .Y(_52_)
);

NAND2X1 _945_ (
    .A(BI[6]),
    .B(_32__bF$buf1),
    .Y(_53_)
);

OAI21X1 _946_ (
    .A(_52_),
    .B(_32__bF$buf0),
    .C(_53_),
    .Y(_7_)
);

INVX4 _947_ (
    .A(ABCmd_i[7]),
    .Y(_54_)
);

NAND2X1 _948_ (
    .A(BI[7]),
    .B(_32__bF$buf3),
    .Y(_55_)
);

OAI21X1 _949_ (
    .A(_54_),
    .B(_32__bF$buf2),
    .C(_55_),
    .Y(_8_)
);

INVX1 _950_ (
    .A(_886_[0]),
    .Y(_56_)
);

INVX1 _951_ (
    .A(AI[0]),
    .Y(_57_)
);

INVX2 _952_ (
    .A(BI_3_bF$buf3),
    .Y(_58_)
);

NOR2X1 _953_ (
    .A(_57_),
    .B(_58_),
    .Y(_59_)
);

AND2X2 _954_ (
    .A(BI_4_bF$buf2),
    .B(AI[1]),
    .Y(_60_)
);

NAND2X1 _955_ (
    .A(_60_),
    .B(_59_),
    .Y(_61_)
);

NAND2X1 _956_ (
    .A(BI_1_bF$buf2),
    .B(AI[2]),
    .Y(_62_)
);

NAND2X1 _957_ (
    .A(BI_0_bF$buf1),
    .B(AI[3]),
    .Y(_63_)
);

OR2X2 _958_ (
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

NAND2X1 _959_ (
    .A(BI[2]),
    .B(AI[1]),
    .Y(_65_)
);

AND2X2 _960_ (
    .A(_62_),
    .B(_63_),
    .Y(_66_)
);

OAI21X1 _961_ (
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

NAND2X1 _962_ (
    .A(BI[2]),
    .B(AI[2]),
    .Y(_68_)
);

INVX1 _963_ (
    .A(_68_),
    .Y(_69_)
);

NAND2X1 _964_ (
    .A(BI_1_bF$buf1),
    .B(AI[3]),
    .Y(_70_)
);

NAND2X1 _965_ (
    .A(BI_0_bF$buf0),
    .B(AI[4]),
    .Y(_71_)
);

OR2X2 _966_ (
    .A(_70_),
    .B(_71_),
    .Y(_72_)
);

INVX1 _967_ (
    .A(BI_0_bF$buf3),
    .Y(_73_)
);

INVX1 _968_ (
    .A(AI[4]),
    .Y(_74_)
);

OAI21X1 _969_ (
    .A(_73_),
    .B(_74_),
    .C(_70_),
    .Y(_75_)
);

NAND3X1 _970_ (
    .A(_75_),
    .B(_69_),
    .C(_72_),
    .Y(_76_)
);

NOR2X1 _971_ (
    .A(_70_),
    .B(_71_),
    .Y(_77_)
);

AND2X2 _972_ (
    .A(_70_),
    .B(_71_),
    .Y(_78_)
);

OAI21X1 _973_ (
    .A(_77_),
    .B(_78_),
    .C(_68_),
    .Y(_79_)
);

NAND3X1 _974_ (
    .A(_79_),
    .B(_67_),
    .C(_76_),
    .Y(_80_)
);

INVX1 _975_ (
    .A(_59_),
    .Y(_81_)
);

NAND2X1 _976_ (
    .A(BI_4_bF$buf1),
    .B(AI[1]),
    .Y(_82_)
);

INVX2 _977_ (
    .A(BI_4_bF$buf0),
    .Y(_83_)
);

NAND2X1 _978_ (
    .A(BI_3_bF$buf2),
    .B(AI[1]),
    .Y(_84_)
);

OAI21X1 _979_ (
    .A(_57_),
    .B(_83_),
    .C(_84_),
    .Y(_85_)
);

OAI21X1 _980_ (
    .A(_82_),
    .B(_81_),
    .C(_85_),
    .Y(_86_)
);

AOI21X1 _981_ (
    .A(_76_),
    .B(_79_),
    .C(_67_),
    .Y(_87_)
);

OAI21X1 _982_ (
    .A(_86_),
    .B(_87_),
    .C(_80_),
    .Y(_88_)
);

OAI21X1 _983_ (
    .A(_68_),
    .B(_78_),
    .C(_72_),
    .Y(_89_)
);

AND2X2 _984_ (
    .A(BI_0_bF$buf2),
    .B(AI_5_bF$buf1),
    .Y(_90_)
);

NAND3X1 _985_ (
    .A(BI_1_bF$buf0),
    .B(AI[4]),
    .C(_90_),
    .Y(_91_)
);

AOI22X1 _986_ (
    .A(BI_0_bF$buf1),
    .B(AI_5_bF$buf0),
    .C(BI_1_bF$buf3),
    .D(AI[4]),
    .Y(_92_)
);

INVX1 _987_ (
    .A(_92_),
    .Y(_93_)
);

NAND2X1 _988_ (
    .A(BI[2]),
    .B(AI[3]),
    .Y(_94_)
);

INVX1 _989_ (
    .A(_94_),
    .Y(_95_)
);

NAND3X1 _990_ (
    .A(_93_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

NAND2X1 _991_ (
    .A(BI_1_bF$buf2),
    .B(AI_5_bF$buf3),
    .Y(_97_)
);

NOR2X1 _992_ (
    .A(_71_),
    .B(_97_),
    .Y(_98_)
);

OAI21X1 _993_ (
    .A(_92_),
    .B(_98_),
    .C(_94_),
    .Y(_99_)
);

NAND3X1 _994_ (
    .A(_96_),
    .B(_99_),
    .C(_89_),
    .Y(_100_)
);

AOI21X1 _995_ (
    .A(_69_),
    .B(_75_),
    .C(_77_),
    .Y(_101_)
);

OAI21X1 _996_ (
    .A(_92_),
    .B(_98_),
    .C(_95_),
    .Y(_102_)
);

NAND3X1 _997_ (
    .A(_93_),
    .B(_94_),
    .C(_91_),
    .Y(_103_)
);

NAND3X1 _998_ (
    .A(_103_),
    .B(_102_),
    .C(_101_),
    .Y(_104_)
);

NAND2X1 _999_ (
    .A(AI[0]),
    .B(BI[5]),
    .Y(_105_)
);

endmodule
