magic
tech scmos
magscale 1 60
timestamp 1709416183
<< checkpaint >>
rect -1200 -1200 381200 381200
<< metal1 >>
rect 89200 183200 96400 196700
rect 287000 180600 290700 199400
<< m2contact >>
rect 88400 183200 89200 196700
rect 290700 180600 291700 199400
<< metal2 >>
rect 119600 291400 120400 291800
rect 94200 290600 120400 291400
rect 88200 259600 93600 260400
rect 88200 232600 92400 233400
rect 88200 227200 91200 228000
rect 90600 211600 91200 227200
rect 91800 217600 92400 232600
rect 93000 233200 93600 259600
rect 94200 237800 94800 290600
rect 146600 289800 147200 291800
rect 114000 289000 147200 289800
rect 114000 286000 114800 289000
rect 173600 288200 174400 291800
rect 127200 287400 174400 288200
rect 127200 286000 128000 287400
rect 200600 286600 201400 291800
rect 227600 291400 228400 291800
rect 154200 285800 201400 286600
rect 217200 290800 228400 291400
rect 217200 285800 217800 290800
rect 254600 290200 255400 291800
rect 221400 289600 255400 290200
rect 221400 286000 222000 289600
rect 281600 289000 282300 291800
rect 228600 288300 282300 289000
rect 228600 285800 229400 288300
rect 230400 286900 291200 287600
rect 230400 285800 231100 286900
rect 236500 285800 290100 286500
rect 288400 206400 289000 258600
rect 289500 233400 290100 285800
rect 290600 260400 291200 286900
rect 290600 259700 291800 260400
rect 289500 232800 291800 233400
rect 288400 205700 291700 206400
rect 90600 152400 91200 170100
rect 88200 151600 91200 152400
rect 92300 147000 92900 178000
rect 88200 146200 92900 147000
rect 93800 120000 94400 176300
rect 88200 119200 94400 120000
rect 99600 89500 100200 96500
rect 102100 91903 102700 96400
rect 102098 91900 102700 91903
rect 102100 90703 102700 91900
rect 104500 91903 105100 96400
rect 108100 93103 108700 96400
rect 117000 94303 117600 96400
rect 132100 95503 132700 96400
rect 132100 95500 232900 95503
rect 132100 94900 233708 95500
rect 117000 93700 206700 94303
rect 108096 93100 179700 93103
rect 108100 92500 179700 93100
rect 104500 91300 152700 91903
rect 102100 90100 125700 90703
rect 98000 88886 100200 89500
rect 98000 88300 98700 88886
rect 125000 88300 125700 90100
rect 152000 88300 152700 91300
rect 179000 88300 179700 92500
rect 206000 88300 206700 93700
rect 233000 89002 233708 94900
rect 232994 88876 233708 89002
rect 232994 88294 233703 88876
<< m3contact >>
rect 94200 236400 94800 237800
rect 288400 258600 289000 259800
rect 93000 231800 93600 233200
rect 91800 216200 92400 217600
rect 90600 210200 91200 211600
rect 92300 178000 92900 179400
rect 90600 170100 91200 171600
rect 93800 176300 94400 177700
<< metal3 >>
rect 284980 259480 288400 259720
rect 94800 236440 98520 236680
rect 93600 231880 98320 232120
rect 92400 216280 98520 216520
rect 91200 210280 98320 210520
rect 92900 179080 98720 179320
rect 94400 177340 97320 177580
rect 91200 171200 97000 171600
<< comment >>
rect 0 0 380000 380000
use PIC  ABCMD_I_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1699925102
transform 1 0 259000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_1
timestamp 1699925102
transform 0 -1 342200 -1 0 229000
box -200 -18300 24200 50600
use PIC  ABCMD_I_2
timestamp 1699925102
transform 0 -1 342200 -1 0 256000
box -200 -18300 24200 50600
use PIC  ABCMD_I_3
timestamp 1699925102
transform 0 -1 342200 -1 0 283000
box -200 -18300 24200 50600
use PIC  ABCMD_I_4
timestamp 1699925102
transform 1 0 232000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_5
timestamp 1699925102
transform 1 0 205000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_6
timestamp 1699925102
transform 1 0 151000 0 -1 342200
box -200 -18300 24200 50600
use PIC  ABCMD_I_7
timestamp 1699925102
transform 1 0 178000 0 -1 342200
box -200 -18300 24200 50600
use POB8  ACC_O_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1699924048
transform 0 1 37800 -1 0 148000
box -200 -18300 24200 50600
use POB8  ACC_O_1
timestamp 1699924048
transform 0 1 37800 -1 0 121000
box -200 -18300 24200 50600
use POB8  ACC_O_2
timestamp 1699924048
transform 0 1 37800 -1 0 229000
box -200 -18300 24200 50600
use POB8  ACC_O_3
timestamp 1699924048
transform 1 0 205000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_4
timestamp 1699924048
transform 1 0 178000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_5
timestamp 1699924048
transform 1 0 151000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_6
timestamp 1699924048
transform 1 0 124000 0 1 37800
box -200 -18300 24200 50600
use POB8  ACC_O_7
timestamp 1699924048
transform 1 0 97000 0 1 37800
box -200 -18300 24200 50600
use ALU_wrapper_Core  ALU_wrapper_Core_0
timestamp 1709017741
transform 1 0 98100 0 1 97000
box -1890 -720 189090 189090
use PIC  CLK
timestamp 1699925102
transform 0 1 37800 -1 0 175000
box -200 -18300 24200 50600
use POB8  DONE_O
timestamp 1699924048
transform 1 0 232000 0 1 37800
box -200 -18300 24200 50600
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 -1 342200 -1 0 175360
box -70 0 2070 50120
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1709081121
transform 1 0 120690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_1
timestamp 1709081121
transform 0 1 37800 -1 0 151309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_2
timestamp 1709081121
transform 1 0 174690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_3
timestamp 1709081121
transform 1 0 147690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_4
timestamp 1709081121
transform 1 0 228690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_5
timestamp 1709081121
transform 1 0 201690 0 1 37800
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_6
timestamp 1709081121
transform 0 1 37800 -1 0 124309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_8
timestamp 1709081121
transform 0 1 37800 -1 0 205309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_9
timestamp 1709081121
transform 0 1 37800 -1 0 178309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_10
timestamp 1709081121
transform 0 1 37800 -1 0 259309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_11
timestamp 1709081121
transform 0 1 37800 -1 0 232309
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_14
timestamp 1709081121
transform 0 -1 342200 -1 0 205305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_15
timestamp 1709081121
transform 0 -1 342200 -1 0 178305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_16
timestamp 1709081121
transform 0 -1 342200 -1 0 259305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_17
timestamp 1709081121
transform 0 -1 342200 -1 0 232305
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_18
timestamp 1709081121
transform 1 0 147690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_19
timestamp 1709081121
transform 1 0 120690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_20
timestamp 1709081121
transform 1 0 201690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_21
timestamp 1709081121
transform 1 0 174690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_22
timestamp 1709081121
transform 1 0 255690 0 -1 342200
box 0 0 3620 50120
use IOFILLER18  IOFILLER18_23
timestamp 1709081121
transform 1 0 228690 0 -1 342200
box 0 0 3620 50120
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 1 0 87287 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_1
timestamp 1692859860
transform 0 1 37800 -1 0 97233
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_2
timestamp 1692859860
transform 1 0 255648 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_3
timestamp 1692859860
transform 0 1 37800 -1 0 292759
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_4
timestamp 1692859860
transform 1 0 87417 0 -1 342200
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_5
timestamp 1692859860
transform 1 0 282662 0 -1 342199
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_6
timestamp 1692859860
transform 0 -1 342200 -1 0 97270
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_7
timestamp 1692859860
transform 0 -1 342200 -1 0 292717
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_8
timestamp 1692859860
transform 0 -1 342200 -1 0 164305
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_9
timestamp 1692859860
transform 0 -1 342200 -1 0 106780
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_10
timestamp 1692859860
transform 0 -1 342200 -1 0 116305
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_11
timestamp 1692859860
transform 0 -1 342200 -1 0 125905
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_12
timestamp 1692859860
transform 0 -1 342200 -1 0 135505
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_13
timestamp 1692859860
transform 0 -1 342200 -1 0 145105
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_14
timestamp 1692859860
transform 0 -1 342200 -1 0 154705
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_15
timestamp 1692859860
transform 0 -1 342200 -1 0 173905
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_16
timestamp 1692859860
transform 1 0 282762 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_17
timestamp 1692859860
transform 1 0 273362 0 1 37800
box -70 0 10070 50120
use IOFILLER50  IOFILLER50_18
timestamp 1692859860
transform 1 0 263968 0 1 37800
box -70 0 10070 50120
use PIC  LOADA_I
timestamp 1699925102
transform 1 0 97000 0 -1 342200
box -200 -18300 24200 50600
use PIC  LOADB_I
timestamp 1699925102
transform 0 1 37800 -1 0 283000
box -200 -18300 24200 50600
use PIC  LOADCMD_I
timestamp 1699925102
transform 1 0 124000 0 -1 342200
box -200 -18300 24200 50600
use MY_LOGO  MY_LOGO_0
timestamp 1700409309
transform 1 0 299100 0 1 21600
box 0 0 40680 14580
use PAD80  PAD80_2 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1709379016
transform 1 0 262500 0 1 19500
box 0 0 17000 17000
use PAD80  PAD80_6
timestamp 1709379016
transform 1 0 343500 0 1 127500
box 0 0 17000 17000
use PAD80  PAD80_7
timestamp 1709379016
transform 1 0 343500 0 1 100500
box 0 0 17000 17000
use PAD80  PAD80_17
timestamp 1709379016
transform 1 0 343500 0 1 154500
box 0 0 17000 17000
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 1 0 37800 0 1 37800
box 0 0 50600 50600
use PCORNER  PCORNER_1
timestamp 1692859860
transform -1 0 342200 0 1 37800
box 0 0 50600 50600
use PCORNER  PCORNER_2
timestamp 1692859860
transform 0 1 37800 -1 0 342200
box 0 0 50600 50600
use PCORNER  PCORNER_3
timestamp 1692859860
transform 0 -1 342200 -1 0 342200
box 0 0 50600 50600
use PVSS  PVSS_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 -1 342200 -1 0 202000
box 0 -18300 24000 50600
use PIC  RESET
timestamp 1699925102
transform 0 1 37800 -1 0 256000
box -200 -18300 24200 50600
use PVDD  VDD_0 ~/ETRI050_DesignKit/devel/Ref_Design/ALU8/chiptop/pads_ETRI050
timestamp 1692859860
transform 0 1 37800 -1 0 202000
box 0 -18300 24000 50600
<< end >>
