/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module ALU_wrapper(
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    output Done_LED,
    output Done_o,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input clk,
    input reset
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire BI_0_bF$buf0 ;
wire BI_0_bF$buf1 ;
wire BI_0_bF$buf2 ;
wire BI_0_bF$buf3 ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire \u_ALU.AI7  ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire ABCmd_i_2_bF$buf0 ;
wire ABCmd_i_2_bF$buf1 ;
wire ABCmd_i_2_bF$buf2 ;
wire ABCmd_i_2_bF$buf3 ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _705__bF$buf0 ;
wire _705__bF$buf1 ;
wire _705__bF$buf2 ;
wire _705__bF$buf3 ;
wire _878_ ;
wire _458_ ;
wire _32__bF$buf0 ;
wire _32__bF$buf1 ;
wire _32__bF$buf2 ;
wire _32__bF$buf3 ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire Done_o ;
wire _740_ ;
wire _320_ ;
wire AI_5_bF$buf0 ;
wire AI_5_bF$buf1 ;
wire AI_5_bF$buf2 ;
wire AI_5_bF$buf3 ;
wire _56_ ;
wire _605_ ;
wire BI_4_bF$buf0 ;
wire BI_4_bF$buf1 ;
wire BI_4_bF$buf2 ;
wire BI_4_bF$buf3 ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire [7:0] _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _713_ ;
wire [6:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire BI_1_bF$buf0 ;
wire BI_1_bF$buf1 ;
wire BI_1_bF$buf2 ;
wire BI_1_bF$buf3 ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [2:0] state ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire [6:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire Done_LED ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire BI_3_bF$buf0 ;
wire BI_3_bF$buf1 ;
wire BI_3_bF$buf2 ;
wire BI_3_bF$buf3 ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire [2:0] _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _0__bF$buf0 ;
wire _0__bF$buf1 ;
wire _0__bF$buf2 ;
wire _0__bF$buf3 ;
wire _0__bF$buf4 ;
wire _22_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_0__1661_ (
);

FILL FILL_2__1679_ (
);

FILL FILL_0__1241_ (
);

FILL FILL_2__1259_ (
);

FILL FILL_1__1822_ (
);

FILL FILL_1__1402_ (
);

OAI21X1 _1677_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .C(_863_),
    .Y(_864_)
);

AOI22X1 _1257_ (
    .A(_321_),
    .B(_324_),
    .C(_358_),
    .D(_359_),
    .Y(_363_)
);

FILL FILL_0__1717_ (
);

FILL FILL_2__1488_ (
);

FILL FILL_0__1470_ (
);

FILL FILL_0__1050_ (
);

FILL FILL_2__1068_ (
);

FILL FILL_3__941_ (
);

FILL FILL_1__1211_ (
);

FILL FILL_3__1137_ (
);

AOI22X1 _1486_ (
    .A(_538_),
    .B(_712_),
    .C(_582_),
    .D(_588_),
    .Y(_12_)
);

NAND3X1 _1066_ (
    .A(_162_),
    .B(_166_),
    .C(_171_),
    .Y(_172_)
);

FILL FILL_2__1700_ (
);

FILL FILL_0__1526_ (
);

FILL FILL_0__1106_ (
);

FILL FILL_2__1297_ (
);

FILL FILL_1__1440_ (
);

FILL FILL_1__1020_ (
);

FILL FILL_3__1786_ (
);

FILL FILL_3__1366_ (
);

FILL FILL94050x82050 (
);

AOI21X1 _1295_ (
    .A(_313_),
    .B(_365_),
    .C(_399_),
    .Y(_400_)
);

FILL FILL_0__1755_ (
);

FILL FILL_0__1335_ (
);

FILL FILL_3__1595_ (
);

FILL FILL_3__1175_ (
);

FILL FILL_0__1564_ (
);

FILL FILL_0__1144_ (
);

FILL FILL_1__1725_ (
);

FILL FILL_1__1305_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_0_BUFX2_insert21 (
);

FILL FILL_0_BUFX2_insert22 (
);

FILL FILL_0_BUFX2_insert23 (
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_0_BUFX2_insert26 (
);

FILL FILL_0_BUFX2_insert27 (
);

FILL FILL_0_BUFX2_insert28 (
);

FILL FILL_0_BUFX2_insert29 (
);

FILL FILL_0__1793_ (
);

FILL FILL_0__1373_ (
);

FILL FILL_1__1534_ (
);

FILL FILL_1__1114_ (
);

NAND2X1 _1389_ (
    .A(AI[6]),
    .B(BI_3_bF$buf0),
    .Y(_493_)
);

FILL FILL_2__1603_ (
);

FILL FILL_0__1429_ (
);

FILL FILL_0__1009_ (
);

FILL FILL_2__958_ (
);

FILL FILL_0__1182_ (
);

NAND2X1 _1601_ (
    .A(AI[4]),
    .B(_705__bF$buf3),
    .Y(_695_)
);

INVX1 _932_ (
    .A(ABCmd_i_2_bF$buf2),
    .Y(_44_)
);

FILL FILL_1__1763_ (
);

FILL FILL_1__1343_ (
);

FILL FILL_3__1689_ (
);

FILL FILL_3__1269_ (
);

OAI21X1 _1198_ (
    .A(_283_),
    .B(_123_),
    .C(_248_),
    .Y(_304_)
);

FILL FILL_2__1412_ (
);

FILL FILL_0__1658_ (
);

FILL FILL_0__1238_ (
);

FILL FILL_1__1819_ (
);

OAI21X1 _1410_ (
    .A(_510_),
    .B(_513_),
    .C(_509_),
    .Y(_514_)
);

FILL FILL_1__1572_ (
);

FILL FILL_1__1152_ (
);

FILL FILL_3__1498_ (
);

FILL FILL_3__1078_ (
);

BUFX2 BUFX2_insert30 (
    .A(BI[4]),
    .Y(BI_4_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .A(BI[4]),
    .Y(BI_4_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .A(BI[4]),
    .Y(BI_4_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .A(BI[4]),
    .Y(BI_4_bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .A(BI[1]),
    .Y(BI_1_bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .A(BI[1]),
    .Y(BI_1_bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .A(BI[1]),
    .Y(BI_1_bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .A(BI[1]),
    .Y(BI_1_bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf3)
);

BUFX2 BUFX2_insert39 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf2)
);

FILL FILL_2__1641_ (
);

FILL FILL_2__1221_ (
);

FILL FILL_0__1467_ (
);

FILL FILL_0__1047_ (
);

FILL FILL_2__996_ (
);

FILL FILL_3__938_ (
);

FILL FILL_3__1710_ (
);

FILL FILL_1__1208_ (
);

NAND3X1 _970_ (
    .A(_75_),
    .B(_69_),
    .C(_72_),
    .Y(_76_)
);

FILL FILL_1__1381_ (
);

FILL FILL_2__1450_ (
);

FILL FILL_2__1030_ (
);

FILL FILL_0__1696_ (
);

FILL FILL_0__1276_ (
);

FILL FILL_1__1437_ (
);

FILL FILL_1__1017_ (
);

FILL FILL_1__1190_ (
);

FILL FILL_3_CLKBUF1_insert11 (
);

FILL FILL_3_CLKBUF1_insert12 (
);

FILL FILL_2__1506_ (
);

FILL FILL_0__1085_ (
);

INVX1 _1504_ (
    .A(_605_),
    .Y(_606_)
);

FILL FILL_3__976_ (
);

FILL FILL_1__1666_ (
);

FILL FILL_1__1246_ (
);

FILL FILL_2__1735_ (
);

FILL FILL_2__1315_ (
);

FILL FILL_3__1804_ (
);

OAI21X1 _1733_ (
    .A(_745_),
    .B(_744_),
    .C(_741_),
    .Y(_746_)
);

AND2X2 _1313_ (
    .A(AI[6]),
    .B(BI_3_bF$buf1),
    .Y(_418_)
);

FILL FILL_1__1475_ (
);

FILL FILL_1__1055_ (
);

FILL FILL_2__1544_ (
);

FILL FILL_2__1124_ (
);

FILL FILL_2__899_ (
);

OAI22X1 _1542_ (
    .A(_592_),
    .B(_167_),
    .C(_423_),
    .D(_597_),
    .Y(_643_)
);

NAND3X1 _1122_ (
    .A(_218_),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

FILL FILL_1__904_ (
);

FILL FILL_1__1284_ (
);

FILL FILL_2__1773_ (
);

FILL FILL_2__1353_ (
);

FILL FILL_0__1599_ (
);

FILL FILL_0__1179_ (
);

FILL FILL_0__926_ (
);

FILL FILL_3__1422_ (
);

INVX1 _929_ (
    .A(ABCmd_i[1]),
    .Y(_42_)
);

OR2X2 _1771_ (
    .A(_761_),
    .B(_844_),
    .Y(_782_)
);

OAI21X1 _1351_ (
    .A(_367_),
    .B(_455_),
    .C(_361_),
    .Y(_456_)
);

FILL FILL_1__1093_ (
);

FILL FILL_0__1811_ (
);

FILL FILL_2__1409_ (
);

FILL FILL_2__920_ (
);

FILL FILL_2__1582_ (
);

FILL FILL_2__1162_ (
);

BUFX2 _1827_ (
    .A(_887_),
    .Y(Done_o)
);

OR2X2 _1407_ (
    .A(_504_),
    .B(_498_),
    .Y(_511_)
);

FILL FILL_3__1651_ (
);

FILL FILL_1__1569_ (
);

FILL FILL_1__1149_ (
);

AOI21X1 _1580_ (
    .A(_677_),
    .B(_679_),
    .C(_712_),
    .Y(_680_)
);

NAND3X1 _1160_ (
    .A(_178_),
    .B(_243_),
    .C(_244_),
    .Y(_266_)
);

FILL FILL_1__942_ (
);

FILL FILL_2__1638_ (
);

FILL FILL_2__1218_ (
);

FILL FILL_0__1200_ (
);

FILL FILL_2__1391_ (
);

FILL FILL_3__1707_ (
);

INVX1 _1636_ (
    .A(ABCmd_i_2_bF$buf0),
    .Y(_824_)
);

AND2X2 _1216_ (
    .A(_318_),
    .B(_317_),
    .Y(_322_)
);

FILL FILL_0__964_ (
);

FILL FILL_3__1040_ (
);

INVX1 _967_ (
    .A(BI_0_bF$buf2),
    .Y(_73_)
);

FILL FILL_1__1798_ (
);

FILL FILL_1__1378_ (
);

FILL FILL_2__1447_ (
);

FILL FILL_2__1027_ (
);

FILL FILL_3__900_ (
);

FILL FILL_3__1516_ (
);

OAI22X1 _1445_ (
    .A(_493_),
    .B(_494_),
    .C(_492_),
    .D(_495_),
    .Y(_548_)
);

NAND2X1 _1025_ (
    .A(BI_0_bF$buf0),
    .B(AI[6]),
    .Y(_131_)
);

FILL FILL_1__1187_ (
);

FILL FILL_1__980_ (
);

FILL FILL_2__1676_ (
);

FILL FILL_2__1256_ (
);

FILL FILL_3__1325_ (
);

NAND2X1 _1674_ (
    .A(_860_),
    .B(_848_),
    .Y(_861_)
);

NAND3X1 _1254_ (
    .A(_359_),
    .B(_358_),
    .C(_357_),
    .Y(_360_)
);

FILL FILL_0__1714_ (
);

FILL FILL_2__1485_ (
);

FILL FILL_2__1065_ (
);

FILL FILL_3__1554_ (
);

NAND2X1 _1483_ (
    .A(ACC[3]),
    .B(_54_),
    .Y(_586_)
);

OAI21X1 _1063_ (
    .A(_84_),
    .B(_150_),
    .C(_111_),
    .Y(_169_)
);

FILL FILL_0__1523_ (
);

FILL FILL_0__1103_ (
);

FILL FILL_2__1294_ (
);

OAI21X1 _1539_ (
    .A(_167_),
    .B(_557_),
    .C(_596_),
    .Y(_640_)
);

NAND3X1 _1119_ (
    .A(_219_),
    .B(_224_),
    .C(_222_),
    .Y(_225_)
);

FILL FILL_3__1783_ (
);

NAND2X1 _1292_ (
    .A(_375_),
    .B(_371_),
    .Y(_397_)
);

FILL FILL_0__1752_ (
);

FILL FILL_0__1332_ (
);

FILL FILL_3__1419_ (
);

AOI21X1 _1768_ (
    .A(_719_),
    .B(_875_),
    .C(_778_),
    .Y(_779_)
);

NAND3X1 _1348_ (
    .A(_401_),
    .B(_452_),
    .C(_451_),
    .Y(_453_)
);

FILL FILL_3__1172_ (
);

FILL FILL_0__1808_ (
);

FILL FILL_2__917_ (
);

FILL FILL_2__1579_ (
);

FILL FILL_0__1561_ (
);

FILL FILL_0__1141_ (
);

FILL FILL_2__1159_ (
);

FILL FILL_1__1722_ (
);

FILL FILL_1__1302_ (
);

OAI21X1 _1577_ (
    .A(_676_),
    .B(_675_),
    .C(ABCmd_i[7]),
    .Y(_677_)
);

OAI21X1 _1157_ (
    .A(_174_),
    .B(_173_),
    .C(_171_),
    .Y(_263_)
);

FILL FILL_1__939_ (
);

FILL FILL_0__1790_ (
);

FILL FILL_2__1388_ (
);

FILL FILL_0__1370_ (
);

FILL FILL_1__1531_ (
);

FILL FILL_1__1111_ (
);

FILL FILL_3__1037_ (
);

NAND2X1 _1386_ (
    .A(_489_),
    .B(_486_),
    .Y(_490_)
);

FILL FILL_2__1600_ (
);

FILL FILL_0__1426_ (
);

FILL FILL_0__1006_ (
);

FILL FILL_2__955_ (
);

FILL FILL_2__1197_ (
);

FILL FILL_1__1760_ (
);

FILL FILL_1__1340_ (
);

FILL FILL_3__1686_ (
);

FILL FILL_3__1266_ (
);

NAND3X1 _1195_ (
    .A(_298_),
    .B(_289_),
    .C(_300_),
    .Y(_301_)
);

FILL FILL_1__977_ (
);

FILL FILL_0__1655_ (
);

FILL FILL_0__1235_ (
);

FILL FILL_1__1816_ (
);

FILL FILL_0__999_ (
);

FILL FILL_3__1495_ (
);

FILL FILL_3__1075_ (
);

FILL FILL_0__1464_ (
);

FILL FILL_0__1044_ (
);

FILL FILL_2__993_ (
);

FILL FILL_1__1205_ (
);

FILL FILL94050x35250 (
);

FILL FILL_0__1693_ (
);

FILL FILL_0__1273_ (
);

FILL FILL_1__1434_ (
);

FILL FILL_1__1014_ (
);

AOI21X1 _1289_ (
    .A(_392_),
    .B(_176_),
    .C(_390_),
    .Y(_394_)
);

FILL FILL_2__1503_ (
);

FILL FILL_0__1749_ (
);

FILL FILL_0__1329_ (
);

FILL FILL_0__1082_ (
);

NAND2X1 _1501_ (
    .A(_602_),
    .B(_600_),
    .Y(_603_)
);

FILL FILL_3__973_ (
);

FILL FILL_1__1663_ (
);

FILL FILL_1__1243_ (
);

FILL FILL_3__1169_ (
);

OAI21X1 _1098_ (
    .A(_83_),
    .B(_149_),
    .C(_198_),
    .Y(_204_)
);

FILL FILL_2__1732_ (
);

FILL FILL_2__1312_ (
);

FILL FILL_0__1558_ (
);

FILL FILL_0__1138_ (
);

FILL FILL94050x7950 (
);

FILL FILL_3__1801_ (
);

FILL FILL_1__1719_ (
);

NAND2X1 _1730_ (
    .A(AI[4]),
    .B(_742_),
    .Y(_743_)
);

FILL FILL94350x74250 (
);

NAND2X1 _1310_ (
    .A(AI[4]),
    .B(BI[5]),
    .Y(_415_)
);

FILL FILL_1__1472_ (
);

FILL FILL_1__1052_ (
);

FILL FILL_3__1398_ (
);

FILL FILL_2__1541_ (
);

FILL FILL_2__1121_ (
);

FILL FILL_0__1787_ (
);

FILL FILL_0__1367_ (
);

FILL FILL_2__896_ (
);

FILL FILL_1__1528_ (
);

FILL FILL_1__1108_ (
);

FILL FILL_1__901_ (
);

FILL FILL_1__1281_ (
);

FILL FILL_2__1770_ (
);

FILL FILL_2__1350_ (
);

FILL FILL_0__1596_ (
);

FILL FILL_0__1176_ (
);

FILL FILL_0__923_ (
);

INVX1 _926_ (
    .A(ABCmd_i[0]),
    .Y(_40_)
);

FILL FILL_1__1757_ (
);

FILL FILL_1__1337_ (
);

FILL FILL_1__1090_ (
);

FILL FILL_2__1826_ (
);

FILL FILL_2__1406_ (
);

BUFX2 _1824_ (
    .A(_886_[6]),
    .Y(ACC_o[6])
);

NAND3X1 _1404_ (
    .A(_502_),
    .B(_507_),
    .C(_479_),
    .Y(_508_)
);

FILL FILL_1__1566_ (
);

FILL FILL_1__1146_ (
);

FILL FILL_2__1215_ (
);

FILL FILL_3__1704_ (
);

DFFSR _1633_ (
    .D(_888_[0]),
    .S(_0__bF$buf1),
    .R(vdd),
    .CLK(clk_bF$buf2),
    .Q(state[0])
);

NAND2X1 _1213_ (
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

FILL FILL_0__961_ (
);

NAND2X1 _964_ (
    .A(BI_1_bF$buf1),
    .B(AI[3]),
    .Y(_70_)
);

FILL FILL_1__1795_ (
);

FILL FILL_1__1375_ (
);

FILL FILL_2__1444_ (
);

FILL FILL_2__1024_ (
);

NAND2X1 _1442_ (
    .A(AI[4]),
    .B(BI[7]),
    .Y(_545_)
);

NAND2X1 _1022_ (
    .A(_90_),
    .B(_127_),
    .Y(_128_)
);

FILL FILL_1__1184_ (
);

FILL FILL_2__1673_ (
);

FILL FILL_2__1253_ (
);

FILL FILL_0__1499_ (
);

FILL FILL_0__1079_ (
);

FILL FILL_3__1322_ (
);

INVX1 _1671_ (
    .A(_857_),
    .Y(_858_)
);

AND2X2 _1251_ (
    .A(_321_),
    .B(_324_),
    .Y(_357_)
);

FILL FILL_0__1711_ (
);

FILL FILL_2__1729_ (
);

FILL FILL_2__1309_ (
);

FILL FILL_2__1482_ (
);

FILL FILL_2__1062_ (
);

OAI21X1 _1727_ (
    .A(_738_),
    .B(_734_),
    .C(_740_),
    .Y(HC)
);

NOR2X1 _1307_ (
    .A(_344_),
    .B(_339_),
    .Y(_412_)
);

FILL FILL_3__1551_ (
);

FILL FILL_1__1469_ (
);

FILL FILL_1__1049_ (
);

NAND2X1 _1480_ (
    .A(_289_),
    .B(_300_),
    .Y(_583_)
);

NAND3X1 _1060_ (
    .A(_164_),
    .B(_165_),
    .C(_163_),
    .Y(_166_)
);

FILL FILL_2__1538_ (
);

FILL FILL_0__1520_ (
);

FILL FILL_2__1118_ (
);

FILL FILL_0__1100_ (
);

FILL FILL_2__1291_ (
);

NAND2X1 _1536_ (
    .A(_622_),
    .B(_624_),
    .Y(_637_)
);

OAI21X1 _1116_ (
    .A(_167_),
    .B(_113_),
    .C(_221_),
    .Y(_222_)
);

FILL FILL_3__1780_ (
);

FILL FILL_1__1698_ (
);

FILL FILL_1__1278_ (
);

FILL FILL_2__1767_ (
);

FILL FILL_2__1347_ (
);

FILL FILL_3__1416_ (
);

FILL FILL94350x62550 (
);

OAI21X1 _1765_ (
    .A(_772_),
    .B(_774_),
    .C(_775_),
    .Y(_776_)
);

NAND3X1 _1345_ (
    .A(_402_),
    .B(_442_),
    .C(_449_),
    .Y(_450_)
);

FILL FILL_1__1087_ (
);

FILL FILL_0__1805_ (
);

FILL FILL_2__914_ (
);

FILL FILL_2__1576_ (
);

FILL FILL_2__1156_ (
);

FILL FILL_3__1225_ (
);

NAND2X1 _1574_ (
    .A(_309_),
    .B(_393_),
    .Y(_674_)
);

NAND3X1 _1154_ (
    .A(_120_),
    .B(_100_),
    .C(_104_),
    .Y(_260_)
);

FILL FILL_1__936_ (
);

FILL FILL_2__1385_ (
);

FILL FILL_0__958_ (
);

FILL FILL_3__1454_ (
);

AND2X2 _1383_ (
    .A(_483_),
    .B(_482_),
    .Y(_487_)
);

FILL FILL_0__1423_ (
);

FILL FILL_0__1003_ (
);

FILL FILL_2__952_ (
);

FILL FILL_2__1194_ (
);

OAI21X1 _1439_ (
    .A(_480_),
    .B(_488_),
    .C(_484_),
    .Y(_542_)
);

AOI21X1 _1019_ (
    .A(_104_),
    .B(_116_),
    .C(_118_),
    .Y(_125_)
);

FILL FILL_3__1683_ (
);

INVX1 _1192_ (
    .A(_297_),
    .Y(_298_)
);

FILL FILL_1__974_ (
);

FILL FILL_0__1652_ (
);

FILL FILL_0__1232_ (
);

FILL FILL_1__1813_ (
);

FILL FILL_3__1739_ (
);

FILL FILL_3__1319_ (
);

OAI21X1 _1668_ (
    .A(_851_),
    .B(_854_),
    .C(_849_),
    .Y(_855_)
);

AOI21X1 _1248_ (
    .A(_342_),
    .B(_345_),
    .C(_338_),
    .Y(_354_)
);

FILL FILL_0__996_ (
);

FILL FILL_3__1072_ (
);

NAND2X1 _999_ (
    .A(AI[0]),
    .B(BI[5]),
    .Y(_105_)
);

FILL FILL_0__1708_ (
);

FILL FILL_2__1479_ (
);

FILL FILL_0__1461_ (
);

FILL FILL_0__1041_ (
);

FILL FILL_2__1059_ (
);

FILL FILL_2__990_ (
);

FILL FILL_1__1202_ (
);

FILL FILL94350x39150 (
);

FILL FILL_3__1548_ (
);

FILL FILL_3__1128_ (
);

INVX1 _1477_ (
    .A(_577_),
    .Y(_580_)
);

OAI21X1 _1057_ (
    .A(_120_),
    .B(_119_),
    .C(_100_),
    .Y(_163_)
);

FILL FILL_0__1517_ (
);

FILL FILL_0__1690_ (
);

FILL FILL_0__1270_ (
);

FILL FILL_2__1288_ (
);

FILL FILL_1__1431_ (
);

FILL FILL_1__1011_ (
);

FILL FILL_3__1777_ (
);

NAND2X1 _1286_ (
    .A(_172_),
    .B(_175_),
    .Y(_391_)
);

FILL FILL_2__1500_ (
);

FILL FILL_0__1746_ (
);

FILL FILL_0__1326_ (
);

FILL FILL_1_BUFX2_insert30 (
);

FILL FILL_1_BUFX2_insert31 (
);

FILL FILL_1_BUFX2_insert32 (
);

FILL FILL_1_BUFX2_insert33 (
);

FILL FILL_1_BUFX2_insert34 (
);

FILL FILL_1_BUFX2_insert35 (
);

FILL FILL_1_BUFX2_insert36 (
);

FILL FILL_1_BUFX2_insert37 (
);

FILL FILL_1_BUFX2_insert38 (
);

FILL FILL_1_BUFX2_insert39 (
);

FILL FILL_0_CLKBUF1_insert10 (
);

FILL FILL_0_CLKBUF1_insert11 (
);

FILL FILL_0_CLKBUF1_insert12 (
);

FILL FILL_2__1097_ (
);

FILL FILL_3__970_ (
);

FILL FILL_1__1660_ (
);

FILL FILL_1__1240_ (
);

FILL FILL_3__1166_ (
);

INVX1 _1095_ (
    .A(_200_),
    .Y(_201_)
);

FILL FILL_0__1555_ (
);

FILL FILL_0__1135_ (
);

FILL FILL_1__1716_ (
);

FILL FILL_0__899_ (
);

FILL FILL_3__1395_ (
);

FILL FILL_0__1784_ (
);

FILL FILL_0__1364_ (
);

FILL FILL_2__893_ (
);

FILL FILL94350x50850 (
);

FILL FILL_1__1525_ (
);

FILL FILL_1__1105_ (
);

FILL FILL_2__949_ (
);

FILL FILL_0__1593_ (
);

FILL FILL_0__1173_ (
);

FILL FILL_0__920_ (
);

AND2X2 _923_ (
    .A(_37_),
    .B(_38_),
    .Y(_39_)
);

FILL FILL_1__1754_ (
);

FILL FILL_1__1334_ (
);

INVX1 _1189_ (
    .A(BI[2]),
    .Y(_295_)
);

FILL FILL_2__1823_ (
);

FILL FILL_2__1403_ (
);

FILL FILL_0__1649_ (
);

FILL FILL_0__1229_ (
);

BUFX2 _1821_ (
    .A(_886_[3]),
    .Y(ACC_o[3])
);

INVX1 _1401_ (
    .A(_498_),
    .Y(_505_)
);

FILL FILL_1__1563_ (
);

FILL FILL_1__1143_ (
);

FILL FILL_3__1069_ (
);

FILL FILL_2__1212_ (
);

FILL FILL_0__1458_ (
);

FILL FILL_0__1038_ (
);

FILL FILL_2__987_ (
);

FILL FILL_3__929_ (
);

FILL FILL_3__1701_ (
);

DFFSR _1630_ (
    .D(_22_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(AI[5])
);

INVX1 _1210_ (
    .A(_315_),
    .Y(_316_)
);

OAI21X1 _961_ (
    .A(_65_),
    .B(_66_),
    .C(_64_),
    .Y(_67_)
);

FILL FILL_1__1792_ (
);

FILL FILL_1__1372_ (
);

FILL FILL_3__1298_ (
);

FILL FILL_2__1441_ (
);

FILL FILL_2__1021_ (
);

FILL FILL_0__1687_ (
);

FILL FILL_0__1267_ (
);

FILL FILL_1__1428_ (
);

FILL FILL_1__1008_ (
);

FILL FILL_1__1181_ (
);

FILL FILL_2__1670_ (
);

FILL FILL_2__1250_ (
);

FILL FILL_0__1496_ (
);

FILL FILL_0__1076_ (
);

FILL FILL94350x27450 (
);

FILL FILL_1_BUFX2_insert0 (
);

FILL FILL_1_BUFX2_insert1 (
);

FILL FILL_1_BUFX2_insert2 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert4 (
);

FILL FILL_3__967_ (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1__1657_ (
);

FILL FILL_1__1237_ (
);

FILL FILL94050x85950 (
);

FILL FILL_2__1726_ (
);

FILL FILL_2__1306_ (
);

NAND2X1 _1724_ (
    .A(ABCmd_i[6]),
    .B(_737_),
    .Y(_738_)
);

OAI22X1 _1304_ (
    .A(_407_),
    .B(_408_),
    .C(_327_),
    .D(_335_),
    .Y(_409_)
);

FILL FILL_1__1466_ (
);

FILL FILL_1__1046_ (
);

FILL FILL_2__1535_ (
);

FILL FILL_2__1115_ (
);

FILL FILL_3__1604_ (
);

AOI22X1 _1533_ (
    .A(_589_),
    .B(_712_),
    .C(_628_),
    .D(_634_),
    .Y(_13_)
);

INVX1 _1113_ (
    .A(_218_),
    .Y(_219_)
);

FILL FILL_1__1695_ (
);

FILL FILL_1__1275_ (
);

FILL FILL_2__1764_ (
);

FILL FILL_2__1344_ (
);

FILL FILL_0__917_ (
);

OAI21X1 _1762_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[6]),
    .C(_825_),
    .Y(_773_)
);

OAI21X1 _1342_ (
    .A(_412_),
    .B(_354_),
    .C(_432_),
    .Y(_447_)
);

FILL FILL_1__1084_ (
);

FILL FILL_0__1802_ (
);

FILL FILL_2__911_ (
);

FILL FILL_2__1573_ (
);

FILL FILL_2__1153_ (
);

FILL FILL93450x4050 (
);

FILL FILL_0__1399_ (
);

BUFX2 _1818_ (
    .A(_886_[0]),
    .Y(ACC_o[0])
);

FILL FILL_3__1222_ (
);

FILL FILL_3_BUFX2_insert0 (
);

FILL FILL_3_BUFX2_insert1 (
);

FILL FILL_3_BUFX2_insert3 (
);

FILL FILL_3_BUFX2_insert4 (
);

FILL FILL_3_BUFX2_insert6 (
);

INVX1 _1571_ (
    .A(_668_),
    .Y(_671_)
);

NAND3X1 _1151_ (
    .A(_252_),
    .B(_253_),
    .C(_254_),
    .Y(_257_)
);

FILL FILL_1__933_ (
);

FILL FILL_2__1209_ (
);

FILL FILL_2__1382_ (
);

DFFSR _1627_ (
    .D(_19_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(AI[2])
);

NAND2X1 _1207_ (
    .A(_226_),
    .B(_233_),
    .Y(_313_)
);

FILL FILL_0__955_ (
);

FILL FILL_3__1451_ (
);

OR2X2 _958_ (
    .A(_62_),
    .B(_63_),
    .Y(_64_)
);

FILL FILL_1__1789_ (
);

FILL FILL_1__1369_ (
);

NAND2X1 _1380_ (
    .A(_482_),
    .B(_483_),
    .Y(_484_)
);

FILL FILL_2__1438_ (
);

FILL FILL_0__1420_ (
);

FILL FILL_0__1000_ (
);

FILL FILL_2__1018_ (
);

FILL FILL_2__1191_ (
);

INVX1 _1436_ (
    .A(AV),
    .Y(_539_)
);

NAND3X1 _1016_ (
    .A(_117_),
    .B(_121_),
    .C(_88_),
    .Y(_122_)
);

FILL FILL_3__1680_ (
);

FILL FILL_1__1598_ (
);

FILL FILL_1__1178_ (
);

FILL FILL_1__971_ (
);

FILL FILL_2__1667_ (
);

FILL FILL_2__1247_ (
);

FILL FILL_1__1810_ (
);

FILL FILL_3__1736_ (
);

FILL FILL_3__1316_ (
);

INVX1 _1665_ (
    .A(BI_1_bF$buf0),
    .Y(_852_)
);

NAND3X1 _1245_ (
    .A(_346_),
    .B(_350_),
    .C(_326_),
    .Y(_351_)
);

FILL FILL_0__993_ (
);

OAI21X1 _996_ (
    .A(_92_),
    .B(_98_),
    .C(_95_),
    .Y(_102_)
);

FILL FILL_0__1705_ (
);

FILL FILL_2__1476_ (
);

FILL FILL_2__1056_ (
);

FILL FILL_3__1545_ (
);

FILL FILL_3__1125_ (
);

NAND2X1 _1474_ (
    .A(_576_),
    .B(_573_),
    .Y(_577_)
);

NAND2X1 _1054_ (
    .A(_152_),
    .B(_155_),
    .Y(_160_)
);

FILL FILL_0__1514_ (
);

FILL FILL_2__1285_ (
);

FILL FILL_3__1354_ (
);

OAI21X1 _1283_ (
    .A(_386_),
    .B(_715_),
    .C(_387_),
    .Y(_388_)
);

FILL FILL_0__1743_ (
);

FILL FILL_0__1323_ (
);

FILL FILL_2__1094_ (
);

AOI22X1 _1759_ (
    .A(_829_),
    .B(BI[6]),
    .C(_769_),
    .D(_830_),
    .Y(_770_)
);

AOI21X1 _1339_ (
    .A(_357_),
    .B(_359_),
    .C(_443_),
    .Y(_444_)
);

FILL FILL_3__1583_ (
);

AND2X2 _1092_ (
    .A(BI_3_bF$buf3),
    .B(AI[4]),
    .Y(_198_)
);

FILL FILL_2__908_ (
);

FILL FILL_0__1552_ (
);

FILL FILL_0__1132_ (
);

FILL FILL_1__1713_ (
);

FILL FILL_3__1639_ (
);

FILL FILL_3__1219_ (
);

XOR2X1 _1568_ (
    .A(_666_),
    .B(_667_),
    .Y(_668_)
);

NAND3X1 _1148_ (
    .A(_68_),
    .B(_75_),
    .C(_72_),
    .Y(_254_)
);

FILL FILL_0__896_ (
);

AOI21X1 _899_ (
    .A(_703_),
    .B(_707_),
    .C(_887_),
    .Y(_708_)
);

FILL FILL_0__1608_ (
);

FILL FILL_2__1799_ (
);

FILL FILL_0__1781_ (
);

FILL FILL_0__1361_ (
);

FILL FILL_2__1379_ (
);

FILL FILL_2__890_ (
);

FILL FILL_1__1522_ (
);

FILL FILL_1__1102_ (
);

FILL FILL_3__1448_ (
);

FILL FILL_3__1028_ (
);

AND2X2 _1797_ (
    .A(_805_),
    .B(_803_),
    .Y(AZ)
);

INVX1 _1377_ (
    .A(_480_),
    .Y(_481_)
);

FILL FILL_0__1417_ (
);

FILL FILL_2__946_ (
);

FILL FILL_0__1590_ (
);

FILL FILL_2__1188_ (
);

FILL FILL_0__1170_ (
);

INVX1 _920_ (
    .A(_32__bF$buf3),
    .Y(_36_)
);

FILL FILL_1__1751_ (
);

FILL FILL_1__1331_ (
);

FILL FILL_3__1677_ (
);

OR2X2 _1186_ (
    .A(_291_),
    .B(_273_),
    .Y(_292_)
);

FILL FILL_1__968_ (
);

FILL FILL_2__1820_ (
);

FILL FILL_2__1400_ (
);

FILL FILL_0__1646_ (
);

FILL FILL_0__1226_ (
);

FILL FILL_1__1807_ (
);

FILL FILL_1__1560_ (
);

FILL FILL_1__1140_ (
);

FILL FILL_3__1066_ (
);

FILL FILL_0__1455_ (
);

FILL FILL_0__1035_ (
);

FILL FILL_2__984_ (
);

FILL FILL_3__926_ (
);

FILL FILL_3__1295_ (
);

FILL FILL_0__1684_ (
);

FILL FILL_0__1264_ (
);

FILL FILL_1__1425_ (
);

FILL FILL_1__1005_ (
);

FILL FILL_0__1493_ (
);

FILL FILL_0__1073_ (
);

FILL FILL_1__1654_ (
);

FILL FILL_1__1234_ (
);

NAND2X1 _1089_ (
    .A(BI[5]),
    .B(AI[2]),
    .Y(_195_)
);

FILL FILL94350x89850 (
);

FILL FILL_2__1723_ (
);

FILL FILL_2__1303_ (
);

FILL FILL_0__1549_ (
);

FILL FILL_0__1129_ (
);

NAND2X1 _1721_ (
    .A(_718_),
    .B(_877_),
    .Y(_735_)
);

NOR2X1 _1301_ (
    .A(_149_),
    .B(_167_),
    .Y(_406_)
);

FILL FILL_1__1463_ (
);

FILL FILL_1__1043_ (
);

FILL FILL_2__1532_ (
);

FILL FILL_2__1112_ (
);

FILL FILL_0__1778_ (
);

FILL FILL_0__1358_ (
);

FILL FILL_3__1601_ (
);

FILL FILL_1__1519_ (
);

NAND2X1 _1530_ (
    .A(ACC[4]),
    .B(_54_),
    .Y(_632_)
);

OAI21X1 _1110_ (
    .A(_194_),
    .B(_191_),
    .C(_211_),
    .Y(_216_)
);

FILL FILL_1__1692_ (
);

FILL FILL_1__1272_ (
);

FILL FILL_3__1198_ (
);

FILL FILL_2__1761_ (
);

FILL FILL_2__1341_ (
);

FILL FILL_0__1587_ (
);

FILL FILL_0__1167_ (
);

FILL FILL_0__914_ (
);

NOR2X1 _917_ (
    .A(LoadB_i),
    .B(_26_),
    .Y(_34_)
);

FILL FILL_1__1748_ (
);

FILL FILL_1__1328_ (
);

FILL FILL_1__1081_ (
);

FILL FILL_2__1817_ (
);

FILL FILL_2__1570_ (
);

FILL FILL_2__1150_ (
);

FILL FILL_0__1396_ (
);

NAND3X1 _1815_ (
    .A(_814_),
    .B(_815_),
    .C(_821_),
    .Y(_822_)
);

FILL FILL_1__1557_ (
);

FILL FILL_1__1137_ (
);

FILL FILL_1__930_ (
);

FILL FILL_2__1206_ (
);

DFFSR _1624_ (
    .D(_16_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf3),
    .Q(_886_[7])
);

AOI21X1 _1204_ (
    .A(_308_),
    .B(_309_),
    .C(_287_),
    .Y(_310_)
);

FILL FILL_0__952_ (
);

NAND2X1 _955_ (
    .A(_60_),
    .B(_59_),
    .Y(_61_)
);

FILL FILL_1__1786_ (
);

FILL FILL_1__1366_ (
);

FILL FILL_2__1435_ (
);

FILL FILL_2__1015_ (
);

FILL FILL_3__1504_ (
);

AOI22X1 _1433_ (
    .A(_534_),
    .B(_536_),
    .C(_530_),
    .D(_532_),
    .Y(_537_)
);

AOI21X1 _1013_ (
    .A(_99_),
    .B(_96_),
    .C(_89_),
    .Y(_119_)
);

FILL FILL_1__1595_ (
);

FILL FILL_1__1175_ (
);

FILL FILL_2__1664_ (
);

FILL FILL_2__1244_ (
);

FILL FILL_3__1733_ (
);

NAND2X1 _1662_ (
    .A(ABCmd_i[5]),
    .B(AI[2]),
    .Y(_849_)
);

NAND2X1 _1242_ (
    .A(_343_),
    .B(_341_),
    .Y(_348_)
);

FILL FILL_0__990_ (
);

OAI21X1 _993_ (
    .A(_92_),
    .B(_98_),
    .C(_94_),
    .Y(_99_)
);

FILL FILL_0__1702_ (
);

FILL FILL_2__1473_ (
);

FILL FILL_2__1053_ (
);

FILL FILL_0__1299_ (
);

OAI21X1 _1718_ (
    .A(_729_),
    .B(_731_),
    .C(_732_),
    .Y(_733_)
);

FILL FILL_3__1122_ (
);

AOI21X1 _1471_ (
    .A(_502_),
    .B(_507_),
    .C(_509_),
    .Y(_574_)
);

OAI21X1 _1051_ (
    .A(_139_),
    .B(_143_),
    .C(_156_),
    .Y(_157_)
);

FILL FILL_0__1511_ (
);

FILL FILL_2__1529_ (
);

FILL FILL_2__1109_ (
);

FILL FILL_2__1282_ (
);

INVX1 _1527_ (
    .A(_303_),
    .Y(_629_)
);

NAND3X1 _1107_ (
    .A(_212_),
    .B(_207_),
    .C(_180_),
    .Y(_213_)
);

FILL FILL_3__999_ (
);

FILL FILL_3__1351_ (
);

FILL FILL_1__1689_ (
);

FILL FILL_1__1269_ (
);

INVX1 _1280_ (
    .A(_886_[1]),
    .Y(_385_)
);

FILL FILL93150x82050 (
);

FILL FILL_0__1740_ (
);

FILL FILL_2__1758_ (
);

FILL FILL_0__1320_ (
);

FILL FILL_2__1338_ (
);

FILL FILL_2__1091_ (
);

FILL FILL_3__1827_ (
);

INVX1 _1756_ (
    .A(\u_ALU.AI7 ),
    .Y(_767_)
);

NAND3X1 _1336_ (
    .A(_438_),
    .B(_440_),
    .C(_439_),
    .Y(_441_)
);

FILL FILL_3__1580_ (
);

FILL FILL_1__1498_ (
);

FILL FILL_1__1078_ (
);

FILL FILL_2__905_ (
);

FILL FILL_2__1567_ (
);

FILL FILL_2__1147_ (
);

FILL FILL_1__1710_ (
);

FILL FILL_3__1636_ (
);

FILL FILL_3__1216_ (
);

NAND2X1 _1565_ (
    .A(_640_),
    .B(_664_),
    .Y(_665_)
);

OAI21X1 _1145_ (
    .A(_73_),
    .B(_149_),
    .C(_62_),
    .Y(_251_)
);

FILL FILL_0__893_ (
);

FILL FILL_1__927_ (
);

NAND2X1 _896_ (
    .A(_702_),
    .B(_704_),
    .Y(_705_)
);

FILL FILL_0__1605_ (
);

FILL FILL_2__1796_ (
);

FILL FILL_2__1376_ (
);

FILL FILL_0__949_ (
);

FILL FILL_3__1445_ (
);

FILL FILL_3__1025_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_2_BUFX2_insert21 (
);

FILL FILL_2_BUFX2_insert22 (
);

FILL FILL_2_BUFX2_insert23 (
);

FILL FILL_2_BUFX2_insert24 (
);

FILL FILL_2_BUFX2_insert25 (
);

FILL FILL_2_BUFX2_insert26 (
);

FILL FILL_2_BUFX2_insert27 (
);

FILL FILL_2_BUFX2_insert28 (
);

FILL FILL_2_BUFX2_insert29 (
);

NOR2X1 _1794_ (
    .A(_802_),
    .B(ACC[4]),
    .Y(_803_)
);

INVX1 _1374_ (
    .A(_477_),
    .Y(_478_)
);

FILL FILL_0__1414_ (
);

FILL FILL_2__943_ (
);

FILL FILL_2__1185_ (
);

FILL FILL_3__1254_ (
);

NAND3X1 _1183_ (
    .A(_59_),
    .B(_277_),
    .C(_288_),
    .Y(_289_)
);

FILL FILL_1__965_ (
);

FILL FILL_0__1643_ (
);

FILL FILL_0__1223_ (
);

FILL FILL_1__1804_ (
);

XOR2X1 _1659_ (
    .A(_846_),
    .B(_828_),
    .Y(ACC[0])
);

NAND2X1 _1239_ (
    .A(_343_),
    .B(_344_),
    .Y(_345_)
);

FILL FILL_0__987_ (
);

FILL FILL_3__1483_ (
);

FILL FILL_0__1452_ (
);

FILL FILL_0__1032_ (
);

FILL FILL_2__981_ (
);

FILL FILL_3__923_ (
);

FILL FILL_3__1119_ (
);

NAND3X1 _1468_ (
    .A(_542_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

OAI21X1 _1048_ (
    .A(_83_),
    .B(_109_),
    .C(_147_),
    .Y(_154_)
);

FILL FILL_0__1508_ (
);

FILL FILL_2__1699_ (
);

FILL FILL_0__1681_ (
);

FILL FILL_2__1279_ (
);

FILL FILL_0__1261_ (
);

FILL FILL_1__1422_ (
);

FILL FILL_1__1002_ (
);

FILL FILL_3__1768_ (
);

FILL FILL_3__1348_ (
);

OAI21X1 _1697_ (
    .A(AI[2]),
    .B(_882_),
    .C(_835_),
    .Y(_883_)
);

OAI21X1 _1277_ (
    .A(_381_),
    .B(_382_),
    .C(_380_),
    .Y(_383_)
);

FILL FILL_0__1737_ (
);

FILL FILL_0__1317_ (
);

FILL FILL_0__1490_ (
);

FILL FILL_2__1088_ (
);

FILL FILL_0__1070_ (
);

FILL FILL_1__1651_ (
);

FILL FILL_1__1231_ (
);

FILL FILL_3__1577_ (
);

OAI21X1 _1086_ (
    .A(_183_),
    .B(_189_),
    .C(_186_),
    .Y(_192_)
);

FILL FILL_2__1720_ (
);

FILL FILL_2__1300_ (
);

FILL FILL_0__1546_ (
);

FILL FILL_0__1126_ (
);

FILL FILL_1__1707_ (
);

FILL FILL_1__1460_ (
);

FILL FILL_1__1040_ (
);

FILL FILL94050x150 (
);

FILL FILL_0__1775_ (
);

FILL FILL_0__1355_ (
);

FILL FILL_1__1516_ (
);

FILL FILL_3__1195_ (
);

FILL FILL_0__1584_ (
);

FILL FILL_0__1164_ (
);

FILL FILL_0__911_ (
);

OAI21X1 _914_ (
    .A(_30_),
    .B(_708_),
    .C(_25_),
    .Y(_31_)
);

FILL FILL_1__1745_ (
);

FILL FILL_1__1325_ (
);

FILL FILL_2__1814_ (
);

FILL FILL_0__1393_ (
);

INVX1 _1812_ (
    .A(_817_),
    .Y(_819_)
);

FILL FILL_1__1554_ (
);

FILL FILL_1__1134_ (
);

FILL FILL_2__1203_ (
);

FILL FILL_0__1449_ (
);

FILL FILL_0__1029_ (
);

FILL FILL_2__978_ (
);

DFFSR _1621_ (
    .D(_13_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf1),
    .Q(_886_[4])
);

NAND3X1 _1201_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_307_)
);

INVX2 _952_ (
    .A(BI_3_bF$buf1),
    .Y(_58_)
);

FILL FILL_1__1783_ (
);

FILL FILL_1__1363_ (
);

FILL FILL_2__1432_ (
);

FILL FILL_2__1012_ (
);

FILL FILL_0__1678_ (
);

FILL FILL_0__1258_ (
);

FILL FILL_3__1501_ (
);

FILL FILL_1__1419_ (
);

OAI21X1 _1430_ (
    .A(_533_),
    .B(_298_),
    .C(ABCmd_i[7]),
    .Y(_534_)
);

AND2X2 _1010_ (
    .A(_115_),
    .B(_111_),
    .Y(_116_)
);

FILL FILL_1__1592_ (
);

FILL FILL_1__1172_ (
);

FILL FILL_3__1098_ (
);

FILL FILL_2__1661_ (
);

FILL FILL_2__1241_ (
);

FILL FILL_0__1487_ (
);

FILL FILL_0__1067_ (
);

FILL FILL_3__1730_ (
);

FILL FILL_1__1648_ (
);

FILL FILL_1__1228_ (
);

NAND3X1 _990_ (
    .A(_93_),
    .B(_95_),
    .C(_91_),
    .Y(_96_)
);

FILL FILL_2__1717_ (
);

FILL FILL_2__1470_ (
);

FILL FILL_2__1050_ (
);

FILL FILL_0__1296_ (
);

OAI21X1 _1715_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_3_bF$buf2),
    .C(_825_),
    .Y(_730_)
);

FILL FILL_1__1457_ (
);

FILL FILL_1__1037_ (
);

FILL FILL_2__1526_ (
);

FILL FILL_2__1106_ (
);

OAI21X1 _1524_ (
    .A(_625_),
    .B(_620_),
    .C(ABCmd_i[7]),
    .Y(_626_)
);

NAND3X1 _1104_ (
    .A(_181_),
    .B(_187_),
    .C(_190_),
    .Y(_210_)
);

FILL FILL_3__996_ (
);

FILL FILL_1__1686_ (
);

FILL FILL_1__1266_ (
);

FILL FILL_2__1755_ (
);

FILL FILL_2__1335_ (
);

FILL FILL_0__908_ (
);

FILL FILL_3__1404_ (
);

XOR2X1 _1753_ (
    .A(_753_),
    .B(_764_),
    .Y(_765_)
);

XOR2X1 _1333_ (
    .A(_410_),
    .B(_405_),
    .Y(_438_)
);

FILL FILL_1__1495_ (
);

FILL FILL_1__1075_ (
);

FILL FILL_2__902_ (
);

FILL FILL_2__1564_ (
);

FILL FILL_2__1144_ (
);

AOI21X1 _1809_ (
    .A(_792_),
    .B(_844_),
    .C(_794_),
    .Y(_816_)
);

OAI21X1 _1562_ (
    .A(_639_),
    .B(_646_),
    .C(_661_),
    .Y(_662_)
);

INVX1 _1142_ (
    .A(_61_),
    .Y(_248_)
);

FILL FILL_0__890_ (
);

FILL FILL_1__924_ (
);

INVX1 _893_ (
    .A(state[0]),
    .Y(_702_)
);

FILL FILL_0__1602_ (
);

FILL FILL_2__1793_ (
);

FILL FILL_2__1373_ (
);

FILL FILL_0__1199_ (
);

DFFSR _1618_ (
    .D(_10_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf1),
    .Q(_886_[1])
);

FILL FILL_0__946_ (
);

FILL FILL_3__1022_ (
);

OAI21X1 _949_ (
    .A(_54_),
    .B(_32__bF$buf3),
    .C(_55_),
    .Y(_8_)
);

NAND2X1 _1791_ (
    .A(_800_),
    .B(_797_),
    .Y(AN)
);

INVX1 _1371_ (
    .A(_474_),
    .Y(_475_)
);

FILL FILL_2__1429_ (
);

FILL FILL_0__1411_ (
);

FILL FILL_2__1009_ (
);

FILL FILL_2__940_ (
);

FILL FILL_2__1182_ (
);

NOR2X1 _1427_ (
    .A(ABCmd_i[7]),
    .B(AZ),
    .Y(_531_)
);

INVX1 _1007_ (
    .A(AI[1]),
    .Y(_113_)
);

FILL FILL_3__899_ (
);

FILL FILL_3__1251_ (
);

FILL FILL_1__1589_ (
);

FILL FILL_1__1169_ (
);

AOI21X1 _1180_ (
    .A(_175_),
    .B(_172_),
    .C(_124_),
    .Y(_286_)
);

FILL FILL_1__962_ (
);

FILL FILL_2__1658_ (
);

FILL FILL_0__1640_ (
);

FILL FILL_2__1238_ (
);

FILL FILL_0__1220_ (
);

FILL FILL_1__1801_ (
);

FILL FILL_3__1727_ (
);

NOR2X1 _1656_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(_825_),
    .Y(_844_)
);

NAND2X1 _1236_ (
    .A(_341_),
    .B(_339_),
    .Y(_342_)
);

FILL FILL_0__984_ (
);

FILL FILL_3__1480_ (
);

INVX1 _987_ (
    .A(_92_),
    .Y(_93_)
);

FILL FILL_1__1398_ (
);

FILL FILL_2__1467_ (
);

FILL FILL_2__1047_ (
);

FILL FILL_3__920_ (
);

FILL FILL_3__1116_ (
);

FILL FILL_3_CLKBUF1_insert8 (
);

FILL FILL_3_CLKBUF1_insert9 (
);

NAND3X1 _1465_ (
    .A(_543_),
    .B(_567_),
    .C(_564_),
    .Y(_568_)
);

OAI21X1 _1045_ (
    .A(_58_),
    .B(_149_),
    .C(_150_),
    .Y(_151_)
);

FILL FILL93150x35250 (
);

FILL FILL_0__1505_ (
);

FILL FILL_2__1696_ (
);

FILL FILL_2__1276_ (
);

FILL FILL_3__1765_ (
);

FILL FILL_3__1345_ (
);

AOI22X1 _1694_ (
    .A(_829_),
    .B(BI[2]),
    .C(_879_),
    .D(_830_),
    .Y(_880_)
);

OAI21X1 _1274_ (
    .A(_54_),
    .B(_377_),
    .C(_379_),
    .Y(_380_)
);

FILL FILL_0__1734_ (
);

FILL FILL_0__1314_ (
);

FILL FILL_2__1085_ (
);

FILL FILL_3__1574_ (
);

FILL FILL_3__1154_ (
);

NOR2X1 _1083_ (
    .A(_131_),
    .B(_188_),
    .Y(_189_)
);

FILL FILL_0__1543_ (
);

FILL FILL_0__1123_ (
);

FILL FILL_1__1704_ (
);

INVX1 _1559_ (
    .A(_658_),
    .Y(_659_)
);

NAND3X1 _1139_ (
    .A(_177_),
    .B(_243_),
    .C(_244_),
    .Y(_245_)
);

FILL FILL_3__1383_ (
);

FILL FILL93450x74250 (
);

FILL FILL_0__1772_ (
);

FILL FILL_0__1352_ (
);

FILL FILL_1__1513_ (
);

FILL FILL_3__1019_ (
);

FILL FILL93450x7950 (
);

NAND2X1 _1788_ (
    .A(_784_),
    .B(_766_),
    .Y(_798_)
);

NOR2X1 _1368_ (
    .A(_471_),
    .B(_470_),
    .Y(_472_)
);

FILL FILL_0__1408_ (
);

FILL FILL_2__937_ (
);

FILL FILL_0__1581_ (
);

FILL FILL_2__1599_ (
);

FILL FILL_2__1179_ (
);

FILL FILL_0__1161_ (
);

AOI22X1 _911_ (
    .A(_712_),
    .B(_713_),
    .C(_28_),
    .D(_711_),
    .Y(_29_)
);

FILL FILL_1__1742_ (
);

FILL FILL_1__1322_ (
);

FILL FILL_3__1668_ (
);

FILL FILL_3__1248_ (
);

NAND2X1 _1597_ (
    .A(AI[2]),
    .B(_705__bF$buf3),
    .Y(_693_)
);

AOI22X1 _1177_ (
    .A(_80_),
    .B(_269_),
    .C(_259_),
    .D(_260_),
    .Y(_283_)
);

FILL FILL_1__959_ (
);

FILL FILL_2__1811_ (
);

FILL FILL_0__1637_ (
);

FILL FILL_0__1217_ (
);

FILL FILL_0__1390_ (
);

FILL FILL_1__1551_ (
);

FILL FILL_1__1131_ (
);

FILL FILL_3__1477_ (
);

FILL FILL_2__1200_ (
);

FILL FILL_0__1446_ (
);

FILL FILL_0__1026_ (
);

FILL FILL_2__975_ (
);

FILL FILL_3__917_ (
);

FILL FILL_1__1607_ (
);

FILL FILL_1__1780_ (
);

FILL FILL_1__1360_ (
);

FILL FILL_1__997_ (
);

FILL FILL_0__1675_ (
);

FILL FILL_0__1255_ (
);

FILL FILL_1__1416_ (
);

FILL FILL_3__1095_ (
);

FILL FILL_0__1484_ (
);

FILL FILL_0__1064_ (
);

FILL FILL_3__955_ (
);

FILL FILL_1__1645_ (
);

FILL FILL_1__1225_ (
);

FILL FILL_2__1714_ (
);

FILL FILL_0__1293_ (
);

AOI22X1 _1712_ (
    .A(_829_),
    .B(BI_3_bF$buf2),
    .C(_726_),
    .D(_830_),
    .Y(_727_)
);

FILL FILL_1__1454_ (
);

FILL FILL_1__1034_ (
);

FILL FILL_2__1523_ (
);

FILL FILL_2__1103_ (
);

FILL FILL_0__1769_ (
);

FILL FILL_0__1349_ (
);

AOI21X1 _1521_ (
    .A(_573_),
    .B(_618_),
    .C(_474_),
    .Y(_623_)
);

OAI21X1 _1101_ (
    .A(_194_),
    .B(_191_),
    .C(_206_),
    .Y(_207_)
);

FILL FILL_1__1683_ (
);

FILL FILL_1__1263_ (
);

FILL FILL_2__1752_ (
);

FILL FILL_2__1332_ (
);

FILL FILL_0__1578_ (
);

FILL FILL_0__1158_ (
);

FILL FILL_0__905_ (
);

FILL FILL_3__1401_ (
);

INVX1 _908_ (
    .A(LoadCmd_i),
    .Y(_26_)
);

FILL FILL_1__1739_ (
);

FILL FILL_1__1319_ (
);

OAI21X1 _1750_ (
    .A(_844_),
    .B(_761_),
    .C(_759_),
    .Y(_762_)
);

OAI21X1 _1330_ (
    .A(_338_),
    .B(_434_),
    .C(_348_),
    .Y(_435_)
);

FILL FILL_1__1492_ (
);

FILL FILL_1__1072_ (
);

FILL FILL_2__1808_ (
);

FILL FILL_2__1561_ (
);

FILL FILL_2__1141_ (
);

FILL FILL_0__1387_ (
);

XOR2X1 _1806_ (
    .A(_813_),
    .B(_810_),
    .Y(_814_)
);

FILL FILL_1__1548_ (
);

FILL FILL_1__1128_ (
);

FILL FILL_1__921_ (
);

NOR2X1 _890_ (
    .A(state[0]),
    .B(_699_),
    .Y(_700_)
);

FILL FILL_2__1790_ (
);

FILL FILL_2__1370_ (
);

FILL FILL_0__1196_ (
);

DFFSR _1615_ (
    .D(_7_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf1),
    .Q(BI[6])
);

FILL FILL_0__943_ (
);

OAI21X1 _946_ (
    .A(_52_),
    .B(_32__bF$buf1),
    .C(_53_),
    .Y(_7_)
);

FILL FILL_1__1777_ (
);

FILL FILL_1__1357_ (
);

FILL FILL_2__1426_ (
);

FILL FILL_2__1006_ (
);

INVX1 _1424_ (
    .A(_524_),
    .Y(_528_)
);

OAI21X1 _1004_ (
    .A(_58_),
    .B(_109_),
    .C(_82_),
    .Y(_110_)
);

FILL FILL_3__896_ (
);

FILL FILL_1__1586_ (
);

FILL FILL_1__1166_ (
);

FILL FILL_2__1655_ (
);

FILL FILL_2__1235_ (
);

FILL FILL_3__1304_ (
);

OAI21X1 _1653_ (
    .A(_834_),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

AOI21X1 _1233_ (
    .A(_184_),
    .B(_186_),
    .C(_189_),
    .Y(_339_)
);

FILL FILL_0__981_ (
);

AND2X2 _984_ (
    .A(BI_0_bF$buf1),
    .B(AI_5_bF$buf3),
    .Y(_90_)
);

FILL FILL_1__1395_ (
);

FILL FILL_2__1464_ (
);

FILL FILL_2__1044_ (
);

NAND2X1 _1709_ (
    .A(ABCmd_i[5]),
    .B(AI[4]),
    .Y(_724_)
);

FILL FILL_3__1533_ (
);

OAI21X1 _1462_ (
    .A(_490_),
    .B(_501_),
    .C(_506_),
    .Y(_565_)
);

NAND2X1 _1042_ (
    .A(_146_),
    .B(_147_),
    .Y(_148_)
);

FILL FILL_0__1502_ (
);

FILL FILL_2__1693_ (
);

FILL FILL_2__1273_ (
);

FILL FILL_0__1099_ (
);

AOI21X1 _1518_ (
    .A(_619_),
    .B(_617_),
    .C(_614_),
    .Y(_620_)
);

FILL FILL_3__1762_ (
);

OAI21X1 _1691_ (
    .A(_876_),
    .B(_871_),
    .C(_872_),
    .Y(_877_)
);

XOR2X1 _1271_ (
    .A(_311_),
    .B(_376_),
    .Y(_377_)
);

FILL FILL_2__1749_ (
);

FILL FILL_0__1731_ (
);

FILL FILL_0__1311_ (
);

FILL FILL_2__1329_ (
);

FILL FILL_2__1082_ (
);

FILL FILL_3__1818_ (
);

OAI21X1 _1747_ (
    .A(_758_),
    .B(_757_),
    .C(_754_),
    .Y(_759_)
);

NAND2X1 _1327_ (
    .A(_431_),
    .B(_427_),
    .Y(_432_)
);

FILL FILL_3__1151_ (
);

FILL FILL_1__1489_ (
);

FILL FILL_1__1069_ (
);

INVX1 _1080_ (
    .A(_185_),
    .Y(_186_)
);

FILL FILL_2__1558_ (
);

FILL FILL_0__1540_ (
);

FILL FILL_0__1120_ (
);

FILL FILL_2__1138_ (
);

FILL FILL_3_BUFX2_insert30 (
);

FILL FILL_3_BUFX2_insert32 (
);

FILL FILL_3_BUFX2_insert33 (
);

FILL FILL_3_BUFX2_insert35 (
);

FILL FILL_3_BUFX2_insert37 (
);

FILL FILL_3_BUFX2_insert38 (
);

FILL FILL_1__1701_ (
);

AOI22X1 _1556_ (
    .A(_635_),
    .B(_712_),
    .C(_651_),
    .D(_656_),
    .Y(_14_)
);

OAI21X1 _1136_ (
    .A(_241_),
    .B(_237_),
    .C(_178_),
    .Y(_242_)
);

FILL FILL_1__918_ (
);

FILL FILL_3__1380_ (
);

FILL FILL93750x78150 (
);

FILL FILL_1__1298_ (
);

FILL FILL_2__1787_ (
);

FILL FILL_2__1367_ (
);

FILL FILL_1__1510_ (
);

FILL FILL_3__1016_ (
);

OAI21X1 _1785_ (
    .A(_844_),
    .B(_794_),
    .C(_792_),
    .Y(_795_)
);

OAI21X1 _1365_ (
    .A(state[0]),
    .B(_699_),
    .C(_886_[2]),
    .Y(_469_)
);

FILL FILL_0__1825_ (
);

FILL FILL_0__1405_ (
);

FILL FILL_2__934_ (
);

FILL FILL_2__1596_ (
);

FILL FILL_2__1176_ (
);

FILL FILL_3__1665_ (
);

FILL FILL_3__1245_ (
);

OAI21X1 _1594_ (
    .A(_40_),
    .B(_705__bF$buf2),
    .C(_691_),
    .Y(_17_)
);

OAI21X1 _1174_ (
    .A(_255_),
    .B(_87_),
    .C(_86_),
    .Y(_280_)
);

FILL FILL_1__956_ (
);

FILL FILL_0__1214_ (
);

FILL FILL_0__978_ (
);

FILL FILL_3__1474_ (
);

FILL FILL_3__1054_ (
);

FILL FILL_0__1443_ (
);

FILL FILL_0__1023_ (
);

FILL FILL_2__972_ (
);

FILL FILL_1__1604_ (
);

INVX1 _1459_ (
    .A(_561_),
    .Y(_562_)
);

INVX1 _1039_ (
    .A(_144_),
    .Y(_145_)
);

FILL FILL_3__1283_ (
);

FILL FILL_1__994_ (
);

FILL FILL_0__1672_ (
);

FILL FILL_0__1252_ (
);

FILL FILL_1__1413_ (
);

FILL FILL_3__1759_ (
);

NAND2X1 _1688_ (
    .A(_874_),
    .B(_861_),
    .Y(_875_)
);

NAND3X1 _1268_ (
    .A(_313_),
    .B(_365_),
    .C(_361_),
    .Y(_374_)
);

FILL FILL_0__1728_ (
);

FILL FILL_0__1308_ (
);

FILL FILL_2__1499_ (
);

FILL FILL_0__1481_ (
);

FILL FILL_0__1061_ (
);

FILL FILL_2__1079_ (
);

FILL FILL_3__952_ (
);

FILL FILL_1__1642_ (
);

FILL FILL_1__1222_ (
);

FILL FILL_3__1148_ (
);

NAND2X1 _1497_ (
    .A(_598_),
    .B(_596_),
    .Y(_599_)
);

AOI22X1 _1077_ (
    .A(BI_0_bF$buf0),
    .B(\u_ALU.AI7 ),
    .C(BI_1_bF$buf3),
    .D(AI[6]),
    .Y(_183_)
);

FILL FILL_2__1711_ (
);

FILL FILL_0__1537_ (
);

FILL FILL_0__1117_ (
);

FILL FILL_0__1290_ (
);

FILL FILL_1__1451_ (
);

FILL FILL_1__1031_ (
);

FILL FILL_3__1377_ (
);

FILL FILL_2__1520_ (
);

FILL FILL_2__1100_ (
);

FILL FILL_0__1766_ (
);

FILL FILL_0__1346_ (
);

FILL FILL_1__1507_ (
);

FILL FILL_1__1680_ (
);

FILL FILL_1__1260_ (
);

FILL FILL_1__897_ (
);

FILL FILL_0__1575_ (
);

FILL FILL_0__1155_ (
);

FILL FILL_0__902_ (
);

INVX1 _905_ (
    .A(LoadB_i),
    .Y(_714_)
);

FILL FILL_1__1736_ (
);

FILL FILL_1__1316_ (
);

FILL FILL_2__1805_ (
);

FILL FILL_0__1384_ (
);

OAI21X1 _1803_ (
    .A(_775_),
    .B(_796_),
    .C(_795_),
    .Y(_811_)
);

FILL FILL_1__1545_ (
);

FILL FILL_1__1125_ (
);

FILL FILL_2__969_ (
);

FILL FILL_0__1193_ (
);

DFFSR _1612_ (
    .D(_4_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf0),
    .Q(BI[3])
);

FILL FILL_0__940_ (
);

OAI21X1 _943_ (
    .A(_50_),
    .B(_32__bF$buf2),
    .C(_51_),
    .Y(_6_)
);

FILL FILL_1__1774_ (
);

FILL FILL_1__1354_ (
);

FILL FILL_2__1423_ (
);

FILL FILL_2__1003_ (
);

FILL FILL_0__1669_ (
);

FILL FILL_0__1249_ (
);

AOI21X1 _1421_ (
    .A(_473_),
    .B(_475_),
    .C(_524_),
    .Y(_525_)
);

AND2X2 _1001_ (
    .A(BI_3_bF$buf3),
    .B(AI[2]),
    .Y(_107_)
);

FILL FILL_1__1583_ (
);

FILL FILL_1__1163_ (
);

FILL FILL_2__1652_ (
);

FILL FILL_2__1232_ (
);

FILL FILL_0__1478_ (
);

FILL FILL_0__1058_ (
);

FILL FILL_3__949_ (
);

FILL FILL_3__1301_ (
);

FILL FILL_1__1639_ (
);

FILL FILL_1__1219_ (
);

OAI21X1 _1650_ (
    .A(ABCmd_i[0]),
    .B(_836_),
    .C(_837_),
    .Y(_838_)
);

INVX1 _1230_ (
    .A(_335_),
    .Y(_336_)
);

AOI21X1 _981_ (
    .A(_76_),
    .B(_79_),
    .C(_67_),
    .Y(_87_)
);

FILL FILL_1__1392_ (
);

FILL FILL_2__1708_ (
);

FILL FILL_2__1461_ (
);

FILL FILL_2__1041_ (
);

FILL FILL_0__1287_ (
);

OAI21X1 _1706_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .C(_720_),
    .Y(_721_)
);

FILL FILL_3__1530_ (
);

FILL FILL_1__1448_ (
);

FILL FILL_1__1028_ (
);

FILL FILL_2__1517_ (
);

FILL FILL_2__1690_ (
);

FILL FILL_2__1270_ (
);

FILL FILL_0__1096_ (
);

NAND3X1 _1515_ (
    .A(_311_),
    .B(_616_),
    .C(_615_),
    .Y(_617_)
);

FILL FILL_1__1677_ (
);

FILL FILL_1__1257_ (
);

FILL FILL_2__1746_ (
);

FILL FILL_2__1326_ (
);

FILL FILL_3__1815_ (
);

NAND2X1 _1744_ (
    .A(AI_5_bF$buf0),
    .B(_755_),
    .Y(_756_)
);

NAND3X1 _1324_ (
    .A(_416_),
    .B(_421_),
    .C(_419_),
    .Y(_429_)
);

FILL FILL_1__1486_ (
);

FILL FILL_1__1066_ (
);

FILL FILL_2__1555_ (
);

FILL FILL_2__1135_ (
);

FILL FILL_3__1204_ (
);

INVX1 _1553_ (
    .A(ACC[5]),
    .Y(_654_)
);

OAI21X1 _1133_ (
    .A(_231_),
    .B(_232_),
    .C(_229_),
    .Y(_239_)
);

FILL FILL_1__915_ (
);

FILL FILL_1__1295_ (
);

FILL FILL_2__1784_ (
);

FILL FILL_2__1364_ (
);

FILL FILL_1_CLKBUF1_insert8 (
);

FILL FILL_1_CLKBUF1_insert9 (
);

DFFSR _1609_ (
    .D(_1_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(BI[0])
);

FILL FILL_0__937_ (
);

FILL FILL94350x4050 (
);

FILL FILL_3__1433_ (
);

OAI21X1 _1782_ (
    .A(_791_),
    .B(_790_),
    .C(_787_),
    .Y(_792_)
);

OAI21X1 _1362_ (
    .A(_466_),
    .B(_464_),
    .C(_465_),
    .Y(_467_)
);

FILL FILL_0__1822_ (
);

FILL FILL_0__1402_ (
);

FILL FILL_2__931_ (
);

FILL FILL_2__1593_ (
);

FILL FILL_2__1173_ (
);

OAI21X1 _1418_ (
    .A(_402_),
    .B(_521_),
    .C(_442_),
    .Y(_522_)
);

FILL FILL_3__1662_ (
);

AOI21X1 _1591_ (
    .A(_689_),
    .B(_703_),
    .C(_712_),
    .Y(_690_)
);

NAND3X1 _1171_ (
    .A(_276_),
    .B(_275_),
    .C(_270_),
    .Y(_277_)
);

FILL FILL_1__953_ (
);

FILL FILL94350x150 (
);

FILL FILL_2__1649_ (
);

FILL FILL_2__1229_ (
);

FILL FILL_0__1211_ (
);

FILL FILL_3__1718_ (
);

INVX2 _1647_ (
    .A(ABCmd_i[5]),
    .Y(_835_)
);

INVX1 _1227_ (
    .A(_327_),
    .Y(_333_)
);

FILL FILL_0__975_ (
);

FILL FILL_3__1051_ (
);

NAND2X1 _978_ (
    .A(BI_3_bF$buf3),
    .B(AI[1]),
    .Y(_84_)
);

FILL FILL_1__1389_ (
);

FILL FILL_2__1458_ (
);

FILL FILL_0__1440_ (
);

FILL FILL_2__1038_ (
);

FILL FILL_0__1020_ (
);

FILL FILL_1__1601_ (
);

FILL FILL_3__1527_ (
);

OAI21X1 _1456_ (
    .A(_423_),
    .B(_558_),
    .C(_494_),
    .Y(_559_)
);

NAND3X1 _1036_ (
    .A(_132_),
    .B(_133_),
    .C(_128_),
    .Y(_142_)
);

FILL FILL_3__1280_ (
);

FILL FILL_1__1198_ (
);

FILL FILL_1__991_ (
);

FILL FILL_2__1687_ (
);

FILL FILL_2__1267_ (
);

FILL FILL_1__1410_ (
);

FILL FILL_3__1756_ (
);

OAI21X1 _1685_ (
    .A(_844_),
    .B(_857_),
    .C(_855_),
    .Y(_872_)
);

OAI21X1 _1265_ (
    .A(_366_),
    .B(_370_),
    .C(_312_),
    .Y(_371_)
);

FILL FILL_0__1725_ (
);

FILL FILL_0__1305_ (
);

FILL FILL_2__1496_ (
);

FILL FILL_2__1076_ (
);

FILL FILL_3__1145_ (
);

OR2X2 _1494_ (
    .A(_595_),
    .B(_593_),
    .Y(_596_)
);

AOI21X1 _1074_ (
    .A(_158_),
    .B(_156_),
    .C(_143_),
    .Y(_180_)
);

FILL FILL_0__1534_ (
);

FILL FILL_0__1114_ (
);

FILL FILL_3__1794_ (
);

FILL FILL_3__1374_ (
);

BUFX2 BUFX2_insert0 (
    .A(BI[3]),
    .Y(BI_3_bF$buf3)
);

BUFX2 BUFX2_insert1 (
    .A(BI[3]),
    .Y(BI_3_bF$buf2)
);

BUFX2 BUFX2_insert2 (
    .A(BI[3]),
    .Y(BI_3_bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .A(BI[3]),
    .Y(BI_3_bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .A(BI[0]),
    .Y(BI_0_bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .A(BI[0]),
    .Y(BI_0_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .A(BI[0]),
    .Y(BI_0_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .A(BI[0]),
    .Y(BI_0_bF$buf0)
);

FILL FILL_0__1763_ (
);

FILL FILL_0__1343_ (
);

FILL FILL_1__1504_ (
);

NAND2X1 _1779_ (
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .Y(_789_)
);

AND2X2 _1359_ (
    .A(_271_),
    .B(_293_),
    .Y(_464_)
);

FILL FILL_3__1183_ (
);

FILL FILL_0__1819_ (
);

FILL FILL_1__894_ (
);

FILL FILL_2__928_ (
);

FILL FILL_0__1572_ (
);

FILL FILL_0__1152_ (
);

INVX1 _902_ (
    .A(LoadA_i),
    .Y(_711_)
);

FILL FILL_1__1733_ (
);

FILL FILL_1__1313_ (
);

FILL FILL_3__1659_ (
);

XNOR2X1 _1588_ (
    .A(_686_),
    .B(_310_),
    .Y(_687_)
);

AOI22X1 _1168_ (
    .A(BI_0_bF$buf2),
    .B(AI[2]),
    .C(BI_1_bF$buf1),
    .D(AI[1]),
    .Y(_274_)
);

FILL FILL_2__1802_ (
);

FILL FILL_0__1208_ (
);

FILL FILL_0__1381_ (
);

FILL FILL_2__1399_ (
);

NAND2X1 _1800_ (
    .A(_806_),
    .B(_807_),
    .Y(_808_)
);

FILL FILL_1__1542_ (
);

FILL FILL_1__1122_ (
);

FILL FILL_3__1048_ (
);

INVX1 _1397_ (
    .A(_500_),
    .Y(_501_)
);

FILL FILL_0__1437_ (
);

FILL FILL_0__1017_ (
);

FILL FILL_2__966_ (
);

FILL FILL_0__1190_ (
);

OAI21X1 _940_ (
    .A(_48_),
    .B(_32__bF$buf0),
    .C(_49_),
    .Y(_5_)
);

FILL FILL_1__1771_ (
);

FILL FILL_1__1351_ (
);

FILL FILL_3__1697_ (
);

FILL FILL_3__1277_ (
);

FILL FILL_1__988_ (
);

FILL FILL_2__1420_ (
);

FILL FILL_2__1000_ (
);

FILL FILL_0__1666_ (
);

FILL FILL_0__1246_ (
);

FILL FILL_1__1827_ (
);

FILL FILL_1__1407_ (
);

FILL FILL_1__1580_ (
);

FILL FILL_1__1160_ (
);

FILL FILL_0__1475_ (
);

FILL FILL_0__1055_ (
);

FILL FILL_3__946_ (
);

FILL FILL_1__1636_ (
);

FILL FILL_1__1216_ (
);

FILL FILL_2__1705_ (
);

FILL FILL_0__1284_ (
);

XOR2X1 _1703_ (
    .A(_877_),
    .B(_718_),
    .Y(_719_)
);

FILL FILL94050x74250 (
);

FILL FILL_1__1445_ (
);

FILL FILL_1__1025_ (
);

FILL FILL_2__1514_ (
);

FILL FILL_0__1093_ (
);

NAND2X1 _1512_ (
    .A(_613_),
    .B(_611_),
    .Y(_614_)
);

FILL FILL_3__984_ (
);

FILL FILL_1__1674_ (
);

FILL FILL_1__1254_ (
);

FILL FILL_2__1743_ (
);

FILL FILL_2__1323_ (
);

FILL FILL_0__1569_ (
);

FILL FILL_0__1149_ (
);

FILL FILL_3__1812_ (
);

AOI21X1 _1741_ (
    .A(HC),
    .B(_751_),
    .C(_752_),
    .Y(_753_)
);

AOI21X1 _1321_ (
    .A(_424_),
    .B(_425_),
    .C(_415_),
    .Y(_426_)
);

FILL FILL_1__1483_ (
);

FILL FILL_1__1063_ (
);

FILL FILL_2__1552_ (
);

FILL FILL_2__1132_ (
);

FILL FILL_0__1798_ (
);

FILL FILL_0__1378_ (
);

FILL FILL_3__1201_ (
);

FILL FILL_1__1539_ (
);

FILL FILL_1__1119_ (
);

NAND3X1 _1550_ (
    .A(_636_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

OAI21X1 _1130_ (
    .A(_231_),
    .B(_232_),
    .C(_235_),
    .Y(_236_)
);

FILL FILL_1__912_ (
);

FILL FILL_1__1292_ (
);

FILL FILL_2__1608_ (
);

FILL FILL_2__1781_ (
);

FILL FILL_2__1361_ (
);

FILL FILL_0__1187_ (
);

OAI21X1 _1606_ (
    .A(_52_),
    .B(_705__bF$buf1),
    .C(_697_),
    .Y(_23_)
);

FILL FILL_0__934_ (
);

FILL FILL_3__1430_ (
);

OAI21X1 _937_ (
    .A(_46_),
    .B(_32__bF$buf1),
    .C(_47_),
    .Y(_4_)
);

FILL FILL_1__1768_ (
);

FILL FILL_1__1348_ (
);

FILL FILL_2__1417_ (
);

FILL FILL_2__1590_ (
);

FILL FILL_2__1170_ (
);

NAND2X1 _1415_ (
    .A(_518_),
    .B(_515_),
    .Y(_519_)
);

FILL FILL_1__1577_ (
);

FILL FILL_1__1157_ (
);

FILL FILL_1__950_ (
);

FILL FILL_2__1646_ (
);

FILL FILL_2__1226_ (
);

FILL FILL_3__1715_ (
);

NAND2X1 _1644_ (
    .A(BI_0_bF$buf3),
    .B(_831_),
    .Y(_832_)
);

AND2X2 _1224_ (
    .A(AI_5_bF$buf3),
    .B(BI_3_bF$buf1),
    .Y(_330_)
);

FILL FILL_0__972_ (
);

INVX1 _975_ (
    .A(_59_),
    .Y(_81_)
);

FILL FILL_1__1386_ (
);

FILL FILL_2__1455_ (
);

FILL FILL_2__1035_ (
);

FILL FILL_3__1524_ (
);

FILL FILL_3__1104_ (
);

NAND2X1 _1453_ (
    .A(\u_ALU.AI7 ),
    .B(BI[5]),
    .Y(_556_)
);

AOI21X1 _1033_ (
    .A(_138_),
    .B(_135_),
    .C(_126_),
    .Y(_139_)
);

FILL FILL_1__1195_ (
);

FILL FILL_2__1684_ (
);

FILL FILL_2__1264_ (
);

NAND3X1 _1509_ (
    .A(_569_),
    .B(_571_),
    .C(_610_),
    .Y(_611_)
);

FILL FILL_3__1333_ (
);

NAND2X1 _1682_ (
    .A(_868_),
    .B(_867_),
    .Y(_869_)
);

NAND3X1 _1262_ (
    .A(_356_),
    .B(_360_),
    .C(_362_),
    .Y(_368_)
);

FILL FILL_0__1722_ (
);

FILL FILL_0__1302_ (
);

FILL FILL_2__1493_ (
);

FILL FILL_2__1073_ (
);

FILL FILL_3__1809_ (
);

FILL FILL94050x62550 (
);

INVX1 _1738_ (
    .A(_750_),
    .Y(_751_)
);

INVX2 _1318_ (
    .A(AI[6]),
    .Y(_423_)
);

FILL FILL_3__1562_ (
);

NAND2X1 _1491_ (
    .A(AI_5_bF$buf1),
    .B(BI[7]),
    .Y(_593_)
);

NAND2X1 _1071_ (
    .A(_168_),
    .B(_169_),
    .Y(_177_)
);

FILL FILL_0__1531_ (
);

FILL FILL_2__1549_ (
);

FILL FILL_2__1129_ (
);

FILL FILL_0__1111_ (
);

NOR2X1 _1547_ (
    .A(_638_),
    .B(_647_),
    .Y(_648_)
);

NAND3X1 _1127_ (
    .A(_219_),
    .B(_227_),
    .C(_226_),
    .Y(_233_)
);

FILL FILL_1__909_ (
);

FILL FILL_3__1791_ (
);

FILL FILL_1__1289_ (
);

FILL FILL_0__1760_ (
);

FILL FILL_2__1778_ (
);

FILL FILL_2__1358_ (
);

FILL FILL_0__1340_ (
);

FILL FILL_1__1501_ (
);

FILL FILL_3__1427_ (
);

OAI21X1 _1776_ (
    .A(_776_),
    .B(_783_),
    .C(_775_),
    .Y(_786_)
);

AND2X2 _1356_ (
    .A(_398_),
    .B(_460_),
    .Y(_461_)
);

FILL FILL_3__1180_ (
);

FILL FILL_1__1098_ (
);

FILL FILL_0__1816_ (
);

FILL FILL_1__891_ (
);

FILL FILL_2__925_ (
);

FILL FILL_2__1587_ (
);

FILL FILL_2__1167_ (
);

FILL FILL_1__1730_ (
);

FILL FILL_1__1310_ (
);

FILL FILL_3__1656_ (
);

NAND2X1 _1585_ (
    .A(_642_),
    .B(_683_),
    .Y(_684_)
);

NAND2X1 _1165_ (
    .A(BI_0_bF$buf1),
    .B(AI[1]),
    .Y(_271_)
);

FILL FILL_1__947_ (
);

FILL FILL_0__1205_ (
);

FILL FILL_2__1396_ (
);

FILL FILL_0__969_ (
);

FILL FILL_3__1045_ (
);

XNOR2X1 _1394_ (
    .A(_497_),
    .B(_492_),
    .Y(_498_)
);

FILL FILL_0__1434_ (
);

FILL FILL_0__1014_ (
);

FILL FILL_2__963_ (
);

FILL FILL_3__905_ (
);

FILL FILL_3__1694_ (
);

FILL FILL_3__1274_ (
);

FILL FILL_1__985_ (
);

FILL FILL_0__1663_ (
);

FILL FILL_0__1243_ (
);

FILL FILL_1__1824_ (
);

FILL FILL_1__1404_ (
);

NAND2X1 _1679_ (
    .A(BI_0_bF$buf2),
    .B(_833_),
    .Y(_866_)
);

OAI21X1 _1259_ (
    .A(_363_),
    .B(_364_),
    .C(_362_),
    .Y(_365_)
);

FILL FILL_3__1083_ (
);

FILL FILL_0__1719_ (
);

FILL FILL_0__1472_ (
);

FILL FILL_0__1052_ (
);

FILL FILL_1__1213_ (
);

FILL FILL_3__1559_ (
);

OAI21X1 _1488_ (
    .A(_545_),
    .B(_550_),
    .C(_549_),
    .Y(_590_)
);

AOI21X1 _1068_ (
    .A(_157_),
    .B(_161_),
    .C(_125_),
    .Y(_174_)
);

FILL FILL_2__1702_ (
);

FILL FILL_0__1528_ (
);

FILL FILL_0__1108_ (
);

FILL FILL_0__1281_ (
);

FILL FILL_2__1299_ (
);

FILL FILL94350x78150 (
);

AOI21X1 _1700_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[2]),
    .C(_885_),
    .Y(_716_)
);

FILL FILL_1__1442_ (
);

FILL FILL_1__1022_ (
);

FILL FILL_3__1788_ (
);

INVX1 _1297_ (
    .A(_401_),
    .Y(_402_)
);

FILL FILL_2__1511_ (
);

FILL FILL_0__1757_ (
);

FILL FILL_0__1337_ (
);

FILL FILL_0__1090_ (
);

FILL FILL_3__981_ (
);

FILL FILL_1__1671_ (
);

FILL FILL_1__1251_ (
);

FILL FILL_3__1177_ (
);

FILL FILL_2__1740_ (
);

FILL FILL_2__1320_ (
);

FILL FILL_0__1566_ (
);

FILL FILL_0__1146_ (
);

FILL FILL_1__1727_ (
);

FILL FILL_1__1307_ (
);

FILL FILL_0_BUFX2_insert40 (
);

FILL FILL_0_BUFX2_insert41 (
);

FILL FILL_1__1480_ (
);

FILL FILL_1__1060_ (
);

FILL FILL_0__1795_ (
);

FILL FILL_0__1375_ (
);

FILL FILL_1__1536_ (
);

FILL FILL_1__1116_ (
);

FILL FILL_2__1605_ (
);

FILL FILL_0__1184_ (
);

NAND2X1 _1603_ (
    .A(AI_5_bF$buf0),
    .B(_705__bF$buf0),
    .Y(_696_)
);

FILL FILL_0__931_ (
);

OAI21X1 _934_ (
    .A(_44_),
    .B(_32__bF$buf3),
    .C(_45_),
    .Y(_3_)
);

FILL FILL_1__1765_ (
);

FILL FILL_1__1345_ (
);

FILL FILL_2__1414_ (
);

NAND3X1 _1412_ (
    .A(_507_),
    .B(_502_),
    .C(_509_),
    .Y(_516_)
);

FILL FILL_1__1574_ (
);

FILL FILL_1__1154_ (
);

FILL FILL_2__1643_ (
);

FILL FILL_2__1223_ (
);

FILL FILL_0__1469_ (
);

FILL FILL_0__1049_ (
);

FILL FILL_2__998_ (
);

FILL FILL_3__1712_ (
);

INVX2 _1641_ (
    .A(ABCmd_i[1]),
    .Y(_829_)
);

NAND2X1 _1221_ (
    .A(BI[5]),
    .B(AI[3]),
    .Y(_327_)
);

AND2X2 _972_ (
    .A(_70_),
    .B(_71_),
    .Y(_78_)
);

FILL FILL_1__1383_ (
);

FILL FILL_2__1452_ (
);

FILL FILL_2__1032_ (
);

FILL FILL_0__1698_ (
);

FILL FILL_0__1278_ (
);

FILL FILL_3__1101_ (
);

FILL FILL_1__1439_ (
);

FILL FILL_1__1019_ (
);

INVX1 _1450_ (
    .A(_549_),
    .Y(_553_)
);

NOR2X1 _1030_ (
    .A(_97_),
    .B(_131_),
    .Y(_136_)
);

FILL FILL_1__1192_ (
);

FILL FILL_2__1508_ (
);

FILL FILL_2__1681_ (
);

FILL FILL_2__1261_ (
);

FILL FILL_0__1087_ (
);

OR2X2 _1506_ (
    .A(_603_),
    .B(_563_),
    .Y(_608_)
);

FILL FILL_3__978_ (
);

FILL FILL_3__1330_ (
);

FILL FILL_1__1668_ (
);

FILL FILL_1__1248_ (
);

FILL FILL_2__1737_ (
);

FILL FILL_2__1317_ (
);

FILL FILL_2__1490_ (
);

FILL FILL_2__1070_ (
);

FILL FILL_3__1806_ (
);

AOI21X1 _1735_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_4_bF$buf0),
    .C(_747_),
    .Y(_748_)
);

AOI22X1 _1315_ (
    .A(AI[6]),
    .B(BI_3_bF$buf1),
    .C(AI_5_bF$buf3),
    .D(BI_4_bF$buf3),
    .Y(_420_)
);

FILL FILL_1__1477_ (
);

FILL FILL_1__1057_ (
);

FILL FILL_2__1546_ (
);

FILL FILL_2__1126_ (
);

XNOR2X1 _1544_ (
    .A(_602_),
    .B(_644_),
    .Y(_645_)
);

NAND3X1 _1124_ (
    .A(_229_),
    .B(_213_),
    .C(_217_),
    .Y(_230_)
);

FILL FILL_1__906_ (
);

FILL FILL_1__1286_ (
);

FILL FILL_2__1775_ (
);

FILL FILL_2__1355_ (
);

FILL FILL_0__928_ (
);

FILL FILL_3__1424_ (
);

FILL FILL_3__1004_ (
);

INVX1 _1773_ (
    .A(_776_),
    .Y(_784_)
);

NAND3X1 _1353_ (
    .A(_402_),
    .B(_452_),
    .C(_451_),
    .Y(_458_)
);

FILL FILL_1__1095_ (
);

FILL FILL_0__1813_ (
);

FILL FILL_2__922_ (
);

FILL FILL_2__1584_ (
);

FILL FILL_2__1164_ (
);

AOI21X1 _1409_ (
    .A(_511_),
    .B(_512_),
    .C(_490_),
    .Y(_513_)
);

FILL FILL_3__1233_ (
);

INVX1 _1582_ (
    .A(_886_[7]),
    .Y(_681_)
);

AOI21X1 _1162_ (
    .A(_267_),
    .B(_266_),
    .C(_265_),
    .Y(_268_)
);

FILL FILL_1__944_ (
);

FILL FILL_0__1202_ (
);

FILL FILL_2__1393_ (
);

FILL FILL_3__1709_ (
);

OAI21X1 _1638_ (
    .A(_824_),
    .B(_825_),
    .C(ABCmd_i[4]),
    .Y(_826_)
);

OAI21X1 _1218_ (
    .A(_323_),
    .B(_322_),
    .C(_315_),
    .Y(_324_)
);

FILL FILL_0__966_ (
);

FILL FILL_3__1462_ (
);

OAI21X1 _969_ (
    .A(_73_),
    .B(_74_),
    .C(_70_),
    .Y(_75_)
);

AOI22X1 _1391_ (
    .A(\u_ALU.AI7 ),
    .B(BI_3_bF$buf0),
    .C(AI[6]),
    .D(BI_4_bF$buf3),
    .Y(_495_)
);

FILL FILL_0__1431_ (
);

FILL FILL_2__1449_ (
);

FILL FILL_2__1029_ (
);

FILL FILL_0__1011_ (
);

FILL FILL_2__960_ (
);

FILL FILL_3__902_ (
);

NOR2X1 _1447_ (
    .A(_547_),
    .B(_548_),
    .Y(_550_)
);

NAND2X1 _1027_ (
    .A(BI[2]),
    .B(AI[4]),
    .Y(_133_)
);

FILL FILL_3__1691_ (
);

FILL FILL_1__1189_ (
);

FILL FILL_1__982_ (
);

FILL FILL_0__1660_ (
);

FILL FILL_2__1678_ (
);

FILL FILL_0__1240_ (
);

FILL FILL_2__1258_ (
);

FILL FILL_1__1821_ (
);

FILL FILL_1__1401_ (
);

FILL FILL_3__1747_ (
);

FILL FILL_3__1327_ (
);

OAI21X1 _1676_ (
    .A(_836_),
    .B(_824_),
    .C(_862_),
    .Y(_863_)
);

AOI21X1 _1256_ (
    .A(_213_),
    .B(_229_),
    .C(_232_),
    .Y(_362_)
);

FILL FILL_3__1080_ (
);

FILL FILL_0__1716_ (
);

FILL FILL_2__1487_ (
);

FILL FILL_2__1067_ (
);

FILL FILL_1__1210_ (
);

FILL FILL_3__1556_ (
);

AOI21X1 _1485_ (
    .A(_587_),
    .B(_703_),
    .C(_712_),
    .Y(_588_)
);

INVX1 _1065_ (
    .A(_170_),
    .Y(_171_)
);

FILL FILL_0__1525_ (
);

FILL FILL_0__1105_ (
);

FILL FILL_2__1296_ (
);

FILL FILL_3__1785_ (
);

INVX1 _1294_ (
    .A(_361_),
    .Y(_399_)
);

FILL FILL_0__1754_ (
);

FILL FILL_0__1334_ (
);

FILL FILL_3__1174_ (
);

FILL FILL_2__919_ (
);

FILL FILL_0__1563_ (
);

FILL FILL_0__1143_ (
);

FILL FILL_1__1724_ (
);

FILL FILL_1__1304_ (
);

FILL FILL_0_BUFX2_insert13 (
);

NOR2X1 _1579_ (
    .A(_678_),
    .B(_25_),
    .Y(_679_)
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

AOI22X1 _1159_ (
    .A(_122_),
    .B(_262_),
    .C(_263_),
    .D(_264_),
    .Y(_265_)
);

FILL FILL_0_BUFX2_insert16 (
);

FILL FILL_0_BUFX2_insert17 (
);

FILL FILL_0_BUFX2_insert18 (
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL94350x7950 (
);

FILL FILL_0__1792_ (
);

FILL FILL_0__1372_ (
);

FILL FILL_1__1533_ (
);

FILL FILL_1__1113_ (
);

FILL FILL_3__1459_ (
);

NAND2X1 _1388_ (
    .A(AI_5_bF$buf1),
    .B(BI[5]),
    .Y(_492_)
);

FILL FILL_2__1602_ (
);

FILL FILL_0__1428_ (
);

FILL FILL_0__1008_ (
);

FILL FILL_2__957_ (
);

FILL FILL_0__1181_ (
);

FILL FILL_2__1199_ (
);

OAI21X1 _1600_ (
    .A(_46_),
    .B(_705__bF$buf0),
    .C(_694_),
    .Y(_20_)
);

OAI21X1 _931_ (
    .A(_42_),
    .B(_32__bF$buf2),
    .C(_43_),
    .Y(_2_)
);

FILL FILL_1__1762_ (
);

FILL FILL_1__1342_ (
);

FILL FILL_3__1688_ (
);

NOR3X1 _1197_ (
    .A(_302_),
    .B(_301_),
    .C(_282_),
    .Y(_303_)
);

FILL FILL_1__979_ (
);

FILL FILL_2__1411_ (
);

FILL FILL_0__1657_ (
);

FILL FILL_0__1237_ (
);

FILL FILL_1__1818_ (
);

FILL FILL_1__1571_ (
);

FILL FILL_1__1151_ (
);

FILL FILL_3__1077_ (
);

BUFX2 BUFX2_insert20 (
    .A(_0_),
    .Y(_0__bF$buf1)
);

BUFX2 BUFX2_insert21 (
    .A(_0_),
    .Y(_0__bF$buf0)
);

BUFX2 BUFX2_insert22 (
    .A(AI[5]),
    .Y(AI_5_bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .A(AI[5]),
    .Y(AI_5_bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .A(AI[5]),
    .Y(AI_5_bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .A(AI[5]),
    .Y(AI_5_bF$buf0)
);

BUFX2 BUFX2_insert26 (
    .A(_32_),
    .Y(_32__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(_32_),
    .Y(_32__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(_32_),
    .Y(_32__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(_32_),
    .Y(_32__bF$buf0)
);

FILL FILL_2__1640_ (
);

FILL FILL_2__1220_ (
);

FILL FILL_0__1466_ (
);

FILL FILL_0__1046_ (
);

FILL FILL_2__995_ (
);

FILL FILL_1__1207_ (
);

FILL FILL_1__1380_ (
);

FILL FILL_0__1695_ (
);

FILL FILL_0__1275_ (
);

FILL FILL_1__1436_ (
);

FILL FILL_1__1016_ (
);

FILL FILL_2__1505_ (
);

FILL FILL_0__1084_ (
);

NAND2X1 _1503_ (
    .A(_563_),
    .B(_603_),
    .Y(_605_)
);

FILL FILL_3__975_ (
);

FILL FILL_1__1665_ (
);

FILL FILL_1__1245_ (
);

FILL FILL_2__1734_ (
);

FILL FILL_2__1314_ (
);

OAI21X1 _1732_ (
    .A(AI[4]),
    .B(_742_),
    .C(_835_),
    .Y(_745_)
);

AND2X2 _1312_ (
    .A(AI_5_bF$buf1),
    .B(BI_4_bF$buf3),
    .Y(_417_)
);

FILL FILL_1__1474_ (
);

FILL FILL_1__1054_ (
);

FILL FILL_2__1543_ (
);

FILL FILL_2__1123_ (
);

FILL FILL_0__1789_ (
);

FILL FILL_0__1369_ (
);

FILL FILL_2__898_ (
);

NAND3X1 _1541_ (
    .A(AI[6]),
    .B(BI[6]),
    .C(_641_),
    .Y(_642_)
);

OAI21X1 _1121_ (
    .A(_167_),
    .B(_113_),
    .C(_220_),
    .Y(_227_)
);

FILL FILL_1__903_ (
);

FILL FILL_1__1283_ (
);

FILL FILL_2__1772_ (
);

FILL FILL_2__1352_ (
);

FILL FILL_0__1598_ (
);

FILL FILL_0__1178_ (
);

FILL FILL_0__925_ (
);

FILL FILL_3__1001_ (
);

OAI21X1 _928_ (
    .A(_40_),
    .B(_32__bF$buf0),
    .C(_41_),
    .Y(_1_)
);

FILL FILL_1__1759_ (
);

FILL FILL_1__1339_ (
);

OAI21X1 _1770_ (
    .A(_750_),
    .B(_780_),
    .C(_749_),
    .Y(_781_)
);

AOI21X1 _1350_ (
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_455_)
);

FILL FILL_1__1092_ (
);

FILL FILL_0__1810_ (
);

FILL FILL_2__1408_ (
);

FILL FILL_2__1581_ (
);

FILL FILL_2__1161_ (
);

BUFX2 _1826_ (
    .A(_887_),
    .Y(Done_LED)
);

AOI22X1 _1406_ (
    .A(_486_),
    .B(_489_),
    .C(_506_),
    .D(_500_),
    .Y(_510_)
);

FILL FILL_3__1230_ (
);

FILL FILL_1__1568_ (
);

FILL FILL_1__1148_ (
);

FILL FILL_1__941_ (
);

FILL FILL_2__1637_ (
);

FILL FILL_2__1217_ (
);

FILL FILL_2__1390_ (
);

FILL FILL_3__1706_ (
);

DFFSR _1635_ (
    .D(_888_[2]),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf2),
    .Q(state[2])
);

NAND3X1 _1215_ (
    .A(_316_),
    .B(_319_),
    .C(_320_),
    .Y(_321_)
);

FILL FILL_0__963_ (
);

FILL FILL_2_CLKBUF1_insert10 (
);

FILL FILL_2_CLKBUF1_insert11 (
);

OR2X2 _966_ (
    .A(_70_),
    .B(_71_),
    .Y(_72_)
);

FILL FILL_2_CLKBUF1_insert12 (
);

FILL FILL_1__1797_ (
);

FILL FILL_1__1377_ (
);

FILL FILL_2__1446_ (
);

FILL FILL_2__1026_ (
);

NOR2X1 _1444_ (
    .A(_130_),
    .B(_167_),
    .Y(_547_)
);

INVX2 _1024_ (
    .A(AI_5_bF$buf1),
    .Y(_130_)
);

FILL FILL_1__1186_ (
);

FILL FILL_2__1675_ (
);

FILL FILL_2__1255_ (
);

FILL FILL94350x19650 (
);

FILL FILL_3__1744_ (
);

FILL FILL_3__1324_ (
);

MUX2X1 _1673_ (
    .A(_859_),
    .B(_858_),
    .S(_855_),
    .Y(_860_)
);

OAI21X1 _1253_ (
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_359_)
);

FILL FILL_0__1713_ (
);

FILL FILL_2__1484_ (
);

FILL FILL_2__1064_ (
);

AND2X2 _1729_ (
    .A(_831_),
    .B(BI_4_bF$buf0),
    .Y(_742_)
);

NAND2X1 _1309_ (
    .A(\u_ALU.AI7 ),
    .B(BI[2]),
    .Y(_414_)
);

FILL FILL_3__1553_ (
);

FILL FILL_3__1133_ (
);

NAND2X1 _1482_ (
    .A(_301_),
    .B(_584_),
    .Y(_585_)
);

NOR2X1 _1062_ (
    .A(_57_),
    .B(_167_),
    .Y(_168_)
);

FILL FILL_0__1522_ (
);

FILL FILL_0__1102_ (
);

FILL FILL_2__1293_ (
);

AOI21X1 _1538_ (
    .A(_590_),
    .B(_605_),
    .C(_604_),
    .Y(_639_)
);

NAND2X1 _1118_ (
    .A(_223_),
    .B(_220_),
    .Y(_224_)
);

FILL FILL_3__1362_ (
);

AOI21X1 _1291_ (
    .A(_395_),
    .B(_389_),
    .C(_246_),
    .Y(_396_)
);

FILL FILL_0__1751_ (
);

FILL FILL_2__1769_ (
);

FILL FILL_0__1331_ (
);

FILL FILL_2__1349_ (
);

INVX1 _1767_ (
    .A(ABCmd_i[6]),
    .Y(_778_)
);

OAI21X1 _1347_ (
    .A(_445_),
    .B(_448_),
    .C(_404_),
    .Y(_452_)
);

FILL FILL_3__1591_ (
);

FILL FILL_1__1089_ (
);

FILL FILL_0__1807_ (
);

FILL FILL_2__916_ (
);

FILL FILL_2__1578_ (
);

FILL FILL_0__1560_ (
);

FILL FILL_0__1140_ (
);

FILL FILL_2__1158_ (
);

FILL FILL_1__1721_ (
);

FILL FILL_1__1301_ (
);

FILL FILL_3__1647_ (
);

FILL FILL_3__1227_ (
);

AOI21X1 _1576_ (
    .A(_393_),
    .B(_309_),
    .C(_308_),
    .Y(_676_)
);

NAND3X1 _1156_ (
    .A(_248_),
    .B(_122_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__938_ (
);

FILL FILL_2__1387_ (
);

FILL FILL_1__1530_ (
);

FILL FILL_1__1110_ (
);

FILL FILL_3__1456_ (
);

OAI21X1 _1385_ (
    .A(_488_),
    .B(_487_),
    .C(_480_),
    .Y(_489_)
);

FILL FILL_0__1425_ (
);

FILL FILL_0__1005_ (
);

FILL FILL_2__954_ (
);

FILL FILL_2__1196_ (
);

FILL FILL_3__1685_ (
);

OAI21X1 _1194_ (
    .A(_278_),
    .B(_299_),
    .C(_81_),
    .Y(_300_)
);

FILL FILL_1__976_ (
);

FILL FILL_0__1654_ (
);

FILL FILL_0__1234_ (
);

FILL FILL_1__1815_ (
);

FILL FILL_0__998_ (
);

FILL FILL_3__1074_ (
);

FILL FILL_0__1463_ (
);

FILL FILL_0__1043_ (
);

FILL FILL_2__992_ (
);

FILL FILL_3__934_ (
);

FILL FILL_1__1204_ (
);

OAI21X1 _1479_ (
    .A(_578_),
    .B(_581_),
    .C(_540_),
    .Y(_582_)
);

OAI21X1 _1059_ (
    .A(_139_),
    .B(_143_),
    .C(_160_),
    .Y(_165_)
);

FILL FILL_0__1519_ (
);

FILL FILL_0__1692_ (
);

FILL FILL_0__1272_ (
);

FILL FILL_1__1433_ (
);

FILL FILL_1__1013_ (
);

FILL FILL_3__1359_ (
);

NAND3X1 _1288_ (
    .A(_176_),
    .B(_390_),
    .C(_392_),
    .Y(_393_)
);

FILL FILL_2__1502_ (
);

FILL FILL_0__1748_ (
);

FILL FILL_0__1328_ (
);

FILL FILL_0__1081_ (
);

FILL FILL_2__1099_ (
);

NAND3X1 _1500_ (
    .A(_601_),
    .B(_598_),
    .C(_596_),
    .Y(_602_)
);

FILL FILL_1__1662_ (
);

FILL FILL_1__1242_ (
);

FILL FILL_3__1588_ (
);

OAI21X1 _1097_ (
    .A(_58_),
    .B(_74_),
    .C(_197_),
    .Y(_203_)
);

FILL FILL_2__1731_ (
);

FILL FILL_2__1311_ (
);

FILL FILL_0__1557_ (
);

FILL FILL_0__1137_ (
);

FILL FILL_1__1718_ (
);

FILL FILL93750x150 (
);

FILL FILL_1__1471_ (
);

FILL FILL_1__1051_ (
);

FILL FILL_2__1540_ (
);

FILL FILL_2__1120_ (
);

FILL FILL_0__1786_ (
);

FILL FILL_0__1366_ (
);

FILL FILL_2__895_ (
);

FILL FILL_1__1527_ (
);

FILL FILL_1__1107_ (
);

FILL FILL_1__900_ (
);

FILL FILL_1__1280_ (
);

FILL FILL_0__1595_ (
);

FILL FILL_0__1175_ (
);

FILL FILL_0__922_ (
);

INVX8 _925_ (
    .A(reset),
    .Y(_0_)
);

FILL FILL_1__1756_ (
);

FILL FILL_1__1336_ (
);

FILL FILL_2__1825_ (
);

FILL FILL_2__1405_ (
);

BUFX2 _1823_ (
    .A(_886_[5]),
    .Y(ACC_o[5])
);

NAND3X1 _1403_ (
    .A(_506_),
    .B(_500_),
    .C(_503_),
    .Y(_507_)
);

FILL FILL_1__1565_ (
);

FILL FILL_1__1145_ (
);

FILL FILL_2__1214_ (
);

FILL FILL_2__989_ (
);

DFFSR _1632_ (
    .D(_24_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf1),
    .Q(\u_ALU.AI7 )
);

OAI21X1 _1212_ (
    .A(_195_),
    .B(_200_),
    .C(_199_),
    .Y(_318_)
);

FILL FILL_0__960_ (
);

INVX1 _963_ (
    .A(_68_),
    .Y(_69_)
);

FILL FILL_1__1794_ (
);

FILL FILL_1__1374_ (
);

FILL FILL_2__1443_ (
);

FILL FILL_2__1023_ (
);

FILL FILL_0__1689_ (
);

FILL FILL_0__1269_ (
);

FILL FILL_3__1512_ (
);

AOI21X1 _1441_ (
    .A(_503_),
    .B(_500_),
    .C(_499_),
    .Y(_544_)
);

AND2X2 _1021_ (
    .A(BI_1_bF$buf3),
    .B(AI[6]),
    .Y(_127_)
);

FILL FILL_1__1183_ (
);

FILL FILL_2__1672_ (
);

FILL FILL_2__1252_ (
);

FILL FILL_0__1498_ (
);

FILL FILL_0__1078_ (
);

FILL FILL_3__1741_ (
);

FILL FILL_1__1659_ (
);

FILL FILL_1__1239_ (
);

AOI21X1 _1670_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI_1_bF$buf2),
    .C(_856_),
    .Y(_857_)
);

NAND3X1 _1250_ (
    .A(_325_),
    .B(_355_),
    .C(_351_),
    .Y(_356_)
);

FILL FILL_0__1710_ (
);

FILL FILL_2__1728_ (
);

FILL FILL_2__1308_ (
);

FILL FILL_2__1481_ (
);

FILL FILL_2__1061_ (
);

INVX1 _1726_ (
    .A(_739_),
    .Y(_740_)
);

XNOR2X1 _1306_ (
    .A(_410_),
    .B(_405_),
    .Y(_411_)
);

FILL FILL_3__1550_ (
);

FILL FILL_3__1130_ (
);

FILL FILL_1__1468_ (
);

FILL FILL_1__1048_ (
);

FILL FILL_2__1537_ (
);

FILL FILL_2__1117_ (
);

FILL FILL_2__1290_ (
);

FILL FILL_3__1606_ (
);

INVX1 _1535_ (
    .A(_387_),
    .Y(_636_)
);

INVX1 _1115_ (
    .A(_220_),
    .Y(_221_)
);

FILL FILL_1__1697_ (
);

FILL FILL_1__1277_ (
);

FILL FILL_2__1766_ (
);

FILL FILL_2__1346_ (
);

FILL FILL_0__919_ (
);

OAI21X1 _1764_ (
    .A(_844_),
    .B(_774_),
    .C(_772_),
    .Y(_775_)
);

OAI21X1 _1344_ (
    .A(_445_),
    .B(_448_),
    .C(_444_),
    .Y(_449_)
);

FILL FILL_1__1086_ (
);

FILL FILL_0__1804_ (
);

FILL FILL_2__913_ (
);

FILL FILL_2__1575_ (
);

FILL FILL_2__1155_ (
);

FILL FILL_3__1644_ (
);

FILL FILL_3__1224_ (
);

NAND3X1 _1573_ (
    .A(_636_),
    .B(_669_),
    .C(_672_),
    .Y(_673_)
);

OAI21X1 _1153_ (
    .A(_118_),
    .B(_119_),
    .C(_116_),
    .Y(_259_)
);

FILL FILL_1__935_ (
);

FILL FILL_2__1384_ (
);

DFFSR _1629_ (
    .D(_21_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(AI[4])
);

NAND2X1 _1209_ (
    .A(BI[7]),
    .B(AI[1]),
    .Y(_315_)
);

FILL FILL_0__957_ (
);

FILL FILL_3__1453_ (
);

FILL FILL_3__1033_ (
);

NAND3X1 _1382_ (
    .A(_481_),
    .B(_484_),
    .C(_485_),
    .Y(_486_)
);

FILL FILL_0__1422_ (
);

FILL FILL_0__1002_ (
);

FILL FILL_2__951_ (
);

FILL FILL_2__1193_ (
);

FILL FILL_3__1509_ (
);

INVX1 _1438_ (
    .A(_523_),
    .Y(_541_)
);

OAI21X1 _1018_ (
    .A(_61_),
    .B(_123_),
    .C(_122_),
    .Y(_124_)
);

FILL FILL_3__1262_ (
);

NAND3X1 _1191_ (
    .A(_294_),
    .B(_296_),
    .C(_292_),
    .Y(_297_)
);

FILL FILL_1__973_ (
);

FILL FILL_2__1669_ (
);

FILL FILL_0__1651_ (
);

FILL FILL_0__1231_ (
);

FILL FILL_2__1249_ (
);

FILL FILL_1__1812_ (
);

FILL FILL_3__1738_ (
);

OAI21X1 _1667_ (
    .A(AI[1]),
    .B(_853_),
    .C(_835_),
    .Y(_854_)
);

AOI22X1 _1247_ (
    .A(_332_),
    .B(_337_),
    .C(_349_),
    .D(_348_),
    .Y(_353_)
);

FILL FILL_0__995_ (
);

FILL FILL_3__1491_ (
);

NAND3X1 _998_ (
    .A(_103_),
    .B(_102_),
    .C(_101_),
    .Y(_104_)
);

FILL FILL_0__1707_ (
);

FILL FILL_2__1478_ (
);

FILL FILL_0__1460_ (
);

FILL FILL_0__1040_ (
);

FILL FILL_2__1058_ (
);

FILL FILL_3__931_ (
);

FILL FILL_1__1201_ (
);

FILL FILL_3__1127_ (
);

AOI21X1 _1476_ (
    .A(_527_),
    .B(_528_),
    .C(_541_),
    .Y(_579_)
);

NAND3X1 _1056_ (
    .A(_161_),
    .B(_125_),
    .C(_157_),
    .Y(_162_)
);

FILL FILL_0__1516_ (
);

FILL FILL_2__1287_ (
);

FILL FILL_1__1430_ (
);

FILL FILL_1__1010_ (
);

FILL FILL_3__1356_ (
);

FILL FILL93150x74250 (
);

INVX1 _1285_ (
    .A(_285_),
    .Y(_390_)
);

FILL FILL_0__1745_ (
);

FILL FILL_0__1325_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_1_BUFX2_insert21 (
);

FILL FILL_1_BUFX2_insert22 (
);

FILL FILL_1_BUFX2_insert23 (
);

FILL FILL_1_BUFX2_insert24 (
);

FILL FILL_1_BUFX2_insert25 (
);

FILL FILL_1_BUFX2_insert26 (
);

FILL FILL_1_BUFX2_insert27 (
);

FILL FILL_1_BUFX2_insert28 (
);

FILL FILL_1_BUFX2_insert29 (
);

FILL FILL_2__1096_ (
);

FILL FILL_3__1585_ (
);

AOI22X1 _1094_ (
    .A(BI_3_bF$buf3),
    .B(AI[4]),
    .C(BI_4_bF$buf1),
    .D(AI[3]),
    .Y(_200_)
);

FILL FILL_0__1554_ (
);

FILL FILL_0__1134_ (
);

FILL FILL_1__1715_ (
);

FILL FILL_0__898_ (
);

FILL FILL_0__1783_ (
);

FILL FILL_0__1363_ (
);

FILL FILL_2__892_ (
);

FILL FILL_1__1524_ (
);

FILL FILL_1__1104_ (
);

NAND2X1 _1799_ (
    .A(_799_),
    .B(_786_),
    .Y(_807_)
);

OAI21X1 _1379_ (
    .A(_415_),
    .B(_420_),
    .C(_419_),
    .Y(_483_)
);

FILL FILL_0__1419_ (
);

FILL FILL_2__948_ (
);

FILL FILL_0__1592_ (
);

FILL FILL_0__1172_ (
);

NAND3X1 _922_ (
    .A(_711_),
    .B(_714_),
    .C(_715_),
    .Y(_38_)
);

FILL FILL_1__1753_ (
);

FILL FILL_1__1333_ (
);

FILL FILL_3__1259_ (
);

NOR2X1 _1188_ (
    .A(_271_),
    .B(_293_),
    .Y(_294_)
);

FILL FILL_2__1822_ (
);

FILL FILL_2__1402_ (
);

FILL FILL_0__1648_ (
);

FILL FILL_0__1228_ (
);

FILL FILL_1__1809_ (
);

BUFX2 _1820_ (
    .A(_886_[2]),
    .Y(ACC_o[2])
);

NAND2X1 _1400_ (
    .A(_491_),
    .B(_431_),
    .Y(_504_)
);

FILL FILL_1__1562_ (
);

FILL FILL_1__1142_ (
);

FILL FILL_3__1488_ (
);

FILL FILL_2__1211_ (
);

FILL FILL_0__1457_ (
);

FILL FILL_0__1037_ (
);

FILL FILL_2__986_ (
);

FILL FILL_3__928_ (
);

AND2X2 _960_ (
    .A(_62_),
    .B(_63_),
    .Y(_66_)
);

FILL FILL_1__1791_ (
);

FILL FILL_1__1371_ (
);

FILL FILL_2__1440_ (
);

FILL FILL_2__1020_ (
);

FILL FILL_0__1686_ (
);

FILL FILL_0__1266_ (
);

FILL FILL_1__1427_ (
);

FILL FILL_1__1007_ (
);

FILL FILL_1__1180_ (
);

FILL FILL_0__1495_ (
);

FILL FILL_0__1075_ (
);

FILL FILL_1__1656_ (
);

FILL FILL_1__1236_ (
);

FILL FILL_2__1725_ (
);

FILL FILL_2__1305_ (
);

NAND3X1 _1723_ (
    .A(_735_),
    .B(_875_),
    .C(_736_),
    .Y(_737_)
);

NAND2X1 _1303_ (
    .A(AI_5_bF$buf2),
    .B(BI_4_bF$buf1),
    .Y(_408_)
);

FILL FILL_1__1465_ (
);

FILL FILL_1__1045_ (
);

FILL FILL_2__1534_ (
);

FILL FILL_2__1114_ (
);

FILL FILL_2__889_ (
);

FILL FILL_3__1603_ (
);

AOI21X1 _1532_ (
    .A(_633_),
    .B(_703_),
    .C(_712_),
    .Y(_634_)
);

NAND2X1 _1112_ (
    .A(AI[0]),
    .B(BI[7]),
    .Y(_218_)
);

FILL FILL_1__1694_ (
);

FILL FILL_1__1274_ (
);

FILL FILL_2__1763_ (
);

FILL FILL_2__1343_ (
);

FILL FILL_0__1589_ (
);

FILL FILL_0__1169_ (
);

FILL FILL_0__916_ (
);

FILL FILL_3__1412_ (
);

OR2X2 _919_ (
    .A(_31_),
    .B(_35_),
    .Y(_888_[1])
);

OAI22X1 _1761_ (
    .A(_835_),
    .B(_767_),
    .C(_771_),
    .D(_770_),
    .Y(_772_)
);

NAND3X1 _1341_ (
    .A(_427_),
    .B(_431_),
    .C(_413_),
    .Y(_446_)
);

FILL FILL_1__1083_ (
);

FILL FILL_2__1819_ (
);

FILL FILL_0__1801_ (
);

FILL FILL_2__910_ (
);

FILL FILL_2__1572_ (
);

FILL FILL_2__1152_ (
);

FILL FILL_0__1398_ (
);

NAND2X1 _1817_ (
    .A(_822_),
    .B(_823_),
    .Y(AV)
);

FILL FILL_3__1641_ (
);

FILL FILL_1__1559_ (
);

FILL FILL_1__1139_ (
);

AOI21X1 _1570_ (
    .A(_619_),
    .B(_617_),
    .C(_658_),
    .Y(_670_)
);

AND2X2 _1150_ (
    .A(_61_),
    .B(_85_),
    .Y(_256_)
);

FILL FILL_1__932_ (
);

FILL FILL_2__1208_ (
);

FILL FILL_2__1381_ (
);

DFFSR _1626_ (
    .D(_18_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(AI[1])
);

AOI21X1 _1206_ (
    .A(_178_),
    .B(_243_),
    .C(_241_),
    .Y(_312_)
);

FILL FILL_0__954_ (
);

FILL FILL_3__1030_ (
);

NAND2X1 _957_ (
    .A(BI_0_bF$buf2),
    .B(AI[3]),
    .Y(_63_)
);

FILL FILL_1__1788_ (
);

FILL FILL_1__1368_ (
);

FILL FILL_2__1437_ (
);

FILL FILL_2__1017_ (
);

FILL FILL_2__1190_ (
);

FILL FILL_3__1506_ (
);

INVX1 _1435_ (
    .A(_886_[3]),
    .Y(_538_)
);

OAI21X1 _1015_ (
    .A(_118_),
    .B(_119_),
    .C(_120_),
    .Y(_121_)
);

FILL FILL_1__1597_ (
);

FILL FILL_1__1177_ (
);

FILL FILL_1__970_ (
);

FILL FILL_2__1666_ (
);

FILL FILL_2__1246_ (
);

FILL FILL_3__1735_ (
);

AOI22X1 _1664_ (
    .A(_829_),
    .B(BI_1_bF$buf2),
    .C(_850_),
    .D(_830_),
    .Y(_851_)
);

NAND3X1 _1244_ (
    .A(_348_),
    .B(_349_),
    .C(_347_),
    .Y(_350_)
);

FILL FILL_0__992_ (
);

AOI21X1 _995_ (
    .A(_69_),
    .B(_75_),
    .C(_77_),
    .Y(_101_)
);

FILL FILL_0__1704_ (
);

FILL FILL_2__1475_ (
);

FILL FILL_2__1055_ (
);

FILL FILL_3__1124_ (
);

NAND3X1 _1473_ (
    .A(_568_),
    .B(_571_),
    .C(_575_),
    .Y(_576_)
);

NAND3X1 _1053_ (
    .A(_126_),
    .B(_135_),
    .C(_138_),
    .Y(_159_)
);

FILL FILL_0__1513_ (
);

FILL FILL_2__1284_ (
);

NAND2X1 _1529_ (
    .A(_630_),
    .B(_629_),
    .Y(_631_)
);

NAND3X1 _1109_ (
    .A(_210_),
    .B(_209_),
    .C(_206_),
    .Y(_215_)
);

FILL FILL_3__1773_ (
);

FILL FILL_3__1353_ (
);

OAI21X1 _1282_ (
    .A(state[1]),
    .B(_712_),
    .C(ABCmd_i[7]),
    .Y(_387_)
);

FILL FILL_0__1742_ (
);

FILL FILL_0__1322_ (
);

FILL FILL_2__1093_ (
);

FILL FILL_3__1409_ (
);

NAND2X1 _1758_ (
    .A(AI[6]),
    .B(_768_),
    .Y(_769_)
);

NOR3X1 _1338_ (
    .A(_353_),
    .B(_354_),
    .C(_326_),
    .Y(_443_)
);

FILL FILL_3__1582_ (
);

FILL FILL_3__1162_ (
);

AND2X2 _1091_ (
    .A(BI_4_bF$buf1),
    .B(AI[3]),
    .Y(_197_)
);

FILL FILL_2__907_ (
);

FILL FILL_2__1569_ (
);

FILL FILL_0__1551_ (
);

FILL FILL_2__1149_ (
);

FILL FILL_0__1131_ (
);

FILL FILL_1__1712_ (
);

FILL FILL_3__1638_ (
);

OAI21X1 _1567_ (
    .A(_423_),
    .B(_167_),
    .C(_641_),
    .Y(_667_)
);

OAI21X1 _1147_ (
    .A(_77_),
    .B(_78_),
    .C(_69_),
    .Y(_253_)
);

FILL FILL_0__895_ (
);

FILL FILL_1__929_ (
);

FILL FILL_3__1391_ (
);

NOR2X1 _898_ (
    .A(state[2]),
    .B(_702_),
    .Y(_707_)
);

FILL FILL_0__1607_ (
);

FILL FILL_2__1798_ (
);

FILL FILL_0__1780_ (
);

FILL FILL_0__1360_ (
);

FILL FILL_2__1378_ (
);

FILL FILL_1__1521_ (
);

FILL FILL_1__1101_ (
);

FILL FILL_3__1027_ (
);

FILL FILL_2_BUFX2_insert40 (
);

FILL FILL_2_BUFX2_insert41 (
);

NOR2X1 _1796_ (
    .A(_804_),
    .B(AN),
    .Y(_805_)
);

NAND2X1 _1376_ (
    .A(AI[3]),
    .B(BI[7]),
    .Y(_480_)
);

FILL FILL_0__1416_ (
);

FILL FILL_2__945_ (
);

FILL FILL_2__1187_ (
);

FILL FILL_1__1750_ (
);

FILL FILL_1__1330_ (
);

FILL FILL_3__1256_ (
);

OAI21X1 _1185_ (
    .A(_62_),
    .B(_271_),
    .C(_290_),
    .Y(_291_)
);

FILL FILL_1__967_ (
);

FILL FILL_0__1645_ (
);

FILL FILL_0__1225_ (
);

FILL FILL_1__1806_ (
);

FILL FILL_0__989_ (
);

FILL FILL_3__1485_ (
);

FILL FILL_0__1454_ (
);

FILL FILL_0__1034_ (
);

FILL FILL_2__983_ (
);

FILL FILL_3__925_ (
);

FILL FILL_0__1683_ (
);

FILL FILL_0__1263_ (
);

FILL FILL_1__1424_ (
);

FILL FILL_1__1004_ (
);

OAI21X1 _1699_ (
    .A(ABCmd_i_2_bF$buf0),
    .B(BI[2]),
    .C(_825_),
    .Y(_885_)
);

OAI21X1 _1279_ (
    .A(_56_),
    .B(_700_),
    .C(_384_),
    .Y(_9_)
);

FILL FILL_0__1739_ (
);

FILL FILL_0__1319_ (
);

FILL FILL_0__1492_ (
);

FILL FILL_0__1072_ (
);

FILL FILL_3__963_ (
);

FILL FILL_1__1653_ (
);

FILL FILL_1__1233_ (
);

FILL FILL_3__1579_ (
);

FILL FILL_3__1159_ (
);

AOI22X1 _1088_ (
    .A(_128_),
    .B(_135_),
    .C(_192_),
    .D(_193_),
    .Y(_194_)
);

FILL FILL_2__1722_ (
);

FILL FILL_2__1302_ (
);

FILL FILL_0__1548_ (
);

FILL FILL_0__1128_ (
);

FILL FILL_1__1709_ (
);

XNOR2X1 _1720_ (
    .A(_723_),
    .B(_733_),
    .Y(_734_)
);

NAND2X1 _1300_ (
    .A(AI[2]),
    .B(BI[7]),
    .Y(_405_)
);

FILL FILL_1__1462_ (
);

FILL FILL_1__1042_ (
);

FILL FILL_3__1388_ (
);

FILL FILL_2__1531_ (
);

FILL FILL_2__1111_ (
);

FILL FILL_0__1777_ (
);

FILL FILL_0__1357_ (
);

FILL FILL_3__1600_ (
);

FILL FILL_1__1518_ (
);

FILL FILL_1__1691_ (
);

FILL FILL_1__1271_ (
);

FILL FILL_2__1760_ (
);

FILL FILL_2__1340_ (
);

FILL FILL_0__1586_ (
);

FILL FILL_0__1166_ (
);

FILL FILL_0__913_ (
);

NOR2X1 _916_ (
    .A(LoadA_i),
    .B(_26_),
    .Y(_33_)
);

FILL FILL_1__1747_ (
);

FILL FILL_1__1327_ (
);

FILL FILL_1__1080_ (
);

FILL FILL_2__1816_ (
);

FILL FILL_0__1395_ (
);

NAND2X1 _1814_ (
    .A(_818_),
    .B(_820_),
    .Y(_821_)
);

FILL FILL_1__1556_ (
);

FILL FILL_1__1136_ (
);

FILL FILL_2__1205_ (
);

DFFSR _1623_ (
    .D(_15_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(_886_[6])
);

OAI21X1 _1203_ (
    .A(_265_),
    .B(_286_),
    .C(_285_),
    .Y(_309_)
);

FILL FILL_0__951_ (
);

AND2X2 _954_ (
    .A(BI_4_bF$buf2),
    .B(AI[1]),
    .Y(_60_)
);

FILL FILL_1__1785_ (
);

FILL FILL_1__1365_ (
);

FILL FILL_2__1434_ (
);

FILL FILL_2__1014_ (
);

FILL FILL_3__1503_ (
);

NOR2X1 _1432_ (
    .A(_535_),
    .B(_25_),
    .Y(_536_)
);

AOI21X1 _1012_ (
    .A(_102_),
    .B(_103_),
    .C(_101_),
    .Y(_118_)
);

FILL FILL_1__1594_ (
);

FILL FILL_1__1174_ (
);

FILL FILL_2__1663_ (
);

FILL FILL_2__1243_ (
);

FILL FILL_0__1489_ (
);

FILL FILL_0__1069_ (
);

FILL FILL_3__1312_ (
);

OAI21X1 _1661_ (
    .A(_828_),
    .B(_847_),
    .C(_845_),
    .Y(_848_)
);

AND2X2 _1241_ (
    .A(_332_),
    .B(_337_),
    .Y(_347_)
);

NOR2X1 _992_ (
    .A(_71_),
    .B(_97_),
    .Y(_98_)
);

FILL FILL_2__1719_ (
);

FILL FILL_0__1701_ (
);

FILL FILL_2__1472_ (
);

FILL FILL_2__1052_ (
);

FILL FILL_0__1298_ (
);

OAI21X1 _1717_ (
    .A(_844_),
    .B(_731_),
    .C(_729_),
    .Y(_732_)
);

FILL FILL_3__1541_ (
);

FILL FILL_1__1459_ (
);

FILL FILL_1__1039_ (
);

NAND3X1 _1470_ (
    .A(_516_),
    .B(_518_),
    .C(_572_),
    .Y(_573_)
);

AND2X2 _1050_ (
    .A(_155_),
    .B(_152_),
    .Y(_156_)
);

FILL FILL_0__1510_ (
);

FILL FILL_2__1528_ (
);

FILL FILL_2__1108_ (
);

FILL FILL_2__1281_ (
);

NAND3X1 _1526_ (
    .A(_25_),
    .B(_627_),
    .C(_626_),
    .Y(_628_)
);

NAND3X1 _1106_ (
    .A(_211_),
    .B(_210_),
    .C(_209_),
    .Y(_212_)
);

FILL FILL_3__1770_ (
);

FILL FILL_1__1688_ (
);

FILL FILL_1__1268_ (
);

FILL FILL_2__1757_ (
);

FILL FILL_2__1337_ (
);

FILL FILL_2__1090_ (
);

FILL FILL_3__1406_ (
);

OAI21X1 _1755_ (
    .A(_763_),
    .B(_753_),
    .C(_762_),
    .Y(_766_)
);

NAND2X1 _1335_ (
    .A(_432_),
    .B(_413_),
    .Y(_440_)
);

FILL FILL_1__1497_ (
);

FILL FILL_1__1077_ (
);

FILL FILL_2__904_ (
);

FILL FILL_2__1566_ (
);

FILL FILL_2__1146_ (
);

INVX1 _1564_ (
    .A(_645_),
    .Y(_664_)
);

INVX1 _1144_ (
    .A(_65_),
    .Y(_250_)
);

FILL FILL_0__892_ (
);

FILL FILL_1__926_ (
);

NOR2X1 _895_ (
    .A(state[2]),
    .B(_703_),
    .Y(_704_)
);

FILL FILL_0__1604_ (
);

FILL FILL_2__1795_ (
);

FILL FILL_2__1375_ (
);

FILL FILL_0__948_ (
);

FILL FILL_3__1024_ (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_2_BUFX2_insert17 (
);

FILL FILL_2_BUFX2_insert18 (
);

FILL FILL_2_BUFX2_insert19 (
);

NAND2X1 _1793_ (
    .A(_734_),
    .B(_801_),
    .Y(_802_)
);

OAI21X1 _1373_ (
    .A(_405_),
    .B(_410_),
    .C(_476_),
    .Y(_477_)
);

FILL FILL_0__1413_ (
);

FILL FILL_2__942_ (
);

FILL FILL_2__1184_ (
);

AOI21X1 _1429_ (
    .A(_292_),
    .B(_296_),
    .C(_294_),
    .Y(_533_)
);

NAND3X1 _1009_ (
    .A(_105_),
    .B(_112_),
    .C(_114_),
    .Y(_115_)
);

FILL FILL_3__1673_ (
);

FILL FILL_3__1253_ (
);

INVX1 _1182_ (
    .A(_278_),
    .Y(_288_)
);

FILL FILL_1__964_ (
);

FILL FILL_0__1642_ (
);

FILL FILL_0__1222_ (
);

FILL FILL_1__1803_ (
);

FILL FILL_3__1309_ (
);

OAI21X1 _1658_ (
    .A(_841_),
    .B(_843_),
    .C(_845_),
    .Y(_846_)
);

XNOR2X1 _1238_ (
    .A(_188_),
    .B(_340_),
    .Y(_344_)
);

FILL FILL_0__986_ (
);

FILL FILL_3__1482_ (
);

FILL FILL_3__1062_ (
);

INVX1 _989_ (
    .A(_94_),
    .Y(_95_)
);

FILL FILL_0__1451_ (
);

FILL FILL_2__1469_ (
);

FILL FILL_0__1031_ (
);

FILL FILL_2__1049_ (
);

FILL FILL_2__980_ (
);

FILL FILL_3__1538_ (
);

OAI21X1 _1467_ (
    .A(_561_),
    .B(_566_),
    .C(_544_),
    .Y(_570_)
);

OAI21X1 _1047_ (
    .A(_58_),
    .B(_149_),
    .C(_146_),
    .Y(_153_)
);

FILL FILL_3__1291_ (
);

FILL FILL_0__1507_ (
);

FILL FILL_2__1698_ (
);

FILL FILL_0__1680_ (
);

FILL FILL_2__1278_ (
);

FILL FILL_0__1260_ (
);

FILL FILL_1__1421_ (
);

FILL FILL_1__1001_ (
);

FILL FILL_3__1767_ (
);

NOR2X1 _1696_ (
    .A(ABCmd_i[0]),
    .B(_881_),
    .Y(_882_)
);

OAI21X1 _1276_ (
    .A(ACC[0]),
    .B(ABCmd_i[7]),
    .C(_715_),
    .Y(_382_)
);

FILL FILL_0__1736_ (
);

FILL FILL_0__1316_ (
);

FILL FILL_2__1087_ (
);

FILL FILL_3__960_ (
);

FILL FILL_1__1650_ (
);

FILL FILL_1__1230_ (
);

FILL FILL_3__1156_ (
);

AOI21X1 _1085_ (
    .A(_190_),
    .B(_187_),
    .C(_181_),
    .Y(_191_)
);

FILL FILL_0__1545_ (
);

FILL FILL_0__1125_ (
);

FILL FILL_1__1706_ (
);

FILL FILL_0__889_ (
);

FILL FILL_3__1385_ (
);

FILL FILL_0__1774_ (
);

FILL FILL_0__1354_ (
);

FILL FILL_1__1515_ (
);

FILL FILL_2__939_ (
);

FILL FILL_0__1583_ (
);

FILL FILL_0__1163_ (
);

FILL FILL_0__910_ (
);

OAI21X1 _913_ (
    .A(LoadA_i),
    .B(LoadB_i),
    .C(_26_),
    .Y(_30_)
);

FILL FILL_1__1744_ (
);

FILL FILL_1__1324_ (
);

NAND2X1 _1599_ (
    .A(AI[3]),
    .B(_705__bF$buf0),
    .Y(_694_)
);

NAND3X1 _1179_ (
    .A(_262_),
    .B(_282_),
    .C(_284_),
    .Y(_285_)
);

FILL FILL_2__1813_ (
);

FILL FILL_0__1639_ (
);

FILL FILL_0__1219_ (
);

FILL FILL_0__1392_ (
);

NAND3X1 _1811_ (
    .A(_800_),
    .B(_817_),
    .C(_797_),
    .Y(_818_)
);

FILL FILL_1__1553_ (
);

FILL FILL_1__1133_ (
);

FILL FILL_3__1479_ (
);

FILL FILL_3__1059_ (
);

FILL FILL_2__1202_ (
);

FILL FILL_0__1448_ (
);

FILL FILL_0__1028_ (
);

FILL FILL_2__977_ (
);

DFFSR _1620_ (
    .D(_12_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf2),
    .Q(_886_[3])
);

NAND3X1 _1200_ (
    .A(_281_),
    .B(_305_),
    .C(_304_),
    .Y(_306_)
);

INVX1 _951_ (
    .A(AI[0]),
    .Y(_57_)
);

FILL FILL_1__1782_ (
);

FILL FILL_1__1362_ (
);

FILL FILL_3__1288_ (
);

FILL FILL_1__999_ (
);

FILL FILL_2__1431_ (
);

FILL FILL_2__1011_ (
);

FILL FILL_0__1677_ (
);

FILL FILL_0__1257_ (
);

FILL FILL_3__1500_ (
);

FILL FILL_1__1418_ (
);

FILL FILL_1__1591_ (
);

FILL FILL_1__1171_ (
);

FILL FILL_2__1660_ (
);

FILL FILL_2__1240_ (
);

FILL FILL_0__1486_ (
);

FILL FILL_0__1066_ (
);

FILL FILL_3__957_ (
);

FILL FILL_1__1647_ (
);

FILL FILL_1__1227_ (
);

FILL FILL_2__1716_ (
);

FILL FILL_0__1295_ (
);

OAI21X1 _1714_ (
    .A(_728_),
    .B(_727_),
    .C(_724_),
    .Y(_729_)
);

FILL FILL_1__1456_ (
);

FILL FILL_1__1036_ (
);

FILL FILL_2__1525_ (
);

FILL FILL_2__1105_ (
);

AOI22X1 _1523_ (
    .A(_611_),
    .B(_613_),
    .C(_624_),
    .D(_622_),
    .Y(_625_)
);

NAND3X1 _1103_ (
    .A(_193_),
    .B(_192_),
    .C(_208_),
    .Y(_209_)
);

FILL FILL_1__1685_ (
);

FILL FILL_1__1265_ (
);

FILL FILL_2__1754_ (
);

FILL FILL_2__1334_ (
);

FILL FILL_0__907_ (
);

FILL FILL_3__1823_ (
);

FILL FILL_3__1403_ (
);

FILL FILL93750x58650 (
);

INVX1 _1752_ (
    .A(_763_),
    .Y(_764_)
);

OAI21X1 _1332_ (
    .A(_436_),
    .B(_433_),
    .C(_411_),
    .Y(_437_)
);

FILL FILL_1__1494_ (
);

FILL FILL_1__1074_ (
);

FILL FILL_2__901_ (
);

FILL FILL_2__1563_ (
);

FILL FILL_2__1143_ (
);

FILL FILL_0__1389_ (
);

NAND3X1 _1808_ (
    .A(ABCmd_i[6]),
    .B(_804_),
    .C(AN),
    .Y(_815_)
);

FILL FILL_3__1212_ (
);

NAND2X1 _1561_ (
    .A(_638_),
    .B(_647_),
    .Y(_661_)
);

INVX1 _1141_ (
    .A(_246_),
    .Y(_247_)
);

FILL FILL_1__923_ (
);

INVX1 _892_ (
    .A(_701_),
    .Y(_887_)
);

FILL FILL_0__1601_ (
);

FILL FILL_2__1792_ (
);

FILL FILL_2__1372_ (
);

FILL FILL_0__1198_ (
);

DFFSR _1617_ (
    .D(_9_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(_886_[0])
);

FILL FILL_0__945_ (
);

FILL FILL_3__1441_ (
);

NAND2X1 _948_ (
    .A(BI[7]),
    .B(_32__bF$buf3),
    .Y(_55_)
);

FILL FILL_1__1779_ (
);

FILL FILL_1__1359_ (
);

NAND3X1 _1790_ (
    .A(_775_),
    .B(_799_),
    .C(_798_),
    .Y(_800_)
);

AOI21X1 _1370_ (
    .A(_375_),
    .B(_459_),
    .C(_470_),
    .Y(_474_)
);

FILL FILL_2__1428_ (
);

FILL FILL_0__1410_ (
);

FILL FILL_2__1008_ (
);

FILL FILL_2__1181_ (
);

OAI21X1 _1426_ (
    .A(_525_),
    .B(_529_),
    .C(ABCmd_i[7]),
    .Y(_530_)
);

OAI21X1 _1006_ (
    .A(_58_),
    .B(_109_),
    .C(_60_),
    .Y(_112_)
);

FILL FILL_3__1670_ (
);

FILL FILL_1__1588_ (
);

FILL FILL_1__1168_ (
);

FILL FILL_1__961_ (
);

FILL FILL_2__1657_ (
);

FILL FILL_2__1237_ (
);

FILL FILL_1__1800_ (
);

FILL FILL_3__1306_ (
);

AOI21X1 _1655_ (
    .A(BI_0_bF$buf3),
    .B(ABCmd_i_2_bF$buf0),
    .C(_842_),
    .Y(_843_)
);

XOR2X1 _1235_ (
    .A(_188_),
    .B(_340_),
    .Y(_341_)
);

FILL FILL_0__983_ (
);

AOI22X1 _986_ (
    .A(BI_0_bF$buf1),
    .B(AI_5_bF$buf3),
    .C(BI_1_bF$buf0),
    .D(AI[4]),
    .Y(_92_)
);

FILL FILL_1__1397_ (
);

FILL FILL_2__1466_ (
);

FILL FILL_2__1046_ (
);

FILL FILL_3__1535_ (
);

OAI21X1 _1464_ (
    .A(_561_),
    .B(_566_),
    .C(_565_),
    .Y(_567_)
);

NAND2X1 _1044_ (
    .A(BI_4_bF$buf2),
    .B(AI[2]),
    .Y(_150_)
);

FILL FILL_0__1504_ (
);

FILL FILL_2__1695_ (
);

FILL FILL_2__1275_ (
);

FILL FILL_3__1764_ (
);

NAND3X1 _1693_ (
    .A(AI[2]),
    .B(BI[2]),
    .C(_831_),
    .Y(_879_)
);

NOR2X1 _1273_ (
    .A(_378_),
    .B(_715_),
    .Y(_379_)
);

FILL FILL_0__1733_ (
);

FILL FILL_0__1313_ (
);

FILL FILL_2__1084_ (
);

AOI21X1 _1749_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[5]),
    .C(_760_),
    .Y(_761_)
);

NOR2X1 _1329_ (
    .A(_343_),
    .B(_341_),
    .Y(_434_)
);

FILL FILL_3__1153_ (
);

FILL FILL94350x43050 (
);

NAND2X1 _1082_ (
    .A(BI_1_bF$buf3),
    .B(\u_ALU.AI7 ),
    .Y(_188_)
);

FILL FILL_0__1542_ (
);

FILL FILL_0__1122_ (
);

FILL FILL_1__1703_ (
);

FILL FILL_3__1209_ (
);

NAND3X1 _1558_ (
    .A(_613_),
    .B(_647_),
    .C(_611_),
    .Y(_658_)
);

NAND3X1 _1138_ (
    .A(_230_),
    .B(_236_),
    .C(_179_),
    .Y(_244_)
);

FILL FILL_3__1382_ (
);

INVX1 _889_ (
    .A(state[2]),
    .Y(_699_)
);

FILL FILL_2__1789_ (
);

FILL FILL_0__1771_ (
);

FILL FILL_2__1369_ (
);

FILL FILL_0__1351_ (
);

FILL FILL_1__1512_ (
);

FILL FILL_3__1438_ (
);

NAND2X1 _1787_ (
    .A(_796_),
    .B(_786_),
    .Y(_797_)
);

AOI22X1 _1367_ (
    .A(_361_),
    .B(_374_),
    .C(_453_),
    .D(_450_),
    .Y(_471_)
);

FILL FILL_3__1191_ (
);

FILL FILL_0__1827_ (
);

FILL FILL_0__1407_ (
);

FILL FILL_2__936_ (
);

FILL FILL_0__1580_ (
);

FILL FILL_2__1598_ (
);

FILL FILL_2__1178_ (
);

FILL FILL_0__1160_ (
);

OAI21X1 _910_ (
    .A(_714_),
    .B(_25_),
    .C(_27_),
    .Y(_28_)
);

FILL FILL_1__1741_ (
);

FILL FILL_1__1321_ (
);

FILL FILL_3__1667_ (
);

OAI21X1 _1596_ (
    .A(_42_),
    .B(_705__bF$buf2),
    .C(_692_),
    .Y(_18_)
);

INVX1 _1176_ (
    .A(_281_),
    .Y(_282_)
);

FILL FILL_1__958_ (
);

FILL FILL_2__1810_ (
);

FILL FILL_0__1636_ (
);

FILL FILL_0__1216_ (
);

FILL FILL_1__1550_ (
);

FILL FILL_1__1130_ (
);

FILL FILL_3__1056_ (
);

FILL FILL_0__1445_ (
);

FILL FILL_0__1025_ (
);

FILL FILL_2__974_ (
);

FILL FILL_1__1606_ (
);

FILL FILL_3__1285_ (
);

FILL FILL_1__996_ (
);

FILL FILL_0__1674_ (
);

FILL FILL_0__1254_ (
);

FILL FILL94050x78150 (
);

FILL FILL_1__1415_ (
);

FILL FILL_0__1483_ (
);

FILL FILL_0__1063_ (
);

FILL FILL_3__954_ (
);

FILL FILL_1__1644_ (
);

FILL FILL_1__1224_ (
);

INVX1 _1499_ (
    .A(_556_),
    .Y(_601_)
);

NAND2X1 _1079_ (
    .A(BI[2]),
    .B(AI_5_bF$buf2),
    .Y(_185_)
);

FILL FILL_2__1713_ (
);

FILL FILL_0__1539_ (
);

FILL FILL_0__1119_ (
);

FILL FILL_0__1292_ (
);

NAND2X1 _1711_ (
    .A(AI[3]),
    .B(_725_),
    .Y(_726_)
);

FILL FILL_1__1453_ (
);

FILL FILL_1__1033_ (
);

FILL FILL_3__1799_ (
);

FILL FILL_3__1379_ (
);

FILL FILL_2__1522_ (
);

FILL FILL_2__1102_ (
);

FILL FILL_0__1768_ (
);

FILL FILL_0__1348_ (
);

FILL FILL_1__1509_ (
);

FILL FILL92850x4050 (
);

OAI21X1 _1520_ (
    .A(_524_),
    .B(_577_),
    .C(_621_),
    .Y(_622_)
);

AND2X2 _1100_ (
    .A(_205_),
    .B(_202_),
    .Y(_206_)
);

FILL FILL_3__992_ (
);

FILL FILL_1__1682_ (
);

FILL FILL_1__1262_ (
);

FILL FILL_3__1188_ (
);

FILL FILL_1__899_ (
);

FILL FILL_2__1751_ (
);

FILL FILL_2__1331_ (
);

FILL FILL_0__1577_ (
);

FILL FILL_0__1157_ (
);

FILL FILL_0__904_ (
);

FILL FILL_3__1820_ (
);

INVX1 _907_ (
    .A(_715_),
    .Y(_25_)
);

FILL FILL_1__1738_ (
);

FILL FILL_1__1318_ (
);

FILL FILL_1__1491_ (
);

FILL FILL_1__1071_ (
);

FILL FILL_2__1807_ (
);

FILL FILL_2__1560_ (
);

FILL FILL_2__1140_ (
);

FILL FILL_0__1386_ (
);

AOI21X1 _1805_ (
    .A(_766_),
    .B(_812_),
    .C(_811_),
    .Y(_813_)
);

FILL FILL_1__1547_ (
);

FILL FILL_1__1127_ (
);

FILL FILL_1__920_ (
);

FILL FILL_0__1195_ (
);

DFFSR _1614_ (
    .D(_6_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(BI[5])
);

FILL FILL_0__942_ (
);

NAND2X1 _945_ (
    .A(BI[6]),
    .B(_32__bF$buf1),
    .Y(_53_)
);

FILL FILL_1__1776_ (
);

FILL FILL_1__1356_ (
);

FILL FILL_2__1425_ (
);

FILL FILL_2__1005_ (
);

OAI21X1 _1423_ (
    .A(_396_),
    .B(_526_),
    .C(_475_),
    .Y(_527_)
);

INVX1 _1003_ (
    .A(AI[2]),
    .Y(_109_)
);

FILL FILL_1__1585_ (
);

FILL FILL_1__1165_ (
);

FILL FILL_2__1654_ (
);

FILL FILL_2__1234_ (
);

FILL FILL_3__1723_ (
);

FILL FILL_3__1303_ (
);

NAND2X1 _1652_ (
    .A(AI[1]),
    .B(ABCmd_i[5]),
    .Y(_840_)
);

NAND2X1 _1232_ (
    .A(_337_),
    .B(_332_),
    .Y(_338_)
);

FILL FILL_0__980_ (
);

OAI21X1 _983_ (
    .A(_68_),
    .B(_78_),
    .C(_72_),
    .Y(_89_)
);

FILL FILL_1__1394_ (
);

FILL FILL_2__1463_ (
);

FILL FILL_2__1043_ (
);

FILL FILL_0__1289_ (
);

AOI22X1 _1708_ (
    .A(_884_),
    .B(_721_),
    .C(_877_),
    .D(_722_),
    .Y(_723_)
);

FILL FILL_3__1532_ (
);

FILL FILL_3__1112_ (
);

NAND3X1 _1461_ (
    .A(_562_),
    .B(_563_),
    .C(_544_),
    .Y(_564_)
);

AND2X2 _1041_ (
    .A(BI_3_bF$buf3),
    .B(AI[3]),
    .Y(_147_)
);

FILL FILL_0__1501_ (
);

FILL FILL_2__1519_ (
);

FILL FILL_2__1692_ (
);

FILL FILL_2__1272_ (
);

FILL FILL_0__1098_ (
);

AOI22X1 _1517_ (
    .A(_573_),
    .B(_618_),
    .C(_616_),
    .D(_474_),
    .Y(_619_)
);

FILL FILL_3__989_ (
);

FILL FILL_3__1341_ (
);

FILL FILL_1__1679_ (
);

FILL FILL_1__1259_ (
);

NOR2X1 _1690_ (
    .A(_857_),
    .B(_855_),
    .Y(_876_)
);

AND2X2 _1270_ (
    .A(_371_),
    .B(_375_),
    .Y(_376_)
);

FILL FILL_2__1748_ (
);

FILL FILL_0__1730_ (
);

FILL FILL_0__1310_ (
);

FILL FILL_2__1328_ (
);

FILL FILL_2__1081_ (
);

FILL FILL_3__1817_ (
);

OAI21X1 _1746_ (
    .A(AI_5_bF$buf0),
    .B(_755_),
    .C(_835_),
    .Y(_758_)
);

NAND3X1 _1326_ (
    .A(_430_),
    .B(_429_),
    .C(_428_),
    .Y(_431_)
);

FILL FILL_3__1570_ (
);

FILL FILL_1__1488_ (
);

FILL FILL_1__1068_ (
);

FILL FILL_2__1557_ (
);

FILL FILL_2__1137_ (
);

FILL FILL_3_BUFX2_insert21 (
);

FILL FILL_3_BUFX2_insert22 (
);

FILL FILL_3_BUFX2_insert24 (
);

FILL FILL_3_BUFX2_insert25 (
);

FILL FILL_3_BUFX2_insert27 (
);

FILL FILL_3_BUFX2_insert29 (
);

FILL FILL_1__1700_ (
);

FILL FILL_3__1206_ (
);

AOI21X1 _1555_ (
    .A(_653_),
    .B(_655_),
    .C(_712_),
    .Y(_656_)
);

AOI21X1 _1135_ (
    .A(_239_),
    .B(_240_),
    .C(_238_),
    .Y(_241_)
);

FILL FILL_1__917_ (
);

FILL FILL_1__1297_ (
);

FILL FILL_2_CLKBUF1_insert8 (
);

FILL FILL_2_CLKBUF1_insert9 (
);

FILL FILL_2__1786_ (
);

FILL FILL_2__1366_ (
);

FILL FILL_0__939_ (
);

FILL FILL_3__1435_ (
);

AOI21X1 _1784_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[7]),
    .C(_793_),
    .Y(_794_)
);

AOI22X1 _1364_ (
    .A(_385_),
    .B(_712_),
    .C(_463_),
    .D(_468_),
    .Y(_10_)
);

FILL FILL_0__1824_ (
);

FILL FILL_0__1404_ (
);

FILL FILL_2__933_ (
);

FILL FILL_2__1595_ (
);

FILL FILL_2__1175_ (
);

FILL FILL_3__1664_ (
);

NAND2X1 _1593_ (
    .A(AI[0]),
    .B(_705__bF$buf2),
    .Y(_691_)
);

OAI21X1 _1173_ (
    .A(_81_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

FILL FILL_1__955_ (
);

FILL FILL_0__1213_ (
);

INVX1 _1649_ (
    .A(AI[0]),
    .Y(_837_)
);

AOI22X1 _1229_ (
    .A(AI_5_bF$buf2),
    .B(BI_3_bF$buf0),
    .C(BI_4_bF$buf1),
    .D(AI[4]),
    .Y(_335_)
);

FILL FILL_0__977_ (
);

FILL FILL_3__1053_ (
);

FILL FILL_0__1442_ (
);

FILL FILL_0__1022_ (
);

FILL FILL_2__971_ (
);

FILL FILL_3__913_ (
);

FILL FILL_1__1603_ (
);

FILL FILL_3__1529_ (
);

FILL FILL_3__1109_ (
);

AOI21X1 _1458_ (
    .A(_552_),
    .B(_554_),
    .C(_560_),
    .Y(_561_)
);

NAND2X1 _1038_ (
    .A(BI[5]),
    .B(AI[1]),
    .Y(_144_)
);

FILL FILL_3__1282_ (
);

FILL FILL_1__993_ (
);

FILL FILL_2__1689_ (
);

FILL FILL_0__1671_ (
);

FILL FILL_0__1251_ (
);

FILL FILL_2__1269_ (
);

FILL FILL_1__1412_ (
);

FILL FILL_3__1338_ (
);

NAND2X1 _1687_ (
    .A(_871_),
    .B(_873_),
    .Y(_874_)
);

NAND3X1 _1267_ (
    .A(_367_),
    .B(_369_),
    .C(_368_),
    .Y(_373_)
);

FILL FILL_3__1091_ (
);

FILL FILL_0__1727_ (
);

FILL FILL_0__1307_ (
);

FILL FILL_2__1498_ (
);

FILL FILL_0__1480_ (
);

FILL FILL_2__1078_ (
);

FILL FILL_0__1060_ (
);

FILL FILL_1__1641_ (
);

FILL FILL_1__1221_ (
);

FILL FILL_3__1567_ (
);

OAI21X1 _1496_ (
    .A(_130_),
    .B(_597_),
    .C(_595_),
    .Y(_598_)
);

NAND3X1 _1076_ (
    .A(BI_0_bF$buf0),
    .B(\u_ALU.AI7 ),
    .C(_127_),
    .Y(_182_)
);

FILL FILL_2__1710_ (
);

FILL FILL_0__1536_ (
);

FILL FILL_0__1116_ (
);

FILL FILL_1__1450_ (
);

FILL FILL_1__1030_ (
);

FILL FILL_3__1796_ (
);

FILL FILL_0__1765_ (
);

FILL FILL_0__1345_ (
);

FILL FILL_1__1506_ (
);

FILL FILL_3__1185_ (
);

FILL FILL_1__896_ (
);

FILL FILL_0__1574_ (
);

FILL FILL_0__1154_ (
);

FILL FILL_0__901_ (
);

OAI21X1 _904_ (
    .A(state[1]),
    .B(state[0]),
    .C(_699_),
    .Y(_713_)
);

FILL FILL_1__1735_ (
);

FILL FILL_1__1315_ (
);

FILL FILL_2__1804_ (
);

FILL FILL_0__1383_ (
);

NOR2X1 _1802_ (
    .A(_837_),
    .B(_835_),
    .Y(_810_)
);

FILL FILL_1__1544_ (
);

FILL FILL_1__1124_ (
);

AND2X2 _1399_ (
    .A(_486_),
    .B(_489_),
    .Y(_503_)
);

FILL FILL_0__1439_ (
);

FILL FILL_0__1019_ (
);

FILL FILL_2__968_ (
);

FILL FILL_0__1192_ (
);

DFFSR _1611_ (
    .D(_3_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf3),
    .Q(BI[2])
);

NAND2X1 _942_ (
    .A(BI[5]),
    .B(_32__bF$buf2),
    .Y(_51_)
);

FILL FILL_1__1773_ (
);

FILL FILL_1__1353_ (
);

FILL FILL_3__1699_ (
);

FILL FILL_3__1279_ (
);

FILL FILL_2__1422_ (
);

FILL FILL_2__1002_ (
);

FILL FILL_0__1668_ (
);

FILL FILL_0__1248_ (
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf1)
);

FILL FILL_1__1409_ (
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf0)
);

NAND2X1 _1420_ (
    .A(_523_),
    .B(_520_),
    .Y(_524_)
);

INVX1 _1000_ (
    .A(_105_),
    .Y(_106_)
);

FILL FILL_3__892_ (
);

FILL FILL_1__1582_ (
);

FILL FILL_1__1162_ (
);

FILL FILL_3__1088_ (
);

FILL FILL_2__1651_ (
);

FILL FILL_2__1231_ (
);

FILL FILL_0__1477_ (
);

FILL FILL_0__1057_ (
);

FILL FILL_3__1720_ (
);

FILL FILL_1__1638_ (
);

FILL FILL_1__1218_ (
);

OAI21X1 _980_ (
    .A(_82_),
    .B(_81_),
    .C(_85_),
    .Y(_86_)
);

FILL FILL_1__1391_ (
);

FILL FILL_2__1707_ (
);

FILL FILL_2__1460_ (
);

FILL FILL_2__1040_ (
);

FILL FILL_0__1286_ (
);

INVX1 _1705_ (
    .A(_716_),
    .Y(_720_)
);

FILL FILL_1__1447_ (
);

FILL FILL_1__1027_ (
);

FILL FILL_2__1516_ (
);

FILL FILL_0__1095_ (
);

NOR2X1 _1514_ (
    .A(_577_),
    .B(_524_),
    .Y(_616_)
);

FILL FILL_3__986_ (
);

FILL FILL_1__1676_ (
);

FILL FILL_1__1256_ (
);

FILL FILL_2__1745_ (
);

FILL FILL_2__1325_ (
);

FILL FILL_3__1814_ (
);

AND2X2 _1743_ (
    .A(_831_),
    .B(BI[5]),
    .Y(_755_)
);

NAND3X1 _1323_ (
    .A(_415_),
    .B(_424_),
    .C(_425_),
    .Y(_428_)
);

FILL FILL_1__1485_ (
);

FILL FILL_1__1065_ (
);

FILL FILL_2__1554_ (
);

FILL FILL_2__1134_ (
);

FILL FILL_3__1203_ (
);

OAI21X1 _1552_ (
    .A(_652_),
    .B(_308_),
    .C(ABCmd_i[7]),
    .Y(_653_)
);

AOI21X1 _1132_ (
    .A(_162_),
    .B(_171_),
    .C(_174_),
    .Y(_238_)
);

FILL FILL_1__914_ (
);

FILL FILL_1__1294_ (
);

FILL FILL_2__1783_ (
);

FILL FILL_2__1363_ (
);

FILL FILL_0__1189_ (
);

OAI21X1 _1608_ (
    .A(_54_),
    .B(_705__bF$buf3),
    .C(_698_),
    .Y(_24_)
);

FILL FILL_0__936_ (
);

FILL FILL_3__1432_ (
);

FILL FILL_3__1012_ (
);

NAND2X1 _939_ (
    .A(BI_4_bF$buf0),
    .B(_32__bF$buf0),
    .Y(_49_)
);

OAI21X1 _1781_ (
    .A(\u_ALU.AI7 ),
    .B(_788_),
    .C(_835_),
    .Y(_791_)
);

OAI21X1 _1361_ (
    .A(_271_),
    .B(_293_),
    .C(ABCmd_i[7]),
    .Y(_466_)
);

FILL FILL_0__1821_ (
);

FILL FILL_2__1419_ (
);

FILL FILL_0__1401_ (
);

FILL FILL_2__930_ (
);

FILL FILL_2__1592_ (
);

FILL FILL_2__1172_ (
);

AOI21X1 _1417_ (
    .A(_437_),
    .B(_441_),
    .C(_404_),
    .Y(_521_)
);

FILL FILL_3__889_ (
);

FILL FILL_3__1241_ (
);

FILL FILL_1__1579_ (
);

FILL FILL_1__1159_ (
);

OAI21X1 _1590_ (
    .A(_54_),
    .B(_687_),
    .C(_688_),
    .Y(_689_)
);

OAI21X1 _1170_ (
    .A(_249_),
    .B(_66_),
    .C(_65_),
    .Y(_276_)
);

FILL FILL_1__952_ (
);

FILL FILL_2__1648_ (
);

FILL FILL_2__1228_ (
);

FILL FILL_0__1210_ (
);

FILL FILL_3__1717_ (
);

AOI22X1 _1646_ (
    .A(BI_0_bF$buf3),
    .B(_833_),
    .C(_830_),
    .D(_832_),
    .Y(_834_)
);

NAND3X1 _1226_ (
    .A(_327_),
    .B(_329_),
    .C(_331_),
    .Y(_332_)
);

FILL FILL_0__974_ (
);

FILL FILL_3__1470_ (
);

INVX2 _977_ (
    .A(BI_4_bF$buf2),
    .Y(_83_)
);

FILL FILL_1__1388_ (
);

FILL FILL_2__1457_ (
);

FILL FILL_2__1037_ (
);

FILL FILL_3__910_ (
);

FILL FILL_1__1600_ (
);

FILL FILL_3__1106_ (
);

INVX1 _1455_ (
    .A(BI[5]),
    .Y(_558_)
);

OAI21X1 _1035_ (
    .A(_137_),
    .B(_136_),
    .C(_134_),
    .Y(_141_)
);

FILL FILL_1__1197_ (
);

FILL FILL_1__990_ (
);

FILL FILL_2__1686_ (
);

FILL FILL_2__1266_ (
);

FILL FILL_3__1335_ (
);

AOI22X1 _1684_ (
    .A(_841_),
    .B(_864_),
    .C(_870_),
    .D(_827_),
    .Y(_871_)
);

AOI21X1 _1264_ (
    .A(_368_),
    .B(_369_),
    .C(_367_),
    .Y(_370_)
);

FILL FILL_0__1724_ (
);

FILL FILL_0__1304_ (
);

FILL FILL94350x58650 (
);

FILL FILL_2__1495_ (
);

FILL FILL_2__1075_ (
);

FILL FILL_3__1564_ (
);

OAI21X1 _1493_ (
    .A(_167_),
    .B(_557_),
    .C(_594_),
    .Y(_595_)
);

OAI21X1 _1073_ (
    .A(_170_),
    .B(_173_),
    .C(_166_),
    .Y(_179_)
);

FILL FILL_0__1533_ (
);

FILL FILL_0__1113_ (
);

OAI21X1 _1549_ (
    .A(_638_),
    .B(_620_),
    .C(_647_),
    .Y(_650_)
);

NAND2X1 _1129_ (
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

FILL FILL_3__1793_ (
);

FILL FILL_0__1762_ (
);

FILL FILL_0__1342_ (
);

FILL FILL_1__1503_ (
);

FILL FILL_3__1429_ (
);

FILL FILL_3__1009_ (
);

AND2X2 _1778_ (
    .A(_831_),
    .B(BI[7]),
    .Y(_788_)
);

OAI21X1 _1358_ (
    .A(_462_),
    .B(_461_),
    .C(_388_),
    .Y(_463_)
);

FILL FILL_3__1182_ (
);

FILL FILL_0__1818_ (
);

FILL FILL_1__893_ (
);

FILL FILL_2__927_ (
);

FILL FILL_2__1589_ (
);

FILL FILL_0__1571_ (
);

FILL FILL_2__1169_ (
);

FILL FILL_0__1151_ (
);

OAI21X1 _901_ (
    .A(_706_),
    .B(_709_),
    .C(LoadB_i),
    .Y(_710_)
);

FILL FILL_1__1732_ (
);

FILL FILL_1__1312_ (
);

FILL FILL_3__1238_ (
);

NAND2X1 _1587_ (
    .A(_389_),
    .B(_247_),
    .Y(_686_)
);

NAND2X1 _1167_ (
    .A(AI[0]),
    .B(BI[2]),
    .Y(_273_)
);

FILL FILL_1__949_ (
);

FILL FILL_2__1801_ (
);

FILL FILL_0__1207_ (
);

FILL FILL_0__1380_ (
);

FILL FILL_2__1398_ (
);

FILL FILL_1__1541_ (
);

FILL FILL_1__1121_ (
);

FILL FILL_3__1467_ (
);

NAND3X1 _1396_ (
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_500_)
);

FILL FILL_0__1436_ (
);

FILL FILL_0__1016_ (
);

FILL FILL_2__965_ (
);

FILL FILL_3__907_ (
);

FILL FILL_1__1770_ (
);

FILL FILL_1__1350_ (
);

FILL FILL_3__1696_ (
);

FILL FILL_1__987_ (
);

FILL FILL_0__1665_ (
);

FILL FILL_0__1245_ (
);

FILL FILL_1__1826_ (
);

FILL FILL_1__1406_ (
);

FILL FILL_3__1085_ (
);

FILL FILL_0__1474_ (
);

FILL FILL_0__1054_ (
);

FILL FILL_1__1215_ (
);

FILL FILL_2__1704_ (
);

FILL FILL_0__1283_ (
);

OAI21X1 _1702_ (
    .A(_884_),
    .B(_716_),
    .C(_717_),
    .Y(_718_)
);

FILL FILL_1__1444_ (
);

FILL FILL_1__1024_ (
);

OAI21X1 _1299_ (
    .A(_325_),
    .B(_403_),
    .C(_358_),
    .Y(_404_)
);

FILL FILL_2__1513_ (
);

FILL FILL_0__1759_ (
);

FILL FILL_0__1339_ (
);

FILL FILL_0__1092_ (
);

NAND3X1 _1511_ (
    .A(_612_),
    .B(_609_),
    .C(_607_),
    .Y(_613_)
);

FILL FILL_3__983_ (
);

FILL FILL_1__1673_ (
);

FILL FILL_1__1253_ (
);

FILL FILL_2__1742_ (
);

FILL FILL_2__1322_ (
);

FILL FILL_0__1568_ (
);

FILL FILL_0__1148_ (
);

FILL FILL_1__1729_ (
);

FILL FILL_1__1309_ (
);

INVX1 _1740_ (
    .A(_749_),
    .Y(_752_)
);

OAI21X1 _1320_ (
    .A(_130_),
    .B(_83_),
    .C(_418_),
    .Y(_425_)
);

FILL FILL_1__1482_ (
);

FILL FILL_1__1062_ (
);

FILL FILL_2__1551_ (
);

FILL FILL_2__1131_ (
);

FILL FILL_0__1797_ (
);

FILL FILL_0__1377_ (
);

FILL FILL_1__1538_ (
);

FILL FILL_1__1118_ (
);

FILL FILL_1__911_ (
);

FILL FILL_1__1291_ (
);

FILL FILL_2__1607_ (
);

FILL FILL_2__1780_ (
);

FILL FILL_2__1360_ (
);

FILL FILL_0__1186_ (
);

NAND2X1 _1605_ (
    .A(AI[6]),
    .B(_705__bF$buf1),
    .Y(_697_)
);

FILL FILL_0__933_ (
);

NAND2X1 _936_ (
    .A(BI_3_bF$buf2),
    .B(_32__bF$buf1),
    .Y(_47_)
);

FILL FILL_1__1767_ (
);

FILL FILL_1__1347_ (
);

FILL FILL_2__1416_ (
);

NAND3X1 _1414_ (
    .A(_477_),
    .B(_516_),
    .C(_517_),
    .Y(_518_)
);

FILL FILL_1__1576_ (
);

FILL FILL_1__1156_ (
);

FILL FILL_2__1645_ (
);

FILL FILL_2__1225_ (
);

FILL FILL_3__1714_ (
);

INVX2 _1643_ (
    .A(ABCmd_i[0]),
    .Y(_831_)
);

OAI21X1 _1223_ (
    .A(_130_),
    .B(_58_),
    .C(_328_),
    .Y(_329_)
);

FILL FILL_0__971_ (
);

NAND3X1 _974_ (
    .A(_79_),
    .B(_67_),
    .C(_76_),
    .Y(_80_)
);

FILL FILL_1__1385_ (
);

FILL FILL_2__1454_ (
);

FILL FILL_2__1034_ (
);

FILL FILL_3__1103_ (
);

NAND2X1 _1452_ (
    .A(AI[6]),
    .B(BI_4_bF$buf3),
    .Y(_555_)
);

OAI21X1 _1032_ (
    .A(_137_),
    .B(_136_),
    .C(_133_),
    .Y(_138_)
);

FILL FILL_0_CLKBUF1_insert8 (
);

FILL FILL_0_CLKBUF1_insert9 (
);

FILL FILL_1__1194_ (
);

FILL FILL_2__1683_ (
);

FILL FILL_2__1263_ (
);

FILL FILL_0__1089_ (
);

NAND2X1 _1508_ (
    .A(_609_),
    .B(_607_),
    .Y(_610_)
);

FILL FILL_3__1752_ (
);

FILL FILL_3__1332_ (
);

AOI21X1 _1681_ (
    .A(_832_),
    .B(_837_),
    .C(ABCmd_i[5]),
    .Y(_868_)
);

INVX1 _1261_ (
    .A(_313_),
    .Y(_367_)
);

FILL FILL_2__1739_ (
);

FILL FILL_0__1721_ (
);

FILL FILL_2__1319_ (
);

FILL FILL_0__1301_ (
);

FILL FILL_2__1492_ (
);

FILL FILL_2__1072_ (
);

OAI21X1 _1737_ (
    .A(_746_),
    .B(_748_),
    .C(_749_),
    .Y(_750_)
);

AOI21X1 _1317_ (
    .A(_419_),
    .B(_421_),
    .C(_416_),
    .Y(_422_)
);

FILL FILL_3__1561_ (
);

FILL FILL_3__1141_ (
);

FILL FILL_1__1479_ (
);

FILL FILL_1__1059_ (
);

INVX1 _1490_ (
    .A(\u_ALU.AI7 ),
    .Y(_592_)
);

NAND3X1 _1070_ (
    .A(_172_),
    .B(_175_),
    .C(_124_),
    .Y(_176_)
);

FILL FILL_0__1530_ (
);

FILL FILL_2__1548_ (
);

FILL FILL_2__1128_ (
);

FILL FILL_0__1110_ (
);

XOR2X1 _1546_ (
    .A(_639_),
    .B(_646_),
    .Y(_647_)
);

AOI21X1 _1126_ (
    .A(_207_),
    .B(_212_),
    .C(_180_),
    .Y(_232_)
);

FILL FILL_1__908_ (
);

FILL FILL_3__1370_ (
);

FILL FILL_1__1288_ (
);

FILL FILL_2__1777_ (
);

FILL FILL_2__1357_ (
);

FILL FILL_1__1500_ (
);

FILL FILL_3__1006_ (
);

NAND2X1 _1775_ (
    .A(_777_),
    .B(_785_),
    .Y(ACC[6])
);

NAND2X1 _1355_ (
    .A(_459_),
    .B(_454_),
    .Y(_460_)
);

FILL FILL_1__1097_ (
);

FILL FILL_0__1815_ (
);

FILL FILL_1__890_ (
);

FILL FILL_2__924_ (
);

FILL FILL_2__1586_ (
);

FILL FILL_2__1166_ (
);

FILL FILL_3__1235_ (
);

NAND3X1 _1584_ (
    .A(_641_),
    .B(_642_),
    .C(_666_),
    .Y(_683_)
);

NAND3X1 _1164_ (
    .A(_251_),
    .B(_250_),
    .C(_64_),
    .Y(_270_)
);

FILL FILL_1__946_ (
);

FILL FILL_0__1204_ (
);

FILL FILL_2__1395_ (
);

FILL FILL_0__968_ (
);

FILL FILL_3__1464_ (
);

OAI21X1 _1393_ (
    .A(_493_),
    .B(_494_),
    .C(_496_),
    .Y(_497_)
);

FILL FILL_0__1433_ (
);

FILL FILL_0__1013_ (
);

FILL FILL_2__962_ (
);

FILL FILL_3__904_ (
);

NAND3X1 _1449_ (
    .A(_546_),
    .B(_549_),
    .C(_551_),
    .Y(_552_)
);

NAND3X1 _1029_ (
    .A(_132_),
    .B(_134_),
    .C(_128_),
    .Y(_135_)
);

FILL FILL_3__1693_ (
);

FILL FILL_1__984_ (
);

FILL FILL_0__1662_ (
);

FILL FILL_0__1242_ (
);

FILL FILL_1__1823_ (
);

FILL FILL_1__1403_ (
);

FILL FILL_3__1749_ (
);

FILL FILL_3__1329_ (
);

MUX2X1 _1678_ (
    .A(ABCmd_i[1]),
    .B(_836_),
    .S(ABCmd_i[0]),
    .Y(_865_)
);

AOI21X1 _1258_ (
    .A(_351_),
    .B(_355_),
    .C(_325_),
    .Y(_364_)
);

FILL FILL_3__1082_ (
);

FILL FILL_0__1718_ (
);

FILL FILL_2__1489_ (
);

FILL FILL_0__1471_ (
);

FILL FILL_2__1069_ (
);

FILL FILL_0__1051_ (
);

FILL FILL_3__942_ (
);

FILL FILL_1__1212_ (
);

FILL FILL_3__1558_ (
);

FILL FILL_3__1138_ (
);

INVX1 _1487_ (
    .A(_886_[4]),
    .Y(_589_)
);

AOI21X1 _1067_ (
    .A(_165_),
    .B(_164_),
    .C(_163_),
    .Y(_173_)
);

FILL FILL_2__1701_ (
);

FILL FILL_0__1527_ (
);

FILL FILL_0__1107_ (
);

FILL FILL_0__1280_ (
);

FILL FILL_2__1298_ (
);

FILL FILL_1__1441_ (
);

FILL FILL_1__1021_ (
);

FILL FILL_3__1367_ (
);

OAI21X1 _1296_ (
    .A(_315_),
    .B(_323_),
    .C(_319_),
    .Y(_401_)
);

FILL FILL_2__1510_ (
);

FILL FILL_0__1756_ (
);

FILL FILL_0__1336_ (
);

FILL FILL_1__1670_ (
);

FILL FILL_1__1250_ (
);

FILL FILL_3__1596_ (
);

FILL FILL_0__1565_ (
);

FILL FILL_0__1145_ (
);

FILL FILL_1__1726_ (
);

FILL FILL_1__1306_ (
);

FILL FILL_0_BUFX2_insert30 (
);

FILL FILL_0_BUFX2_insert31 (
);

FILL FILL_0_BUFX2_insert32 (
);

FILL FILL_0_BUFX2_insert33 (
);

FILL FILL_0_BUFX2_insert34 (
);

FILL FILL_0_BUFX2_insert35 (
);

FILL FILL_0_BUFX2_insert36 (
);

FILL FILL_0_BUFX2_insert37 (
);

FILL FILL92850x58650 (
);

FILL FILL_0_BUFX2_insert38 (
);

FILL FILL_0_BUFX2_insert39 (
);

FILL FILL_0__1794_ (
);

FILL FILL_0__1374_ (
);

FILL FILL_1__1535_ (
);

FILL FILL_1__1115_ (
);

FILL FILL_2__1604_ (
);

FILL FILL_2__959_ (
);

FILL FILL_0__1183_ (
);

OAI21X1 _1602_ (
    .A(_48_),
    .B(_705__bF$buf3),
    .C(_695_),
    .Y(_21_)
);

FILL FILL_0__930_ (
);

NAND2X1 _933_ (
    .A(BI[2]),
    .B(_32__bF$buf0),
    .Y(_45_)
);

FILL FILL_1__1764_ (
);

FILL FILL_1__1344_ (
);

NAND3X1 _1199_ (
    .A(_61_),
    .B(_122_),
    .C(_261_),
    .Y(_305_)
);

FILL FILL_2__1413_ (
);

FILL FILL_0__1659_ (
);

FILL FILL_0__1239_ (
);

NAND3X1 _1411_ (
    .A(_478_),
    .B(_514_),
    .C(_508_),
    .Y(_515_)
);

FILL FILL_1__1573_ (
);

FILL FILL_1__1153_ (
);

BUFX2 BUFX2_insert40 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf1)
);

BUFX2 BUFX2_insert41 (
    .A(ABCmd_i[2]),
    .Y(ABCmd_i_2_bF$buf0)
);

FILL FILL_2__1642_ (
);

FILL FILL_2__1222_ (
);

FILL FILL_0__1468_ (
);

FILL FILL_0__1048_ (
);

FILL FILL_2__997_ (
);

FILL FILL_3__939_ (
);

FILL FILL_1__1209_ (
);

INVX1 _1640_ (
    .A(_827_),
    .Y(_828_)
);

AOI21X1 _1220_ (
    .A(_206_),
    .B(_209_),
    .C(_194_),
    .Y(_326_)
);

NOR2X1 _971_ (
    .A(_70_),
    .B(_71_),
    .Y(_77_)
);

FILL FILL_1__1382_ (
);

FILL FILL_2__1451_ (
);

FILL FILL_2__1031_ (
);

FILL FILL_0__1697_ (
);

FILL FILL_0__1277_ (
);

FILL FILL_3__1520_ (
);

FILL FILL_1__1438_ (
);

FILL FILL_1__1018_ (
);

FILL FILL_1__1191_ (
);

FILL FILL_2__1507_ (
);

FILL FILL_2__1680_ (
);

FILL FILL_2__1260_ (
);

FILL FILL_0__1086_ (
);

OAI21X1 _1505_ (
    .A(_604_),
    .B(_606_),
    .C(_591_),
    .Y(_607_)
);

FILL FILL_1__1667_ (
);

FILL FILL_1__1247_ (
);

FILL FILL_2__1736_ (
);

FILL FILL_2__1316_ (
);

OAI21X1 _1734_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_4_bF$buf0),
    .C(_825_),
    .Y(_747_)
);

NAND2X1 _1314_ (
    .A(_417_),
    .B(_418_),
    .Y(_419_)
);

FILL FILL_1__1476_ (
);

FILL FILL_1__1056_ (
);

FILL FILL_2__1545_ (
);

FILL FILL_2__1125_ (
);

NAND2X1 _1543_ (
    .A(_643_),
    .B(_642_),
    .Y(_644_)
);

NAND2X1 _1123_ (
    .A(_228_),
    .B(_225_),
    .Y(_229_)
);

FILL FILL_1__905_ (
);

FILL FILL_1__1285_ (
);

FILL FILL_2__1774_ (
);

FILL FILL_2__1354_ (
);

FILL FILL_0__927_ (
);

FILL FILL_3__1003_ (
);

AOI22X1 _1772_ (
    .A(_759_),
    .B(_782_),
    .C(_781_),
    .D(_764_),
    .Y(_783_)
);

NAND3X1 _1352_ (
    .A(_401_),
    .B(_442_),
    .C(_449_),
    .Y(_457_)
);

FILL FILL_1__1094_ (
);

FILL FILL_0__1812_ (
);

FILL FILL_2__921_ (
);

FILL FILL_2__1583_ (
);

FILL FILL_2__1163_ (
);

NAND2X1 _1408_ (
    .A(_498_),
    .B(_504_),
    .Y(_512_)
);

FILL FILL_3__1652_ (
);

FILL FILL_3__1232_ (
);

AOI22X1 _1581_ (
    .A(_657_),
    .B(_712_),
    .C(_673_),
    .D(_680_),
    .Y(_15_)
);

OAI21X1 _1161_ (
    .A(_241_),
    .B(_237_),
    .C(_177_),
    .Y(_267_)
);

FILL FILL_1__943_ (
);

FILL FILL_2__1639_ (
);

FILL FILL_0__1201_ (
);

FILL FILL_2__1219_ (
);

FILL FILL93750x82050 (
);

FILL FILL_2__1392_ (
);

INVX4 _1637_ (
    .A(ABCmd_i[3]),
    .Y(_825_)
);

NOR2X1 _1217_ (
    .A(_317_),
    .B(_318_),
    .Y(_323_)
);

FILL FILL_0__965_ (
);

FILL FILL_3__1461_ (
);

FILL FILL_3__1041_ (
);

INVX1 _968_ (
    .A(AI[4]),
    .Y(_74_)
);

FILL FILL_1__1799_ (
);

FILL FILL_1__1379_ (
);

NAND2X1 _1390_ (
    .A(\u_ALU.AI7 ),
    .B(BI_4_bF$buf3),
    .Y(_494_)
);

FILL FILL_2__1448_ (
);

FILL FILL_0__1430_ (
);

FILL FILL_2__1028_ (
);

FILL FILL_0__1010_ (
);

FILL FILL_3__1517_ (
);

NAND2X1 _1446_ (
    .A(_547_),
    .B(_548_),
    .Y(_549_)
);

OAI21X1 _1026_ (
    .A(_129_),
    .B(_130_),
    .C(_131_),
    .Y(_132_)
);

FILL FILL_3__1270_ (
);

FILL FILL_1__1188_ (
);

FILL FILL_1__981_ (
);

FILL FILL_2__1677_ (
);

FILL FILL_2__1257_ (
);

FILL FILL_1__1820_ (
);

FILL FILL_1__1400_ (
);

FILL FILL_3__1746_ (
);

INVX1 _1675_ (
    .A(_842_),
    .Y(_862_)
);

NAND3X1 _1255_ (
    .A(_356_),
    .B(_360_),
    .C(_314_),
    .Y(_361_)
);

FILL FILL_0__1715_ (
);

FILL FILL_2__1486_ (
);

FILL FILL_2__1066_ (
);

FILL FILL_3__1135_ (
);

OAI21X1 _1484_ (
    .A(_54_),
    .B(_585_),
    .C(_586_),
    .Y(_587_)
);

XNOR2X1 _1064_ (
    .A(_169_),
    .B(_168_),
    .Y(_170_)
);

FILL FILL_0__1524_ (
);

FILL FILL_0__1104_ (
);

FILL FILL_2__1295_ (
);

FILL FILL_3__1364_ (
);

OAI21X1 _1293_ (
    .A(_397_),
    .B(_396_),
    .C(_375_),
    .Y(_398_)
);

FILL FILL_0__1753_ (
);

FILL FILL_0__1333_ (
);

AOI21X1 _1769_ (
    .A(_779_),
    .B(ACC[3]),
    .C(_739_),
    .Y(_780_)
);

NAND3X1 _1349_ (
    .A(_450_),
    .B(_453_),
    .C(_400_),
    .Y(_454_)
);

FILL FILL_3__1593_ (
);

FILL FILL_0__1809_ (
);

FILL FILL_2__918_ (
);

FILL FILL_0__1562_ (
);

FILL FILL_0__1142_ (
);

FILL FILL_1__1723_ (
);

FILL FILL_1__1303_ (
);

FILL FILL_3__1649_ (
);

FILL FILL_3__1229_ (
);

NOR2X1 _1578_ (
    .A(ABCmd_i[7]),
    .B(ACC[6]),
    .Y(_678_)
);

NAND3X1 _1158_ (
    .A(_170_),
    .B(_162_),
    .C(_166_),
    .Y(_264_)
);

FILL FILL_0__1791_ (
);

FILL FILL_0__1371_ (
);

FILL FILL_2__1389_ (
);

FILL FILL_1__1532_ (
);

FILL FILL_1__1112_ (
);

FILL FILL_3__1458_ (
);

FILL FILL_3__1038_ (
);

OR2X2 _1387_ (
    .A(_188_),
    .B(_340_),
    .Y(_491_)
);

FILL FILL_2__1601_ (
);

FILL FILL_0__1427_ (
);

FILL FILL_0__1007_ (
);

FILL FILL_2__956_ (
);

FILL FILL_0__1180_ (
);

FILL FILL_2__1198_ (
);

NAND2X1 _930_ (
    .A(BI_1_bF$buf2),
    .B(_32__bF$buf2),
    .Y(_43_)
);

FILL FILL_1__1761_ (
);

FILL FILL_1__1341_ (
);

FILL FILL_3__1267_ (
);

AOI21X1 _1196_ (
    .A(_280_),
    .B(_269_),
    .C(_279_),
    .Y(_302_)
);

FILL FILL_1__978_ (
);

FILL FILL_2__1410_ (
);

FILL FILL_0__1656_ (
);

FILL FILL_0__1236_ (
);

FILL FILL_1__1817_ (
);

FILL FILL_1__1570_ (
);

FILL FILL_1__1150_ (
);

FILL FILL_3__1496_ (
);

BUFX2 BUFX2_insert13 (
    .A(_705_),
    .Y(_705__bF$buf3)
);

BUFX2 BUFX2_insert14 (
    .A(_705_),
    .Y(_705__bF$buf2)
);

BUFX2 BUFX2_insert15 (
    .A(_705_),
    .Y(_705__bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .A(_705_),
    .Y(_705__bF$buf0)
);

BUFX2 BUFX2_insert17 (
    .A(_0_),
    .Y(_0__bF$buf4)
);

BUFX2 BUFX2_insert18 (
    .A(_0_),
    .Y(_0__bF$buf3)
);

BUFX2 BUFX2_insert19 (
    .A(_0_),
    .Y(_0__bF$buf2)
);

FILL FILL_0__1465_ (
);

FILL FILL_0__1045_ (
);

FILL FILL_2__994_ (
);

FILL FILL_3__936_ (
);

FILL FILL_1__1206_ (
);

FILL FILL_0__1694_ (
);

FILL FILL_0__1274_ (
);

FILL FILL_1__1435_ (
);

FILL FILL_1__1015_ (
);

FILL FILL_2__1504_ (
);

FILL FILL_0__1083_ (
);

NOR2X1 _1502_ (
    .A(_563_),
    .B(_603_),
    .Y(_604_)
);

FILL FILL_1__1664_ (
);

FILL FILL_1__1244_ (
);

NAND3X1 _1099_ (
    .A(_195_),
    .B(_203_),
    .C(_204_),
    .Y(_205_)
);

FILL FILL_2__1733_ (
);

FILL FILL_2__1313_ (
);

FILL FILL_0__1559_ (
);

FILL FILL_0__1139_ (
);

FILL FILL_3__1802_ (
);

AOI22X1 _1731_ (
    .A(_829_),
    .B(BI_4_bF$buf0),
    .C(_743_),
    .D(_830_),
    .Y(_744_)
);

INVX1 _1311_ (
    .A(_415_),
    .Y(_416_)
);

FILL FILL93750x4050 (
);

FILL FILL_1__1473_ (
);

FILL FILL_1__1053_ (
);

FILL FILL_3__1399_ (
);

FILL FILL_2__1542_ (
);

FILL FILL_2__1122_ (
);

FILL FILL_0__1788_ (
);

FILL FILL_0__1368_ (
);

FILL FILL_2__897_ (
);

FILL FILL_1__1529_ (
);

FILL FILL_1__1109_ (
);

NOR2X1 _1540_ (
    .A(_592_),
    .B(_597_),
    .Y(_641_)
);

NAND2X1 _1120_ (
    .A(_223_),
    .B(_221_),
    .Y(_226_)
);

FILL FILL_1__902_ (
);

FILL FILL_1__1282_ (
);

FILL FILL_2__1771_ (
);

FILL FILL_2__1351_ (
);

FILL FILL_0__1597_ (
);

FILL FILL_0__1177_ (
);

FILL FILL_0__924_ (
);

FILL FILL_3__1420_ (
);

NAND2X1 _927_ (
    .A(BI_0_bF$buf1),
    .B(_32__bF$buf2),
    .Y(_41_)
);

FILL FILL_1__1758_ (
);

FILL FILL_1__1338_ (
);

FILL FILL_1__1091_ (
);

FILL FILL_2__1827_ (
);

FILL FILL_2__1407_ (
);

FILL FILL_2__1580_ (
);

FILL FILL_2__1160_ (
);

BUFX2 _1825_ (
    .A(_886_[7]),
    .Y(ACC_o[7])
);

OAI21X1 _1405_ (
    .A(_411_),
    .B(_436_),
    .C(_439_),
    .Y(_509_)
);

FILL FILL_1__1567_ (
);

FILL FILL_1__1147_ (
);

FILL FILL_1__940_ (
);

FILL FILL_2__1636_ (
);

FILL FILL_2__1216_ (
);

DFFSR _1634_ (
    .D(_888_[1]),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf2),
    .Q(state[1])
);

OR2X2 _1214_ (
    .A(_318_),
    .B(_317_),
    .Y(_320_)
);

FILL FILL_0__962_ (
);

NAND2X1 _965_ (
    .A(BI_0_bF$buf2),
    .B(AI[4]),
    .Y(_71_)
);

FILL FILL_1__1796_ (
);

FILL FILL_1__1376_ (
);

FILL FILL_2__1445_ (
);

FILL FILL_2__1025_ (
);

FILL FILL_3__1514_ (
);

INVX1 _1443_ (
    .A(_545_),
    .Y(_546_)
);

INVX1 _1023_ (
    .A(BI_1_bF$buf3),
    .Y(_129_)
);

FILL FILL_1__1185_ (
);

FILL FILL_2__1674_ (
);

FILL FILL_2__1254_ (
);

FILL FILL_3__1743_ (
);

OAI21X1 _1672_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(_825_),
    .C(_858_),
    .Y(_859_)
);

NAND3X1 _1252_ (
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_358_)
);

FILL FILL_0__1712_ (
);

FILL FILL_2__1483_ (
);

FILL FILL_2__1063_ (
);

NAND2X1 _1728_ (
    .A(ABCmd_i[5]),
    .B(AI_5_bF$buf0),
    .Y(_741_)
);

AOI21X1 _1308_ (
    .A(_347_),
    .B(_349_),
    .C(_412_),
    .Y(_413_)
);

FILL FILL_3__1132_ (
);

NAND2X1 _1481_ (
    .A(_297_),
    .B(_583_),
    .Y(_584_)
);

INVX4 _1061_ (
    .A(BI[6]),
    .Y(_167_)
);

FILL FILL_0__1521_ (
);

FILL FILL_2__1539_ (
);

FILL FILL_0__1101_ (
);

FILL FILL_2__1119_ (
);

FILL FILL_2__1292_ (
);

FILL FILL_3__1608_ (
);

INVX1 _1537_ (
    .A(_613_),
    .Y(_638_)
);

NOR2X1 _1117_ (
    .A(_167_),
    .B(_113_),
    .Y(_223_)
);

FILL FILL_3__1781_ (
);

FILL FILL_3__1361_ (
);

FILL FILL_1__1699_ (
);

FILL FILL_1__1279_ (
);

OAI21X1 _1290_ (
    .A(_307_),
    .B(_394_),
    .C(_393_),
    .Y(_395_)
);

FILL FILL_0__1750_ (
);

FILL FILL_2__1768_ (
);

FILL FILL_0__1330_ (
);

FILL FILL_2__1348_ (
);

FILL FILL_3__1417_ (
);

NAND2X1 _1766_ (
    .A(_776_),
    .B(_766_),
    .Y(_777_)
);

NAND3X1 _1346_ (
    .A(_437_),
    .B(_441_),
    .C(_444_),
    .Y(_451_)
);

FILL FILL_3__1590_ (
);

FILL FILL_3__1170_ (
);

FILL FILL_1__1088_ (
);

FILL FILL_0__1806_ (
);

FILL FILL93750x35250 (
);

FILL FILL_2__915_ (
);

FILL FILL_2__1577_ (
);

FILL FILL_2__1157_ (
);

FILL FILL_1_CLKBUF1_insert10 (
);

FILL FILL_1_CLKBUF1_insert11 (
);

FILL FILL_1__1720_ (
);

FILL FILL_1_CLKBUF1_insert12 (
);

FILL FILL_1__1300_ (
);

FILL FILL_3__1646_ (
);

NOR2X1 _1575_ (
    .A(_307_),
    .B(_674_),
    .Y(_675_)
);

NAND3X1 _1155_ (
    .A(_260_),
    .B(_259_),
    .C(_258_),
    .Y(_261_)
);

FILL FILL_1__937_ (
);

FILL FILL_2__1386_ (
);

FILL FILL_0__959_ (
);

FILL FILL_3__1035_ (
);

NOR2X1 _1384_ (
    .A(_482_),
    .B(_483_),
    .Y(_488_)
);

FILL FILL_0__1424_ (
);

FILL FILL_0__1004_ (
);

FILL FILL_2__953_ (
);

FILL FILL_2__1195_ (
);

FILL FILL_3__1264_ (
);

INVX1 _1193_ (
    .A(_277_),
    .Y(_299_)
);

FILL FILL_1__975_ (
);

FILL FILL_0__1653_ (
);

FILL FILL_0__1233_ (
);

FILL FILL_1__1814_ (
);

OAI21X1 _1669_ (
    .A(ABCmd_i_2_bF$buf1),
    .B(BI_1_bF$buf2),
    .C(_825_),
    .Y(_856_)
);

OAI21X1 _1249_ (
    .A(_353_),
    .B(_354_),
    .C(_352_),
    .Y(_355_)
);

FILL FILL_0__997_ (
);

FILL FILL_3__1493_ (
);

FILL FILL_0__1709_ (
);

FILL FILL_0__1462_ (
);

FILL FILL_0__1042_ (
);

FILL FILL_2__991_ (
);

FILL FILL_3__933_ (
);

FILL FILL_1__1203_ (
);

OAI21X1 _1478_ (
    .A(_580_),
    .B(_579_),
    .C(ABCmd_i[7]),
    .Y(_581_)
);

NAND3X1 _1058_ (
    .A(_159_),
    .B(_158_),
    .C(_156_),
    .Y(_164_)
);

FILL FILL_0__1518_ (
);

FILL FILL_0__1691_ (
);

FILL FILL_0__1271_ (
);

FILL FILL_2__1289_ (
);

FILL FILL_1__1432_ (
);

FILL FILL_1__1012_ (
);

FILL FILL_3__1778_ (
);

FILL FILL_3__1358_ (
);

NAND3X1 _1287_ (
    .A(_122_),
    .B(_262_),
    .C(_391_),
    .Y(_392_)
);

FILL FILL_2__1501_ (
);

FILL FILL_0__1747_ (
);

FILL FILL_0__1327_ (
);

FILL FILL_1_BUFX2_insert40 (
);

FILL FILL_1_BUFX2_insert41 (
);

FILL FILL_0__1080_ (
);

FILL FILL_2__1098_ (
);

FILL FILL_3__971_ (
);

FILL FILL_1__1661_ (
);

FILL FILL_1__1241_ (
);

FILL FILL_3__1587_ (
);

FILL FILL_3__1167_ (
);

NAND3X1 _1096_ (
    .A(_196_),
    .B(_201_),
    .C(_199_),
    .Y(_202_)
);

FILL FILL_2__1730_ (
);

FILL FILL_2__1310_ (
);

FILL FILL_0__1556_ (
);

FILL FILL_0__1136_ (
);

FILL FILL_1__1717_ (
);

FILL FILL_1__1470_ (
);

FILL FILL_1__1050_ (
);

FILL FILL_3__1396_ (
);

FILL FILL_0__1785_ (
);

FILL FILL_0__1365_ (
);

FILL FILL_2__894_ (
);

FILL FILL_1__1526_ (
);

FILL FILL_1__1106_ (
);

FILL FILL_0__1594_ (
);

FILL FILL_0__1174_ (
);

FILL FILL_0__921_ (
);

OAI21X1 _924_ (
    .A(_26_),
    .B(_708_),
    .C(_39_),
    .Y(_888_[2])
);

FILL FILL_1__1755_ (
);

FILL FILL_1__1335_ (
);

FILL FILL_2__1824_ (
);

FILL FILL_2__1404_ (
);

BUFX2 _1822_ (
    .A(_886_[4]),
    .Y(ACC_o[4])
);

NAND2X1 _1402_ (
    .A(_504_),
    .B(_505_),
    .Y(_506_)
);

FILL FILL_1__1564_ (
);

FILL FILL_1__1144_ (
);

FILL FILL_2__1213_ (
);

FILL FILL_0__1459_ (
);

FILL FILL_0__1039_ (
);

FILL FILL_2__988_ (
);

FILL FILL_3__1702_ (
);

DFFSR _1631_ (
    .D(_23_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf1),
    .Q(AI[6])
);

NOR2X1 _1211_ (
    .A(_109_),
    .B(_167_),
    .Y(_317_)
);

NAND2X1 _962_ (
    .A(BI[2]),
    .B(AI[2]),
    .Y(_68_)
);

FILL FILL_1__1793_ (
);

FILL FILL_1__1373_ (
);

FILL FILL_3__1299_ (
);

FILL FILL_2__1442_ (
);

FILL FILL_2__1022_ (
);

FILL FILL_0__1688_ (
);

FILL FILL_0__1268_ (
);

FILL FILL_3__1511_ (
);

FILL FILL_1__1429_ (
);

FILL FILL_1__1009_ (
);

INVX1 _1440_ (
    .A(_542_),
    .Y(_543_)
);

OAI21X1 _1020_ (
    .A(_92_),
    .B(_94_),
    .C(_91_),
    .Y(_126_)
);

FILL FILL_1__1182_ (
);

FILL FILL_2__1671_ (
);

FILL FILL_2__1251_ (
);

FILL FILL_0__1497_ (
);

FILL FILL_0__1077_ (
);

FILL FILL_3__968_ (
);

FILL FILL_3__1320_ (
);

FILL FILL_1__1658_ (
);

FILL FILL_1__1238_ (
);

FILL FILL_2__1727_ (
);

FILL FILL_2__1307_ (
);

FILL FILL_2__1480_ (
);

FILL FILL_2__1060_ (
);

FILL FILL93450x58650 (
);

OAI21X1 _1725_ (
    .A(_733_),
    .B(_723_),
    .C(_732_),
    .Y(_739_)
);

XNOR2X1 _1305_ (
    .A(_409_),
    .B(_406_),
    .Y(_410_)
);

FILL FILL_1__1467_ (
);

FILL FILL_1__1047_ (
);

FILL FILL_2__1536_ (
);

FILL FILL_2__1116_ (
);

INVX1 _1534_ (
    .A(_886_[5]),
    .Y(_635_)
);

AOI22X1 _1114_ (
    .A(_107_),
    .B(_197_),
    .C(_151_),
    .D(_145_),
    .Y(_220_)
);

FILL FILL_1__1696_ (
);

FILL FILL_1__1276_ (
);

FILL FILL_2__1765_ (
);

FILL FILL_2__1345_ (
);

FILL FILL_0__918_ (
);

FILL FILL_3__1414_ (
);

AOI21X1 _1763_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[6]),
    .C(_773_),
    .Y(_774_)
);

AOI21X1 _1343_ (
    .A(_446_),
    .B(_447_),
    .C(_411_),
    .Y(_448_)
);

FILL FILL_1__1085_ (
);

FILL FILL_0__1803_ (
);

FILL FILL_2__912_ (
);

FILL FILL_2__1574_ (
);

FILL FILL_2__1154_ (
);

BUFX2 _1819_ (
    .A(_886_[1]),
    .Y(ACC_o[1])
);

FILL FILL_3__1643_ (
);

OAI21X1 _1572_ (
    .A(_662_),
    .B(_670_),
    .C(_671_),
    .Y(_672_)
);

AOI21X1 _1152_ (
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

FILL FILL_1__934_ (
);

FILL FILL_2__1383_ (
);

DFFSR _1628_ (
    .D(_20_),
    .S(vdd),
    .R(_0__bF$buf0),
    .CLK(clk_bF$buf4),
    .Q(AI[3])
);

OAI21X1 _1208_ (
    .A(_235_),
    .B(_231_),
    .C(_217_),
    .Y(_314_)
);

FILL FILL_0__956_ (
);

FILL FILL_3__1032_ (
);

NAND2X1 _959_ (
    .A(BI[2]),
    .B(AI[1]),
    .Y(_65_)
);

OR2X2 _1381_ (
    .A(_483_),
    .B(_482_),
    .Y(_485_)
);

FILL FILL_0__1421_ (
);

FILL FILL_2__1439_ (
);

FILL FILL_0__1001_ (
);

FILL FILL_2__1019_ (
);

FILL FILL_2__950_ (
);

FILL FILL_2__1192_ (
);

FILL FILL_3__1508_ (
);

OAI21X1 _1437_ (
    .A(_539_),
    .B(_715_),
    .C(_387_),
    .Y(_540_)
);

AOI21X1 _1017_ (
    .A(_121_),
    .B(_117_),
    .C(_88_),
    .Y(_123_)
);

FILL FILL_3__1681_ (
);

FILL FILL_3__1261_ (
);

FILL FILL_1__1599_ (
);

FILL FILL_1__1179_ (
);

OAI21X1 _1190_ (
    .A(_57_),
    .B(_295_),
    .C(_291_),
    .Y(_296_)
);

FILL FILL_1__972_ (
);

FILL FILL_2__1668_ (
);

FILL FILL_0__1650_ (
);

FILL FILL_0__1230_ (
);

FILL FILL_2__1248_ (
);

FILL FILL_1__1811_ (
);

FILL FILL_3__1317_ (
);

NOR2X1 _1666_ (
    .A(ABCmd_i[0]),
    .B(_852_),
    .Y(_853_)
);

OAI21X1 _1246_ (
    .A(_211_),
    .B(_191_),
    .C(_210_),
    .Y(_352_)
);

FILL FILL_0__994_ (
);

FILL FILL_3__1490_ (
);

FILL FILL_3__1070_ (
);

NAND3X1 _997_ (
    .A(_93_),
    .B(_94_),
    .C(_91_),
    .Y(_103_)
);

FILL FILL_0__1706_ (
);

FILL FILL_2__1477_ (
);

FILL FILL_2__1057_ (
);

FILL FILL_1__1200_ (
);

FILL FILL_3__1546_ (
);

NOR3X1 _1475_ (
    .A(_541_),
    .B(_577_),
    .C(_525_),
    .Y(_578_)
);

NAND3X1 _1055_ (
    .A(_160_),
    .B(_159_),
    .C(_158_),
    .Y(_161_)
);

FILL FILL_0__1515_ (
);

FILL FILL_2__1286_ (
);

FILL FILL_3__1775_ (
);

NAND3X1 _1284_ (
    .A(_176_),
    .B(_245_),
    .C(_242_),
    .Y(_389_)
);

FILL FILL_0__1744_ (
);

FILL FILL_0__1324_ (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_1_BUFX2_insert18 (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_2__1095_ (
);

FILL FILL_3__1164_ (
);

NAND2X1 _1093_ (
    .A(_197_),
    .B(_198_),
    .Y(_199_)
);

FILL FILL_2__909_ (
);

FILL FILL_0__1553_ (
);

FILL FILL_0__1133_ (
);

FILL FILL_1__1714_ (
);

NAND3X1 _1569_ (
    .A(_668_),
    .B(_663_),
    .C(_660_),
    .Y(_669_)
);

AOI21X1 _1149_ (
    .A(_254_),
    .B(_253_),
    .C(_252_),
    .Y(_255_)
);

FILL FILL_0__897_ (
);

FILL FILL94350x82050 (
);

FILL FILL_3__1393_ (
);

FILL FILL_0__1782_ (
);

FILL FILL_0__1362_ (
);

FILL FILL_2__891_ (
);

FILL FILL_1__1523_ (
);

FILL FILL_1__1103_ (
);

FILL FILL_3__1449_ (
);

NAND3X1 _1798_ (
    .A(_775_),
    .B(_796_),
    .C(_798_),
    .Y(_806_)
);

NOR2X1 _1378_ (
    .A(_74_),
    .B(_167_),
    .Y(_482_)
);

FILL FILL_0__1418_ (
);

FILL FILL_2__947_ (
);

FILL FILL_0__1591_ (
);

FILL FILL_2__1189_ (
);

FILL FILL_0__1171_ (
);

FILL FILL93750x85950 (
);

AOI22X1 _921_ (
    .A(_36_),
    .B(_33_),
    .C(_706_),
    .D(_34_),
    .Y(_37_)
);

FILL FILL_1__1752_ (
);

FILL FILL_1__1332_ (
);

FILL FILL_3__1678_ (
);

FILL FILL_3__1258_ (
);

NAND2X1 _1187_ (
    .A(AI[0]),
    .B(BI_1_bF$buf0),
    .Y(_293_)
);

FILL FILL_1__969_ (
);

FILL FILL_2__1821_ (
);

FILL FILL_2__1401_ (
);

FILL FILL_0__1647_ (
);

FILL FILL_0__1227_ (
);

FILL FILL_1__1808_ (
);

FILL FILL_1__1561_ (
);

FILL FILL_1__1141_ (
);

FILL FILL_3__1487_ (
);

FILL FILL_3__1067_ (
);

FILL FILL_2__1210_ (
);

FILL FILL_0__1456_ (
);

FILL FILL_0__1036_ (
);

FILL FILL_2__985_ (
);

FILL FILL_1__1790_ (
);

FILL FILL_1__1370_ (
);

FILL FILL_3__1296_ (
);

FILL FILL_0__1685_ (
);

FILL FILL_0__1265_ (
);

FILL FILL_1__1426_ (
);

FILL FILL_1__1006_ (
);

FILL FILL_0__1494_ (
);

FILL FILL_0__1074_ (
);

FILL FILL_3__965_ (
);

FILL FILL_1__1655_ (
);

FILL FILL_1__1235_ (
);

FILL FILL_2__1724_ (
);

FILL FILL_2__1304_ (
);

NAND3X1 _1722_ (
    .A(_872_),
    .B(_722_),
    .C(_861_),
    .Y(_736_)
);

NAND2X1 _1302_ (
    .A(BI_3_bF$buf0),
    .B(AI[4]),
    .Y(_407_)
);

FILL FILL_1__1464_ (
);

FILL FILL_1__1044_ (
);

FILL FILL_2__1533_ (
);

FILL FILL_2__1113_ (
);

FILL FILL_0__1779_ (
);

FILL FILL_0__1359_ (
);

OAI21X1 _1531_ (
    .A(_54_),
    .B(_631_),
    .C(_632_),
    .Y(_633_)
);

NAND3X1 _1111_ (
    .A(_215_),
    .B(_214_),
    .C(_216_),
    .Y(_217_)
);

FILL FILL_1__1693_ (
);

FILL FILL_1__1273_ (
);

FILL FILL_3__1199_ (
);

FILL FILL_2__1762_ (
);

FILL FILL_2__1342_ (
);

FILL FILL_0__1588_ (
);

FILL FILL_0__1168_ (
);

FILL FILL_0__915_ (
);

FILL FILL_3__1411_ (
);

OAI22X1 _918_ (
    .A(_33_),
    .B(_32__bF$buf3),
    .C(_705__bF$buf1),
    .D(_34_),
    .Y(_35_)
);

FILL FILL_1__1749_ (
);

FILL FILL_1__1329_ (
);

OAI21X1 _1760_ (
    .A(AI[6]),
    .B(_768_),
    .C(_835_),
    .Y(_771_)
);

AOI21X1 _1340_ (
    .A(_439_),
    .B(_440_),
    .C(_438_),
    .Y(_445_)
);

FILL FILL_1__1082_ (
);

FILL FILL_2__1818_ (
);

FILL FILL_0__1800_ (
);

FILL FILL_2__1571_ (
);

FILL FILL_2__1151_ (
);

FILL FILL_0__1397_ (
);

NAND3X1 _1816_ (
    .A(_818_),
    .B(_820_),
    .C(CO),
    .Y(_823_)
);

FILL FILL_3__1220_ (
);

FILL FILL_1__1558_ (
);

FILL FILL_1__1138_ (
);

FILL FILL_1__931_ (
);

FILL FILL_2__1207_ (
);

FILL FILL_2__1380_ (
);

DFFSR _1625_ (
    .D(_17_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf4),
    .Q(AI[0])
);

OAI21X1 _1205_ (
    .A(_268_),
    .B(_310_),
    .C(_247_),
    .Y(_311_)
);

FILL FILL_0__953_ (
);

NAND2X1 _956_ (
    .A(BI_1_bF$buf1),
    .B(AI[2]),
    .Y(_62_)
);

FILL FILL_1__1787_ (
);

FILL FILL_1__1367_ (
);

FILL FILL_2__1436_ (
);

FILL FILL_2__1016_ (
);

OAI21X1 _1434_ (
    .A(_712_),
    .B(_537_),
    .C(_469_),
    .Y(_11_)
);

NAND2X1 _1014_ (
    .A(_111_),
    .B(_115_),
    .Y(_120_)
);

FILL FILL_1__1596_ (
);

FILL FILL_1__1176_ (
);

FILL FILL_2__1665_ (
);

FILL FILL_2__1245_ (
);

FILL FILL_3__1314_ (
);

NAND3X1 _1663_ (
    .A(AI[1]),
    .B(BI_1_bF$buf2),
    .C(_831_),
    .Y(_850_)
);

NAND2X1 _1243_ (
    .A(_344_),
    .B(_339_),
    .Y(_349_)
);

FILL FILL_0__991_ (
);

NAND3X1 _994_ (
    .A(_96_),
    .B(_99_),
    .C(_89_),
    .Y(_100_)
);

FILL FILL_0__1703_ (
);

FILL FILL_2__1474_ (
);

FILL FILL_2__1054_ (
);

XOR2X1 _1719_ (
    .A(_723_),
    .B(_733_),
    .Y(ACC[3])
);

FILL FILL_3__1543_ (
);

OAI21X1 _1472_ (
    .A(_478_),
    .B(_574_),
    .C(_516_),
    .Y(_575_)
);

NAND3X1 _1052_ (
    .A(_142_),
    .B(_141_),
    .C(_140_),
    .Y(_158_)
);

FILL FILL_0__1512_ (
);

FILL FILL_2__1283_ (
);

OAI21X1 _1528_ (
    .A(_302_),
    .B(_282_),
    .C(_301_),
    .Y(_630_)
);

OAI21X1 _1108_ (
    .A(_160_),
    .B(_139_),
    .C(_159_),
    .Y(_214_)
);

FILL FILL_3__1772_ (
);

INVX1 _1281_ (
    .A(AN),
    .Y(_386_)
);

FILL FILL93750x7950 (
);

FILL FILL_0__1741_ (
);

FILL FILL_2__1759_ (
);

FILL FILL_0__1321_ (
);

FILL FILL_2__1339_ (
);

FILL FILL_2__1092_ (
);

FILL FILL_3__1408_ (
);

AND2X2 _1757_ (
    .A(_831_),
    .B(BI[6]),
    .Y(_768_)
);

NAND3X1 _1337_ (
    .A(_441_),
    .B(_437_),
    .C(_404_),
    .Y(_442_)
);

FILL FILL_3__1161_ (
);

FILL FILL_1__1499_ (
);

FILL FILL_1__1079_ (
);

FILL FILL93150x4050 (
);

INVX1 _1090_ (
    .A(_195_),
    .Y(_196_)
);

FILL FILL_2__906_ (
);

FILL FILL_0__1550_ (
);

FILL FILL_2__1568_ (
);

FILL FILL_2__1148_ (
);

FILL FILL_0__1130_ (
);

FILL FILL_1__1711_ (
);

FILL FILL_3__1217_ (
);

OAI21X1 _1566_ (
    .A(_602_),
    .B(_644_),
    .C(_665_),
    .Y(_666_)
);

AOI21X1 _1146_ (
    .A(_250_),
    .B(_251_),
    .C(_249_),
    .Y(_252_)
);

FILL FILL_0__894_ (
);

FILL FILL_1__928_ (
);

FILL FILL_3__1390_ (
);

INVX1 _897_ (
    .A(_705__bF$buf1),
    .Y(_706_)
);

FILL FILL_0__1606_ (
);

FILL FILL_2__1797_ (
);

FILL FILL_2__1377_ (
);

FILL FILL_1__1520_ (
);

FILL FILL_1__1100_ (
);

FILL FILL_3__1446_ (
);

FILL FILL_2_BUFX2_insert30 (
);

FILL FILL_2_BUFX2_insert31 (
);

FILL FILL_2_BUFX2_insert32 (
);

FILL FILL_2_BUFX2_insert33 (
);

FILL FILL_2_BUFX2_insert34 (
);

FILL FILL_2_BUFX2_insert35 (
);

FILL FILL_2_BUFX2_insert36 (
);

FILL FILL_2_BUFX2_insert37 (
);

FILL FILL_2_BUFX2_insert38 (
);

FILL FILL_2_BUFX2_insert39 (
);

NAND3X1 _1795_ (
    .A(_765_),
    .B(_777_),
    .C(_785_),
    .Y(_804_)
);

AOI21X1 _1375_ (
    .A(_438_),
    .B(_440_),
    .C(_433_),
    .Y(_479_)
);

FILL FILL_0__1415_ (
);

FILL FILL_2__944_ (
);

FILL FILL_2__1186_ (
);

FILL FILL_3__1675_ (
);

INVX1 _1184_ (
    .A(_274_),
    .Y(_290_)
);

FILL FILL_1__966_ (
);

FILL FILL_0__1644_ (
);

FILL FILL_0__1224_ (
);

FILL FILL_1__1805_ (
);

FILL FILL_0__988_ (
);

FILL FILL_3__1064_ (
);

FILL FILL_0__1453_ (
);

FILL FILL_0__1033_ (
);

FILL FILL_2__982_ (
);

NAND2X1 _1469_ (
    .A(_571_),
    .B(_568_),
    .Y(_572_)
);

NAND3X1 _1049_ (
    .A(_144_),
    .B(_153_),
    .C(_154_),
    .Y(_155_)
);

FILL FILL_3__1293_ (
);

FILL FILL_0__1509_ (
);

FILL FILL_0__1682_ (
);

FILL FILL_0__1262_ (
);

FILL FILL_1__1423_ (
);

FILL FILL_1__1003_ (
);

FILL FILL_3__1349_ (
);

OAI21X1 _1698_ (
    .A(_880_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

NAND2X1 _1278_ (
    .A(_700_),
    .B(_383_),
    .Y(_384_)
);

FILL FILL_0__1738_ (
);

FILL FILL_0__1318_ (
);

FILL FILL_0__1491_ (
);

FILL FILL_2__1089_ (
);

FILL FILL_0__1071_ (
);

FILL FILL_3__962_ (
);

FILL FILL_1__1652_ (
);

FILL FILL_1__1232_ (
);

FILL FILL94350x35250 (
);

FILL FILL_3__1158_ (
);

NAND3X1 _1087_ (
    .A(_184_),
    .B(_185_),
    .C(_182_),
    .Y(_193_)
);

FILL FILL_2__1721_ (
);

FILL FILL_2__1301_ (
);

FILL FILL_0__1547_ (
);

FILL FILL_0__1127_ (
);

FILL FILL_1__1708_ (
);

FILL FILL_1__1461_ (
);

FILL FILL_1__1041_ (
);

FILL FILL_3__1387_ (
);

FILL FILL_2__1530_ (
);

FILL FILL_2__1110_ (
);

FILL FILL_0__1776_ (
);

FILL FILL_0__1356_ (
);

FILL FILL_1__1517_ (
);

FILL FILL_1__1690_ (
);

FILL FILL_1__1270_ (
);

FILL FILL_3__1196_ (
);

FILL FILL_0__1585_ (
);

FILL FILL_0__1165_ (
);

FILL FILL_0__912_ (
);

NAND2X1 _915_ (
    .A(state[1]),
    .B(_707_),
    .Y(_32_)
);

FILL FILL_1__1746_ (
);

FILL FILL_1__1326_ (
);

FILL FILL_2__1815_ (
);

FILL FILL_0__1394_ (
);

NAND3X1 _1813_ (
    .A(_806_),
    .B(_819_),
    .C(_807_),
    .Y(_820_)
);

FILL FILL_1__1555_ (
);

FILL FILL_1__1135_ (
);

FILL FILL_2__1204_ (
);

FILL FILL_2__979_ (
);

DFFSR _1622_ (
    .D(_14_),
    .S(vdd),
    .R(_0__bF$buf1),
    .CLK(clk_bF$buf2),
    .Q(_886_[5])
);

INVX1 _1202_ (
    .A(_307_),
    .Y(_308_)
);

FILL FILL_0__950_ (
);

NOR2X1 _953_ (
    .A(_57_),
    .B(_58_),
    .Y(_59_)
);

FILL FILL_1__1784_ (
);

FILL FILL_1__1364_ (
);

FILL FILL_2__1433_ (
);

FILL FILL_2__1013_ (
);

FILL FILL_0__1679_ (
);

FILL FILL_0__1259_ (
);

NOR2X1 _1431_ (
    .A(ABCmd_i[7]),
    .B(ACC[2]),
    .Y(_535_)
);

NAND3X1 _1011_ (
    .A(_100_),
    .B(_104_),
    .C(_116_),
    .Y(_117_)
);

FILL FILL_1__1593_ (
);

FILL FILL_1__1173_ (
);

FILL FILL_3__1099_ (
);

FILL FILL_2__1662_ (
);

FILL FILL_2__1242_ (
);

FILL FILL_0__1488_ (
);

FILL FILL_0__1068_ (
);

FILL FILL_3__959_ (
);

FILL FILL_3__1731_ (
);

FILL FILL_3__1311_ (
);

FILL FILL_1__1649_ (
);

FILL FILL_1__1229_ (
);

NOR2X1 _1660_ (
    .A(_843_),
    .B(_841_),
    .Y(_847_)
);

NAND3X1 _1240_ (
    .A(_345_),
    .B(_338_),
    .C(_342_),
    .Y(_346_)
);

NAND2X1 _991_ (
    .A(BI_1_bF$buf0),
    .B(AI_5_bF$buf3),
    .Y(_97_)
);

FILL FILL_2__1718_ (
);

FILL FILL_0__1700_ (
);

FILL FILL_2__1471_ (
);

FILL FILL_2__1051_ (
);

FILL FILL_0__1297_ (
);

AOI21X1 _1716_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI_3_bF$buf2),
    .C(_730_),
    .Y(_731_)
);

FILL FILL_3__1540_ (
);

FILL FILL_3__1120_ (
);

FILL FILL_1__1458_ (
);

FILL FILL_1__1038_ (
);

FILL FILL_2__1527_ (
);

FILL FILL_2__1107_ (
);

FILL FILL_2__1280_ (
);

OR2X2 _1525_ (
    .A(ABCmd_i[7]),
    .B(CO),
    .Y(_627_)
);

NAND2X1 _1105_ (
    .A(_202_),
    .B(_205_),
    .Y(_211_)
);

FILL FILL_3__997_ (
);

FILL FILL_1__1687_ (
);

FILL FILL_1__1267_ (
);

FILL FILL_2__1756_ (
);

FILL FILL_2__1336_ (
);

FILL FILL_0__909_ (
);

FILL FILL_3__1825_ (
);

INVX1 _1754_ (
    .A(_765_),
    .Y(ACC[5])
);

NAND3X1 _1334_ (
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_439_)
);

FILL FILL_1__1496_ (
);

FILL FILL_1__1076_ (
);

FILL FILL_2__903_ (
);

FILL FILL_2__1565_ (
);

FILL FILL_2__1145_ (
);

FILL FILL_3__1214_ (
);

INVX1 _1563_ (
    .A(_662_),
    .Y(_663_)
);

NOR2X1 _1143_ (
    .A(_62_),
    .B(_63_),
    .Y(_249_)
);

FILL FILL_0__891_ (
);

FILL FILL_1__925_ (
);

INVX2 _894_ (
    .A(state[1]),
    .Y(_703_)
);

FILL FILL_0__1603_ (
);

FILL FILL_2__1794_ (
);

FILL FILL_2__1374_ (
);

DFFSR _1619_ (
    .D(_11_),
    .S(vdd),
    .R(_0__bF$buf2),
    .CLK(clk_bF$buf3),
    .Q(_886_[2])
);

FILL FILL_0__947_ (
);

FILL FILL_3__1443_ (
);

NOR2X1 _1792_ (
    .A(ACC[0]),
    .B(_737_),
    .Y(_801_)
);

NAND2X1 _1372_ (
    .A(_406_),
    .B(_409_),
    .Y(_476_)
);

FILL FILL_0__1412_ (
);

FILL FILL_2__941_ (
);

FILL FILL_2__1183_ (
);

NOR2X1 _1428_ (
    .A(_531_),
    .B(_715_),
    .Y(_532_)
);

OAI21X1 _1008_ (
    .A(_83_),
    .B(_113_),
    .C(_107_),
    .Y(_114_)
);

FILL FILL_3__1672_ (
);

NOR3X1 _1181_ (
    .A(_285_),
    .B(_265_),
    .C(_286_),
    .Y(_287_)
);

FILL FILL_1__963_ (
);

FILL FILL_2__1659_ (
);

FILL FILL_0__1641_ (
);

FILL FILL_0__1221_ (
);

FILL FILL_2__1239_ (
);

FILL FILL_1__1802_ (
);

FILL FILL_3__1728_ (
);

FILL FILL_3__1308_ (
);

OAI21X1 _1657_ (
    .A(_844_),
    .B(_843_),
    .C(_841_),
    .Y(_845_)
);

OAI21X1 _1237_ (
    .A(_183_),
    .B(_185_),
    .C(_182_),
    .Y(_343_)
);

FILL FILL_0__985_ (
);

FILL FILL_3__1061_ (
);

NAND2X1 _988_ (
    .A(BI[2]),
    .B(AI[3]),
    .Y(_94_)
);

FILL FILL_1__1399_ (
);

FILL FILL94050x58650 (
);

FILL FILL_0__1450_ (
);

FILL FILL_2__1468_ (
);

FILL FILL_0__1030_ (
);

FILL FILL_2__1048_ (
);

FILL FILL_3__921_ (
);

FILL FILL_3__1537_ (
);

FILL FILL_3__1117_ (
);

NAND3X1 _1466_ (
    .A(_563_),
    .B(_562_),
    .C(_565_),
    .Y(_569_)
);

NAND3X1 _1046_ (
    .A(_151_),
    .B(_145_),
    .C(_148_),
    .Y(_152_)
);

FILL FILL_3__1290_ (
);

FILL FILL_0__1506_ (
);

FILL FILL_2__1697_ (
);

FILL FILL_2__1277_ (
);

FILL FILL_1__1420_ (
);

FILL FILL_1__1000_ (
);

FILL FILL_3__1346_ (
);

INVX1 _1695_ (
    .A(BI[2]),
    .Y(_881_)
);

AOI21X1 _1275_ (
    .A(BI_0_bF$buf1),
    .B(AI[0]),
    .C(_54_),
    .Y(_381_)
);

FILL FILL_0__1735_ (
);

FILL FILL_0__1315_ (
);

FILL FILL_2__1086_ (
);

FILL FILL_3__1575_ (
);

OAI21X1 _1084_ (
    .A(_183_),
    .B(_189_),
    .C(_185_),
    .Y(_190_)
);

FILL FILL_0__1544_ (
);

FILL FILL_0__1124_ (
);

FILL FILL_1__1705_ (
);

FILL FILL94350x11850 (
);

FILL FILL_0__1773_ (
);

FILL FILL_0__1353_ (
);

FILL FILL_1__1514_ (
);

INVX1 _1789_ (
    .A(_796_),
    .Y(_799_)
);

NAND3X1 _1369_ (
    .A(_376_),
    .B(_472_),
    .C(_311_),
    .Y(_473_)
);

FILL FILL_3__1193_ (
);

FILL FILL_0__1409_ (
);

FILL FILL_2__938_ (
);

FILL FILL_0__1582_ (
);

FILL FILL_0__1162_ (
);

NAND2X1 _912_ (
    .A(_29_),
    .B(_710_),
    .Y(_888_[0])
);

FILL FILL_1__1743_ (
);

FILL FILL_1__1323_ (
);

FILL FILL_3__1249_ (
);

OAI21X1 _1598_ (
    .A(_44_),
    .B(_705__bF$buf3),
    .C(_693_),
    .Y(_19_)
);

OAI21X1 _1178_ (
    .A(_283_),
    .B(_123_),
    .C(_61_),
    .Y(_284_)
);

FILL FILL_2__1812_ (
);

FILL FILL_0__1638_ (
);

FILL FILL_0__1218_ (
);

FILL FILL_0__1391_ (
);

XOR2X1 _1810_ (
    .A(_816_),
    .B(_767_),
    .Y(_817_)
);

FILL FILL_1__1552_ (
);

FILL FILL_1__1132_ (
);

FILL FILL_3__1058_ (
);

FILL FILL_2__1201_ (
);

FILL FILL_0__1447_ (
);

FILL FILL_0__1027_ (
);

FILL FILL_2__976_ (
);

FILL FILL_3__918_ (
);

FILL FILL_1__1608_ (
);

INVX1 _950_ (
    .A(_886_[0]),
    .Y(_56_)
);

FILL FILL_1__1781_ (
);

FILL FILL_1__1361_ (
);

FILL FILL_3__1287_ (
);

FILL FILL_1__998_ (
);

FILL FILL_2__1430_ (
);

FILL FILL_2__1010_ (
);

FILL FILL_0__1676_ (
);

FILL FILL_0__1256_ (
);

FILL FILL_1__1417_ (
);

FILL FILL_1__1590_ (
);

FILL FILL_1__1170_ (
);

FILL FILL_3__1096_ (
);

FILL FILL_0__1485_ (
);

FILL FILL_0__1065_ (
);

FILL FILL_1__1646_ (
);

FILL FILL_1__1226_ (
);

FILL FILL_2__1715_ (
);

FILL FILL_0__1294_ (
);

OAI21X1 _1713_ (
    .A(AI[3]),
    .B(_725_),
    .C(_835_),
    .Y(_728_)
);

FILL FILL_1__1455_ (
);

FILL FILL_1__1035_ (
);

FILL FILL_2__1524_ (
);

FILL FILL_2__1104_ (
);

OAI21X1 _1522_ (
    .A(_396_),
    .B(_526_),
    .C(_623_),
    .Y(_624_)
);

AOI21X1 _1102_ (
    .A(_132_),
    .B(_134_),
    .C(_136_),
    .Y(_208_)
);

FILL FILL_3__994_ (
);

FILL FILL_1__1684_ (
);

FILL FILL_1__1264_ (
);

FILL FILL94350x85950 (
);

FILL FILL_2__1753_ (
);

FILL FILL_2__1333_ (
);

FILL FILL_0__1579_ (
);

FILL FILL_0__1159_ (
);

FILL FILL_0__906_ (
);

FILL FILL_3__1822_ (
);

OAI21X1 _909_ (
    .A(_707_),
    .B(_887_),
    .C(_26_),
    .Y(_27_)
);

OAI21X1 _1751_ (
    .A(_759_),
    .B(_761_),
    .C(_762_),
    .Y(_763_)
);

AOI21X1 _1331_ (
    .A(_427_),
    .B(_431_),
    .C(_435_),
    .Y(_436_)
);

FILL FILL_1__1493_ (
);

FILL FILL_1__1073_ (
);

FILL FILL_2__1809_ (
);

FILL FILL_2__900_ (
);

FILL FILL_2__1562_ (
);

FILL FILL_2__1142_ (
);

FILL FILL_0__1388_ (
);

OAI21X1 _1807_ (
    .A(_809_),
    .B(_808_),
    .C(_814_),
    .Y(CO)
);

FILL FILL_3__1211_ (
);

FILL FILL_1__1549_ (
);

FILL FILL_1__1129_ (
);

NAND3X1 _1560_ (
    .A(_622_),
    .B(_659_),
    .C(_624_),
    .Y(_660_)
);

AOI21X1 _1140_ (
    .A(_242_),
    .B(_245_),
    .C(_176_),
    .Y(_246_)
);

FILL FILL_1__922_ (
);

NAND2X1 _891_ (
    .A(state[1]),
    .B(_700_),
    .Y(_701_)
);

FILL FILL_0__1600_ (
);

FILL FILL_2__1791_ (
);

FILL FILL_2__1371_ (
);

FILL FILL_0__1197_ (
);

DFFSR _1616_ (
    .D(_8_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf3),
    .Q(BI[7])
);

FILL FILL_0__944_ (
);

FILL FILL_3__1440_ (
);

FILL FILL_3__1020_ (
);

INVX4 _947_ (
    .A(ABCmd_i[7]),
    .Y(_54_)
);

FILL FILL_1__1778_ (
);

FILL FILL_1__1358_ (
);

FILL FILL_2__1427_ (
);

FILL FILL_2__1007_ (
);

FILL FILL_2__1180_ (
);

NOR2X1 _1425_ (
    .A(_528_),
    .B(_527_),
    .Y(_529_)
);

NAND3X1 _1005_ (
    .A(_110_),
    .B(_106_),
    .C(_108_),
    .Y(_111_)
);

FILL FILL_3__897_ (
);

FILL FILL_1__1587_ (
);

FILL FILL_1__1167_ (
);

FILL FILL_1__960_ (
);

FILL FILL_2__1656_ (
);

FILL FILL_2__1236_ (
);

FILL FILL_3__1725_ (
);

OAI21X1 _1654_ (
    .A(BI_0_bF$buf3),
    .B(ABCmd_i_2_bF$buf0),
    .C(_825_),
    .Y(_842_)
);

NAND2X1 _1234_ (
    .A(BI[2]),
    .B(AI[6]),
    .Y(_340_)
);

FILL FILL_0__982_ (
);

NAND3X1 _985_ (
    .A(BI_1_bF$buf1),
    .B(AI[4]),
    .C(_90_),
    .Y(_91_)
);

FILL FILL_1__1396_ (
);

FILL FILL_2__1465_ (
);

FILL FILL_2__1045_ (
);

FILL FILL_3__1114_ (
);

INVX1 _1463_ (
    .A(_563_),
    .Y(_566_)
);

INVX2 _1043_ (
    .A(AI[3]),
    .Y(_149_)
);

FILL FILL_0__1503_ (
);

FILL FILL_2__1694_ (
);

FILL FILL_2__1274_ (
);

NAND2X1 _1519_ (
    .A(_573_),
    .B(_618_),
    .Y(_621_)
);

FILL FILL_3__1343_ (
);

NAND2X1 _1692_ (
    .A(ABCmd_i[5]),
    .B(AI[3]),
    .Y(_878_)
);

NOR2X1 _1272_ (
    .A(ABCmd_i[7]),
    .B(HC),
    .Y(_378_)
);

FILL FILL_0__1732_ (
);

FILL FILL_0__1312_ (
);

FILL FILL_2__1083_ (
);

OAI21X1 _1748_ (
    .A(ABCmd_i_2_bF$buf2),
    .B(BI[5]),
    .C(_825_),
    .Y(_760_)
);

NOR2X1 _1328_ (
    .A(_432_),
    .B(_413_),
    .Y(_433_)
);

FILL FILL_3__1572_ (
);

NAND3X1 _1081_ (
    .A(_184_),
    .B(_186_),
    .C(_182_),
    .Y(_187_)
);

FILL FILL_2__1559_ (
);

FILL FILL_0__1541_ (
);

FILL FILL_0__1121_ (
);

FILL FILL_2__1139_ (
);

FILL FILL_3_BUFX2_insert40 (
);

FILL FILL_3_BUFX2_insert41 (
);

FILL FILL_1__1702_ (
);

FILL FILL_3__1208_ (
);

INVX1 _1557_ (
    .A(_886_[6]),
    .Y(_657_)
);

NAND3X1 _1137_ (
    .A(_240_),
    .B(_239_),
    .C(_238_),
    .Y(_243_)
);

FILL FILL_1__919_ (
);

FILL FILL_1__1299_ (
);

FILL FILL_2__1788_ (
);

FILL FILL_0__1770_ (
);

FILL FILL_2__1368_ (
);

FILL FILL_0__1350_ (
);

FILL FILL_1__1511_ (
);

FILL FILL_3__1437_ (
);

FILL FILL_3__1017_ (
);

OAI21X1 _1786_ (
    .A(_792_),
    .B(_794_),
    .C(_795_),
    .Y(_796_)
);

AOI21X1 _1366_ (
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_470_)
);

FILL FILL_3__1190_ (
);

FILL FILL_0__1826_ (
);

FILL FILL_0__1406_ (
);

FILL FILL_2__935_ (
);

FILL FILL_2__1597_ (
);

FILL FILL_2__1177_ (
);

FILL FILL_1__1740_ (
);

FILL FILL_1__1320_ (
);

FILL FILL_3__1246_ (
);

NAND2X1 _1595_ (
    .A(AI[1]),
    .B(_705__bF$buf2),
    .Y(_692_)
);

NAND3X1 _1175_ (
    .A(_269_),
    .B(_279_),
    .C(_280_),
    .Y(_281_)
);

FILL FILL_1__957_ (
);

FILL FILL_0__1215_ (
);

FILL FILL_0__979_ (
);

FILL FILL_3__1475_ (
);

FILL FILL_0__1444_ (
);

FILL FILL_0__1024_ (
);

FILL FILL_2__973_ (
);

FILL FILL_3__915_ (
);

FILL FILL_1__1605_ (
);

FILL FILL_1__995_ (
);

FILL FILL_0__1673_ (
);

FILL FILL_0__1253_ (
);

FILL FILL_1__1414_ (
);

INVX1 _1689_ (
    .A(_875_),
    .Y(ACC[1])
);

NAND3X1 _1269_ (
    .A(_373_),
    .B(_374_),
    .C(_372_),
    .Y(_375_)
);

FILL FILL_3__1093_ (
);

FILL FILL_0__1729_ (
);

FILL FILL_0__1309_ (
);

FILL FILL_0__1482_ (
);

FILL FILL_0__1062_ (
);

FILL FILL_1__1643_ (
);

FILL FILL_1__1223_ (
);

FILL FILL_3__1569_ (
);

FILL FILL_3__1149_ (
);

OAI21X1 _1498_ (
    .A(_592_),
    .B(_558_),
    .C(_599_),
    .Y(_600_)
);

INVX1 _1078_ (
    .A(_183_),
    .Y(_184_)
);

FILL FILL_2__1712_ (
);

FILL FILL_0__1538_ (
);

FILL FILL_0__1118_ (
);

FILL FILL_0__1291_ (
);

AND2X2 _1710_ (
    .A(_831_),
    .B(BI_3_bF$buf2),
    .Y(_725_)
);

FILL FILL92550x58650 (
);

FILL FILL_1__1452_ (
);

FILL FILL_1__1032_ (
);

FILL FILL_3__1798_ (
);

FILL FILL_2__1521_ (
);

FILL FILL_2__1101_ (
);

FILL FILL_0__1767_ (
);

FILL FILL_0__1347_ (
);

FILL FILL93150x7950 (
);

FILL FILL_1__1508_ (
);

FILL FILL_3__991_ (
);

FILL FILL_1__1681_ (
);

FILL FILL_1__1261_ (
);

FILL FILL_3__1187_ (
);

FILL FILL_1__898_ (
);

FILL FILL_2__1750_ (
);

FILL FILL_2__1330_ (
);

FILL FILL_0__1576_ (
);

FILL FILL_0__1156_ (
);

FILL FILL_0__903_ (
);

NOR2X1 _906_ (
    .A(state[1]),
    .B(_712_),
    .Y(_715_)
);

FILL FILL_1__1737_ (
);

FILL FILL_1__1317_ (
);

FILL FILL_1__1490_ (
);

FILL FILL_1__1070_ (
);

FILL FILL_2__1806_ (
);

FILL FILL_0__1385_ (
);

NOR2X1 _1804_ (
    .A(_796_),
    .B(_776_),
    .Y(_812_)
);

FILL FILL_1__1546_ (
);

FILL FILL_1__1126_ (
);

FILL FILL_0__1194_ (
);

DFFSR _1613_ (
    .D(_5_),
    .S(vdd),
    .R(_0__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(BI[4])
);

FILL FILL_0__941_ (
);

INVX1 _944_ (
    .A(ABCmd_i[6]),
    .Y(_52_)
);

FILL FILL_1__1775_ (
);

FILL FILL_1__1355_ (
);

FILL FILL_2__1424_ (
);

FILL FILL_2__1004_ (
);

NAND2X1 _1422_ (
    .A(_376_),
    .B(_472_),
    .Y(_526_)
);

NAND2X1 _1002_ (
    .A(_60_),
    .B(_107_),
    .Y(_108_)
);

FILL FILL_3__894_ (
);

FILL FILL_1__1584_ (
);

FILL FILL_1__1164_ (
);

FILL FILL_2__1653_ (
);

FILL FILL_2__1233_ (
);

FILL FILL_0__1479_ (
);

FILL FILL_0__1059_ (
);

FILL FILL_3__1722_ (
);

NAND2X1 _1651_ (
    .A(_835_),
    .B(_838_),
    .Y(_839_)
);

NAND3X1 _1231_ (
    .A(_333_),
    .B(_336_),
    .C(_334_),
    .Y(_337_)
);

OAI21X1 _982_ (
    .A(_86_),
    .B(_87_),
    .C(_80_),
    .Y(_88_)
);

FILL FILL_1__1393_ (
);

FILL FILL_2__1709_ (
);

FILL FILL_2__1462_ (
);

FILL FILL_2__1042_ (
);

FILL FILL_0__1288_ (
);

INVX1 _1707_ (
    .A(_718_),
    .Y(_722_)
);

FILL FILL_3__1111_ (
);

FILL FILL_1__1449_ (
);

FILL FILL_1__1029_ (
);

NAND3X1 _1460_ (
    .A(_560_),
    .B(_554_),
    .C(_552_),
    .Y(_563_)
);

AND2X2 _1040_ (
    .A(BI_4_bF$buf2),
    .B(AI[2]),
    .Y(_146_)
);

FILL FILL_2__1518_ (
);

FILL FILL_0__1500_ (
);

FILL FILL_2__1691_ (
);

FILL FILL_2__1271_ (
);

FILL FILL_0__1097_ (
);

NAND2X1 _1516_ (
    .A(_576_),
    .B(_523_),
    .Y(_618_)
);

FILL FILL_3__988_ (
);

FILL FILL_3__1760_ (
);

FILL FILL_3__1340_ (
);

FILL FILL_1__1678_ (
);

FILL FILL_1__1258_ (
);

FILL FILL_2__1747_ (
);

FILL FILL_2__1327_ (
);

FILL FILL_2__1080_ (
);

AOI22X1 _1745_ (
    .A(_829_),
    .B(BI[5]),
    .C(_756_),
    .D(_830_),
    .Y(_757_)
);

NOR2X1 _1325_ (
    .A(_414_),
    .B(_127_),
    .Y(_430_)
);

FILL FILL_1__1487_ (
);

FILL FILL_1__1067_ (
);

FILL FILL_2__1556_ (
);

FILL FILL_2__1136_ (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_3_BUFX2_insert19 (
);

AOI21X1 _1554_ (
    .A(_54_),
    .B(_654_),
    .C(state[1]),
    .Y(_655_)
);

NAND3X1 _1134_ (
    .A(_235_),
    .B(_213_),
    .C(_217_),
    .Y(_240_)
);

FILL FILL_1__916_ (
);

FILL FILL_1__1296_ (
);

FILL FILL93450x82050 (
);

FILL FILL_2__1785_ (
);

FILL FILL_2__1365_ (
);

FILL FILL_0__938_ (
);

FILL FILL_3__1014_ (
);

OAI21X1 _1783_ (
    .A(ABCmd_i_2_bF$buf3),
    .B(BI[7]),
    .C(_825_),
    .Y(_793_)
);

AOI21X1 _1363_ (
    .A(_467_),
    .B(_703_),
    .C(_712_),
    .Y(_468_)
);

FILL FILL_0__1823_ (
);

FILL FILL_0__1403_ (
);

FILL FILL_2__932_ (
);

FILL FILL_2__1594_ (
);

FILL FILL_2__1174_ (
);

NAND3X1 _1419_ (
    .A(_515_),
    .B(_518_),
    .C(_522_),
    .Y(_523_)
);

FILL FILL_3__1243_ (
);

AOI22X1 _1592_ (
    .A(_681_),
    .B(_712_),
    .C(_685_),
    .D(_690_),
    .Y(_16_)
);

AOI21X1 _1172_ (
    .A(_270_),
    .B(_276_),
    .C(_275_),
    .Y(_278_)
);

FILL FILL_1__954_ (
);

FILL FILL_0__1212_ (
);

INVX1 _1648_ (
    .A(BI_0_bF$buf3),
    .Y(_836_)
);

NAND2X1 _1228_ (
    .A(_328_),
    .B(_330_),
    .Y(_334_)
);

FILL FILL_0__976_ (
);

FILL FILL_3__1472_ (
);

OAI21X1 _979_ (
    .A(_57_),
    .B(_83_),
    .C(_84_),
    .Y(_85_)
);

FILL FILL_2__1459_ (
);

FILL FILL_0__1441_ (
);

FILL FILL_0__1021_ (
);

FILL FILL_2__1039_ (
);

FILL FILL_2__970_ (
);

FILL FILL_3__912_ (
);

FILL FILL_1__1602_ (
);

FILL FILL_3__1108_ (
);

AND2X2 _1457_ (
    .A(_557_),
    .B(_559_),
    .Y(_560_)
);

AOI21X1 _1037_ (
    .A(_141_),
    .B(_142_),
    .C(_140_),
    .Y(_143_)
);

FILL FILL_1__1199_ (
);

FILL FILL_1__992_ (
);

FILL FILL_2__1688_ (
);

FILL FILL_0__1670_ (
);

FILL FILL_2__1268_ (
);

FILL FILL_0__1250_ (
);

FILL FILL_1__1411_ (
);

FILL FILL_3__1757_ (
);

FILL FILL_3__1337_ (
);

OAI21X1 _1686_ (
    .A(_855_),
    .B(_857_),
    .C(_872_),
    .Y(_873_)
);

OAI21X1 _1266_ (
    .A(_177_),
    .B(_237_),
    .C(_244_),
    .Y(_372_)
);

FILL FILL_3__1090_ (
);

FILL FILL_0__1726_ (
);

FILL FILL_0__1306_ (
);

FILL FILL_2__1497_ (
);

FILL FILL_2__1077_ (
);

FILL FILL_3__950_ (
);

FILL FILL_1__1640_ (
);

FILL FILL_1__1220_ (
);

FILL FILL_3__1566_ (
);

FILL FILL_3__1146_ (
);

INVX1 _1495_ (
    .A(BI[7]),
    .Y(_597_)
);

OAI21X1 _1075_ (
    .A(_137_),
    .B(_133_),
    .C(_128_),
    .Y(_181_)
);

FILL FILL_0__1535_ (
);

FILL FILL_0__1115_ (
);

FILL FILL_3__1375_ (
);

FILL FILL_0__1764_ (
);

FILL FILL_0__1344_ (
);

FILL FILL_1__1505_ (
);

FILL FILL_1__895_ (
);

FILL FILL_2__929_ (
);

FILL FILL_0__1573_ (
);

FILL FILL_0__1153_ (
);

FILL FILL_0__900_ (
);

INVX4 _903_ (
    .A(_700_),
    .Y(_712_)
);

FILL FILL_1__1734_ (
);

FILL FILL_1__1314_ (
);

NAND2X1 _1589_ (
    .A(AN),
    .B(_54_),
    .Y(_688_)
);

OAI21X1 _1169_ (
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(_275_)
);

FILL FILL_2__1803_ (
);

FILL FILL_0__1209_ (
);

FILL FILL_0__1382_ (
);

NAND2X1 _1801_ (
    .A(ABCmd_i[6]),
    .B(_804_),
    .Y(_809_)
);

FILL FILL_1__1543_ (
);

FILL FILL_1__1123_ (
);

FILL FILL_3__1469_ (
);

FILL FILL_3__1049_ (
);

OAI21X1 _1398_ (
    .A(_499_),
    .B(_501_),
    .C(_490_),
    .Y(_502_)
);

FILL FILL_0__1438_ (
);

FILL FILL_0__1018_ (
);

FILL FILL_2__967_ (
);

FILL FILL_3__909_ (
);

FILL FILL_0__1191_ (
);

DFFSR _1610_ (
    .D(_2_),
    .S(vdd),
    .R(_0__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(BI[1])
);

INVX1 _941_ (
    .A(ABCmd_i[5]),
    .Y(_50_)
);

FILL FILL_1__1772_ (
);

FILL FILL_1__1352_ (
);

FILL FILL_1__989_ (
);

FILL FILL_2__1421_ (
);

FILL FILL_2__1001_ (
);

FILL FILL_0__1667_ (
);

FILL FILL_0__1247_ (
);

FILL FILL_1__1408_ (
);

FILL FILL_3__891_ (
);

FILL FILL_1__1581_ (
);

FILL FILL_1__1161_ (
);

FILL FILL_3__1087_ (
);

FILL FILL_2__1650_ (
);

FILL FILL_2__1230_ (
);

FILL FILL_0__1476_ (
);

FILL FILL_0__1056_ (
);

FILL FILL_3__947_ (
);

FILL FILL_1__1637_ (
);

FILL FILL_1__1217_ (
);

FILL FILL_1__1390_ (
);

FILL FILL_2__1706_ (
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert2 (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_0_BUFX2_insert4 (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0__1285_ (
);

INVX1 _1704_ (
    .A(_719_),
    .Y(ACC[2])
);

FILL FILL_1__1446_ (
);

FILL FILL_1__1026_ (
);

FILL FILL_2__1515_ (
);

FILL FILL_0__1094_ (
);

NOR2X1 _1513_ (
    .A(_397_),
    .B(_460_),
    .Y(_615_)
);

FILL FILL_1__1675_ (
);

FILL FILL_1__1255_ (
);

FILL FILL_2__1744_ (
);

FILL FILL_2__1324_ (
);

NAND2X1 _1742_ (
    .A(ABCmd_i[5]),
    .B(AI[6]),
    .Y(_754_)
);

OAI22X1 _1322_ (
    .A(_127_),
    .B(_414_),
    .C(_422_),
    .D(_426_),
    .Y(_427_)
);

FILL FILL_1__1484_ (
);

FILL FILL_1__1064_ (
);

FILL FILL_2__1553_ (
);

FILL FILL_2__1133_ (
);

FILL FILL_0__1799_ (
);

FILL FILL_0__1379_ (
);

AOI21X1 _1551_ (
    .A(_285_),
    .B(_306_),
    .C(_303_),
    .Y(_652_)
);

AOI21X1 _1131_ (
    .A(_236_),
    .B(_230_),
    .C(_179_),
    .Y(_237_)
);

FILL FILL_1__913_ (
);

FILL FILL_1__1293_ (
);

FILL FILL_2_BUFX2_insert0 (
);

FILL FILL_2_BUFX2_insert1 (
);

FILL FILL_2_BUFX2_insert2 (
);

FILL FILL_2_BUFX2_insert3 (
);

FILL FILL_2_BUFX2_insert4 (
);

FILL FILL_2_BUFX2_insert5 (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_2__1782_ (
);

FILL FILL_2__1362_ (
);

FILL FILL_0__1188_ (
);

NAND2X1 _1607_ (
    .A(\u_ALU.AI7 ),
    .B(_705__bF$buf0),
    .Y(_698_)
);

FILL FILL_0__935_ (
);

FILL FILL_3__1011_ (
);

INVX1 _938_ (
    .A(ABCmd_i[4]),
    .Y(_48_)
);

FILL FILL_1__1769_ (
);

FILL FILL_1__1349_ (
);

AOI22X1 _1780_ (
    .A(_829_),
    .B(BI[7]),
    .C(_789_),
    .D(_830_),
    .Y(_790_)
);

NAND2X1 _1360_ (
    .A(ACC[1]),
    .B(_54_),
    .Y(_465_)
);

FILL FILL_0__1820_ (
);

FILL FILL_0__1400_ (
);

FILL FILL_2__1418_ (
);

FILL FILL_2__1591_ (
);

FILL FILL_2__1171_ (
);

NAND3X1 _1416_ (
    .A(_442_),
    .B(_457_),
    .C(_519_),
    .Y(_520_)
);

FILL FILL_3__1660_ (
);

FILL FILL_3__1240_ (
);

FILL FILL_1__1578_ (
);

FILL FILL_1__1158_ (
);

FILL FILL_1__951_ (
);

FILL FILL_2__1647_ (
);

FILL FILL_2__1227_ (
);

NAND2X1 _1645_ (
    .A(AI[0]),
    .B(ABCmd_i[1]),
    .Y(_833_)
);

OAI21X1 _1225_ (
    .A(_83_),
    .B(_74_),
    .C(_330_),
    .Y(_331_)
);

FILL FILL_0__973_ (
);

NAND2X1 _976_ (
    .A(BI_4_bF$buf2),
    .B(AI[1]),
    .Y(_82_)
);

FILL FILL_1__1387_ (
);

FILL FILL_2__1456_ (
);

FILL FILL_2__1036_ (
);

FILL FILL_3__1525_ (
);

OR2X2 _1454_ (
    .A(_555_),
    .B(_556_),
    .Y(_557_)
);

AOI21X1 _1034_ (
    .A(_93_),
    .B(_95_),
    .C(_98_),
    .Y(_140_)
);

FILL FILL_1__1196_ (
);

FILL FILL_2__1685_ (
);

FILL FILL_2__1265_ (
);

FILL FILL_3__1754_ (
);

NAND3X1 _1683_ (
    .A(_840_),
    .B(_863_),
    .C(_869_),
    .Y(_870_)
);

OAI21X1 _1263_ (
    .A(_363_),
    .B(_364_),
    .C(_314_),
    .Y(_369_)
);

FILL FILL_0__1723_ (
);

FILL FILL_0__1303_ (
);

FILL FILL_2__1494_ (
);

FILL FILL_2__1074_ (
);

XOR2X1 _1739_ (
    .A(HC),
    .B(_751_),
    .Y(ACC[4])
);

OAI21X1 _1319_ (
    .A(_423_),
    .B(_58_),
    .C(_417_),
    .Y(_424_)
);

FILL FILL_3__1143_ (
);

OAI21X1 _1492_ (
    .A(_423_),
    .B(_167_),
    .C(_557_),
    .Y(_594_)
);

INVX1 _1072_ (
    .A(_177_),
    .Y(_178_)
);

FILL FILL93450x35250 (
);

FILL FILL_0__1532_ (
);

FILL FILL_0__1112_ (
);

OAI21X1 _1548_ (
    .A(_614_),
    .B(_637_),
    .C(_648_),
    .Y(_649_)
);

NAND3X1 _1128_ (
    .A(_218_),
    .B(_224_),
    .C(_222_),
    .Y(_234_)
);

FILL FILL_3__1372_ (
);

FILL FILL94050x4050 (
);

FILL FILL_0__1761_ (
);

FILL FILL_2__1779_ (
);

FILL FILL_2__1359_ (
);

FILL FILL_0__1341_ (
);

FILL FILL_1__1502_ (
);

FILL FILL_3__1008_ (
);

NAND2X1 _1777_ (
    .A(ABCmd_i[5]),
    .B(ABCmd_i[4]),
    .Y(_787_)
);

OAI21X1 _1357_ (
    .A(_460_),
    .B(_398_),
    .C(ABCmd_i[7]),
    .Y(_462_)
);

FILL FILL_1__1099_ (
);

FILL FILL_0__1817_ (
);

FILL FILL_1__892_ (
);

FILL FILL_2__926_ (
);

FILL FILL_0__1570_ (
);

FILL FILL_2__1588_ (
);

FILL FILL_2__1168_ (
);

FILL FILL_0__1150_ (
);

NOR2X1 _900_ (
    .A(LoadCmd_i),
    .B(_708_),
    .Y(_709_)
);

FILL FILL_1__1731_ (
);

FILL FILL_1__1311_ (
);

FILL FILL_3__1657_ (
);

FILL FILL_3__1237_ (
);

OAI21X1 _1586_ (
    .A(_684_),
    .B(_682_),
    .C(_636_),
    .Y(_685_)
);

OR2X2 _1166_ (
    .A(_62_),
    .B(_271_),
    .Y(_272_)
);

FILL FILL_1__948_ (
);

FILL FILL93750x74250 (
);

FILL FILL_2__1800_ (
);

FILL FILL_0__1206_ (
);

FILL FILL_2__1397_ (
);

FILL FILL_1__1540_ (
);

FILL FILL_1__1120_ (
);

FILL FILL_3__1466_ (
);

FILL FILL_3__1046_ (
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf3)
);

AOI21X1 _1395_ (
    .A(_491_),
    .B(_431_),
    .C(_498_),
    .Y(_499_)
);

FILL FILL_0__1435_ (
);

FILL FILL_0__1015_ (
);

FILL FILL_2__964_ (
);

FILL FILL_3__1275_ (
);

FILL FILL_1__986_ (
);

FILL FILL_0__1664_ (
);

FILL FILL_0__1244_ (
);

FILL FILL_1__1825_ (
);

FILL FILL_1__1405_ (
);

FILL FILL_0__1473_ (
);

FILL FILL_0__1053_ (
);

FILL FILL_3__944_ (
);

FILL FILL_1__1214_ (
);

INVX1 _1489_ (
    .A(_590_),
    .Y(_591_)
);

OAI21X1 _1069_ (
    .A(_174_),
    .B(_173_),
    .C(_170_),
    .Y(_175_)
);

FILL FILL_2__1703_ (
);

FILL FILL_0__1529_ (
);

FILL FILL_0__1109_ (
);

FILL FILL_0__1282_ (
);

OAI21X1 _1701_ (
    .A(_844_),
    .B(_716_),
    .C(_884_),
    .Y(_717_)
);

FILL FILL_1__1443_ (
);

FILL FILL_1__1023_ (
);

FILL FILL_3__1789_ (
);

FILL FILL_3__1369_ (
);

AOI21X1 _1298_ (
    .A(_346_),
    .B(_350_),
    .C(_352_),
    .Y(_403_)
);

FILL FILL_2__1512_ (
);

FILL FILL_0__1758_ (
);

FILL FILL_0__1338_ (
);

FILL FILL_0__1091_ (
);

NAND2X1 _1510_ (
    .A(_569_),
    .B(_571_),
    .Y(_612_)
);

FILL FILL_1__1672_ (
);

FILL FILL_1__1252_ (
);

FILL FILL_3__1598_ (
);

FILL FILL_3__1178_ (
);

FILL FILL_1__889_ (
);

FILL FILL_2__1741_ (
);

FILL FILL_2__1321_ (
);

FILL FILL_0__1567_ (
);

FILL FILL_0__1147_ (
);

FILL FILL_3__1810_ (
);

FILL FILL_1__1728_ (
);

FILL FILL_1__1308_ (
);

FILL FILL_1__1481_ (
);

FILL FILL_1__1061_ (
);

FILL FILL_2__1550_ (
);

FILL FILL_2__1130_ (
);

FILL FILL_0__1796_ (
);

FILL FILL_0__1376_ (
);

FILL FILL_1__1537_ (
);

FILL FILL_1__1117_ (
);

FILL FILL_1__910_ (
);

FILL FILL_1__1290_ (
);

FILL FILL_2__1606_ (
);

FILL FILL_0__1185_ (
);

OAI21X1 _1604_ (
    .A(_50_),
    .B(_705__bF$buf2),
    .C(_696_),
    .Y(_22_)
);

FILL FILL_0__932_ (
);

INVX1 _935_ (
    .A(ABCmd_i[3]),
    .Y(_46_)
);

FILL FILL_1__1766_ (
);

FILL FILL_1__1346_ (
);

FILL FILL93750x62550 (
);

FILL FILL_2__1415_ (
);

OAI21X1 _1413_ (
    .A(_510_),
    .B(_513_),
    .C(_479_),
    .Y(_517_)
);

FILL FILL_1__1575_ (
);

FILL FILL_1__1155_ (
);

FILL FILL_2__1644_ (
);

FILL FILL_2__1224_ (
);

FILL FILL_2__999_ (
);

NAND2X1 _1642_ (
    .A(ABCmd_i[0]),
    .B(_829_),
    .Y(_830_)
);

AND2X2 _1222_ (
    .A(BI_4_bF$buf1),
    .B(AI[4]),
    .Y(_328_)
);

FILL FILL_0__970_ (
);

OAI21X1 _973_ (
    .A(_77_),
    .B(_78_),
    .C(_68_),
    .Y(_79_)
);

FILL FILL_1__1384_ (
);

FILL FILL_2__1453_ (
);

FILL FILL_2__1033_ (
);

FILL FILL_0__1699_ (
);

FILL FILL_0__1279_ (
);

FILL FILL93150x58650 (
);

FILL FILL_3__1522_ (
);

OAI21X1 _1451_ (
    .A(_550_),
    .B(_553_),
    .C(_545_),
    .Y(_554_)
);

AOI22X1 _1031_ (
    .A(BI_0_bF$buf0),
    .B(AI[6]),
    .C(BI_1_bF$buf3),
    .D(AI_5_bF$buf2),
    .Y(_137_)
);

FILL FILL_1__1193_ (
);

FILL FILL_2__1509_ (
);

FILL FILL_2__1682_ (
);

FILL FILL_2__1262_ (
);

FILL FILL_0__1088_ (
);

NAND3X1 _1507_ (
    .A(_590_),
    .B(_605_),
    .C(_608_),
    .Y(_609_)
);

FILL FILL_3__979_ (
);

FILL FILL_3__1751_ (
);

FILL FILL_1__1669_ (
);

FILL FILL_1__1249_ (
);

NAND2X1 _1680_ (
    .A(_866_),
    .B(_865_),
    .Y(_867_)
);

AOI21X1 _1260_ (
    .A(_361_),
    .B(_365_),
    .C(_313_),
    .Y(_366_)
);

FILL FILL_2__1738_ (
);

FILL FILL_0__1720_ (
);

FILL FILL_2__1318_ (
);

FILL FILL_0__1300_ (
);

FILL FILL_2__1491_ (
);

FILL FILL_2__1071_ (
);

FILL FILL_3__1807_ (
);

OAI21X1 _1736_ (
    .A(_844_),
    .B(_748_),
    .C(_746_),
    .Y(_749_)
);

INVX1 _1316_ (
    .A(_420_),
    .Y(_421_)
);

FILL FILL_3__1140_ (
);

FILL FILL_1__1478_ (
);

FILL FILL_1__1058_ (
);

FILL FILL_2__1547_ (
);

FILL FILL_2__1127_ (
);

XOR2X1 _1545_ (
    .A(_645_),
    .B(_640_),
    .Y(_646_)
);

AOI21X1 _1125_ (
    .A(_216_),
    .B(_215_),
    .C(_214_),
    .Y(_231_)
);

FILL FILL_1__907_ (
);

FILL FILL_1__1287_ (
);

FILL FILL_2__1776_ (
);

FILL FILL_2__1356_ (
);

FILL FILL_0__929_ (
);

FILL FILL_3__1425_ (
);

NAND2X1 _1774_ (
    .A(_784_),
    .B(_783_),
    .Y(_785_)
);

NAND3X1 _1354_ (
    .A(_457_),
    .B(_458_),
    .C(_456_),
    .Y(_459_)
);

FILL FILL_1__1096_ (
);

FILL FILL_0__1814_ (
);

FILL FILL_2__923_ (
);

FILL FILL_2__1585_ (
);

FILL FILL_2__1165_ (
);

FILL FILL_3__1654_ (
);

AOI21X1 _1583_ (
    .A(_660_),
    .B(_663_),
    .C(_668_),
    .Y(_682_)
);

NAND3X1 _1163_ (
    .A(_256_),
    .B(_257_),
    .C(_80_),
    .Y(_269_)
);

FILL FILL_1__945_ (
);

FILL FILL_0__1203_ (
);

FILL FILL_2__1394_ (
);

NOR2X1 _1639_ (
    .A(ABCmd_i[5]),
    .B(_826_),
    .Y(_827_)
);

NAND2X1 _1219_ (
    .A(_324_),
    .B(_321_),
    .Y(_325_)
);

FILL FILL_0__967_ (
);

FILL FILL_3__1043_ (
);

INVX1 _1392_ (
    .A(_495_),
    .Y(_496_)
);

FILL FILL_0__1432_ (
);

FILL FILL_0__1012_ (
);

FILL FILL_2__961_ (
);

FILL FILL_3__1519_ (
);

INVX1 _1448_ (
    .A(_550_),
    .Y(_551_)
);

INVX1 _1028_ (
    .A(_133_),
    .Y(_134_)
);

FILL FILL_3__1272_ (
);

FILL FILL_1__983_ (
);

endmodule
