magic
tech scmos
magscale 1 2
timestamp 1715667437
<< metal1 >>
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 527 6137 593 6143
rect 5827 6137 5853 6143
rect 907 6123 920 6127
rect 907 6113 923 6123
rect 1347 6117 1373 6123
rect 5387 6117 5413 6123
rect 917 6083 923 6113
rect 917 6080 943 6083
rect 917 6077 947 6080
rect 933 6067 947 6077
rect 1607 6077 1633 6083
rect 907 6046 920 6047
rect 907 6033 913 6046
rect 6323 5998 6383 6258
rect 6290 5982 6383 5998
rect 1907 5917 1933 5923
rect 5547 5917 5613 5923
rect 840 5903 853 5907
rect 837 5893 853 5903
rect 5247 5903 5260 5907
rect 5247 5893 5263 5903
rect 837 5867 843 5893
rect 5257 5867 5263 5893
rect 827 5857 843 5867
rect 827 5853 840 5857
rect 5247 5857 5263 5867
rect 5247 5853 5260 5857
rect 147 5837 173 5843
rect 1347 5817 1413 5823
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 367 5617 393 5623
rect 3707 5617 3753 5623
rect 4647 5617 4673 5623
rect 4687 5617 4713 5623
rect 187 5593 213 5607
rect 780 5603 793 5607
rect 777 5593 793 5603
rect 2800 5603 2813 5607
rect 2797 5593 2813 5603
rect 2947 5597 2973 5603
rect 3827 5603 3840 5607
rect 4080 5603 4093 5607
rect 3827 5593 3843 5603
rect 197 5567 203 5593
rect 777 5567 783 5593
rect 197 5557 213 5567
rect 200 5553 213 5557
rect 767 5557 783 5567
rect 2797 5563 2803 5593
rect 3837 5567 3843 5593
rect 2757 5557 2803 5563
rect 767 5553 780 5557
rect 2757 5547 2763 5557
rect 3827 5557 3843 5567
rect 4077 5593 4093 5603
rect 4077 5567 4083 5593
rect 4077 5557 4093 5567
rect 3827 5553 3840 5557
rect 4080 5553 4093 5557
rect 2327 5537 2373 5543
rect 193 5527 207 5533
rect 2607 5537 2653 5543
rect 2740 5545 2763 5547
rect 2747 5537 2763 5545
rect 2747 5533 2760 5537
rect 2787 5537 2853 5543
rect 193 5526 220 5527
rect 193 5520 213 5526
rect 197 5517 213 5520
rect 200 5513 213 5517
rect 1807 5517 1853 5523
rect 2633 5503 2647 5513
rect 2633 5500 2673 5503
rect 2637 5497 2673 5500
rect 6323 5478 6383 5982
rect 6290 5462 6383 5478
rect 3460 5383 3473 5387
rect 3457 5373 3473 5383
rect 3587 5383 3600 5387
rect 3587 5373 3603 5383
rect 3827 5383 3840 5387
rect 4373 5383 4387 5393
rect 3827 5373 3843 5383
rect 4373 5380 4413 5383
rect 4377 5377 4413 5380
rect 3457 5347 3463 5373
rect 3457 5337 3473 5347
rect 3460 5333 3473 5337
rect 147 5317 173 5323
rect 187 5317 213 5323
rect 227 5317 293 5323
rect 747 5317 773 5323
rect 3597 5326 3603 5373
rect 3837 5327 3843 5373
rect 3837 5326 3860 5327
rect 3427 5317 3513 5323
rect 3837 5317 3853 5326
rect 3840 5313 3853 5317
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 2107 5097 2233 5103
rect 2560 5103 2573 5107
rect 2557 5093 2573 5103
rect 2747 5097 2793 5103
rect 4053 5103 4067 5113
rect 4053 5100 4153 5103
rect 4057 5097 4153 5100
rect 5167 5097 5213 5103
rect 5307 5097 5373 5103
rect 5927 5097 6013 5103
rect 620 5083 633 5087
rect 617 5073 633 5083
rect 760 5083 773 5087
rect 757 5073 773 5083
rect 900 5083 913 5087
rect 897 5073 913 5083
rect 2007 5083 2020 5087
rect 2557 5083 2563 5093
rect 2007 5073 2023 5083
rect 107 5017 173 5023
rect 617 5023 623 5073
rect 757 5047 763 5073
rect 897 5047 903 5073
rect 757 5037 773 5047
rect 760 5033 773 5037
rect 887 5037 903 5047
rect 2017 5043 2023 5073
rect 2537 5077 2563 5083
rect 2407 5063 2420 5067
rect 2407 5053 2423 5063
rect 2417 5047 2423 5053
rect 2537 5047 2543 5077
rect 2657 5047 2663 5093
rect 2940 5083 2953 5087
rect 2937 5073 2953 5083
rect 4080 5083 4093 5087
rect 4077 5073 4093 5083
rect 4220 5083 4233 5087
rect 4217 5073 4233 5083
rect 2937 5047 2943 5073
rect 2017 5037 2053 5043
rect 887 5033 900 5037
rect 2417 5037 2433 5047
rect 2420 5033 2433 5037
rect 2537 5037 2553 5047
rect 2540 5033 2553 5037
rect 2647 5037 2663 5047
rect 2647 5033 2660 5037
rect 2927 5037 2943 5047
rect 4077 5047 4083 5073
rect 4217 5047 4223 5073
rect 4077 5037 4093 5047
rect 2927 5033 2940 5037
rect 4080 5033 4093 5037
rect 4217 5037 4233 5047
rect 4220 5033 4233 5037
rect 5127 5037 5173 5043
rect 617 5017 653 5023
rect 5287 5017 5373 5023
rect 5807 5017 5853 5023
rect 6323 4958 6383 5462
rect 6290 4942 6383 4958
rect 4893 4903 4907 4913
rect 4893 4900 4973 4903
rect 4897 4897 4973 4900
rect 5027 4897 5053 4903
rect 1893 4883 1907 4893
rect 1877 4880 1907 4883
rect 1877 4877 1903 4880
rect 787 4857 813 4863
rect 1877 4863 1883 4877
rect 1947 4877 1993 4883
rect 2020 4883 2033 4887
rect 2017 4873 2033 4883
rect 4867 4877 4953 4883
rect 6067 4877 6093 4883
rect 2017 4863 2023 4873
rect 1857 4857 1883 4863
rect 1977 4857 2023 4863
rect 2093 4863 2107 4873
rect 2093 4860 2133 4863
rect 2097 4857 2133 4860
rect 747 4797 813 4803
rect 1087 4797 1133 4803
rect 1307 4797 1373 4803
rect 1857 4803 1863 4857
rect 1977 4827 1983 4857
rect 2247 4863 2260 4867
rect 2247 4853 2263 4863
rect 2687 4857 2723 4863
rect 1967 4817 1983 4827
rect 2257 4827 2263 4853
rect 2717 4827 2723 4857
rect 2257 4817 2273 4827
rect 1967 4813 1980 4817
rect 2260 4813 2273 4817
rect 2717 4817 2733 4827
rect 2720 4813 2733 4817
rect 3577 4823 3583 4873
rect 3577 4817 3613 4823
rect 1857 4797 1893 4803
rect 5247 4797 5273 4803
rect 5287 4797 5373 4803
rect 5447 4797 5513 4803
rect 2087 4777 2173 4783
rect 5567 4777 5613 4783
rect 2687 4757 2713 4763
rect 4587 4757 4613 4763
rect 2833 4723 2847 4733
rect 2833 4720 2893 4723
rect 2837 4717 2893 4720
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 1287 4637 1313 4643
rect 2757 4637 2793 4643
rect 2757 4607 2763 4637
rect 2747 4597 2763 4607
rect 2747 4593 2760 4597
rect 547 4577 613 4583
rect 827 4577 893 4583
rect 1307 4577 1353 4583
rect 1847 4583 1860 4587
rect 2800 4583 2813 4587
rect 1847 4574 1863 4583
rect 1840 4573 1863 4574
rect 1300 4563 1313 4567
rect 1297 4553 1313 4563
rect 1447 4563 1460 4567
rect 1447 4553 1463 4563
rect 1297 4503 1303 4553
rect 1247 4497 1303 4503
rect 1457 4503 1463 4553
rect 1857 4506 1863 4573
rect 2797 4573 2813 4583
rect 3977 4577 4033 4583
rect 1887 4557 1913 4563
rect 2020 4563 2033 4567
rect 2017 4553 2033 4563
rect 2797 4563 2803 4573
rect 2777 4557 2803 4563
rect 2017 4523 2023 4553
rect 2777 4527 2783 4557
rect 2017 4520 2043 4523
rect 2017 4517 2047 4520
rect 2777 4517 2793 4527
rect 2033 4507 2047 4517
rect 2780 4513 2793 4517
rect 1427 4497 1463 4503
rect 3977 4506 3983 4577
rect 4000 4563 4013 4567
rect 3997 4553 4013 4563
rect 5940 4563 5953 4567
rect 5937 4553 5953 4563
rect 6047 4563 6060 4567
rect 6047 4553 6063 4563
rect 3997 4527 4003 4553
rect 3997 4517 4013 4527
rect 4000 4513 4013 4517
rect 5647 4517 5673 4523
rect 5937 4523 5943 4553
rect 5907 4517 5943 4523
rect 6057 4503 6063 4553
rect 6027 4497 6063 4503
rect 3867 4477 3913 4483
rect 6323 4438 6383 4942
rect 6290 4422 6383 4438
rect 767 4377 793 4383
rect 787 4357 833 4363
rect 907 4337 953 4343
rect 1080 4343 1093 4347
rect 1077 4333 1093 4343
rect 4580 4343 4593 4347
rect 4577 4333 4593 4343
rect 1077 4307 1083 4333
rect 1077 4297 1093 4307
rect 1080 4293 1093 4297
rect 3247 4297 3293 4303
rect 3993 4303 4007 4313
rect 4577 4307 4583 4333
rect 3993 4300 4033 4303
rect 3997 4297 4033 4300
rect 4567 4297 4583 4307
rect 4567 4293 4580 4297
rect 5327 4297 5373 4303
rect 427 4277 473 4283
rect 3987 4277 4013 4283
rect 4427 4277 4473 4283
rect 5887 4277 5953 4283
rect 6207 4277 6253 4283
rect -63 4162 30 4178
rect 3307 4173 3310 4187
rect -63 3658 -3 4162
rect 3867 4137 3913 4143
rect 4777 4143 4783 4163
rect 4747 4137 4783 4143
rect 167 4077 213 4083
rect 1387 4077 1453 4083
rect 147 4057 173 4063
rect 267 4057 333 4063
rect 347 4057 393 4063
rect 2767 4057 2873 4063
rect 4187 4057 4233 4063
rect 4487 4057 4553 4063
rect 5247 4057 5333 4063
rect 60 4043 73 4047
rect 57 4033 73 4043
rect 467 4037 503 4043
rect 57 4007 63 4033
rect 497 4007 503 4037
rect 597 4007 603 4053
rect 727 4043 740 4047
rect 1120 4043 1133 4047
rect 727 4033 743 4043
rect 737 4007 743 4033
rect 1117 4033 1133 4043
rect 1247 4043 1260 4047
rect 1247 4033 1263 4043
rect 1407 4037 1443 4043
rect 1117 4007 1123 4033
rect 1257 4007 1263 4033
rect 57 3997 73 4007
rect 60 3993 73 3997
rect 497 3997 513 4007
rect 500 3993 513 3997
rect 587 3997 603 4007
rect 587 3993 600 3997
rect 1107 3997 1123 4007
rect 1107 3993 1120 3997
rect 1247 3997 1263 4007
rect 1437 4007 1443 4037
rect 1567 4043 1580 4047
rect 1880 4043 1893 4047
rect 1567 4033 1583 4043
rect 1577 4007 1583 4033
rect 1877 4033 1893 4043
rect 1967 4043 1980 4047
rect 2240 4043 2253 4047
rect 1967 4033 1983 4043
rect 1437 3997 1453 4007
rect 1247 3993 1260 3997
rect 1440 3993 1453 3997
rect 1567 3997 1583 4007
rect 1567 3993 1580 3997
rect 1877 4003 1883 4033
rect 1847 3997 1883 4003
rect 1977 4007 1983 4033
rect 2237 4033 2253 4043
rect 4060 4043 4073 4047
rect 4057 4033 4073 4043
rect 4360 4043 4373 4047
rect 4357 4033 4373 4043
rect 5720 4043 5733 4047
rect 5717 4033 5733 4043
rect 5807 4043 5820 4047
rect 5807 4033 5823 4043
rect 1977 3997 1993 4007
rect 1980 3993 1993 3997
rect 2237 4003 2243 4033
rect 4057 4007 4063 4033
rect 4357 4007 4363 4033
rect 5717 4007 5723 4033
rect 5817 4007 5823 4033
rect 2217 3997 2243 4003
rect 2217 3987 2223 3997
rect 2787 3997 2833 4003
rect 4057 3997 4073 4007
rect 4060 3993 4073 3997
rect 4357 3997 4373 4007
rect 4360 3993 4373 3997
rect 5717 3997 5733 4007
rect 5720 3993 5733 3997
rect 5807 3997 5823 4007
rect 5807 3993 5820 3997
rect 1687 3977 1773 3983
rect 2207 3977 2223 3987
rect 2207 3973 2220 3977
rect 6087 3977 6233 3983
rect 5787 3957 5833 3963
rect 5687 3937 5733 3943
rect 6323 3918 6383 4422
rect 6290 3902 6383 3918
rect 3867 3857 3933 3863
rect 307 3837 333 3843
rect 1327 3843 1340 3847
rect 1327 3833 1343 3843
rect 457 3787 463 3833
rect 567 3817 603 3823
rect 447 3777 463 3787
rect 597 3787 603 3817
rect 1307 3823 1320 3827
rect 1307 3813 1323 3823
rect 597 3777 613 3787
rect 447 3773 460 3777
rect 600 3773 613 3777
rect 853 3783 867 3793
rect 827 3780 867 3783
rect 827 3777 863 3780
rect 987 3777 1013 3783
rect 267 3757 333 3763
rect 847 3757 893 3763
rect 1317 3763 1323 3813
rect 1337 3787 1343 3833
rect 3747 3837 3793 3843
rect 5087 3837 5133 3843
rect 5520 3823 5533 3827
rect 2987 3820 3023 3823
rect 2987 3817 3027 3820
rect 1337 3777 1353 3787
rect 1340 3773 1353 3777
rect 1833 3783 1847 3793
rect 2137 3787 2143 3813
rect 3013 3807 3027 3817
rect 5517 3813 5533 3823
rect 1833 3780 1873 3783
rect 1837 3777 1873 3780
rect 2127 3777 2143 3787
rect 2677 3780 2713 3783
rect 2673 3777 2713 3780
rect 2127 3773 2140 3777
rect 1287 3757 1323 3763
rect 1467 3740 1503 3743
rect 1467 3737 1507 3740
rect 1493 3727 1507 3737
rect 1517 3727 1523 3773
rect 2673 3766 2687 3777
rect 3887 3757 3933 3763
rect 4367 3757 4413 3763
rect 5367 3757 5453 3763
rect 5517 3763 5523 3813
rect 5517 3757 5553 3763
rect 5647 3757 5733 3763
rect 1506 3720 1507 3727
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 2687 3617 2733 3623
rect 2687 3560 2763 3563
rect 2687 3557 2767 3560
rect 2753 3548 2767 3557
rect 547 3537 603 3543
rect 597 3483 603 3537
rect 1427 3537 1453 3543
rect 1857 3537 1893 3543
rect 727 3523 740 3527
rect 860 3523 873 3527
rect 727 3513 743 3523
rect 737 3487 743 3513
rect 857 3513 873 3523
rect 987 3523 1000 3527
rect 1020 3523 1033 3527
rect 987 3513 1003 3523
rect 857 3487 863 3513
rect 597 3477 623 3483
rect 737 3477 753 3487
rect 397 3460 453 3463
rect 393 3457 453 3460
rect 393 3447 407 3457
rect 617 3463 623 3477
rect 740 3473 753 3477
rect 857 3477 873 3487
rect 860 3473 873 3477
rect 617 3457 653 3463
rect 997 3463 1003 3513
rect 1017 3513 1033 3523
rect 1267 3523 1280 3527
rect 1267 3513 1283 3523
rect 1687 3523 1700 3527
rect 1687 3513 1703 3523
rect 1807 3523 1820 3527
rect 1857 3523 1863 3537
rect 4527 3537 4593 3543
rect 5887 3537 5913 3543
rect 5927 3537 5973 3543
rect 1807 3513 1823 3523
rect 1017 3487 1023 3513
rect 1277 3487 1283 3513
rect 1697 3487 1703 3513
rect 1817 3487 1823 3513
rect 1017 3477 1033 3487
rect 1020 3473 1033 3477
rect 1267 3477 1283 3487
rect 1517 3477 1553 3483
rect 1267 3473 1280 3477
rect 997 3457 1053 3463
rect 1517 3443 1523 3477
rect 1697 3477 1713 3487
rect 1700 3473 1713 3477
rect 1807 3477 1823 3487
rect 1837 3517 1863 3523
rect 1837 3487 1843 3517
rect 2087 3523 2100 3527
rect 2720 3523 2733 3527
rect 2087 3513 2103 3523
rect 2097 3487 2103 3513
rect 1837 3477 1853 3487
rect 1807 3473 1820 3477
rect 1840 3473 1853 3477
rect 2087 3477 2103 3487
rect 2717 3513 2733 3523
rect 4427 3523 4440 3527
rect 4427 3513 4443 3523
rect 4847 3523 4860 3527
rect 4847 3513 4863 3523
rect 5007 3523 5020 3527
rect 5007 3513 5023 3523
rect 2087 3473 2100 3477
rect 2717 3483 2723 3513
rect 2687 3477 2723 3483
rect 4437 3487 4443 3513
rect 4437 3477 4453 3487
rect 4440 3473 4453 3477
rect 4857 3483 4863 3513
rect 4837 3480 4863 3483
rect 4833 3477 4863 3480
rect 5017 3487 5023 3513
rect 5017 3477 5033 3487
rect 4833 3467 4847 3477
rect 5020 3473 5033 3477
rect 5107 3457 5133 3463
rect 6147 3457 6173 3463
rect 1517 3437 1553 3443
rect 6323 3398 6383 3902
rect 6290 3382 6383 3398
rect 1967 3337 1993 3343
rect 927 3317 953 3323
rect 2207 3317 2253 3323
rect 3227 3317 3293 3323
rect 4240 3323 4253 3327
rect 4237 3313 4253 3323
rect 4847 3317 4933 3323
rect 5727 3323 5740 3327
rect 5727 3313 5743 3323
rect 317 3297 353 3303
rect 317 3267 323 3297
rect 447 3297 473 3303
rect 1173 3303 1187 3313
rect 1700 3303 1713 3307
rect 1173 3300 1223 3303
rect 1177 3297 1223 3300
rect 307 3257 323 3267
rect 1217 3263 1223 3297
rect 1697 3293 1713 3303
rect 2120 3303 2133 3307
rect 2117 3293 2133 3303
rect 4047 3297 4083 3303
rect 1697 3267 1703 3293
rect 2117 3267 2123 3293
rect 1217 3257 1243 3263
rect 1697 3257 1713 3267
rect 307 3253 320 3257
rect 427 3237 553 3243
rect 887 3237 973 3243
rect 1237 3243 1243 3257
rect 1700 3253 1713 3257
rect 2107 3257 2123 3267
rect 4077 3267 4083 3297
rect 4077 3257 4093 3267
rect 2107 3253 2120 3257
rect 4080 3253 4093 3257
rect 4237 3263 4243 3313
rect 5737 3303 5743 3313
rect 5737 3297 5763 3303
rect 5757 3267 5763 3297
rect 6047 3303 6060 3307
rect 6047 3293 6063 3303
rect 4207 3257 4243 3263
rect 5747 3257 5763 3267
rect 5747 3253 5760 3257
rect 5907 3257 5933 3263
rect 1237 3237 1293 3243
rect 2527 3237 2613 3243
rect 4847 3237 4953 3243
rect 5487 3237 5533 3243
rect 5787 3237 5833 3243
rect 6057 3243 6063 3293
rect 6187 3257 6213 3263
rect 6027 3237 6063 3243
rect 6227 3237 6253 3243
rect 767 3217 813 3223
rect 2207 3217 2293 3223
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 2897 3107 2903 3123
rect 2887 3097 2903 3107
rect 2887 3093 2900 3097
rect 1547 3037 1633 3043
rect 5307 3037 5373 3043
rect 567 3017 593 3023
rect 1657 3017 1693 3023
rect 320 3006 340 3007
rect 320 3003 333 3006
rect 317 2993 333 3003
rect 317 2967 323 2993
rect 940 3003 953 3007
rect 937 2993 953 3003
rect 1607 3003 1620 3007
rect 1657 3003 1663 3017
rect 1887 3017 1933 3023
rect 2747 3017 2773 3023
rect 5347 3017 5413 3023
rect 5497 3017 5553 3023
rect 2933 3003 2947 3013
rect 3200 3003 3213 3007
rect 1607 2993 1623 3003
rect 187 2957 213 2963
rect 317 2957 333 2967
rect 320 2953 333 2957
rect 937 2963 943 2993
rect 1617 2963 1623 2993
rect 907 2957 943 2963
rect 1597 2960 1623 2963
rect 1593 2957 1623 2960
rect 1637 2997 1663 3003
rect 2917 3000 2947 3003
rect 2917 2997 2943 3000
rect 1637 2967 1643 2997
rect 2917 2967 2923 2997
rect 3197 2993 3213 3003
rect 3927 3003 3940 3007
rect 3927 2993 3943 3003
rect 4867 3003 4880 3007
rect 5060 3003 5073 3007
rect 4867 2993 4883 3003
rect 1637 2957 1653 2967
rect 1593 2947 1607 2957
rect 1640 2953 1653 2957
rect 2917 2957 2933 2967
rect 2920 2953 2933 2957
rect 3197 2963 3203 2993
rect 3937 2967 3943 2993
rect 4877 2967 4883 2993
rect 3167 2957 3203 2963
rect 3927 2957 3943 2967
rect 3927 2953 3940 2957
rect 4867 2957 4883 2967
rect 5057 2993 5073 3003
rect 5180 3003 5193 3007
rect 5177 2993 5193 3003
rect 5497 3003 5503 3017
rect 5807 3017 5833 3023
rect 5957 3017 5993 3023
rect 5477 2997 5503 3003
rect 5057 2967 5063 2993
rect 5177 2967 5183 2993
rect 5477 2967 5483 2997
rect 5607 3003 5620 3007
rect 5640 3003 5653 3007
rect 5607 2993 5623 3003
rect 5057 2957 5073 2967
rect 4867 2953 4880 2957
rect 5060 2953 5073 2957
rect 5177 2957 5193 2967
rect 5180 2953 5193 2957
rect 5467 2957 5483 2967
rect 5467 2953 5480 2957
rect 5617 2947 5623 2993
rect 5637 2993 5653 3003
rect 5767 3003 5780 3007
rect 5957 3003 5963 3017
rect 6147 3017 6233 3023
rect 5767 2993 5783 3003
rect 5637 2967 5643 2993
rect 5637 2957 5653 2967
rect 5640 2953 5653 2957
rect 5777 2963 5783 2993
rect 5937 2997 5963 3003
rect 5937 2967 5943 2997
rect 6207 3003 6220 3007
rect 6207 2993 6223 3003
rect 5777 2957 5813 2963
rect 5937 2957 5953 2967
rect 5940 2953 5953 2957
rect 6217 2947 6223 2993
rect 4207 2937 4253 2943
rect 6323 2878 6383 3382
rect 6290 2862 6383 2878
rect 1387 2797 1453 2803
rect 1667 2797 1693 2803
rect 2467 2783 2480 2787
rect 2467 2773 2483 2783
rect 3207 2783 3220 2787
rect 3240 2783 3253 2787
rect 3207 2773 3223 2783
rect 3237 2780 3253 2783
rect 2477 2747 2483 2773
rect 2467 2737 2483 2747
rect 3217 2743 3223 2773
rect 3233 2773 3253 2780
rect 3387 2783 3400 2787
rect 3420 2783 3433 2787
rect 3387 2773 3403 2783
rect 3233 2766 3247 2773
rect 3397 2747 3403 2773
rect 3197 2737 3223 2743
rect 2467 2733 2480 2737
rect 2827 2717 2953 2723
rect 3197 2723 3203 2737
rect 3387 2737 3403 2747
rect 3417 2773 3433 2783
rect 3540 2783 3553 2787
rect 3537 2773 3553 2783
rect 3667 2777 3703 2783
rect 3417 2747 3423 2773
rect 3537 2747 3543 2773
rect 3697 2747 3703 2777
rect 6177 2777 6213 2783
rect 6177 2747 6183 2777
rect 3417 2737 3433 2747
rect 3387 2733 3400 2737
rect 3420 2733 3433 2737
rect 3537 2737 3553 2747
rect 3540 2733 3553 2737
rect 3697 2737 3713 2747
rect 3700 2733 3713 2737
rect 6167 2737 6183 2747
rect 6167 2733 6180 2737
rect 3167 2717 3203 2723
rect 3507 2717 3573 2723
rect 3907 2717 3953 2723
rect 4647 2717 4713 2723
rect 5147 2717 5233 2723
rect 5987 2717 6033 2723
rect 5567 2697 5633 2703
rect 3907 2677 3973 2683
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 2887 2537 2953 2543
rect 2887 2517 2913 2523
rect 987 2497 1013 2503
rect 1587 2497 1653 2503
rect 3367 2497 3433 2503
rect 4087 2497 4173 2503
rect 5607 2497 5653 2503
rect 6167 2497 6233 2503
rect 2180 2483 2193 2487
rect 2177 2473 2193 2483
rect 2307 2483 2320 2487
rect 2307 2473 2323 2483
rect 3387 2483 3400 2487
rect 3387 2473 3403 2483
rect 3807 2483 3820 2487
rect 5780 2483 5793 2487
rect 3807 2473 3823 2483
rect 2177 2447 2183 2473
rect 2177 2437 2193 2447
rect 2180 2433 2193 2437
rect 1467 2417 1493 2423
rect 2317 2423 2323 2473
rect 3397 2447 3403 2473
rect 3240 2443 3253 2447
rect 3237 2433 3253 2443
rect 3397 2437 3413 2447
rect 3400 2433 3413 2437
rect 3237 2427 3243 2433
rect 2247 2417 2323 2423
rect 3227 2417 3243 2427
rect 3227 2413 3240 2417
rect 3817 2407 3823 2473
rect 5777 2473 5793 2483
rect 5940 2483 5953 2487
rect 5937 2473 5953 2483
rect 6067 2483 6080 2487
rect 6067 2473 6083 2483
rect 5777 2443 5783 2473
rect 5747 2437 5783 2443
rect 5937 2447 5943 2473
rect 5937 2437 5953 2447
rect 5940 2433 5953 2437
rect 6077 2443 6083 2473
rect 6077 2437 6113 2443
rect 3817 2406 3840 2407
rect 3817 2397 3833 2406
rect 3820 2393 3833 2397
rect 6267 2397 6293 2403
rect 6323 2358 6383 2862
rect 6290 2342 6383 2358
rect 3887 2297 3953 2303
rect 1287 2277 1353 2283
rect 2267 2277 2313 2283
rect 3820 2283 3833 2287
rect 3817 2274 3833 2283
rect 3817 2273 3840 2274
rect 2967 2257 3003 2263
rect 2997 2226 3003 2257
rect 3127 2257 3153 2263
rect 3253 2263 3267 2273
rect 3253 2260 3293 2263
rect 3257 2257 3293 2260
rect 3537 2223 3543 2273
rect 3817 2263 3823 2273
rect 5280 2263 5293 2267
rect 3797 2257 3823 2263
rect 3797 2227 3803 2257
rect 5277 2253 5293 2263
rect 6060 2263 6073 2267
rect 6057 2253 6073 2263
rect 6200 2263 6213 2267
rect 6197 2253 6213 2263
rect 5277 2227 5283 2253
rect 3537 2217 3563 2223
rect 3797 2217 3813 2227
rect 1987 2197 2013 2203
rect 2207 2197 2233 2203
rect 2247 2197 2273 2203
rect 3367 2197 3433 2203
rect 3557 2203 3563 2217
rect 3800 2213 3813 2217
rect 5267 2217 5283 2227
rect 6057 2227 6063 2253
rect 6057 2217 6073 2227
rect 5267 2213 5280 2217
rect 6060 2213 6073 2217
rect 6197 2223 6203 2253
rect 6167 2217 6203 2223
rect 3557 2197 3593 2203
rect 4507 2197 4593 2203
rect 5087 2197 5193 2203
rect 5407 2197 5513 2203
rect 6027 2197 6093 2203
rect 967 2177 1013 2183
rect 1027 2177 1093 2183
rect 5607 2177 5673 2183
rect 2967 2157 2993 2163
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 2847 2017 2893 2023
rect 197 1977 253 1983
rect 197 1866 203 1977
rect 467 1977 493 1983
rect 507 1977 573 1983
rect 2347 1977 2373 1983
rect 2477 1977 2533 1983
rect 760 1963 773 1967
rect 757 1953 773 1963
rect 907 1963 920 1967
rect 907 1953 923 1963
rect 1767 1963 1780 1967
rect 1767 1953 1783 1963
rect 633 1927 647 1933
rect 627 1920 647 1927
rect 757 1927 763 1953
rect 917 1927 923 1953
rect 1777 1927 1783 1953
rect 2157 1957 2193 1963
rect 2157 1927 2163 1957
rect 627 1917 643 1920
rect 757 1917 773 1927
rect 627 1913 640 1917
rect 760 1913 773 1917
rect 907 1917 923 1927
rect 907 1913 920 1917
rect 1307 1917 1333 1923
rect 1767 1917 1783 1927
rect 1767 1913 1780 1917
rect 2147 1917 2163 1927
rect 2147 1913 2160 1917
rect 2477 1906 2483 1977
rect 5867 1977 5933 1983
rect 5947 1977 5973 1983
rect 6080 1983 6093 1987
rect 6077 1973 6093 1983
rect 6147 1977 6183 1983
rect 3760 1963 3773 1967
rect 3757 1953 3773 1963
rect 6077 1963 6083 1973
rect 6057 1957 6083 1963
rect 6177 1963 6183 1977
rect 6177 1957 6203 1963
rect 3757 1923 3763 1953
rect 6057 1927 6063 1957
rect 6197 1927 6203 1957
rect 3727 1917 3763 1923
rect 5367 1917 5393 1923
rect 6047 1917 6063 1927
rect 6047 1913 6060 1917
rect 6187 1917 6203 1927
rect 6187 1913 6200 1917
rect 4587 1897 4613 1903
rect 6323 1838 6383 2342
rect 6290 1822 6383 1838
rect 1667 1757 1713 1763
rect 4447 1757 4493 1763
rect 4847 1757 4913 1763
rect 5707 1757 5753 1763
rect 187 1743 200 1747
rect 187 1733 203 1743
rect 1307 1743 1320 1747
rect 1460 1743 1473 1747
rect 1307 1733 1323 1743
rect 197 1707 203 1733
rect 187 1697 203 1707
rect 1317 1703 1323 1733
rect 1297 1697 1323 1703
rect 1457 1733 1473 1743
rect 1720 1743 1733 1747
rect 1717 1733 1733 1743
rect 3840 1743 3853 1747
rect 3837 1733 3853 1743
rect 5447 1737 5473 1743
rect 6100 1743 6113 1747
rect 6097 1733 6113 1743
rect 6240 1743 6253 1747
rect 6237 1733 6253 1743
rect 1457 1707 1463 1733
rect 1717 1707 1723 1733
rect 3837 1727 3843 1733
rect 3820 1726 3843 1727
rect 3827 1717 3843 1726
rect 3827 1713 3840 1717
rect 6077 1707 6083 1733
rect 1457 1697 1473 1707
rect 187 1693 200 1697
rect 1297 1687 1303 1697
rect 1460 1693 1473 1697
rect 1717 1697 1733 1707
rect 1720 1693 1733 1697
rect 6067 1697 6083 1707
rect 6097 1707 6103 1733
rect 6237 1707 6243 1733
rect 6097 1697 6113 1707
rect 6067 1693 6080 1697
rect 6100 1693 6113 1697
rect 6237 1697 6253 1707
rect 6240 1693 6253 1697
rect 407 1677 433 1683
rect 1287 1677 1303 1687
rect 1287 1673 1300 1677
rect 2187 1677 2273 1683
rect 3667 1677 3733 1683
rect 4587 1677 4613 1683
rect 5567 1677 5613 1683
rect 5907 1657 6013 1663
rect 2007 1597 2033 1603
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 2047 1537 2093 1543
rect 1773 1467 1787 1473
rect 787 1457 893 1463
rect 1773 1460 1793 1467
rect 1777 1457 1793 1460
rect 1780 1453 1793 1457
rect 1867 1457 1953 1463
rect 2587 1457 2633 1463
rect 4667 1457 4773 1463
rect 4847 1457 4873 1463
rect 5007 1457 5073 1463
rect 1400 1443 1413 1447
rect 1397 1433 1413 1443
rect 1540 1443 1553 1447
rect 1537 1433 1553 1443
rect 2047 1443 2060 1447
rect 3480 1443 3493 1447
rect 2047 1433 2063 1443
rect 1397 1407 1403 1433
rect 1537 1407 1543 1433
rect 2057 1407 2063 1433
rect 3477 1433 3493 1443
rect 4160 1443 4173 1447
rect 4157 1433 4173 1443
rect 4267 1443 4280 1447
rect 4540 1443 4553 1447
rect 4267 1433 4283 1443
rect 1397 1397 1413 1407
rect 1400 1393 1413 1397
rect 1527 1397 1543 1407
rect 1527 1393 1540 1397
rect 2047 1397 2063 1407
rect 2047 1393 2060 1397
rect 3477 1403 3483 1433
rect 3447 1397 3483 1403
rect 4157 1407 4163 1433
rect 4157 1397 4173 1407
rect 4160 1393 4173 1397
rect 4277 1403 4283 1433
rect 4537 1433 4553 1443
rect 4687 1437 4713 1443
rect 5720 1443 5733 1447
rect 5717 1433 5733 1443
rect 5847 1443 5860 1447
rect 5880 1443 5893 1447
rect 5847 1433 5863 1443
rect 4537 1403 4543 1433
rect 5717 1407 5723 1433
rect 5857 1407 5863 1433
rect 4277 1400 4303 1403
rect 4277 1397 4307 1400
rect 4537 1397 4563 1403
rect 5717 1397 5733 1407
rect 4293 1387 4307 1397
rect 3827 1377 3853 1383
rect 4007 1377 4053 1383
rect 4557 1383 4563 1397
rect 5720 1393 5733 1397
rect 5847 1397 5863 1407
rect 5877 1433 5893 1443
rect 6020 1443 6033 1447
rect 6017 1433 6033 1443
rect 5877 1403 5883 1433
rect 6017 1407 6023 1433
rect 5877 1397 5903 1403
rect 6017 1397 6033 1407
rect 5847 1393 5860 1397
rect 4557 1377 4593 1383
rect 5897 1363 5903 1397
rect 6020 1393 6033 1397
rect 6157 1387 6163 1473
rect 6147 1377 6163 1387
rect 6147 1373 6160 1377
rect 5867 1357 5903 1363
rect 6323 1318 6383 1822
rect 6290 1302 6383 1318
rect 2397 1260 2453 1263
rect 2393 1257 2453 1260
rect 207 1237 273 1243
rect 347 1223 360 1227
rect 347 1213 363 1223
rect 1227 1223 1240 1227
rect 1227 1213 1243 1223
rect 1387 1217 1413 1223
rect 1967 1223 1980 1227
rect 1967 1213 1983 1223
rect 357 1187 363 1213
rect 347 1177 363 1187
rect 347 1173 360 1177
rect 207 1157 273 1163
rect 1237 1163 1243 1213
rect 1977 1183 1983 1213
rect 2297 1223 2303 1253
rect 2393 1247 2407 1257
rect 2787 1237 2853 1243
rect 4607 1237 4653 1243
rect 4967 1237 5013 1243
rect 2247 1217 2303 1223
rect 2567 1223 2580 1227
rect 2700 1223 2713 1227
rect 2567 1213 2583 1223
rect 2577 1187 2583 1213
rect 2697 1213 2713 1223
rect 3020 1223 3033 1227
rect 3017 1213 3033 1223
rect 3320 1223 3333 1227
rect 3317 1213 3333 1223
rect 3880 1223 3893 1227
rect 3877 1213 3893 1223
rect 5600 1223 5613 1227
rect 5287 1217 5323 1223
rect 1957 1177 1983 1183
rect 1957 1167 1963 1177
rect 2567 1177 2583 1187
rect 2567 1173 2580 1177
rect 2697 1183 2703 1213
rect 2667 1177 2703 1183
rect 3017 1187 3023 1213
rect 3317 1187 3323 1213
rect 3017 1177 3033 1187
rect 3020 1173 3033 1177
rect 3307 1177 3323 1187
rect 3877 1187 3883 1213
rect 3877 1177 3893 1187
rect 3307 1173 3320 1177
rect 3880 1173 3893 1177
rect 4987 1177 5033 1183
rect 5317 1183 5323 1217
rect 5597 1213 5613 1223
rect 5760 1223 5773 1227
rect 5757 1213 5773 1223
rect 5597 1187 5603 1213
rect 5317 1180 5343 1183
rect 5317 1177 5347 1180
rect 5333 1167 5347 1177
rect 5587 1177 5603 1187
rect 5757 1187 5763 1213
rect 6037 1187 6043 1233
rect 6200 1223 6213 1227
rect 6197 1213 6213 1223
rect 6197 1187 6203 1213
rect 5757 1177 5773 1187
rect 5587 1173 5600 1177
rect 5760 1173 5773 1177
rect 6037 1177 6053 1187
rect 6040 1173 6053 1177
rect 6197 1177 6213 1187
rect 6200 1173 6213 1177
rect 1237 1157 1293 1163
rect 1787 1157 1873 1163
rect 1940 1165 1963 1167
rect 1947 1157 1963 1165
rect 1947 1153 1960 1157
rect 2407 1157 2493 1163
rect 2687 1157 2713 1163
rect 3127 1157 3153 1163
rect 3547 1157 3653 1163
rect 4847 1157 4913 1163
rect 5027 1157 5053 1163
rect 5827 1157 5893 1163
rect 1847 1137 1893 1143
rect 4967 1137 5033 1143
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 5487 1017 5513 1023
rect 5167 977 5233 983
rect 207 937 293 943
rect 447 937 533 943
rect 1667 937 1753 943
rect 1827 937 1853 943
rect 2247 943 2260 947
rect 2247 933 2263 943
rect 220 923 233 927
rect 217 913 233 923
rect 380 923 393 927
rect 377 913 393 923
rect 2257 923 2263 933
rect 2827 937 2893 943
rect 3087 937 3173 943
rect 3957 937 4013 943
rect 2460 923 2473 927
rect 2257 917 2283 923
rect 217 883 223 913
rect 187 877 223 883
rect 377 887 383 913
rect 377 877 393 887
rect 380 873 393 877
rect 2153 867 2167 873
rect 2140 866 2167 867
rect 2147 860 2167 866
rect 2147 857 2163 860
rect 2147 853 2160 857
rect 2277 863 2283 917
rect 2457 913 2473 923
rect 2967 917 3013 923
rect 3127 923 3140 927
rect 3957 923 3963 937
rect 5697 937 5733 943
rect 5697 923 5703 937
rect 6127 937 6173 943
rect 6187 937 6233 943
rect 3127 920 3143 923
rect 3127 913 3147 920
rect 2457 887 2463 913
rect 3133 906 3147 913
rect 3937 917 3963 923
rect 5677 917 5703 923
rect 2457 877 2473 887
rect 2460 873 2473 877
rect 2867 877 2893 883
rect 3937 883 3943 917
rect 3907 877 3943 883
rect 5677 883 5683 917
rect 5967 923 5980 927
rect 6180 923 6193 927
rect 5967 913 5983 923
rect 5977 883 5983 913
rect 5647 877 5683 883
rect 5957 877 5983 883
rect 6177 913 6193 923
rect 6177 887 6183 913
rect 6177 877 6193 887
rect 2247 857 2283 863
rect 2447 857 2493 863
rect 4387 857 4453 863
rect 5957 847 5963 877
rect 6180 873 6193 877
rect 5987 857 6033 863
rect 2247 837 2313 843
rect 5957 846 5980 847
rect 5957 837 5973 846
rect 5960 833 5973 837
rect 1347 817 1393 823
rect 6323 798 6383 1302
rect 6290 782 6383 798
rect 1527 757 1573 763
rect 5907 714 5913 727
rect 5907 713 5920 714
rect 767 697 793 703
rect 940 703 953 707
rect 937 693 953 703
rect 1847 697 1873 703
rect 2007 703 2020 707
rect 2007 693 2023 703
rect 2707 703 2720 707
rect 2707 693 2723 703
rect 4647 703 4660 707
rect 4647 693 4663 703
rect 5087 697 5123 703
rect 937 667 943 693
rect 927 657 943 667
rect 2017 663 2023 693
rect 2717 666 2723 693
rect 4657 667 4663 693
rect 1997 660 2023 663
rect 1993 657 2023 660
rect 927 653 940 657
rect 1993 647 2007 657
rect 4647 657 4663 667
rect 5117 667 5123 697
rect 5227 697 5253 703
rect 5540 703 5553 707
rect 5537 693 5553 703
rect 5687 697 5713 703
rect 5537 667 5543 693
rect 5117 657 5133 667
rect 4647 653 4660 657
rect 5120 653 5133 657
rect 5537 657 5553 667
rect 5540 653 5553 657
rect 187 637 253 643
rect 887 637 933 643
rect 1287 637 1333 643
rect 1707 637 1773 643
rect 1827 637 1953 643
rect 2647 637 2753 643
rect 3787 637 3873 643
rect 4287 637 4353 643
rect 5667 637 5713 643
rect -63 522 30 538
rect -63 18 -3 522
rect 1047 457 1073 463
rect 127 417 233 423
rect 1027 417 1073 423
rect 1837 417 1893 423
rect 1207 403 1220 407
rect 1837 403 1843 417
rect 1947 417 1993 423
rect 2047 417 2173 423
rect 3007 417 3113 423
rect 4047 417 4073 423
rect 5867 417 5893 423
rect 6027 417 6073 423
rect 2400 403 2413 407
rect 1207 393 1223 403
rect 1217 367 1223 393
rect 1817 397 1843 403
rect 1817 363 1823 397
rect 2397 393 2413 403
rect 2880 403 2893 407
rect 2877 393 2893 403
rect 3327 403 3340 407
rect 3660 403 3673 407
rect 3327 393 3343 403
rect 2397 367 2403 393
rect 2853 367 2867 373
rect 1787 357 1823 363
rect 2387 357 2403 367
rect 2387 353 2400 357
rect 2847 360 2867 367
rect 2877 367 2883 393
rect 3337 367 3343 393
rect 3657 393 3673 403
rect 4487 397 4513 403
rect 5767 403 5780 407
rect 5767 393 5783 403
rect 2847 357 2863 360
rect 2877 357 2893 367
rect 2847 353 2860 357
rect 2880 353 2893 357
rect 3327 357 3343 367
rect 3327 353 3340 357
rect 3657 363 3663 393
rect 3627 357 3663 363
rect 3747 357 3773 363
rect 5777 366 5783 393
rect 5327 337 5393 343
rect 3747 297 3773 303
rect 6323 278 6383 782
rect 6290 262 6383 278
rect 3127 217 3173 223
rect 197 197 253 203
rect 197 147 203 197
rect 507 197 573 203
rect 1067 197 1133 203
rect 4087 197 4113 203
rect 4227 197 4333 203
rect 1187 177 1223 183
rect 187 137 203 147
rect 1217 147 1223 177
rect 1507 177 1533 183
rect 1733 183 1747 193
rect 1733 180 1783 183
rect 1737 177 1783 180
rect 1353 147 1367 153
rect 1777 147 1783 177
rect 2067 183 2080 187
rect 2220 183 2233 187
rect 2067 173 2083 183
rect 2077 147 2083 173
rect 2217 173 2233 183
rect 4067 177 4093 183
rect 2217 147 2223 173
rect 1217 137 1233 147
rect 187 133 200 137
rect 1220 133 1233 137
rect 1353 140 1373 147
rect 1357 137 1373 140
rect 1360 133 1373 137
rect 1777 137 1793 147
rect 1780 133 1793 137
rect 2077 137 2093 147
rect 2080 133 2093 137
rect 2207 137 2223 147
rect 2207 133 2220 137
rect 207 117 273 123
rect 427 117 493 123
rect 987 117 1053 123
rect 1367 117 1413 123
rect 1527 117 1593 123
rect 1867 117 1933 123
rect 2007 117 2153 123
rect 2327 117 2373 123
rect 2387 117 2433 123
rect 2927 117 3073 123
rect 3327 117 3393 123
rect 3947 117 3973 123
rect 5267 117 5333 123
rect 5467 117 5513 123
rect 2487 97 2533 103
rect 3307 97 3353 103
rect 4407 93 4413 107
rect 5407 97 5493 103
rect 2347 57 2373 63
rect 1487 37 1513 43
rect -63 2 30 18
rect 6323 2 6383 262
<< m2contact >>
rect 2653 6253 2667 6267
rect 3253 6253 3267 6267
rect 3433 6253 3447 6267
rect 4033 6253 4047 6267
rect 5133 6253 5147 6267
rect 513 6133 527 6147
rect 593 6133 607 6147
rect 5813 6133 5827 6147
rect 5853 6133 5867 6147
rect 893 6113 907 6127
rect 1333 6113 1347 6127
rect 1373 6113 1387 6127
rect 5373 6113 5387 6127
rect 5413 6113 5427 6127
rect 1593 6073 1607 6087
rect 1633 6073 1647 6087
rect 933 6053 947 6067
rect 893 6033 907 6047
rect 913 6032 927 6046
rect 1893 5913 1907 5927
rect 1933 5913 1947 5927
rect 5533 5913 5547 5927
rect 5613 5914 5627 5928
rect 853 5893 867 5907
rect 5233 5893 5247 5907
rect 813 5853 827 5867
rect 5233 5853 5247 5867
rect 133 5833 147 5847
rect 173 5833 187 5847
rect 1333 5813 1347 5827
rect 1413 5813 1427 5827
rect 3433 5713 3447 5727
rect 3973 5713 3987 5727
rect 4833 5713 4847 5727
rect 6093 5713 6107 5727
rect 353 5613 367 5627
rect 393 5613 407 5627
rect 3693 5613 3707 5627
rect 3753 5613 3767 5627
rect 4633 5613 4647 5627
rect 4673 5613 4687 5627
rect 4713 5613 4727 5627
rect 173 5593 187 5607
rect 213 5593 227 5607
rect 793 5593 807 5607
rect 2813 5593 2827 5607
rect 2933 5593 2947 5607
rect 2973 5593 2987 5607
rect 3813 5593 3827 5607
rect 213 5553 227 5567
rect 753 5553 767 5567
rect 3813 5553 3827 5567
rect 4093 5593 4107 5607
rect 4093 5553 4107 5567
rect 193 5533 207 5547
rect 2313 5533 2327 5547
rect 2373 5532 2387 5546
rect 2593 5533 2607 5547
rect 2653 5533 2667 5547
rect 2733 5531 2747 5545
rect 2773 5533 2787 5547
rect 2853 5531 2867 5545
rect 213 5512 227 5526
rect 1793 5513 1807 5527
rect 1853 5513 1867 5527
rect 2633 5513 2647 5527
rect 2673 5493 2687 5507
rect 4373 5393 4387 5407
rect 3473 5373 3487 5387
rect 3573 5373 3587 5387
rect 3813 5373 3827 5387
rect 4413 5373 4427 5387
rect 3473 5333 3487 5347
rect 133 5313 147 5327
rect 173 5313 187 5327
rect 213 5313 227 5327
rect 293 5313 307 5327
rect 733 5313 747 5327
rect 773 5313 787 5327
rect 3413 5313 3427 5327
rect 3513 5311 3527 5325
rect 3593 5312 3607 5326
rect 3853 5312 3867 5326
rect 2913 5193 2927 5207
rect 4493 5193 4507 5207
rect 5493 5193 5507 5207
rect 5633 5193 5647 5207
rect 4053 5113 4067 5127
rect 2093 5093 2107 5107
rect 2233 5093 2247 5107
rect 2573 5093 2587 5107
rect 2653 5093 2667 5107
rect 2733 5093 2747 5107
rect 2793 5093 2807 5107
rect 4153 5093 4167 5107
rect 5153 5093 5167 5107
rect 5213 5094 5227 5108
rect 5293 5093 5307 5107
rect 5373 5093 5387 5107
rect 5913 5093 5927 5107
rect 6013 5093 6027 5107
rect 633 5073 647 5087
rect 773 5073 787 5087
rect 913 5073 927 5087
rect 1993 5073 2007 5087
rect 93 5013 107 5027
rect 173 5013 187 5027
rect 773 5033 787 5047
rect 873 5033 887 5047
rect 2393 5053 2407 5067
rect 2953 5073 2967 5087
rect 4093 5073 4107 5087
rect 4233 5073 4247 5087
rect 2053 5033 2067 5047
rect 2433 5033 2447 5047
rect 2553 5033 2567 5047
rect 2633 5033 2647 5047
rect 2913 5033 2927 5047
rect 4093 5033 4107 5047
rect 4233 5033 4247 5047
rect 5113 5033 5127 5047
rect 5173 5033 5187 5047
rect 653 5013 667 5027
rect 5273 5013 5287 5027
rect 5373 5013 5387 5027
rect 5793 5013 5807 5027
rect 5853 5013 5867 5027
rect 4893 4913 4907 4927
rect 1893 4893 1907 4907
rect 4973 4893 4987 4907
rect 5013 4893 5027 4907
rect 5053 4893 5067 4907
rect 773 4853 787 4867
rect 813 4853 827 4867
rect 1933 4873 1947 4887
rect 1993 4873 2007 4887
rect 2033 4873 2047 4887
rect 2093 4873 2107 4887
rect 3573 4873 3587 4887
rect 4853 4873 4867 4887
rect 4953 4873 4967 4887
rect 6053 4873 6067 4887
rect 6093 4873 6107 4887
rect 733 4791 747 4805
rect 813 4793 827 4807
rect 1073 4793 1087 4807
rect 1133 4793 1147 4807
rect 1293 4793 1307 4807
rect 1373 4793 1387 4807
rect 2133 4852 2147 4866
rect 2233 4853 2247 4867
rect 2673 4853 2687 4867
rect 1953 4813 1967 4827
rect 2273 4813 2287 4827
rect 2733 4813 2747 4827
rect 3613 4813 3627 4827
rect 1893 4793 1907 4807
rect 5233 4791 5247 4805
rect 5273 4793 5287 4807
rect 5373 4793 5387 4807
rect 5433 4793 5447 4807
rect 5513 4791 5527 4805
rect 2073 4773 2087 4787
rect 2173 4773 2187 4787
rect 5553 4773 5567 4787
rect 5613 4773 5627 4787
rect 2673 4753 2687 4767
rect 2713 4752 2727 4766
rect 4573 4753 4587 4767
rect 4613 4753 4627 4767
rect 2833 4733 2847 4747
rect 2893 4713 2907 4727
rect 2593 4673 2607 4687
rect 3333 4673 3347 4687
rect 3653 4673 3667 4687
rect 1273 4632 1287 4646
rect 1313 4633 1327 4647
rect 2793 4633 2807 4647
rect 2733 4593 2747 4607
rect 533 4573 547 4587
rect 613 4573 627 4587
rect 813 4573 827 4587
rect 893 4573 907 4587
rect 1293 4573 1307 4587
rect 1353 4573 1367 4587
rect 1833 4574 1847 4588
rect 1313 4553 1327 4567
rect 1433 4553 1447 4567
rect 1233 4493 1247 4507
rect 1413 4493 1427 4507
rect 2813 4573 2827 4587
rect 1873 4553 1887 4567
rect 1913 4553 1927 4567
rect 2033 4553 2047 4567
rect 2793 4513 2807 4527
rect 1853 4492 1867 4506
rect 2033 4493 2047 4507
rect 4033 4573 4047 4587
rect 4013 4553 4027 4567
rect 5953 4553 5967 4567
rect 6033 4553 6047 4567
rect 4013 4513 4027 4527
rect 5633 4513 5647 4527
rect 5673 4513 5687 4527
rect 5893 4513 5907 4527
rect 3973 4492 3987 4506
rect 6013 4493 6027 4507
rect 3853 4473 3867 4487
rect 3913 4473 3927 4487
rect 753 4373 767 4387
rect 793 4373 807 4387
rect 773 4353 787 4367
rect 833 4353 847 4367
rect 893 4333 907 4347
rect 953 4333 967 4347
rect 1093 4333 1107 4347
rect 4593 4333 4607 4347
rect 3993 4313 4007 4327
rect 1093 4293 1107 4307
rect 3233 4293 3247 4307
rect 3293 4293 3307 4307
rect 4033 4293 4047 4307
rect 4553 4293 4567 4307
rect 5313 4293 5327 4307
rect 5373 4293 5387 4307
rect 413 4273 427 4287
rect 473 4273 487 4287
rect 3973 4273 3987 4287
rect 4013 4272 4027 4286
rect 4413 4273 4427 4287
rect 4473 4273 4487 4287
rect 5873 4273 5887 4287
rect 5953 4273 5967 4287
rect 6193 4273 6207 4287
rect 6253 4273 6267 4287
rect 3293 4173 3307 4187
rect 2513 4153 2527 4167
rect 2773 4153 2787 4167
rect 3873 4153 3887 4167
rect 3893 4153 3907 4167
rect 4473 4153 4487 4167
rect 3853 4133 3867 4147
rect 3913 4133 3927 4147
rect 4733 4133 4747 4147
rect 153 4073 167 4087
rect 213 4073 227 4087
rect 1373 4073 1387 4087
rect 1453 4073 1467 4087
rect 133 4053 147 4067
rect 173 4052 187 4066
rect 253 4054 267 4068
rect 333 4053 347 4067
rect 393 4052 407 4066
rect 593 4053 607 4067
rect 2753 4053 2767 4067
rect 2873 4054 2887 4068
rect 4173 4053 4187 4067
rect 4233 4053 4247 4067
rect 4473 4053 4487 4067
rect 4553 4054 4567 4068
rect 5233 4053 5247 4067
rect 5333 4053 5347 4067
rect 73 4033 87 4047
rect 453 4033 467 4047
rect 713 4033 727 4047
rect 1133 4033 1147 4047
rect 1233 4033 1247 4047
rect 1393 4033 1407 4047
rect 73 3993 87 4007
rect 513 3993 527 4007
rect 573 3993 587 4007
rect 733 3993 747 4007
rect 1093 3993 1107 4007
rect 1233 3993 1247 4007
rect 1553 4033 1567 4047
rect 1893 4033 1907 4047
rect 1953 4033 1967 4047
rect 1453 3993 1467 4007
rect 1553 3993 1567 4007
rect 1833 3993 1847 4007
rect 2253 4033 2267 4047
rect 4073 4033 4087 4047
rect 4373 4033 4387 4047
rect 5733 4033 5747 4047
rect 5793 4033 5807 4047
rect 1993 3993 2007 4007
rect 2773 3993 2787 4007
rect 2833 3993 2847 4007
rect 4073 3993 4087 4007
rect 4373 3993 4387 4007
rect 5733 3993 5747 4007
rect 5793 3993 5807 4007
rect 1673 3973 1687 3987
rect 1773 3973 1787 3987
rect 2193 3973 2207 3987
rect 6073 3971 6087 3985
rect 6233 3973 6247 3987
rect 5773 3952 5787 3966
rect 5833 3953 5847 3967
rect 5673 3933 5687 3947
rect 5733 3933 5747 3947
rect 3853 3853 3867 3867
rect 3933 3853 3947 3867
rect 293 3833 307 3847
rect 333 3833 347 3847
rect 453 3833 467 3847
rect 1313 3833 1327 3847
rect 553 3813 567 3827
rect 433 3773 447 3787
rect 1293 3813 1307 3827
rect 853 3793 867 3807
rect 613 3773 627 3787
rect 813 3773 827 3787
rect 973 3773 987 3787
rect 1013 3773 1027 3787
rect 253 3753 267 3767
rect 333 3753 347 3767
rect 833 3753 847 3767
rect 893 3753 907 3767
rect 1273 3751 1287 3765
rect 3733 3832 3747 3846
rect 3793 3833 3807 3847
rect 5073 3833 5087 3847
rect 5133 3833 5147 3847
rect 2133 3813 2147 3827
rect 2973 3813 2987 3827
rect 1833 3793 1847 3807
rect 1353 3773 1367 3787
rect 1513 3773 1527 3787
rect 3013 3793 3027 3807
rect 5533 3813 5547 3827
rect 1873 3773 1887 3787
rect 2113 3773 2127 3787
rect 1453 3733 1467 3747
rect 2713 3773 2727 3787
rect 2673 3752 2687 3766
rect 3873 3753 3887 3767
rect 3933 3753 3947 3767
rect 4353 3753 4367 3767
rect 4413 3753 4427 3767
rect 5353 3753 5367 3767
rect 5453 3753 5467 3767
rect 5553 3753 5567 3767
rect 5633 3753 5647 3767
rect 5733 3753 5747 3767
rect 1492 3713 1506 3727
rect 1513 3713 1527 3727
rect 2673 3613 2687 3627
rect 2733 3613 2747 3627
rect 2673 3553 2687 3567
rect 533 3533 547 3547
rect 1413 3533 1427 3547
rect 1453 3533 1467 3547
rect 713 3513 727 3527
rect 873 3513 887 3527
rect 973 3513 987 3527
rect 453 3453 467 3467
rect 753 3473 767 3487
rect 873 3473 887 3487
rect 653 3453 667 3467
rect 1033 3513 1047 3527
rect 1253 3513 1267 3527
rect 1673 3513 1687 3527
rect 1793 3513 1807 3527
rect 1893 3533 1907 3547
rect 2753 3534 2767 3548
rect 4513 3533 4527 3547
rect 4593 3533 4607 3547
rect 5873 3533 5887 3547
rect 5913 3533 5927 3547
rect 5973 3533 5987 3547
rect 1033 3473 1047 3487
rect 1253 3473 1267 3487
rect 1053 3451 1067 3465
rect 393 3433 407 3447
rect 1553 3473 1567 3487
rect 1713 3473 1727 3487
rect 1793 3473 1807 3487
rect 2073 3513 2087 3527
rect 1853 3473 1867 3487
rect 2073 3473 2087 3487
rect 2733 3513 2747 3527
rect 4413 3513 4427 3527
rect 4833 3513 4847 3527
rect 4993 3513 5007 3527
rect 2673 3472 2687 3486
rect 4453 3473 4467 3487
rect 5033 3473 5047 3487
rect 4833 3453 4847 3467
rect 5093 3452 5107 3466
rect 5133 3453 5147 3467
rect 6133 3453 6147 3467
rect 6173 3452 6187 3466
rect 1553 3433 1567 3447
rect 1953 3333 1967 3347
rect 1993 3333 2007 3347
rect 913 3313 927 3327
rect 953 3313 967 3327
rect 1173 3313 1187 3327
rect 2193 3313 2207 3327
rect 2253 3313 2267 3327
rect 3213 3313 3227 3327
rect 3293 3313 3307 3327
rect 4253 3313 4267 3327
rect 4833 3313 4847 3327
rect 4933 3313 4947 3327
rect 5713 3313 5727 3327
rect 353 3293 367 3307
rect 433 3293 447 3307
rect 473 3293 487 3307
rect 293 3253 307 3267
rect 1713 3293 1727 3307
rect 2133 3293 2147 3307
rect 4033 3293 4047 3307
rect 413 3233 427 3247
rect 553 3233 567 3247
rect 873 3233 887 3247
rect 973 3233 987 3247
rect 1713 3253 1727 3267
rect 2093 3253 2107 3267
rect 4093 3253 4107 3267
rect 4193 3253 4207 3267
rect 6033 3293 6047 3307
rect 5733 3253 5747 3267
rect 5893 3253 5907 3267
rect 5933 3253 5947 3267
rect 1293 3233 1307 3247
rect 2513 3231 2527 3245
rect 2613 3233 2627 3247
rect 4833 3233 4847 3247
rect 4953 3233 4967 3247
rect 5473 3233 5487 3247
rect 5533 3233 5547 3247
rect 5773 3233 5787 3247
rect 5833 3233 5847 3247
rect 6013 3233 6027 3247
rect 6173 3253 6187 3267
rect 6213 3253 6227 3267
rect 6213 3232 6227 3246
rect 6253 3233 6267 3247
rect 753 3213 767 3227
rect 813 3213 827 3227
rect 2193 3213 2207 3227
rect 2293 3213 2307 3227
rect 2473 3113 2487 3127
rect 3293 3113 3307 3127
rect 2873 3093 2887 3107
rect 1533 3033 1547 3047
rect 1633 3033 1647 3047
rect 5293 3033 5307 3047
rect 5373 3032 5387 3046
rect 553 3013 567 3027
rect 593 3013 607 3027
rect 333 2992 347 3006
rect 953 2993 967 3007
rect 1593 2993 1607 3007
rect 1693 3013 1707 3027
rect 1873 3013 1887 3027
rect 1933 3013 1947 3027
rect 2733 3013 2747 3027
rect 2773 3013 2787 3027
rect 2933 3013 2947 3027
rect 5333 3013 5347 3027
rect 5413 3013 5427 3027
rect 173 2953 187 2967
rect 213 2953 227 2967
rect 333 2953 347 2967
rect 893 2953 907 2967
rect 3213 2993 3227 3007
rect 3913 2993 3927 3007
rect 4853 2993 4867 3007
rect 1653 2953 1667 2967
rect 2933 2953 2947 2967
rect 3153 2952 3167 2966
rect 3913 2953 3927 2967
rect 4853 2953 4867 2967
rect 5073 2993 5087 3007
rect 5193 2993 5207 3007
rect 5553 3013 5567 3027
rect 5793 3013 5807 3027
rect 5833 3013 5847 3027
rect 5593 2993 5607 3007
rect 5073 2953 5087 2967
rect 5193 2953 5207 2967
rect 5453 2953 5467 2967
rect 5653 2993 5667 3007
rect 5753 2993 5767 3007
rect 5993 3013 6007 3027
rect 6133 3013 6147 3027
rect 6233 3013 6247 3027
rect 5653 2953 5667 2967
rect 6193 2993 6207 3007
rect 5813 2953 5827 2967
rect 5953 2953 5967 2967
rect 1593 2933 1607 2947
rect 4193 2931 4207 2945
rect 4253 2933 4267 2947
rect 5613 2933 5627 2947
rect 6213 2933 6227 2947
rect 1373 2793 1387 2807
rect 1453 2793 1467 2807
rect 1653 2793 1667 2807
rect 1693 2793 1707 2807
rect 2453 2773 2467 2787
rect 3193 2773 3207 2787
rect 2453 2733 2467 2747
rect 3253 2773 3267 2787
rect 3373 2773 3387 2787
rect 3233 2752 3247 2766
rect 2813 2713 2827 2727
rect 2953 2713 2967 2727
rect 3153 2713 3167 2727
rect 3373 2733 3387 2747
rect 3433 2773 3447 2787
rect 3553 2773 3567 2787
rect 3653 2773 3667 2787
rect 6213 2773 6227 2787
rect 3433 2733 3447 2747
rect 3553 2733 3567 2747
rect 3713 2733 3727 2747
rect 6153 2733 6167 2747
rect 3493 2713 3507 2727
rect 3573 2713 3587 2727
rect 3893 2711 3907 2725
rect 3953 2713 3967 2727
rect 4633 2713 4647 2727
rect 4713 2713 4727 2727
rect 5133 2713 5147 2727
rect 5233 2713 5247 2727
rect 5973 2713 5987 2727
rect 6033 2713 6047 2727
rect 5553 2693 5567 2707
rect 5633 2693 5647 2707
rect 3893 2673 3907 2687
rect 3973 2673 3987 2687
rect 2873 2533 2887 2547
rect 2953 2533 2967 2547
rect 2873 2512 2887 2526
rect 2913 2513 2927 2527
rect 973 2493 987 2507
rect 1013 2493 1027 2507
rect 1573 2493 1587 2507
rect 1653 2493 1667 2507
rect 3353 2493 3367 2507
rect 3433 2493 3447 2507
rect 4073 2493 4087 2507
rect 4173 2493 4187 2507
rect 5593 2493 5607 2507
rect 5653 2493 5667 2507
rect 6153 2492 6167 2506
rect 6233 2493 6247 2507
rect 2193 2473 2207 2487
rect 2293 2473 2307 2487
rect 3373 2473 3387 2487
rect 3793 2473 3807 2487
rect 2193 2433 2207 2447
rect 1453 2413 1467 2427
rect 1493 2413 1507 2427
rect 2233 2413 2247 2427
rect 3253 2433 3267 2447
rect 3413 2433 3427 2447
rect 3213 2413 3227 2427
rect 5793 2473 5807 2487
rect 5953 2473 5967 2487
rect 6053 2473 6067 2487
rect 5733 2433 5747 2447
rect 5953 2433 5967 2447
rect 6113 2433 6127 2447
rect 3833 2392 3847 2406
rect 6253 2393 6267 2407
rect 6293 2392 6307 2406
rect 3873 2293 3887 2307
rect 3953 2293 3967 2307
rect 1273 2273 1287 2287
rect 1353 2273 1367 2287
rect 2253 2273 2267 2287
rect 2313 2274 2327 2288
rect 3253 2273 3267 2287
rect 3533 2273 3547 2287
rect 3833 2274 3847 2288
rect 2953 2253 2967 2267
rect 3113 2252 3127 2266
rect 3153 2253 3167 2267
rect 3293 2253 3307 2267
rect 2993 2212 3007 2226
rect 5293 2253 5307 2267
rect 6073 2253 6087 2267
rect 6213 2253 6227 2267
rect 1973 2193 1987 2207
rect 2013 2193 2027 2207
rect 2193 2193 2207 2207
rect 2233 2193 2247 2207
rect 2273 2193 2287 2207
rect 3353 2193 3367 2207
rect 3433 2193 3447 2207
rect 3813 2213 3827 2227
rect 5253 2213 5267 2227
rect 6073 2213 6087 2227
rect 6153 2213 6167 2227
rect 3593 2193 3607 2207
rect 4493 2193 4507 2207
rect 4593 2193 4607 2207
rect 5073 2191 5087 2205
rect 5193 2193 5207 2207
rect 5393 2193 5407 2207
rect 5513 2193 5527 2207
rect 6013 2193 6027 2207
rect 6093 2193 6107 2207
rect 953 2173 967 2187
rect 1013 2173 1027 2187
rect 1093 2173 1107 2187
rect 5593 2173 5607 2187
rect 5673 2173 5687 2187
rect 2953 2152 2967 2166
rect 2993 2153 3007 2167
rect 2833 2013 2847 2027
rect 2893 2013 2907 2027
rect 253 1973 267 1987
rect 453 1973 467 1987
rect 493 1973 507 1987
rect 573 1973 587 1987
rect 2333 1973 2347 1987
rect 2373 1973 2387 1987
rect 773 1953 787 1967
rect 893 1953 907 1967
rect 1753 1953 1767 1967
rect 633 1933 647 1947
rect 613 1913 627 1927
rect 2193 1953 2207 1967
rect 773 1913 787 1927
rect 893 1913 907 1927
rect 1293 1913 1307 1927
rect 1333 1913 1347 1927
rect 1753 1913 1767 1927
rect 2133 1913 2147 1927
rect 2533 1973 2547 1987
rect 5853 1973 5867 1987
rect 5933 1973 5947 1987
rect 5973 1973 5987 1987
rect 6093 1973 6107 1987
rect 6133 1974 6147 1988
rect 3773 1953 3787 1967
rect 3713 1913 3727 1927
rect 5353 1913 5367 1927
rect 5393 1913 5407 1927
rect 6033 1913 6047 1927
rect 6173 1913 6187 1927
rect 2473 1892 2487 1906
rect 4573 1893 4587 1907
rect 4613 1893 4627 1907
rect 193 1852 207 1866
rect 1653 1753 1667 1767
rect 1713 1753 1727 1767
rect 4433 1753 4447 1767
rect 4493 1753 4507 1767
rect 4833 1753 4847 1767
rect 4913 1753 4927 1767
rect 5693 1753 5707 1767
rect 5753 1753 5767 1767
rect 173 1733 187 1747
rect 1293 1733 1307 1747
rect 173 1693 187 1707
rect 1473 1733 1487 1747
rect 1733 1733 1747 1747
rect 3853 1733 3867 1747
rect 5433 1733 5447 1747
rect 5473 1733 5487 1747
rect 6073 1733 6087 1747
rect 6113 1733 6127 1747
rect 6253 1733 6267 1747
rect 3813 1712 3827 1726
rect 1473 1693 1487 1707
rect 1733 1693 1747 1707
rect 6053 1693 6067 1707
rect 6113 1693 6127 1707
rect 6253 1693 6267 1707
rect 393 1673 407 1687
rect 433 1671 447 1685
rect 1273 1673 1287 1687
rect 2173 1673 2187 1687
rect 2273 1673 2287 1687
rect 3653 1673 3667 1687
rect 3733 1673 3747 1687
rect 4573 1673 4587 1687
rect 4613 1673 4627 1687
rect 5553 1671 5567 1685
rect 5613 1673 5627 1687
rect 5893 1653 5907 1667
rect 6013 1653 6027 1667
rect 1993 1592 2007 1606
rect 2033 1593 2047 1607
rect 2033 1533 2047 1547
rect 2093 1533 2107 1547
rect 1773 1473 1787 1487
rect 6153 1473 6167 1487
rect 773 1453 787 1467
rect 893 1453 907 1467
rect 1793 1453 1807 1467
rect 1853 1453 1867 1467
rect 1953 1453 1967 1467
rect 2573 1453 2587 1467
rect 2633 1453 2647 1467
rect 4653 1453 4667 1467
rect 4773 1453 4787 1467
rect 4833 1453 4847 1467
rect 4873 1453 4887 1467
rect 4993 1453 5007 1467
rect 5073 1453 5087 1467
rect 1413 1433 1427 1447
rect 1553 1433 1567 1447
rect 2033 1433 2047 1447
rect 3493 1433 3507 1447
rect 4173 1433 4187 1447
rect 4253 1433 4267 1447
rect 1413 1393 1427 1407
rect 1513 1393 1527 1407
rect 2033 1393 2047 1407
rect 3433 1393 3447 1407
rect 4173 1393 4187 1407
rect 4553 1433 4567 1447
rect 4673 1433 4687 1447
rect 4713 1433 4727 1447
rect 5733 1433 5747 1447
rect 5833 1433 5847 1447
rect 3813 1373 3827 1387
rect 3853 1373 3867 1387
rect 3993 1373 4007 1387
rect 4053 1373 4067 1387
rect 4293 1373 4307 1387
rect 5733 1393 5747 1407
rect 5833 1393 5847 1407
rect 5893 1433 5907 1447
rect 6033 1433 6047 1447
rect 4593 1373 4607 1387
rect 5853 1353 5867 1367
rect 6033 1393 6047 1407
rect 6133 1373 6147 1387
rect 2293 1253 2307 1267
rect 193 1233 207 1247
rect 273 1233 287 1247
rect 333 1213 347 1227
rect 1213 1213 1227 1227
rect 1373 1213 1387 1227
rect 1413 1213 1427 1227
rect 1953 1213 1967 1227
rect 333 1173 347 1187
rect 193 1153 207 1167
rect 273 1153 287 1167
rect 2233 1212 2247 1226
rect 2453 1253 2467 1267
rect 2393 1233 2407 1247
rect 2773 1233 2787 1247
rect 2853 1233 2867 1247
rect 4593 1233 4607 1247
rect 4653 1233 4667 1247
rect 4953 1233 4967 1247
rect 5013 1233 5027 1247
rect 6033 1233 6047 1247
rect 2553 1213 2567 1227
rect 2713 1213 2727 1227
rect 3033 1213 3047 1227
rect 3333 1213 3347 1227
rect 3893 1213 3907 1227
rect 5273 1213 5287 1227
rect 2553 1173 2567 1187
rect 2653 1173 2667 1187
rect 3033 1173 3047 1187
rect 3293 1173 3307 1187
rect 3893 1173 3907 1187
rect 4973 1173 4987 1187
rect 5033 1173 5047 1187
rect 5613 1213 5627 1227
rect 5773 1213 5787 1227
rect 5573 1173 5587 1187
rect 6213 1213 6227 1227
rect 5773 1173 5787 1187
rect 6053 1173 6067 1187
rect 6213 1173 6227 1187
rect 1293 1153 1307 1167
rect 1773 1153 1787 1167
rect 1873 1153 1887 1167
rect 1933 1151 1947 1165
rect 2393 1153 2407 1167
rect 2493 1153 2507 1167
rect 2673 1153 2687 1167
rect 2713 1153 2727 1167
rect 3113 1153 3127 1167
rect 3153 1153 3167 1167
rect 3533 1153 3547 1167
rect 3653 1153 3667 1167
rect 4833 1153 4847 1167
rect 4913 1151 4927 1165
rect 5013 1152 5027 1166
rect 5053 1153 5067 1167
rect 5333 1153 5347 1167
rect 5813 1151 5827 1165
rect 5893 1153 5907 1167
rect 1833 1132 1847 1146
rect 1893 1133 1907 1147
rect 4953 1133 4967 1147
rect 5033 1132 5047 1146
rect 5473 1013 5487 1027
rect 5513 1013 5527 1027
rect 5153 973 5167 987
rect 5233 973 5247 987
rect 193 933 207 947
rect 293 933 307 947
rect 433 933 447 947
rect 533 933 547 947
rect 1653 932 1667 946
rect 1753 933 1767 947
rect 1813 933 1827 947
rect 1853 933 1867 947
rect 2233 933 2247 947
rect 233 913 247 927
rect 393 913 407 927
rect 2813 932 2827 946
rect 2893 933 2907 947
rect 3073 933 3087 947
rect 3173 934 3187 948
rect 173 873 187 887
rect 393 873 407 887
rect 2153 873 2167 887
rect 2133 852 2147 866
rect 2233 853 2247 867
rect 2473 913 2487 927
rect 2953 913 2967 927
rect 3013 913 3027 927
rect 3113 913 3127 927
rect 4013 933 4027 947
rect 5733 933 5747 947
rect 6113 933 6127 947
rect 6173 933 6187 947
rect 6233 933 6247 947
rect 3133 892 3147 906
rect 2473 873 2487 887
rect 2853 873 2867 887
rect 2893 873 2907 887
rect 3893 873 3907 887
rect 5633 873 5647 887
rect 5953 913 5967 927
rect 6193 913 6207 927
rect 2433 853 2447 867
rect 2493 853 2507 867
rect 4373 853 4387 867
rect 4453 853 4467 867
rect 6193 873 6207 887
rect 5973 853 5987 867
rect 6033 853 6047 867
rect 2233 832 2247 846
rect 2313 833 2327 847
rect 5973 832 5987 846
rect 1333 813 1347 827
rect 1393 813 1407 827
rect 1513 753 1527 767
rect 1573 753 1587 767
rect 5893 713 5907 727
rect 5913 714 5927 728
rect 753 693 767 707
rect 793 693 807 707
rect 953 693 967 707
rect 1833 693 1847 707
rect 1873 693 1887 707
rect 1993 693 2007 707
rect 2693 693 2707 707
rect 4633 693 4647 707
rect 5073 693 5087 707
rect 913 653 927 667
rect 2713 652 2727 666
rect 4633 653 4647 667
rect 5213 693 5227 707
rect 5253 693 5267 707
rect 5553 693 5567 707
rect 5673 693 5687 707
rect 5713 693 5727 707
rect 5133 653 5147 667
rect 5553 653 5567 667
rect 173 633 187 647
rect 253 633 267 647
rect 873 633 887 647
rect 933 633 947 647
rect 1273 633 1287 647
rect 1333 633 1347 647
rect 1693 633 1707 647
rect 1773 631 1787 645
rect 1813 631 1827 645
rect 1953 633 1967 647
rect 1993 633 2007 647
rect 2633 633 2647 647
rect 2753 633 2767 647
rect 3773 633 3787 647
rect 3873 633 3887 647
rect 4273 631 4287 645
rect 4353 633 4367 647
rect 5653 633 5667 647
rect 5713 633 5727 647
rect 1033 453 1047 467
rect 1073 453 1087 467
rect 113 413 127 427
rect 233 413 247 427
rect 1013 413 1027 427
rect 1073 413 1087 427
rect 1193 393 1207 407
rect 1893 413 1907 427
rect 1933 413 1947 427
rect 1993 413 2007 427
rect 2033 413 2047 427
rect 2173 413 2187 427
rect 2993 413 3007 427
rect 3113 414 3127 428
rect 4033 413 4047 427
rect 4073 413 4087 427
rect 5853 414 5867 428
rect 5893 413 5907 427
rect 6013 413 6027 427
rect 6073 413 6087 427
rect 1213 353 1227 367
rect 1773 353 1787 367
rect 2413 393 2427 407
rect 2893 393 2907 407
rect 3313 393 3327 407
rect 2853 373 2867 387
rect 2373 353 2387 367
rect 2833 353 2847 367
rect 3673 393 3687 407
rect 4473 393 4487 407
rect 4513 393 4527 407
rect 5753 393 5767 407
rect 2893 353 2907 367
rect 3313 353 3327 367
rect 3613 353 3627 367
rect 3733 353 3747 367
rect 3773 353 3787 367
rect 5773 352 5787 366
rect 5313 333 5327 347
rect 5393 333 5407 347
rect 3733 293 3747 307
rect 3773 293 3787 307
rect 3113 212 3127 226
rect 3173 213 3187 227
rect 253 193 267 207
rect 493 193 507 207
rect 573 193 587 207
rect 1053 193 1067 207
rect 1133 193 1147 207
rect 1733 193 1747 207
rect 4073 193 4087 207
rect 4113 193 4127 207
rect 4213 193 4227 207
rect 4333 193 4347 207
rect 1173 173 1187 187
rect 173 133 187 147
rect 1493 173 1507 187
rect 1533 173 1547 187
rect 1353 153 1367 167
rect 2053 173 2067 187
rect 2233 173 2247 187
rect 4053 173 4067 187
rect 4093 173 4107 187
rect 1233 133 1247 147
rect 1373 133 1387 147
rect 1793 133 1807 147
rect 2093 133 2107 147
rect 2193 133 2207 147
rect 193 112 207 126
rect 273 113 287 127
rect 413 113 427 127
rect 493 113 507 127
rect 973 113 987 127
rect 1053 113 1067 127
rect 1353 113 1367 127
rect 1413 113 1427 127
rect 1513 113 1527 127
rect 1593 113 1607 127
rect 1853 111 1867 125
rect 1933 113 1947 127
rect 1993 113 2007 127
rect 2153 113 2167 127
rect 2313 113 2327 127
rect 2373 113 2387 127
rect 2433 111 2447 125
rect 2913 113 2927 127
rect 3073 113 3087 127
rect 3313 113 3327 127
rect 3393 113 3407 127
rect 3933 113 3947 127
rect 3973 113 3987 127
rect 5253 113 5267 127
rect 5333 113 5347 127
rect 5453 113 5467 127
rect 5513 113 5527 127
rect 2473 93 2487 107
rect 2533 93 2547 107
rect 3293 93 3307 107
rect 3353 92 3367 106
rect 4393 93 4407 107
rect 4413 93 4427 107
rect 5393 93 5407 107
rect 5493 92 5507 106
rect 2333 53 2347 67
rect 2373 53 2387 67
rect 1473 33 1487 47
rect 1513 33 1527 47
<< metal2 >>
rect 1696 6267 1703 6303
rect 116 6116 123 6173
rect 196 6116 223 6123
rect 96 5947 103 6083
rect 196 6063 203 6116
rect 316 6076 343 6083
rect 196 6056 223 6063
rect 96 5896 103 5933
rect 216 5896 223 6056
rect 116 5847 123 5863
rect 116 5836 133 5847
rect 120 5833 133 5836
rect 156 5807 163 5853
rect 176 5847 183 5894
rect 276 5856 303 5863
rect 276 5608 283 5813
rect 296 5787 303 5856
rect 160 5603 173 5607
rect 156 5596 173 5603
rect 160 5593 173 5596
rect 96 5527 103 5563
rect 196 5547 203 5594
rect 227 5603 240 5607
rect 227 5596 243 5603
rect 227 5593 240 5596
rect 316 5607 323 5852
rect 213 5547 227 5553
rect 156 5447 163 5533
rect 116 5376 123 5433
rect 16 4767 23 5374
rect 196 5346 203 5512
rect 96 5340 103 5343
rect 136 5340 143 5343
rect 93 5327 107 5340
rect 133 5327 147 5340
rect 36 5007 43 5074
rect 16 4347 23 4653
rect 36 4507 43 4933
rect 56 4807 63 5032
rect 76 5027 83 5043
rect 76 5016 93 5027
rect 80 5013 93 5016
rect 116 4856 123 4993
rect 156 4868 163 5033
rect 176 5027 183 5313
rect 196 4823 203 5332
rect 216 5327 223 5512
rect 256 5507 263 5563
rect 296 5560 303 5563
rect 293 5547 307 5560
rect 316 5507 323 5553
rect 336 5523 343 6076
rect 356 6027 363 6114
rect 376 6047 383 6153
rect 513 6128 527 6133
rect 593 6120 607 6133
rect 596 6116 603 6120
rect 436 5947 443 6083
rect 476 6027 483 6083
rect 356 5807 363 5853
rect 436 5827 443 5933
rect 356 5687 363 5793
rect 456 5727 463 6013
rect 516 5896 523 6114
rect 656 6107 663 6153
rect 596 6027 603 6053
rect 616 5967 623 6083
rect 676 6007 683 6133
rect 716 6128 723 6173
rect 753 6120 767 6133
rect 756 6116 763 6120
rect 816 6107 823 6153
rect 880 6123 893 6127
rect 876 6116 893 6123
rect 880 6113 893 6116
rect 1236 6116 1243 6153
rect 736 6047 743 6083
rect 576 5867 583 5933
rect 636 5896 643 5993
rect 496 5827 503 5863
rect 496 5787 503 5813
rect 616 5727 623 5863
rect 656 5747 663 5863
rect 716 5863 723 5993
rect 856 5987 863 6083
rect 916 6067 923 6114
rect 933 6067 947 6072
rect 887 6033 893 6047
rect 920 6046 940 6047
rect 927 6033 933 6046
rect 1016 6027 1023 6083
rect 1056 6047 1063 6114
rect 1256 6080 1263 6083
rect 1253 6067 1267 6080
rect 1336 6007 1343 6113
rect 1356 6027 1363 6133
rect 1387 6114 1393 6127
rect 1433 6120 1447 6133
rect 1436 6116 1443 6120
rect 1387 6113 1400 6114
rect 1476 6087 1483 6193
rect 1580 6083 1593 6087
rect 1376 6007 1383 6072
rect 1536 6027 1543 6083
rect 1576 6076 1593 6083
rect 1580 6073 1593 6076
rect 1616 6067 1623 6114
rect 1636 6087 1643 6213
rect 1676 6116 1683 6153
rect 1716 6116 1723 6193
rect 1616 6027 1623 6053
rect 856 5907 863 5973
rect 896 5896 903 5973
rect 936 5896 943 5993
rect 1467 5956 1493 5963
rect 716 5856 763 5863
rect 396 5627 403 5713
rect 696 5687 703 5853
rect 356 5547 363 5613
rect 393 5600 407 5613
rect 396 5596 403 5600
rect 436 5596 443 5633
rect 496 5587 503 5673
rect 596 5608 603 5633
rect 696 5596 703 5673
rect 736 5608 743 5813
rect 796 5807 803 5863
rect 816 5783 823 5853
rect 836 5847 843 5893
rect 996 5866 1003 5953
rect 1047 5916 1073 5923
rect 1116 5866 1123 5933
rect 1316 5896 1323 5953
rect 1476 5896 1483 5933
rect 1256 5866 1263 5893
rect 916 5860 923 5863
rect 913 5847 927 5860
rect 796 5776 823 5783
rect 796 5607 803 5776
rect 1036 5747 1043 5813
rect 1056 5787 1063 5833
rect 1156 5827 1163 5863
rect 1336 5843 1343 5852
rect 1376 5847 1383 5893
rect 1536 5866 1543 5933
rect 1596 5896 1603 5993
rect 1696 5896 1703 6083
rect 1727 5956 1753 5963
rect 1736 5908 1743 5933
rect 1316 5836 1343 5843
rect 456 5527 463 5563
rect 336 5516 363 5523
rect 273 5388 287 5393
rect 316 5376 323 5413
rect 296 5340 303 5343
rect 293 5327 307 5340
rect 356 5327 363 5516
rect 516 5523 523 5594
rect 576 5560 583 5563
rect 573 5547 587 5560
rect 516 5516 533 5523
rect 476 5416 483 5453
rect 376 5346 383 5413
rect 236 5076 243 5273
rect 256 4967 263 5043
rect 216 4827 223 4854
rect 96 4787 103 4823
rect 136 4807 143 4823
rect 176 4816 203 4823
rect 56 4063 63 4713
rect 76 4568 83 4613
rect 96 4607 103 4773
rect 36 4056 63 4063
rect 16 3567 23 3853
rect 36 3786 43 4056
rect 76 4047 83 4493
rect 136 4427 143 4793
rect 156 4527 163 4593
rect 136 4227 143 4303
rect 136 4067 143 4173
rect 176 4087 183 4816
rect 236 4787 243 4893
rect 296 4887 303 5273
rect 316 5043 323 5313
rect 396 5287 403 5374
rect 336 5088 343 5133
rect 536 5127 543 5513
rect 556 5287 563 5473
rect 616 5403 623 5563
rect 656 5487 663 5594
rect 756 5467 763 5553
rect 776 5427 783 5594
rect 876 5527 883 5563
rect 976 5527 983 5563
rect 1036 5543 1043 5733
rect 1316 5647 1323 5836
rect 1416 5827 1423 5863
rect 1456 5860 1463 5863
rect 1453 5847 1467 5860
rect 1336 5687 1343 5813
rect 1476 5787 1483 5813
rect 1616 5767 1623 5863
rect 1716 5827 1723 5863
rect 1756 5767 1763 5863
rect 1796 5767 1803 6253
rect 1836 6116 1843 6213
rect 1916 6086 1923 6173
rect 1956 6123 1963 6303
rect 2116 6296 2143 6303
rect 2856 6296 2883 6303
rect 1956 6116 1973 6123
rect 2036 6116 2063 6123
rect 1996 6027 2003 6083
rect 1893 5900 1907 5913
rect 1896 5896 1903 5900
rect 1176 5596 1203 5603
rect 1016 5536 1043 5543
rect 1056 5563 1063 5593
rect 1196 5567 1203 5596
rect 1056 5556 1083 5563
rect 607 5396 623 5403
rect 593 5380 607 5393
rect 596 5376 603 5380
rect 636 5376 643 5413
rect 796 5376 803 5513
rect 616 5323 623 5343
rect 656 5340 663 5343
rect 653 5327 667 5340
rect 716 5327 723 5374
rect 856 5346 863 5413
rect 913 5380 927 5393
rect 916 5376 923 5380
rect 776 5340 783 5343
rect 773 5327 787 5340
rect 976 5343 983 5374
rect 1016 5347 1023 5536
rect 1056 5427 1063 5556
rect 1256 5543 1263 5563
rect 1256 5536 1283 5543
rect 1116 5376 1123 5413
rect 616 5316 643 5323
rect 316 5036 343 5043
rect 296 4856 323 4863
rect 316 4667 323 4856
rect 336 4703 343 5036
rect 356 5023 363 5043
rect 356 5016 383 5023
rect 356 4727 363 4993
rect 376 4987 383 5016
rect 376 4863 383 4973
rect 456 4903 463 5074
rect 496 4967 503 5043
rect 536 5027 543 5043
rect 527 5016 543 5027
rect 527 5013 540 5016
rect 447 4896 463 4903
rect 376 4856 393 4863
rect 436 4856 443 4893
rect 556 4856 563 5013
rect 576 4987 583 5033
rect 596 5027 603 5113
rect 616 4967 623 5273
rect 636 5267 643 5316
rect 736 5267 743 5313
rect 636 5087 643 5153
rect 696 5076 703 5113
rect 736 5087 743 5253
rect 676 5023 683 5043
rect 667 5016 683 5023
rect 416 4767 423 4823
rect 476 4787 483 4854
rect 336 4696 363 4703
rect 216 4556 223 4593
rect 196 4267 203 4513
rect 236 4363 243 4512
rect 296 4423 303 4593
rect 356 4556 363 4696
rect 376 4487 383 4523
rect 296 4416 323 4423
rect 276 4363 283 4393
rect 216 4356 243 4363
rect 256 4356 283 4363
rect 216 4127 223 4356
rect 256 4336 263 4356
rect 56 3828 63 4034
rect 133 4040 147 4053
rect 156 4047 163 4073
rect 136 4036 143 4040
rect 76 3947 83 3993
rect 16 3347 23 3553
rect 16 3266 23 3333
rect 36 3107 43 3633
rect 56 3527 63 3814
rect 156 3787 163 3933
rect 176 3867 183 4052
rect 216 4036 223 4073
rect 236 4067 243 4303
rect 296 4300 303 4303
rect 293 4287 307 4300
rect 316 4187 323 4416
rect 336 4207 343 4413
rect 396 4336 403 4453
rect 416 4387 423 4753
rect 436 4527 443 4773
rect 576 4767 583 4823
rect 476 4607 483 4733
rect 496 4583 503 4673
rect 476 4576 503 4583
rect 476 4556 483 4576
rect 516 4556 523 4753
rect 656 4727 663 5013
rect 756 5003 763 5313
rect 773 5307 787 5313
rect 896 5307 903 5343
rect 956 5336 983 5343
rect 1176 5346 1183 5433
rect 1056 5340 1063 5343
rect 1053 5327 1067 5340
rect 776 5087 783 5113
rect 793 5088 807 5093
rect 836 5076 843 5153
rect 896 5147 903 5173
rect 773 5027 787 5033
rect 756 4996 783 5003
rect 736 4883 743 4933
rect 736 4876 763 4883
rect 756 4868 763 4876
rect 776 4867 783 4996
rect 796 4907 803 4953
rect 876 4947 883 5033
rect 896 4907 903 5133
rect 916 5087 923 5193
rect 956 5076 963 5113
rect 836 4868 843 4893
rect 936 4868 943 5032
rect 1036 5027 1043 5113
rect 1056 5043 1063 5273
rect 1196 5103 1203 5393
rect 1233 5380 1247 5393
rect 1276 5388 1283 5536
rect 1336 5527 1343 5673
rect 1876 5647 1883 5863
rect 1936 5827 1943 5913
rect 1976 5896 1983 5953
rect 2016 5896 2023 5953
rect 2056 5947 2063 6116
rect 2116 6116 2123 6296
rect 2076 5967 2083 6114
rect 2316 6100 2323 6103
rect 2313 6087 2327 6100
rect 2356 6103 2363 6193
rect 2356 6096 2383 6103
rect 2656 6103 2663 6253
rect 2656 6096 2683 6103
rect 2076 5867 2083 5894
rect 2136 5647 2143 5863
rect 1436 5596 1443 5633
rect 1816 5608 1823 5633
rect 1636 5566 1643 5593
rect 1536 5388 1543 5563
rect 1647 5556 1663 5563
rect 1787 5513 1793 5527
rect 1816 5447 1823 5594
rect 1976 5596 1983 5633
rect 2036 5596 2063 5603
rect 1856 5527 1863 5563
rect 1896 5560 1903 5563
rect 1893 5547 1907 5560
rect 1956 5527 1963 5593
rect 1236 5376 1243 5380
rect 1576 5376 1583 5433
rect 1816 5376 1823 5433
rect 1976 5376 1983 5533
rect 2056 5527 2063 5596
rect 2196 5607 2203 5953
rect 2256 5896 2263 5933
rect 2236 5787 2243 5852
rect 2336 5827 2343 6093
rect 2456 5896 2463 5993
rect 2476 5860 2483 5863
rect 2256 5767 2263 5813
rect 2216 5707 2223 5753
rect 2156 5487 2163 5563
rect 1336 5347 1343 5374
rect 1256 5287 1263 5343
rect 1296 5147 1303 5332
rect 1396 5287 1403 5343
rect 1196 5096 1223 5103
rect 1056 5036 1103 5043
rect 1136 5040 1143 5043
rect 1133 5027 1147 5040
rect 1036 4856 1063 4863
rect 536 4587 543 4613
rect 576 4563 583 4713
rect 616 4587 623 4633
rect 576 4556 603 4563
rect 633 4560 647 4573
rect 636 4556 643 4560
rect 676 4556 683 4813
rect 696 4787 703 4823
rect 720 4805 740 4807
rect 720 4802 733 4805
rect 716 4793 733 4802
rect 696 4567 703 4673
rect 496 4427 503 4523
rect 536 4427 543 4523
rect 507 4416 523 4423
rect 376 4187 383 4303
rect 416 4300 423 4303
rect 413 4287 427 4300
rect 456 4267 463 4373
rect 516 4336 523 4416
rect 556 4336 563 4433
rect 576 4387 583 4513
rect 596 4447 603 4556
rect 716 4523 723 4793
rect 696 4516 723 4523
rect 596 4347 603 4393
rect 396 4087 403 4213
rect 436 4127 443 4253
rect 476 4247 483 4273
rect 536 4227 543 4303
rect 576 4283 583 4303
rect 556 4276 583 4283
rect 496 4147 503 4193
rect 236 4058 253 4067
rect 240 4054 253 4058
rect 240 4053 260 4054
rect 276 3996 303 4003
rect 276 3787 283 3953
rect 296 3947 303 3996
rect 316 3967 323 4013
rect 336 3847 343 4053
rect 416 4063 423 4113
rect 416 4056 443 4063
rect 393 4040 407 4052
rect 436 4047 443 4056
rect 396 4036 403 4040
rect 436 4036 453 4047
rect 440 4033 453 4036
rect 376 3927 383 4003
rect 416 3947 423 4003
rect 236 3780 243 3783
rect 133 3520 147 3533
rect 136 3516 143 3520
rect 56 3127 63 3373
rect 116 3323 123 3483
rect 156 3447 163 3483
rect 196 3387 203 3772
rect 233 3767 247 3780
rect 266 3773 267 3780
rect 253 3767 267 3773
rect 296 3767 303 3833
rect 353 3820 367 3833
rect 356 3816 363 3820
rect 396 3816 403 3853
rect 436 3827 443 3893
rect 456 3847 463 3993
rect 476 3828 483 4073
rect 496 3843 503 4133
rect 536 4048 543 4173
rect 556 4067 563 4276
rect 596 4067 603 4293
rect 616 4187 623 4473
rect 636 4306 643 4453
rect 696 4336 703 4516
rect 736 4427 743 4693
rect 756 4627 763 4733
rect 776 4556 783 4773
rect 796 4687 803 4853
rect 816 4807 823 4853
rect 836 4707 843 4854
rect 936 4807 943 4854
rect 996 4820 1003 4823
rect 896 4727 903 4773
rect 796 4587 803 4673
rect 956 4647 963 4812
rect 993 4807 1007 4820
rect 813 4560 827 4573
rect 856 4567 863 4593
rect 816 4556 823 4560
rect 796 4387 803 4523
rect 756 4343 763 4373
rect 736 4336 763 4343
rect 776 4306 783 4353
rect 816 4343 823 4373
rect 836 4367 843 4512
rect 876 4487 883 4633
rect 893 4567 907 4573
rect 796 4336 823 4343
rect 853 4340 867 4353
rect 896 4347 903 4553
rect 856 4336 863 4340
rect 716 4227 723 4303
rect 796 4223 803 4336
rect 916 4327 923 4633
rect 976 4587 983 4673
rect 1056 4667 1063 4856
rect 1076 4807 1083 4953
rect 1096 4767 1103 5013
rect 1176 4923 1183 5033
rect 1196 4967 1203 5074
rect 1216 5046 1223 5096
rect 1273 5088 1287 5093
rect 1296 4987 1303 5043
rect 1176 4916 1203 4923
rect 1156 4856 1163 4893
rect 1196 4868 1203 4916
rect 1136 4820 1143 4823
rect 1133 4807 1147 4820
rect 996 4556 1003 4633
rect 956 4447 963 4523
rect 996 4367 1003 4393
rect 787 4216 803 4223
rect 636 4036 643 4073
rect 716 4047 723 4113
rect 776 4067 783 4213
rect 816 4127 823 4153
rect 556 4000 563 4003
rect 516 3927 523 3993
rect 553 3987 567 4000
rect 576 3963 583 3993
rect 556 3956 583 3963
rect 556 3867 563 3956
rect 596 3907 603 4032
rect 616 3907 623 3973
rect 656 3887 663 4003
rect 496 3836 513 3843
rect 456 3816 473 3823
rect 336 3780 343 3783
rect 333 3767 347 3780
rect 416 3727 423 3772
rect 436 3647 443 3773
rect 216 3447 223 3513
rect 276 3480 283 3483
rect 273 3467 287 3480
rect 96 3316 123 3323
rect 96 3296 103 3316
rect 136 3296 143 3333
rect 216 3328 223 3433
rect 316 3427 323 3613
rect 256 3296 263 3353
rect 116 3207 123 3263
rect 16 2967 23 3033
rect 16 2787 23 2913
rect 36 2607 43 3053
rect 93 3000 107 3013
rect 136 3008 143 3093
rect 176 3027 183 3293
rect 280 3263 293 3267
rect 236 3260 243 3263
rect 233 3247 247 3260
rect 276 3256 293 3263
rect 280 3253 293 3256
rect 316 3247 323 3313
rect 276 3027 283 3053
rect 96 2996 103 3000
rect 176 2967 183 3013
rect 273 3000 287 3013
rect 276 2996 283 3000
rect 196 2967 203 2994
rect 316 2967 323 3212
rect 336 3027 343 3593
rect 456 3587 463 3816
rect 513 3820 527 3833
rect 553 3827 567 3832
rect 516 3816 523 3820
rect 576 3786 583 3873
rect 496 3780 503 3783
rect 493 3767 507 3780
rect 536 3707 543 3783
rect 396 3476 423 3483
rect 356 3307 363 3473
rect 393 3447 407 3453
rect 416 3447 423 3476
rect 436 3307 443 3533
rect 456 3467 463 3573
rect 496 3547 503 3633
rect 536 3547 543 3573
rect 496 3516 503 3533
rect 536 3516 543 3533
rect 576 3523 583 3772
rect 596 3727 603 3853
rect 676 3816 683 3973
rect 696 3967 703 4003
rect 716 3867 723 3913
rect 616 3567 623 3773
rect 736 3783 743 3993
rect 756 3827 763 3973
rect 776 3967 783 4003
rect 836 3967 843 4173
rect 856 3987 863 4253
rect 936 4227 943 4353
rect 1016 4336 1023 4653
rect 956 4306 963 4333
rect 916 4063 923 4153
rect 976 4087 983 4303
rect 916 4056 943 4063
rect 936 4036 943 4056
rect 776 3816 783 3873
rect 856 3820 903 3823
rect 853 3816 903 3820
rect 696 3776 743 3783
rect 696 3647 703 3776
rect 800 3783 813 3787
rect 796 3776 813 3783
rect 800 3773 813 3776
rect 576 3516 603 3523
rect 516 3447 523 3483
rect 416 3256 443 3263
rect 376 3067 383 3252
rect 413 3227 427 3233
rect 436 3147 443 3256
rect 456 3207 463 3373
rect 536 3296 543 3353
rect 556 3327 563 3472
rect 596 3303 603 3516
rect 676 3516 683 3613
rect 716 3587 723 3673
rect 716 3527 723 3552
rect 656 3480 663 3483
rect 696 3480 703 3483
rect 653 3467 667 3480
rect 693 3467 707 3480
rect 676 3387 683 3413
rect 636 3307 643 3353
rect 596 3296 623 3303
rect 476 3187 483 3293
rect 507 3263 520 3267
rect 507 3253 523 3263
rect 556 3260 563 3263
rect 456 3023 463 3153
rect 496 3047 503 3193
rect 516 3087 523 3253
rect 553 3247 567 3260
rect 436 3016 463 3023
rect 340 3006 360 3007
rect 347 3003 360 3006
rect 347 2996 363 3003
rect 347 2993 360 2996
rect 76 2743 83 2952
rect 176 2776 183 2913
rect 216 2788 223 2953
rect 256 2887 263 2963
rect 336 2907 343 2953
rect 276 2776 283 2813
rect 76 2736 103 2743
rect 216 2727 223 2774
rect 396 2776 403 2893
rect 436 2787 443 3016
rect 516 2996 523 3052
rect 553 3000 567 3013
rect 576 3007 583 3233
rect 616 3167 623 3296
rect 676 3296 683 3373
rect 736 3367 743 3753
rect 756 3607 763 3773
rect 836 3767 843 3814
rect 853 3807 867 3816
rect 956 3827 963 3992
rect 996 3943 1003 4253
rect 1036 4247 1043 4573
rect 1056 4567 1063 4613
rect 1056 4167 1063 4513
rect 1076 4487 1083 4523
rect 1096 4347 1103 4433
rect 1116 4387 1123 4513
rect 1136 4507 1143 4554
rect 1156 4403 1163 4753
rect 1176 4687 1183 4812
rect 1196 4667 1203 4713
rect 1216 4627 1223 4733
rect 1236 4707 1243 4973
rect 1276 4856 1283 4953
rect 1356 4867 1363 5133
rect 1433 5080 1447 5093
rect 1436 5076 1443 5080
rect 1376 5047 1383 5074
rect 1296 4820 1303 4823
rect 1293 4807 1307 4820
rect 1336 4787 1343 4823
rect 1256 4667 1263 4753
rect 1336 4727 1343 4773
rect 1313 4647 1327 4653
rect 1260 4646 1280 4647
rect 1267 4633 1273 4646
rect 1196 4556 1203 4593
rect 1216 4583 1223 4613
rect 1216 4576 1243 4583
rect 1236 4556 1243 4576
rect 1147 4396 1163 4403
rect 1136 4336 1143 4393
rect 1176 4336 1183 4453
rect 1196 4427 1203 4493
rect 1216 4387 1223 4523
rect 1236 4347 1243 4493
rect 1016 4047 1023 4073
rect 1056 4063 1063 4153
rect 1036 4056 1063 4063
rect 1036 4036 1043 4056
rect 1076 4048 1083 4333
rect 1096 4247 1103 4293
rect 1116 4227 1123 4303
rect 1233 4303 1247 4312
rect 1196 4300 1247 4303
rect 1196 4296 1243 4300
rect 1256 4287 1263 4373
rect 1276 4347 1283 4593
rect 1296 4523 1303 4573
rect 1316 4567 1323 4612
rect 1356 4587 1363 4813
rect 1376 4807 1383 4893
rect 1396 4823 1403 4933
rect 1416 4887 1423 5032
rect 1456 5007 1463 5043
rect 1516 4987 1523 5074
rect 1536 4947 1543 5293
rect 1556 5167 1563 5343
rect 1636 5127 1643 5374
rect 1636 5007 1643 5043
rect 1636 4967 1643 4993
rect 1456 4896 1493 4903
rect 1456 4883 1463 4896
rect 1436 4876 1463 4883
rect 1436 4856 1443 4876
rect 1473 4860 1487 4873
rect 1476 4856 1483 4860
rect 1596 4856 1603 4893
rect 1396 4816 1423 4823
rect 1416 4803 1423 4816
rect 1416 4796 1443 4803
rect 1436 4567 1443 4796
rect 1456 4607 1463 4823
rect 1496 4803 1503 4823
rect 1476 4796 1503 4803
rect 1296 4516 1323 4523
rect 1316 4336 1323 4516
rect 1356 4447 1363 4523
rect 1396 4467 1403 4523
rect 1296 4300 1303 4303
rect 1293 4287 1307 4300
rect 1133 4047 1147 4053
rect 1116 4007 1123 4034
rect 1193 4040 1207 4053
rect 1236 4047 1243 4133
rect 1196 4036 1203 4040
rect 1096 3967 1103 3993
rect 976 3936 1003 3943
rect 976 3787 983 3936
rect 1027 3923 1040 3927
rect 1027 3920 1043 3923
rect 1027 3913 1047 3920
rect 1033 3907 1047 3913
rect 776 3567 783 3713
rect 856 3687 863 3772
rect 916 3763 923 3783
rect 996 3786 1003 3853
rect 1016 3847 1023 3873
rect 1056 3816 1063 3953
rect 916 3756 943 3763
rect 893 3747 907 3753
rect 893 3740 913 3747
rect 896 3736 913 3740
rect 900 3733 913 3736
rect 936 3727 943 3756
rect 847 3676 863 3687
rect 847 3673 860 3676
rect 796 3516 803 3633
rect 836 3486 843 3593
rect 876 3527 883 3673
rect 916 3607 923 3693
rect 756 3303 763 3473
rect 776 3427 783 3483
rect 856 3467 863 3514
rect 976 3527 983 3553
rect 856 3367 863 3453
rect 876 3447 883 3473
rect 756 3296 783 3303
rect 556 2996 563 3000
rect 456 2967 463 2994
rect 576 2887 583 2953
rect 596 2867 603 3013
rect 636 2996 643 3073
rect 696 3067 703 3263
rect 736 3256 763 3263
rect 756 3227 763 3256
rect 716 3087 723 3113
rect 673 3000 687 3013
rect 676 2996 683 3000
rect 696 2960 703 2963
rect 693 2947 707 2960
rect 636 2788 643 2873
rect 256 2740 263 2743
rect 253 2727 267 2740
rect 36 1607 43 2513
rect 76 2476 103 2483
rect 156 2476 183 2483
rect 76 2407 83 2476
rect 76 2223 83 2393
rect 136 2268 143 2313
rect 176 2283 183 2476
rect 196 2467 203 2573
rect 316 2527 323 2773
rect 576 2743 583 2773
rect 696 2746 703 2893
rect 736 2847 743 3133
rect 756 2987 763 3213
rect 776 3107 783 3296
rect 796 3247 803 3353
rect 916 3327 923 3433
rect 936 3427 943 3483
rect 893 3300 907 3313
rect 896 3296 903 3300
rect 876 3247 883 3263
rect 796 3207 803 3233
rect 827 3213 833 3227
rect 876 3187 883 3233
rect 916 3227 923 3253
rect 793 3008 807 3013
rect 876 2996 883 3093
rect 916 3067 923 3153
rect 816 2887 823 2963
rect 856 2867 863 2952
rect 896 2903 903 2953
rect 876 2896 903 2903
rect 496 2707 503 2743
rect 536 2736 583 2743
rect 316 2483 323 2513
rect 356 2488 363 2613
rect 296 2476 323 2483
rect 416 2476 423 2573
rect 276 2367 283 2443
rect 276 2307 283 2353
rect 176 2276 203 2283
rect 76 2216 103 2223
rect 156 2220 163 2223
rect 96 2007 103 2216
rect 153 2207 167 2220
rect 96 1887 103 1923
rect 136 1920 143 1923
rect 133 1907 147 1920
rect 156 1867 163 1913
rect 176 1907 183 2254
rect 196 2226 203 2276
rect 316 2256 323 2293
rect 196 1887 203 1993
rect 256 1987 263 2191
rect 296 2127 303 2212
rect 356 2047 363 2474
rect 396 2407 403 2443
rect 436 2440 443 2443
rect 433 2427 447 2440
rect 376 2267 383 2293
rect 456 1987 463 2293
rect 476 2227 483 2433
rect 496 2267 503 2693
rect 656 2627 663 2743
rect 716 2667 723 2774
rect 756 2643 763 2743
rect 716 2636 763 2643
rect 516 2476 543 2483
rect 516 2427 523 2476
rect 516 2287 523 2413
rect 556 2367 563 2443
rect 536 2256 543 2313
rect 596 2226 603 2273
rect 656 2256 663 2513
rect 716 2488 723 2636
rect 756 2476 763 2613
rect 776 2487 783 2653
rect 796 2627 803 2743
rect 876 2723 883 2896
rect 916 2843 923 2994
rect 936 2947 943 3392
rect 976 3387 983 3472
rect 996 3427 1003 3593
rect 1016 3407 1023 3773
rect 1076 3727 1083 3783
rect 1036 3527 1043 3553
rect 1076 3516 1083 3573
rect 1116 3527 1123 3773
rect 1136 3687 1143 3993
rect 1216 3967 1223 4003
rect 956 3007 963 3313
rect 976 3307 983 3373
rect 1036 3307 1043 3473
rect 1060 3465 1080 3467
rect 1067 3462 1080 3465
rect 1067 3460 1083 3462
rect 1067 3453 1087 3460
rect 1073 3447 1087 3453
rect 1016 3260 1023 3263
rect 1013 3247 1027 3260
rect 976 3187 983 3233
rect 1016 3027 1023 3233
rect 1036 3107 1043 3253
rect 1036 3003 1043 3093
rect 1016 2996 1043 3003
rect 1056 2987 1063 3413
rect 1096 3367 1103 3483
rect 1116 3323 1123 3473
rect 1136 3367 1143 3533
rect 1156 3527 1163 3853
rect 1216 3847 1223 3913
rect 1236 3843 1243 3993
rect 1256 3863 1263 4153
rect 1336 4036 1343 4173
rect 1376 4087 1383 4173
rect 1396 4167 1403 4453
rect 1416 4147 1423 4493
rect 1456 4487 1463 4554
rect 1476 4527 1483 4796
rect 1516 4767 1523 4812
rect 1536 4767 1543 4854
rect 1576 4803 1583 4812
rect 1616 4803 1623 4823
rect 1576 4796 1603 4803
rect 1616 4796 1643 4803
rect 1536 4627 1543 4753
rect 1556 4556 1563 4733
rect 1576 4707 1583 4773
rect 1596 4467 1603 4796
rect 1616 4568 1623 4613
rect 1636 4607 1643 4796
rect 1676 4747 1683 5253
rect 1696 5207 1703 5233
rect 1756 5187 1763 5273
rect 1836 5207 1843 5343
rect 1956 5207 1963 5343
rect 1696 4823 1703 5074
rect 1716 5047 1723 5113
rect 1856 5047 1863 5153
rect 1876 5007 1883 5193
rect 1936 5076 1943 5113
rect 1996 5087 2003 5343
rect 2076 5243 2083 5343
rect 2156 5307 2163 5413
rect 2216 5388 2223 5693
rect 2236 5467 2243 5633
rect 2236 5407 2243 5432
rect 2256 5387 2263 5533
rect 2276 5527 2283 5563
rect 2326 5552 2327 5560
rect 2313 5547 2327 5552
rect 2176 5347 2183 5374
rect 2276 5346 2283 5473
rect 2336 5376 2343 5553
rect 2356 5487 2363 5852
rect 2473 5847 2487 5860
rect 2456 5596 2463 5713
rect 2496 5607 2503 5773
rect 2376 5567 2383 5594
rect 2376 5507 2383 5532
rect 2056 5236 2083 5243
rect 1773 4900 1787 4913
rect 1776 4896 1783 4900
rect 1836 4863 1843 4953
rect 1896 4907 1903 4953
rect 1956 4927 1963 5043
rect 1816 4856 1843 4863
rect 1696 4816 1723 4823
rect 1696 4763 1703 4816
rect 1696 4756 1723 4763
rect 1636 4556 1643 4593
rect 1716 4523 1723 4756
rect 1473 4340 1487 4353
rect 1476 4336 1483 4340
rect 1536 4306 1543 4453
rect 1636 4348 1643 4493
rect 1656 4487 1663 4523
rect 1696 4516 1723 4523
rect 1456 4300 1463 4303
rect 1436 4263 1443 4293
rect 1453 4287 1467 4300
rect 1496 4267 1503 4303
rect 1616 4267 1623 4303
rect 1436 4256 1463 4263
rect 1436 4123 1443 4233
rect 1456 4207 1463 4256
rect 1476 4187 1483 4253
rect 1416 4116 1443 4123
rect 1373 4048 1387 4052
rect 1396 4047 1403 4113
rect 1276 4007 1283 4034
rect 1316 4000 1323 4003
rect 1313 3987 1327 4000
rect 1416 4003 1423 4116
rect 1467 4073 1473 4087
rect 1516 4036 1523 4073
rect 1556 4047 1563 4133
rect 1436 4007 1443 4034
rect 1396 3996 1423 4003
rect 1256 3860 1283 3863
rect 1256 3856 1287 3860
rect 1273 3847 1287 3856
rect 1236 3836 1263 3843
rect 1216 3816 1223 3833
rect 1256 3816 1263 3836
rect 1296 3827 1303 3953
rect 1316 3847 1323 3973
rect 1396 3967 1403 3996
rect 1456 3967 1463 3993
rect 1316 3786 1323 3812
rect 1336 3787 1343 3953
rect 1416 3887 1423 3913
rect 1416 3816 1423 3873
rect 1496 3827 1503 4003
rect 1576 4006 1583 4053
rect 1613 4040 1627 4053
rect 1616 4036 1623 4040
rect 1656 4036 1663 4293
rect 1676 4067 1683 4493
rect 1696 4307 1703 4516
rect 1736 4507 1743 4733
rect 1756 4567 1763 4653
rect 1776 4556 1783 4593
rect 1836 4588 1843 4833
rect 1856 4703 1863 4873
rect 1876 4867 1883 4893
rect 1893 4860 1907 4872
rect 1933 4860 1947 4873
rect 1956 4867 1963 4913
rect 1896 4856 1903 4860
rect 1936 4856 1943 4860
rect 1856 4696 1883 4703
rect 1716 4427 1723 4473
rect 1736 4336 1743 4393
rect 1756 4387 1763 4553
rect 1856 4527 1863 4673
rect 1876 4567 1883 4696
rect 1796 4447 1803 4512
rect 1876 4507 1883 4532
rect 1840 4506 1860 4507
rect 1840 4503 1853 4506
rect 1836 4493 1853 4503
rect 1796 4303 1803 4373
rect 1716 4267 1723 4303
rect 1776 4296 1803 4303
rect 1736 4048 1743 4073
rect 1516 3787 1523 3873
rect 1556 3867 1563 3993
rect 1636 3967 1643 4003
rect 1676 4000 1683 4003
rect 1673 3987 1687 4000
rect 1576 3867 1583 3893
rect 1593 3860 1607 3873
rect 1596 3856 1603 3860
rect 1636 3816 1663 3823
rect 1196 3727 1203 3783
rect 1236 3762 1243 3783
rect 1236 3755 1273 3762
rect 1196 3627 1203 3713
rect 1193 3520 1207 3533
rect 1196 3516 1203 3520
rect 1236 3516 1243 3593
rect 1256 3527 1263 3713
rect 1276 3487 1283 3713
rect 1296 3707 1303 3753
rect 1356 3627 1363 3773
rect 1396 3763 1403 3772
rect 1436 3763 1443 3783
rect 1376 3756 1403 3763
rect 1416 3756 1443 3763
rect 1316 3516 1323 3593
rect 1356 3516 1363 3573
rect 1376 3567 1383 3756
rect 1416 3687 1423 3756
rect 1447 3733 1453 3747
rect 1476 3727 1483 3772
rect 1493 3727 1507 3733
rect 1506 3720 1507 3727
rect 1527 3713 1533 3727
rect 1396 3527 1403 3633
rect 1496 3547 1503 3692
rect 1176 3387 1183 3483
rect 1107 3316 1123 3323
rect 1096 3296 1103 3313
rect 1173 3307 1187 3313
rect 1196 3267 1203 3453
rect 1236 3403 1243 3433
rect 1256 3427 1263 3473
rect 1336 3447 1343 3483
rect 1416 3447 1423 3533
rect 1453 3520 1467 3533
rect 1500 3523 1513 3527
rect 1456 3516 1463 3520
rect 1496 3516 1513 3523
rect 1500 3513 1513 3516
rect 1236 3396 1273 3403
rect 1427 3403 1440 3407
rect 1427 3393 1443 3403
rect 1216 3327 1223 3353
rect 896 2836 923 2843
rect 896 2827 903 2836
rect 896 2743 903 2813
rect 953 2780 967 2793
rect 956 2776 963 2780
rect 896 2736 923 2743
rect 976 2727 983 2933
rect 1076 2887 1083 3253
rect 1116 3047 1123 3263
rect 1156 3187 1163 3263
rect 1216 3266 1223 3313
rect 1276 3296 1283 3333
rect 1296 3260 1303 3263
rect 1293 3247 1307 3260
rect 1176 3167 1183 3213
rect 1176 2966 1183 2993
rect 1176 2907 1183 2952
rect 1196 2927 1203 3113
rect 1256 2996 1263 3153
rect 1356 3127 1363 3333
rect 1416 3296 1423 3353
rect 1436 3347 1443 3393
rect 1516 3267 1523 3473
rect 1536 3327 1543 3533
rect 1556 3487 1563 3673
rect 1656 3647 1663 3816
rect 1676 3787 1683 3933
rect 1576 3527 1583 3613
rect 1660 3523 1673 3527
rect 1656 3516 1673 3523
rect 1660 3513 1673 3516
rect 1436 3207 1443 3263
rect 1556 3187 1563 3433
rect 1636 3367 1643 3483
rect 1676 3427 1683 3473
rect 1676 3287 1683 3353
rect 1656 3256 1683 3263
rect 1316 3047 1323 3113
rect 1376 3067 1383 3133
rect 1516 3107 1523 3133
rect 1316 2966 1323 3033
rect 1396 2996 1403 3053
rect 1496 3008 1503 3093
rect 1527 3033 1533 3047
rect 1596 3007 1603 3113
rect 1616 3107 1623 3133
rect 1476 2967 1483 2994
rect 1416 2927 1423 2963
rect 1593 2947 1607 2952
rect 1016 2816 1053 2823
rect 1016 2787 1023 2816
rect 1033 2780 1047 2793
rect 1036 2776 1043 2780
rect 876 2716 903 2723
rect 856 2476 863 2673
rect 696 2407 703 2443
rect 896 2443 903 2716
rect 973 2480 987 2493
rect 976 2476 983 2480
rect 876 2436 903 2443
rect 516 2027 523 2212
rect 556 2067 563 2223
rect 636 2187 643 2223
rect 696 2007 703 2313
rect 776 2256 783 2432
rect 836 2407 843 2432
rect 796 2187 803 2223
rect 856 2207 863 2254
rect 876 2223 883 2436
rect 1016 2407 1023 2493
rect 1036 2447 1043 2713
rect 1076 2707 1083 2743
rect 1096 2667 1103 2793
rect 1176 2776 1183 2813
rect 1216 2776 1223 2873
rect 1196 2687 1203 2743
rect 1236 2740 1243 2743
rect 1233 2727 1247 2740
rect 1116 2476 1163 2483
rect 936 2256 943 2393
rect 996 2226 1003 2313
rect 1156 2287 1163 2476
rect 1196 2327 1203 2673
rect 1256 2587 1263 2733
rect 1256 2327 1263 2443
rect 1296 2347 1303 2873
rect 1373 2780 1387 2793
rect 1416 2788 1423 2833
rect 1376 2776 1383 2780
rect 1416 2747 1423 2774
rect 1356 2627 1363 2743
rect 1396 2707 1403 2733
rect 1376 2607 1383 2653
rect 1336 2547 1343 2593
rect 1196 2276 1273 2283
rect 1113 2260 1127 2273
rect 1196 2268 1203 2276
rect 1116 2256 1123 2260
rect 876 2216 903 2223
rect 696 1983 703 1993
rect 256 1956 263 1973
rect 156 1767 163 1853
rect 196 1767 203 1852
rect 160 1743 173 1747
rect 156 1736 173 1743
rect 56 1667 63 1734
rect 160 1733 173 1736
rect 216 1743 223 1913
rect 236 1867 243 1923
rect 276 1867 283 1923
rect 336 1867 343 1954
rect 476 1923 483 1954
rect 496 1926 503 1973
rect 573 1960 587 1973
rect 676 1976 703 1983
rect 576 1956 583 1960
rect 676 1956 683 1976
rect 633 1947 647 1954
rect 207 1736 223 1743
rect 76 1696 103 1703
rect 76 1647 83 1696
rect 76 1436 83 1633
rect 176 1443 183 1693
rect 196 1627 203 1732
rect 336 1706 343 1773
rect 376 1767 383 1893
rect 436 1827 443 1923
rect 456 1916 483 1923
rect 456 1736 463 1916
rect 156 1436 183 1443
rect 196 1436 203 1533
rect 236 1448 243 1573
rect 156 1247 163 1436
rect 276 1407 283 1613
rect 336 1436 343 1493
rect 356 1487 363 1733
rect 496 1707 503 1773
rect 396 1700 403 1703
rect 376 1647 383 1693
rect 393 1687 407 1700
rect 393 1667 407 1673
rect 433 1667 447 1671
rect 356 1383 363 1403
rect 336 1376 363 1383
rect 160 1223 173 1227
rect 156 1216 173 1223
rect 36 667 43 1214
rect 160 1213 173 1216
rect 96 1127 103 1183
rect 136 1087 143 1183
rect 196 1167 203 1233
rect 56 827 63 914
rect 160 883 173 887
rect 156 876 173 883
rect 160 873 173 876
rect 116 723 123 872
rect 196 827 203 933
rect 216 928 223 1233
rect 273 1220 287 1233
rect 276 1216 283 1220
rect 336 1227 343 1376
rect 416 1247 423 1473
rect 436 1447 443 1613
rect 476 1436 483 1593
rect 516 1507 523 1893
rect 556 1867 563 1923
rect 596 1867 603 1923
rect 616 1787 623 1913
rect 573 1740 587 1753
rect 576 1736 583 1740
rect 596 1487 603 1573
rect 616 1463 623 1773
rect 636 1547 643 1912
rect 656 1847 663 1893
rect 696 1887 703 1923
rect 756 1887 763 1993
rect 776 1967 783 2013
rect 836 1956 843 2113
rect 896 2067 903 2216
rect 916 2167 923 2223
rect 956 2187 963 2223
rect 1016 2223 1023 2254
rect 1016 2216 1043 2223
rect 976 2127 983 2193
rect 876 1956 883 2013
rect 896 1967 903 2053
rect 916 1927 923 2093
rect 976 1956 983 2113
rect 996 1967 1003 2033
rect 696 1767 703 1873
rect 756 1847 763 1873
rect 656 1706 663 1753
rect 716 1736 723 1793
rect 776 1748 783 1913
rect 856 1887 863 1923
rect 736 1587 743 1703
rect 796 1667 803 1793
rect 896 1747 903 1913
rect 1016 1907 1023 2173
rect 1036 2167 1043 2216
rect 1096 2187 1103 2223
rect 1156 2203 1163 2252
rect 1296 2226 1303 2273
rect 1136 2196 1163 2203
rect 1036 1927 1043 2153
rect 596 1456 623 1463
rect 596 1436 603 1456
rect 556 1407 563 1434
rect 416 1216 423 1233
rect 456 1216 463 1253
rect 356 1187 363 1214
rect 256 1047 263 1172
rect 276 1067 283 1153
rect 236 927 243 973
rect 293 920 307 933
rect 336 927 343 1173
rect 296 916 303 920
rect 356 887 363 1113
rect 316 876 343 883
rect 253 723 267 733
rect 96 716 123 723
rect 236 720 267 723
rect 236 716 263 720
rect 96 696 103 716
rect 236 696 243 716
rect 76 403 83 652
rect 116 567 123 663
rect 176 647 183 693
rect 316 666 323 853
rect 336 767 343 876
rect 376 727 383 1073
rect 396 1067 403 1183
rect 396 927 403 1053
rect 436 1047 443 1183
rect 496 1127 503 1403
rect 596 1216 603 1333
rect 616 1247 623 1392
rect 676 1387 683 1533
rect 736 1436 743 1473
rect 816 1467 823 1733
rect 847 1703 860 1707
rect 847 1696 863 1703
rect 847 1693 860 1696
rect 836 1627 843 1693
rect 896 1467 903 1693
rect 773 1448 787 1453
rect 916 1448 923 1753
rect 936 1587 943 1873
rect 1076 1867 1083 1923
rect 976 1736 983 1813
rect 1036 1667 1043 1793
rect 1076 1736 1083 1853
rect 1116 1736 1123 1893
rect 1136 1807 1143 2196
rect 1216 2167 1223 2223
rect 1156 1743 1163 2013
rect 1296 1927 1303 2153
rect 1236 1827 1243 1923
rect 1196 1747 1203 1813
rect 1256 1767 1263 1853
rect 1276 1807 1283 1913
rect 1246 1753 1247 1760
rect 1156 1736 1183 1743
rect 1136 1667 1143 1703
rect 756 1327 763 1403
rect 836 1347 843 1434
rect 516 987 523 1214
rect 620 1183 633 1187
rect 616 1176 633 1183
rect 620 1173 633 1176
rect 576 1127 583 1172
rect 656 1167 663 1253
rect 696 1228 703 1273
rect 736 1216 743 1253
rect 536 947 543 1073
rect 616 1007 623 1153
rect 716 1127 723 1183
rect 756 1167 763 1183
rect 433 920 447 933
rect 436 916 443 920
rect 533 923 547 933
rect 533 920 563 923
rect 536 916 563 920
rect 616 916 623 993
rect 256 660 263 663
rect 253 647 267 660
rect 253 627 267 633
rect 116 427 123 553
rect 76 396 103 403
rect 233 400 247 413
rect 236 396 243 400
rect 276 396 283 473
rect 116 360 123 363
rect 113 347 127 360
rect 156 267 163 394
rect 216 360 223 363
rect 213 347 227 360
rect 256 327 263 363
rect 156 176 163 253
rect 253 188 267 193
rect 296 176 303 353
rect 316 347 323 652
rect 336 487 343 713
rect 396 696 403 873
rect 416 827 423 883
rect 456 747 463 872
rect 596 827 603 883
rect 596 747 603 813
rect 536 696 543 733
rect 416 567 423 663
rect 476 627 483 694
rect 596 663 603 693
rect 396 408 403 433
rect 196 147 203 174
rect 336 147 343 313
rect 376 307 383 363
rect 396 176 403 273
rect 436 188 443 313
rect 456 287 463 573
rect 516 567 523 663
rect 576 656 603 663
rect 476 307 483 473
rect 516 408 523 493
rect 596 483 603 593
rect 616 547 623 653
rect 596 476 623 483
rect 616 367 623 476
rect 636 408 643 933
rect 656 707 663 993
rect 716 916 723 973
rect 756 967 763 1153
rect 796 1027 803 1253
rect 816 1087 823 1313
rect 896 1247 903 1403
rect 916 1216 923 1313
rect 956 1186 963 1333
rect 976 1228 983 1433
rect 996 1407 1003 1653
rect 1033 1440 1047 1453
rect 1036 1436 1043 1440
rect 1076 1436 1083 1533
rect 1016 1216 1023 1273
rect 1056 1247 1063 1403
rect 1116 1383 1123 1473
rect 1156 1436 1163 1613
rect 1176 1607 1183 1736
rect 1233 1740 1247 1753
rect 1236 1736 1243 1740
rect 1296 1747 1303 1892
rect 1116 1376 1133 1383
rect 1076 1223 1083 1253
rect 1056 1216 1083 1223
rect 996 1180 1003 1183
rect 856 1147 863 1172
rect 993 1167 1007 1180
rect 1036 1147 1043 1183
rect 696 787 703 883
rect 667 696 683 703
rect 716 696 723 813
rect 736 767 743 872
rect 796 707 803 953
rect 836 928 843 973
rect 876 916 883 953
rect 936 887 943 1133
rect 896 723 903 872
rect 876 716 903 723
rect 696 627 703 663
rect 756 647 763 693
rect 776 607 783 694
rect 876 696 883 716
rect 816 567 823 652
rect 856 647 863 663
rect 896 660 903 663
rect 893 647 907 660
rect 856 636 873 647
rect 860 633 873 636
rect 696 396 703 433
rect 496 327 503 353
rect 536 343 543 363
rect 516 336 543 343
rect 516 267 523 336
rect 96 140 103 143
rect 93 127 107 140
rect 136 123 143 143
rect 173 127 187 133
rect 136 116 163 123
rect 156 103 163 116
rect 193 103 207 112
rect 236 107 243 132
rect 273 127 287 132
rect 156 100 207 103
rect 156 96 203 100
rect 356 87 363 173
rect 416 140 423 143
rect 413 127 427 140
rect 496 127 503 193
rect 516 147 523 253
rect 573 188 587 193
rect 616 176 623 233
rect 636 188 643 394
rect 776 367 783 553
rect 876 507 883 553
rect 856 447 863 473
rect 836 396 843 433
rect 876 396 883 493
rect 676 307 683 363
rect 656 296 673 303
rect 656 167 663 296
rect 753 180 767 193
rect 756 176 763 180
rect 796 167 803 333
rect 816 307 823 363
rect 916 267 923 653
rect 936 647 943 753
rect 956 707 963 1073
rect 1016 947 1023 1053
rect 973 920 987 933
rect 976 916 983 920
rect 1056 887 1063 1153
rect 1096 827 1103 1233
rect 1116 928 1123 1333
rect 1136 1227 1143 1373
rect 1176 1327 1183 1403
rect 1176 1228 1183 1253
rect 1216 1227 1223 1593
rect 1156 1180 1163 1183
rect 1153 1167 1167 1180
rect 1196 1163 1203 1183
rect 1176 1156 1203 1163
rect 1176 1143 1183 1156
rect 1156 1136 1183 1143
rect 1156 947 1163 1136
rect 1127 916 1143 923
rect 1176 916 1183 1053
rect 1216 887 1223 1173
rect 1236 1147 1243 1653
rect 1276 1547 1283 1673
rect 1296 1667 1303 1693
rect 1316 1647 1323 2513
rect 1356 2488 1363 2553
rect 1376 2367 1383 2443
rect 1436 2407 1443 2933
rect 1616 2923 1623 2994
rect 1596 2916 1623 2923
rect 1456 2807 1463 2893
rect 1516 2776 1523 2913
rect 1536 2847 1543 2873
rect 1596 2787 1603 2916
rect 1636 2803 1643 3033
rect 1656 3007 1663 3213
rect 1676 3107 1683 3256
rect 1696 3227 1703 3973
rect 1736 3947 1743 4034
rect 1756 3987 1763 4273
rect 1776 4247 1783 4296
rect 1816 4187 1823 4493
rect 1836 4147 1843 4493
rect 1876 4336 1883 4453
rect 1896 4363 1903 4793
rect 1916 4747 1923 4823
rect 1936 4556 1943 4673
rect 1956 4607 1963 4813
rect 1976 4787 1983 4993
rect 1996 4887 2003 5013
rect 2016 4907 2023 5173
rect 2056 5087 2063 5236
rect 2236 5107 2243 5343
rect 2356 5267 2363 5343
rect 2036 5047 2043 5074
rect 2093 5080 2107 5093
rect 2096 5076 2103 5080
rect 2176 5047 2183 5074
rect 2056 4927 2063 5033
rect 2116 4967 2123 5043
rect 2156 4967 2163 4993
rect 2047 4883 2060 4887
rect 2047 4873 2063 4883
rect 1916 4387 1923 4553
rect 1976 4447 1983 4523
rect 1996 4467 2003 4873
rect 2056 4856 2063 4873
rect 2093 4867 2107 4873
rect 1896 4356 1923 4363
rect 1916 4348 1923 4356
rect 1896 4300 1903 4303
rect 1893 4287 1907 4300
rect 1820 4004 1833 4007
rect 1773 3987 1787 3993
rect 1816 3993 1833 4004
rect 1736 3816 1743 3893
rect 1776 3816 1783 3973
rect 1816 3827 1823 3993
rect 1836 3883 1843 3972
rect 1856 3907 1863 4273
rect 1876 4187 1883 4213
rect 1876 4007 1883 4133
rect 1916 4063 1923 4253
rect 1936 4247 1943 4303
rect 1896 4060 1923 4063
rect 1893 4056 1923 4060
rect 1893 4047 1907 4056
rect 1956 4047 1963 4293
rect 1976 4127 1983 4433
rect 1996 4043 2003 4373
rect 2016 4367 2023 4813
rect 2036 4687 2043 4823
rect 2076 4787 2083 4823
rect 2033 4567 2047 4573
rect 2056 4556 2063 4593
rect 2076 4583 2083 4773
rect 2096 4687 2103 4753
rect 2116 4747 2123 4913
rect 2136 4887 2143 4933
rect 2196 4856 2203 4893
rect 2236 4867 2243 5032
rect 2296 4927 2303 5133
rect 2376 5076 2383 5133
rect 2396 5067 2403 5173
rect 2136 4827 2143 4852
rect 2256 4787 2263 4913
rect 2276 4867 2283 4893
rect 2316 4856 2323 4973
rect 2356 4887 2363 4913
rect 2356 4856 2363 4873
rect 2187 4773 2193 4787
rect 2276 4763 2283 4813
rect 2336 4767 2343 4823
rect 2256 4756 2283 4763
rect 2076 4576 2103 4583
rect 2096 4556 2103 4576
rect 2196 4547 2203 4752
rect 2033 4507 2047 4512
rect 2116 4487 2123 4512
rect 2107 4476 2123 4487
rect 2107 4473 2120 4476
rect 2136 4367 2143 4453
rect 2156 4447 2163 4543
rect 2216 4427 2223 4543
rect 2256 4447 2263 4756
rect 2396 4647 2403 5032
rect 2416 4927 2423 5374
rect 2436 5343 2443 5563
rect 2476 5560 2483 5563
rect 2473 5547 2487 5560
rect 2516 5547 2523 5894
rect 2536 5867 2543 5913
rect 2596 5896 2603 5973
rect 2576 5860 2583 5863
rect 2573 5847 2587 5860
rect 2656 5847 2663 6073
rect 2716 5896 2723 6013
rect 2756 6007 2763 6134
rect 2876 6116 2883 6296
rect 2896 6296 2923 6303
rect 2896 6107 2903 6296
rect 3336 6267 3343 6303
rect 3916 6296 3943 6303
rect 2836 5987 2843 6083
rect 2856 5907 2863 6013
rect 2916 5987 2923 6103
rect 2956 6103 2963 6193
rect 2956 6096 2983 6103
rect 2816 5863 2823 5894
rect 2936 5896 2943 6093
rect 2696 5827 2703 5863
rect 2736 5860 2743 5863
rect 2733 5847 2747 5860
rect 2736 5767 2743 5793
rect 2636 5587 2643 5653
rect 2596 5547 2603 5563
rect 2656 5547 2663 5613
rect 2716 5596 2723 5653
rect 2576 5536 2593 5543
rect 2496 5376 2503 5453
rect 2536 5376 2543 5453
rect 2436 5336 2463 5343
rect 2456 5307 2463 5336
rect 2476 5127 2483 5343
rect 2516 5247 2523 5343
rect 2447 5043 2460 5047
rect 2447 5036 2463 5043
rect 2447 5033 2460 5036
rect 2436 4903 2443 5033
rect 2536 5027 2543 5313
rect 2556 5087 2563 5333
rect 2576 5107 2583 5536
rect 2633 5507 2647 5513
rect 2596 5187 2603 5493
rect 2656 5427 2663 5512
rect 2633 5380 2647 5393
rect 2636 5376 2643 5380
rect 2676 5376 2683 5493
rect 2696 5387 2703 5563
rect 2776 5547 2783 5863
rect 2796 5856 2823 5863
rect 2796 5563 2803 5856
rect 2856 5727 2863 5893
rect 2896 5860 2903 5863
rect 2893 5847 2907 5860
rect 2827 5603 2840 5607
rect 2827 5596 2843 5603
rect 2876 5596 2883 5733
rect 2896 5627 2903 5753
rect 2827 5593 2840 5596
rect 2936 5607 2943 5673
rect 2796 5556 2823 5563
rect 2733 5527 2747 5531
rect 2656 5107 2663 5343
rect 2716 5327 2723 5433
rect 2816 5376 2823 5556
rect 2756 5207 2763 5343
rect 2796 5323 2803 5343
rect 2796 5316 2823 5323
rect 2696 5076 2703 5133
rect 2796 5107 2803 5253
rect 2816 5247 2823 5316
rect 2816 5147 2823 5233
rect 2856 5187 2863 5531
rect 2936 5407 2943 5553
rect 2956 5383 2963 5693
rect 2976 5647 2983 6096
rect 3256 6103 3263 6253
rect 3256 6096 3283 6103
rect 2996 5947 3003 6094
rect 3436 6103 3443 6253
rect 3416 6096 3443 6103
rect 3036 5863 3043 5993
rect 3276 5987 3283 6073
rect 3296 6007 3303 6093
rect 3676 6067 3683 6253
rect 3716 6100 3723 6103
rect 3713 6087 3727 6100
rect 3776 6067 3783 6103
rect 3107 5936 3123 5943
rect 3096 5896 3103 5933
rect 3036 5856 3063 5863
rect 3116 5847 3123 5936
rect 3216 5896 3223 5973
rect 3296 5956 3333 5963
rect 3136 5827 3143 5894
rect 3296 5866 3303 5956
rect 3316 5908 3323 5933
rect 2976 5566 2983 5593
rect 2976 5427 2983 5473
rect 2936 5376 2963 5383
rect 2876 5307 2883 5373
rect 2916 5267 2923 5343
rect 2936 5247 2943 5313
rect 2733 5080 2747 5093
rect 2736 5076 2743 5080
rect 2567 5043 2580 5047
rect 2620 5043 2633 5047
rect 2567 5033 2583 5043
rect 2616 5036 2633 5043
rect 2620 5033 2633 5036
rect 2416 4896 2443 4903
rect 2416 4867 2423 4896
rect 2456 4883 2463 4933
rect 2496 4887 2503 4913
rect 2436 4876 2463 4883
rect 2436 4856 2443 4876
rect 2456 4747 2463 4812
rect 2536 4747 2543 4893
rect 2576 4867 2583 5033
rect 2596 4856 2603 4913
rect 2636 4856 2643 5012
rect 2656 4883 2663 5072
rect 2776 4987 2783 5093
rect 2796 5047 2803 5093
rect 2876 5076 2883 5153
rect 2916 5087 2923 5193
rect 2956 5087 2963 5253
rect 3016 5227 3023 5473
rect 3036 5356 3043 5493
rect 3056 5467 3063 5513
rect 3076 5487 3083 5793
rect 3096 5707 3103 5753
rect 3096 5566 3103 5693
rect 3136 5596 3143 5773
rect 3196 5747 3203 5863
rect 3356 5860 3363 5863
rect 3353 5847 3367 5860
rect 3256 5603 3263 5633
rect 3256 5596 3283 5603
rect 3196 5567 3203 5594
rect 3176 5467 3183 5533
rect 3256 5507 3263 5596
rect 3256 5467 3263 5493
rect 3276 5487 3283 5533
rect 3080 5463 3093 5467
rect 3076 5453 3093 5463
rect 3076 5407 3083 5453
rect 2900 5043 2913 5047
rect 2856 5040 2863 5043
rect 2853 5027 2867 5040
rect 2896 5036 2913 5043
rect 2900 5033 2913 5036
rect 2656 4880 2683 4883
rect 2656 4876 2687 4880
rect 2673 4867 2687 4876
rect 2556 4807 2563 4853
rect 2616 4820 2623 4823
rect 2613 4807 2627 4820
rect 2626 4800 2627 4807
rect 2393 4540 2407 4553
rect 2396 4536 2403 4540
rect 2296 4376 2303 4433
rect 1976 4036 2003 4043
rect 2016 4036 2023 4292
rect 2076 4247 2083 4293
rect 2096 4167 2103 4353
rect 2236 4336 2263 4343
rect 2136 4267 2143 4303
rect 2056 4036 2063 4153
rect 1896 3996 1923 4003
rect 1896 3947 1903 3996
rect 1836 3876 1863 3883
rect 1836 3807 1843 3853
rect 1716 3527 1723 3773
rect 1756 3707 1763 3783
rect 1796 3607 1803 3783
rect 1796 3527 1803 3593
rect 1727 3483 1740 3487
rect 1727 3473 1743 3483
rect 1716 3307 1723 3433
rect 1736 3367 1743 3473
rect 1756 3407 1763 3453
rect 1776 3323 1783 3483
rect 1793 3467 1807 3473
rect 1816 3403 1823 3533
rect 1767 3316 1783 3323
rect 1796 3396 1823 3403
rect 1753 3300 1767 3313
rect 1756 3296 1763 3300
rect 1713 3247 1727 3253
rect 1676 3027 1683 3053
rect 1693 3000 1707 3013
rect 1696 2996 1703 3000
rect 1656 2927 1663 2953
rect 1776 2947 1783 2994
rect 1616 2796 1643 2803
rect 1616 2776 1623 2796
rect 1653 2780 1667 2793
rect 1656 2776 1663 2780
rect 1696 2747 1703 2793
rect 1456 2427 1463 2733
rect 1536 2723 1543 2743
rect 1516 2716 1543 2723
rect 1496 2476 1503 2553
rect 1516 2547 1523 2716
rect 1716 2607 1723 2913
rect 1796 2887 1803 3396
rect 1836 3387 1843 3772
rect 1856 3667 1863 3876
rect 1896 3847 1903 3933
rect 1916 3816 1923 3973
rect 1956 3863 1963 3993
rect 1976 3887 1983 4036
rect 1993 3987 2007 3993
rect 2036 3867 2043 4003
rect 2096 3927 2103 4113
rect 2116 4003 2123 4053
rect 2156 4036 2163 4093
rect 2176 4087 2183 4303
rect 2196 4247 2203 4293
rect 2236 4267 2243 4336
rect 2436 4323 2443 4413
rect 2476 4327 2483 4433
rect 2436 4316 2463 4323
rect 2356 4296 2383 4303
rect 2376 4243 2383 4296
rect 2356 4236 2383 4243
rect 2196 4187 2203 4233
rect 2196 4036 2203 4173
rect 2116 3996 2143 4003
rect 1956 3856 1983 3863
rect 1876 3647 1883 3773
rect 1916 3687 1923 3713
rect 1936 3707 1943 3783
rect 1976 3727 1983 3856
rect 2076 3827 2083 3853
rect 1996 3747 2003 3814
rect 2116 3803 2123 3933
rect 2136 3827 2143 3996
rect 2156 3947 2163 3973
rect 2196 3816 2203 3973
rect 2116 3796 2143 3803
rect 2056 3687 2063 3783
rect 1956 3627 1963 3673
rect 1893 3528 1907 3533
rect 1936 3516 1943 3593
rect 1856 3447 1863 3473
rect 1816 3266 1823 3313
rect 1856 3308 1863 3353
rect 1896 3296 1903 3453
rect 1916 3427 1923 3483
rect 1976 3427 1983 3653
rect 2076 3527 2083 3773
rect 2096 3487 2103 3794
rect 2113 3767 2127 3773
rect 1996 3347 2003 3393
rect 2036 3387 2043 3483
rect 1947 3333 1953 3347
rect 1916 3260 1923 3263
rect 1913 3247 1927 3260
rect 1816 3007 1823 3093
rect 1836 2996 1843 3053
rect 1876 3027 1883 3173
rect 1873 3000 1887 3013
rect 1876 2996 1883 3000
rect 1856 2960 1863 2963
rect 1853 2947 1867 2960
rect 1896 2907 1903 2953
rect 1916 2927 1923 3212
rect 1936 3107 1943 3253
rect 1956 3227 1963 3273
rect 1976 3266 1983 3333
rect 2036 3296 2043 3352
rect 2076 3347 2083 3473
rect 2116 3367 2123 3713
rect 2136 3307 2143 3796
rect 2156 3528 2163 3751
rect 2216 3587 2223 3973
rect 2236 3867 2243 4093
rect 2256 4047 2263 4113
rect 2316 4048 2323 4093
rect 2356 4087 2363 4236
rect 2296 3967 2303 4003
rect 2276 3787 2283 3853
rect 2316 3803 2323 3973
rect 2336 3947 2343 4003
rect 2376 3987 2383 4193
rect 2396 4087 2403 4233
rect 2436 4207 2443 4316
rect 2476 4067 2483 4273
rect 2496 4127 2503 4633
rect 2556 4576 2563 4613
rect 2516 4487 2523 4543
rect 2596 4487 2603 4673
rect 2616 4427 2623 4753
rect 2636 4467 2643 4793
rect 2696 4787 2703 4913
rect 2716 4787 2723 4973
rect 2813 4860 2827 4873
rect 2816 4856 2823 4860
rect 2747 4823 2760 4827
rect 2747 4816 2763 4823
rect 2796 4820 2803 4823
rect 2747 4813 2760 4816
rect 2793 4807 2807 4820
rect 2806 4800 2807 4807
rect 2720 4766 2733 4767
rect 2676 4727 2683 4753
rect 2727 4753 2733 4766
rect 2676 4607 2683 4673
rect 2696 4556 2703 4693
rect 2796 4647 2803 4713
rect 2733 4607 2747 4613
rect 2796 4563 2803 4612
rect 2816 4587 2823 4793
rect 2833 4727 2847 4733
rect 2836 4627 2843 4692
rect 2856 4687 2863 4893
rect 2876 4807 2883 4973
rect 2876 4603 2883 4733
rect 2896 4727 2903 4913
rect 2936 4887 2943 5074
rect 3016 5076 3023 5213
rect 3056 5108 3063 5273
rect 3076 5207 3083 5354
rect 3316 5327 3323 5813
rect 3356 5443 3363 5713
rect 3336 5436 3363 5443
rect 3336 5356 3343 5436
rect 3356 5367 3363 5413
rect 3376 5407 3383 5894
rect 3396 5608 3403 6053
rect 3776 6027 3783 6053
rect 3416 5907 3423 6013
rect 3456 5896 3463 5953
rect 3573 5908 3587 5913
rect 3713 5900 3727 5913
rect 3716 5896 3723 5900
rect 3836 5896 3843 6094
rect 3876 5947 3883 6133
rect 3936 6116 3943 6296
rect 4576 6296 4603 6303
rect 4736 6296 4763 6303
rect 4876 6296 4903 6303
rect 4036 6103 4043 6253
rect 4016 6096 4043 6103
rect 4296 6096 4323 6103
rect 4296 6087 4303 6096
rect 3896 6080 3903 6083
rect 3893 6067 3907 6080
rect 3656 5867 3663 5894
rect 3596 5807 3603 5863
rect 3916 5866 3923 5893
rect 3656 5827 3663 5853
rect 3427 5713 3433 5727
rect 3656 5608 3663 5733
rect 3696 5707 3703 5863
rect 3696 5627 3703 5693
rect 3436 5527 3443 5594
rect 3753 5600 3767 5613
rect 3756 5596 3763 5600
rect 3816 5607 3823 5863
rect 3856 5807 3863 5863
rect 3856 5647 3863 5793
rect 3936 5667 3943 5933
rect 3996 5896 4003 5993
rect 4056 5866 4063 5913
rect 4116 5896 4123 5973
rect 4236 5876 4263 5883
rect 4096 5827 4103 5863
rect 3856 5623 3863 5633
rect 3836 5616 3863 5623
rect 3396 5367 3403 5513
rect 3576 5487 3583 5593
rect 3413 5327 3427 5333
rect 3216 5147 3223 5313
rect 3376 5287 3383 5312
rect 3436 5207 3443 5413
rect 3487 5383 3500 5387
rect 3487 5376 3503 5383
rect 3536 5376 3543 5473
rect 3576 5387 3583 5452
rect 3487 5373 3500 5376
rect 3456 5326 3463 5373
rect 3596 5347 3603 5593
rect 3776 5543 3783 5552
rect 3776 5536 3803 5543
rect 3656 5376 3663 5413
rect 3476 5267 3483 5333
rect 3513 5307 3527 5311
rect 3236 5167 3243 5193
rect 3216 5107 3223 5133
rect 2956 5007 2963 5033
rect 2956 4727 2963 4823
rect 2867 4596 2883 4603
rect 2796 4556 2823 4563
rect 2856 4556 2863 4593
rect 2896 4576 2903 4713
rect 2916 4607 2923 4673
rect 2716 4487 2723 4523
rect 2776 4487 2783 4553
rect 2936 4540 2943 4543
rect 2796 4427 2803 4513
rect 2466 4053 2467 4060
rect 2453 4048 2467 4053
rect 2296 3796 2323 3803
rect 2256 3547 2263 3733
rect 2216 3483 2223 3513
rect 2216 3476 2243 3483
rect 2196 3463 2203 3472
rect 2196 3456 2223 3463
rect 2180 3323 2193 3327
rect 2176 3313 2193 3323
rect 2056 3243 2063 3263
rect 2036 3236 2063 3243
rect 1976 3107 1983 3133
rect 1816 2747 1823 2774
rect 1807 2723 1820 2727
rect 1807 2713 1823 2723
rect 1536 2476 1543 2513
rect 1656 2507 1663 2533
rect 1573 2480 1587 2493
rect 1576 2476 1583 2480
rect 1516 2440 1523 2443
rect 1513 2427 1527 2440
rect 1353 2260 1367 2273
rect 1356 2256 1363 2260
rect 1416 2256 1423 2333
rect 1436 2287 1443 2313
rect 1476 2223 1483 2273
rect 1396 2220 1403 2223
rect 1376 2187 1383 2213
rect 1393 2207 1407 2220
rect 1456 2216 1483 2223
rect 1376 1987 1383 2053
rect 1373 1960 1387 1973
rect 1376 1956 1383 1960
rect 1336 1627 1343 1913
rect 1356 1887 1363 1923
rect 1416 1847 1423 2113
rect 1436 1923 1443 2193
rect 1496 2107 1503 2413
rect 1516 2167 1523 2333
rect 1536 2047 1543 2293
rect 1556 2267 1563 2411
rect 1596 2256 1603 2393
rect 1616 2307 1623 2493
rect 1656 2476 1683 2483
rect 1736 2476 1743 2533
rect 1636 2327 1643 2373
rect 1556 2147 1563 2213
rect 1576 2187 1583 2223
rect 1656 2087 1663 2476
rect 1776 2403 1783 2473
rect 1796 2446 1803 2653
rect 1816 2647 1823 2713
rect 1836 2707 1843 2793
rect 1896 2776 1903 2893
rect 1936 2847 1943 3013
rect 1956 2996 1983 3003
rect 2036 2996 2043 3236
rect 2096 3067 2103 3253
rect 2116 3043 2123 3294
rect 2176 3296 2183 3313
rect 2216 3307 2223 3456
rect 2196 3227 2203 3263
rect 2196 3127 2203 3213
rect 2096 3036 2123 3043
rect 1956 2947 1963 2996
rect 2096 2967 2103 3036
rect 2216 3003 2223 3173
rect 2196 2996 2223 3003
rect 2136 2960 2143 2963
rect 2133 2947 2147 2960
rect 1916 2736 1943 2743
rect 1876 2567 1883 2732
rect 1856 2436 1883 2443
rect 1756 2396 1783 2403
rect 1507 1956 1523 1963
rect 1436 1916 1463 1923
rect 1376 1736 1383 1793
rect 1296 1483 1303 1553
rect 1276 1476 1303 1483
rect 1276 1436 1283 1476
rect 1316 1436 1323 1533
rect 1296 1216 1303 1353
rect 1336 1347 1343 1403
rect 1376 1227 1383 1613
rect 1256 1127 1263 1214
rect 1396 1183 1403 1633
rect 1436 1567 1443 1734
rect 1456 1607 1463 1893
rect 1476 1747 1483 1853
rect 1516 1787 1523 1956
rect 1536 1867 1543 2033
rect 1616 1956 1623 2073
rect 1636 1920 1643 1923
rect 1633 1907 1647 1920
rect 1487 1703 1500 1707
rect 1487 1696 1503 1703
rect 1487 1693 1500 1696
rect 1536 1607 1543 1703
rect 1416 1447 1423 1493
rect 1436 1436 1443 1513
rect 1516 1447 1523 1553
rect 1416 1347 1423 1393
rect 1496 1396 1513 1403
rect 1476 1216 1483 1333
rect 1496 1287 1503 1373
rect 1496 1247 1503 1273
rect 1516 1216 1523 1393
rect 1536 1367 1543 1453
rect 1556 1447 1563 1613
rect 1576 1467 1583 1833
rect 1596 1747 1603 1793
rect 1616 1736 1623 1833
rect 1676 1763 1683 2313
rect 1713 2260 1727 2273
rect 1756 2267 1763 2396
rect 1716 2256 1723 2260
rect 1696 1967 1703 2133
rect 1756 1967 1763 2213
rect 1776 2167 1783 2353
rect 1876 2347 1883 2436
rect 1736 1956 1753 1963
rect 1716 1887 1723 1923
rect 1676 1756 1703 1763
rect 1653 1740 1667 1753
rect 1656 1736 1663 1740
rect 1636 1403 1643 1653
rect 1656 1487 1663 1673
rect 1696 1667 1703 1756
rect 1756 1763 1763 1913
rect 1796 1827 1803 2293
rect 1856 2268 1863 2313
rect 1896 2307 1903 2453
rect 1916 2387 1923 2713
rect 1936 2703 1943 2736
rect 1956 2727 1963 2873
rect 1976 2787 1983 2853
rect 2016 2827 2023 2931
rect 2236 2907 2243 3476
rect 2256 3407 2263 3493
rect 2256 3266 2263 3313
rect 2276 3307 2283 3773
rect 2336 3763 2343 3912
rect 2436 3907 2443 4003
rect 2516 3987 2523 4153
rect 2593 4040 2607 4053
rect 2636 4043 2643 4323
rect 2736 4167 2743 4393
rect 2776 4167 2783 4273
rect 2596 4036 2603 4040
rect 2636 4036 2663 4043
rect 2316 3756 2343 3763
rect 2316 3547 2323 3756
rect 2576 3647 2583 4003
rect 2596 3796 2603 3973
rect 2656 3967 2663 4036
rect 2676 4007 2683 4153
rect 2753 4040 2767 4053
rect 2756 4036 2763 4040
rect 2616 3807 2623 3833
rect 2676 3787 2683 3893
rect 2640 3763 2653 3767
rect 2636 3753 2653 3763
rect 2336 3503 2343 3573
rect 2296 3496 2343 3503
rect 2576 3487 2583 3612
rect 2636 3536 2643 3753
rect 2676 3703 2683 3752
rect 2656 3700 2683 3703
rect 2653 3696 2683 3700
rect 2653 3687 2667 3696
rect 2696 3687 2703 4033
rect 2776 4007 2783 4132
rect 2796 3927 2803 4153
rect 2816 4007 2823 4213
rect 2836 4107 2843 4453
rect 2856 4147 2863 4413
rect 2876 4068 2883 4453
rect 2916 4367 2923 4533
rect 2933 4527 2947 4540
rect 2936 4336 2943 4373
rect 2956 4363 2963 4692
rect 2976 4687 2983 4953
rect 2996 4826 3003 5043
rect 3076 4856 3083 4973
rect 3116 4947 3123 5093
rect 3356 4967 3363 5073
rect 3416 5063 3423 5113
rect 3396 5056 3423 5063
rect 3456 5027 3463 5063
rect 3116 4887 3123 4912
rect 3113 4860 3127 4873
rect 3216 4868 3223 4953
rect 3116 4856 3123 4860
rect 3356 4856 3363 4932
rect 3096 4820 3103 4823
rect 3093 4807 3107 4820
rect 3416 4823 3423 5013
rect 3436 4826 3443 4973
rect 3476 4967 3483 5153
rect 3496 4856 3503 5293
rect 3536 5167 3543 5253
rect 3556 5207 3563 5343
rect 3716 5346 3723 5433
rect 3776 5376 3783 5493
rect 3796 5403 3803 5536
rect 3816 5507 3823 5553
rect 3796 5400 3823 5403
rect 3796 5396 3827 5400
rect 3813 5387 3827 5396
rect 3836 5347 3843 5616
rect 3976 5587 3983 5713
rect 4016 5596 4023 5813
rect 4096 5607 4103 5693
rect 4236 5667 4243 5876
rect 4296 5747 4303 6073
rect 4376 6067 4383 6103
rect 4396 6087 4403 6173
rect 4576 6116 4583 6296
rect 4756 6116 4763 6296
rect 4376 6007 4383 6053
rect 4576 5887 4583 5933
rect 4616 5887 4623 6083
rect 4536 5876 4563 5883
rect 4536 5847 4543 5876
rect 4256 5687 4263 5733
rect 4196 5616 4203 5653
rect 3856 5347 3863 5373
rect 3616 5336 3643 5343
rect 3576 5167 3583 5293
rect 3596 5127 3603 5312
rect 3616 5267 3623 5336
rect 3516 4887 3523 5063
rect 3556 5063 3563 5113
rect 3556 5056 3583 5063
rect 3536 4923 3543 5053
rect 3536 4916 3563 4923
rect 3536 4856 3543 4893
rect 3556 4867 3563 4916
rect 3576 4887 3583 5013
rect 3596 4987 3603 5033
rect 3396 4816 3423 4823
rect 3036 4543 3043 4573
rect 3056 4567 3063 4713
rect 3036 4536 3063 4543
rect 2956 4360 2983 4363
rect 2956 4356 2987 4360
rect 2973 4347 2987 4356
rect 2916 4247 2923 4303
rect 2916 4187 2923 4233
rect 2896 4067 2903 4113
rect 2916 4036 2923 4133
rect 2936 4047 2943 4273
rect 2996 4147 3003 4373
rect 3016 4127 3023 4353
rect 3073 4340 3087 4353
rect 3076 4336 3083 4340
rect 3096 4327 3103 4433
rect 3036 4300 3043 4303
rect 3033 4286 3047 4300
rect 3036 4147 3043 4193
rect 2716 3787 2723 3853
rect 2773 3820 2787 3833
rect 2776 3816 2783 3820
rect 2816 3816 2823 3853
rect 2836 3827 2843 3993
rect 2856 3967 2863 4003
rect 2896 3947 2903 4003
rect 2796 3780 2803 3783
rect 2793 3767 2807 3780
rect 2856 3767 2863 3913
rect 2956 3907 2963 4023
rect 2896 3816 2903 3853
rect 2933 3820 2947 3833
rect 2976 3827 2983 4013
rect 2936 3816 2943 3820
rect 2716 3727 2723 3752
rect 2696 3683 2713 3687
rect 2676 3676 2713 3683
rect 2676 3663 2683 3676
rect 2700 3673 2713 3676
rect 2656 3656 2683 3663
rect 2656 3547 2663 3656
rect 2673 3627 2687 3633
rect 2676 3507 2683 3553
rect 2296 3327 2303 3453
rect 2316 3296 2323 3473
rect 2360 3303 2373 3307
rect 2356 3296 2373 3303
rect 2360 3293 2373 3296
rect 2387 3296 2403 3303
rect 2016 2776 2023 2813
rect 2076 2746 2083 2893
rect 2113 2780 2127 2793
rect 2116 2776 2123 2780
rect 1936 2696 1963 2703
rect 1936 2407 1943 2593
rect 1956 2587 1963 2696
rect 1956 2507 1963 2573
rect 1996 2503 2003 2673
rect 2016 2647 2023 2713
rect 2036 2547 2043 2732
rect 2136 2707 2143 2743
rect 1996 2496 2023 2503
rect 2016 2446 2023 2496
rect 1956 2347 1963 2432
rect 2013 2383 2027 2393
rect 2013 2380 2043 2383
rect 2016 2376 2043 2380
rect 1896 2256 1903 2293
rect 1996 2287 2003 2333
rect 2036 2287 2043 2376
rect 1936 2226 1943 2273
rect 2056 2256 2063 2633
rect 2116 2476 2123 2613
rect 2176 2467 2183 2793
rect 2276 2776 2283 3193
rect 2296 2996 2303 3213
rect 2336 2887 2343 2963
rect 2356 2807 2363 3173
rect 2376 2967 2383 3253
rect 2396 3167 2403 3296
rect 2416 3227 2423 3313
rect 2496 3296 2503 3393
rect 2476 3260 2483 3263
rect 2473 3247 2487 3260
rect 2436 3107 2443 3133
rect 2476 3127 2483 3212
rect 2396 2943 2403 3033
rect 2456 2996 2463 3073
rect 2396 2936 2423 2943
rect 2416 2776 2423 2936
rect 2456 2787 2463 2833
rect 2196 2487 2203 2774
rect 2236 2476 2243 2693
rect 2256 2627 2263 2743
rect 2296 2740 2303 2743
rect 2293 2727 2307 2740
rect 2280 2483 2293 2487
rect 2276 2476 2293 2483
rect 2280 2473 2293 2476
rect 2136 2440 2143 2443
rect 2133 2427 2147 2440
rect 2207 2443 2220 2447
rect 2207 2436 2223 2443
rect 2256 2440 2263 2443
rect 2207 2433 2220 2436
rect 2253 2427 2267 2440
rect 2096 2226 2103 2333
rect 2176 2256 2183 2413
rect 1836 2187 1843 2223
rect 1996 2220 2003 2223
rect 1993 2207 2007 2220
rect 2116 2223 2123 2253
rect 2116 2216 2163 2223
rect 2196 2220 2203 2223
rect 1976 2127 1983 2193
rect 1856 1967 1863 2113
rect 1876 1956 1883 2093
rect 1936 1956 1943 2053
rect 1836 1916 1853 1923
rect 1856 1847 1863 1913
rect 1816 1807 1823 1833
rect 1736 1760 1763 1763
rect 1733 1756 1763 1760
rect 1716 1667 1723 1753
rect 1733 1747 1747 1756
rect 1716 1627 1723 1653
rect 1736 1567 1743 1693
rect 1796 1647 1803 1703
rect 1676 1436 1683 1493
rect 1716 1436 1723 1493
rect 1756 1447 1763 1613
rect 1796 1527 1803 1633
rect 1773 1487 1787 1493
rect 1796 1483 1803 1513
rect 1816 1507 1823 1653
rect 1796 1476 1823 1483
rect 1636 1396 1663 1403
rect 1536 1227 1543 1313
rect 1296 1047 1303 1153
rect 1316 1147 1323 1183
rect 1356 1180 1363 1183
rect 1353 1167 1367 1180
rect 1376 1176 1403 1183
rect 1336 1087 1343 1153
rect 1036 696 1043 793
rect 1076 666 1083 773
rect 1156 747 1163 883
rect 1236 863 1243 1013
rect 1256 916 1263 973
rect 1316 916 1323 973
rect 1336 867 1343 1033
rect 1356 947 1363 993
rect 1236 856 1263 863
rect 976 607 983 663
rect 1096 567 1103 733
rect 1196 696 1203 733
rect 1136 587 1143 663
rect 1236 627 1243 694
rect 1256 663 1263 856
rect 1336 767 1343 813
rect 1356 807 1363 893
rect 1376 783 1383 1176
rect 1396 923 1403 973
rect 1416 947 1423 1213
rect 1456 1127 1463 1183
rect 1556 1167 1563 1293
rect 1613 1220 1627 1233
rect 1616 1216 1623 1220
rect 1656 1216 1663 1396
rect 1473 1087 1487 1093
rect 1467 1080 1487 1087
rect 1467 1076 1483 1080
rect 1467 1073 1480 1076
rect 1496 1007 1503 1113
rect 1396 916 1423 923
rect 1393 807 1407 813
rect 1376 776 1403 783
rect 1356 696 1363 772
rect 1396 687 1403 776
rect 1256 656 1273 663
rect 1273 647 1287 653
rect 1296 627 1303 663
rect 1336 660 1343 663
rect 1333 647 1347 660
rect 936 407 943 473
rect 976 396 983 513
rect 1087 453 1093 467
rect 1033 447 1047 453
rect 1073 427 1087 432
rect 1013 400 1027 413
rect 1016 396 1023 400
rect 1136 396 1143 513
rect 1176 487 1183 613
rect 1316 587 1323 633
rect 1196 447 1203 493
rect 1196 407 1203 433
rect 1356 407 1363 593
rect 1396 463 1403 673
rect 1416 667 1423 853
rect 1436 747 1443 883
rect 1453 700 1467 713
rect 1456 696 1463 700
rect 1496 696 1503 833
rect 1516 767 1523 893
rect 1536 827 1543 953
rect 1556 927 1563 1073
rect 1636 1007 1643 1183
rect 1656 963 1663 1153
rect 1696 1087 1703 1233
rect 1716 1227 1723 1373
rect 1736 1247 1743 1403
rect 1776 1367 1783 1452
rect 1793 1447 1807 1453
rect 1816 1436 1823 1476
rect 1836 1467 1843 1734
rect 1856 1627 1863 1833
rect 1876 1667 1883 1793
rect 1896 1787 1903 1873
rect 1956 1867 1963 1993
rect 1976 1887 1983 2013
rect 1996 1807 2003 2152
rect 2016 2127 2023 2193
rect 2016 1926 2023 1973
rect 2056 1968 2063 2193
rect 2087 1983 2100 1987
rect 2087 1973 2103 1983
rect 2096 1956 2103 1973
rect 2136 1967 2143 2216
rect 2193 2207 2207 2220
rect 2236 2207 2243 2413
rect 2316 2288 2323 2693
rect 2336 2647 2343 2774
rect 2356 2607 2363 2733
rect 2396 2707 2403 2743
rect 2436 2740 2443 2743
rect 2433 2727 2447 2740
rect 2396 2587 2403 2633
rect 2436 2488 2443 2533
rect 2356 2476 2383 2483
rect 2356 2347 2363 2476
rect 2256 2226 2263 2273
rect 2356 2256 2363 2293
rect 2376 2267 2383 2413
rect 2116 1920 2123 1923
rect 1976 1707 1983 1773
rect 1896 1647 1903 1703
rect 1916 1623 1923 1673
rect 1896 1616 1923 1623
rect 1853 1440 1867 1453
rect 1856 1436 1863 1440
rect 1796 1228 1803 1293
rect 1647 956 1663 963
rect 1636 916 1643 953
rect 1653 927 1667 932
rect 1676 886 1683 933
rect 1696 923 1703 1033
rect 1716 947 1723 1173
rect 1776 1180 1783 1183
rect 1736 1067 1743 1172
rect 1773 1167 1787 1180
rect 1696 916 1723 923
rect 1753 920 1767 933
rect 1796 923 1803 993
rect 1816 947 1823 1173
rect 1836 1167 1843 1353
rect 1896 1347 1903 1616
rect 1916 1267 1923 1573
rect 1956 1567 1963 1703
rect 1996 1627 2003 1793
rect 2016 1687 2023 1912
rect 2113 1907 2127 1920
rect 2056 1736 2063 1833
rect 2136 1743 2143 1913
rect 2116 1736 2143 1743
rect 2156 1736 2163 1973
rect 2176 1907 2183 2093
rect 2196 1967 2203 2013
rect 2233 1960 2247 1973
rect 2276 1968 2283 2193
rect 2336 2067 2343 2223
rect 2396 2127 2403 2443
rect 2456 2387 2463 2733
rect 2476 2727 2483 2793
rect 2496 2687 2503 3093
rect 2516 2887 2523 3231
rect 2536 3007 2543 3053
rect 2556 3047 2563 3373
rect 2576 3367 2583 3413
rect 2596 3327 2603 3503
rect 2616 3387 2623 3493
rect 2676 3407 2683 3472
rect 2696 3447 2703 3653
rect 2747 3613 2753 3627
rect 2576 3266 2583 3293
rect 2616 3260 2623 3263
rect 2613 3247 2627 3260
rect 2656 3247 2663 3252
rect 2647 3236 2663 3247
rect 2647 3233 2660 3236
rect 2616 3207 2623 3233
rect 2576 3047 2583 3073
rect 2576 2996 2583 3033
rect 2696 3008 2703 3353
rect 2716 3227 2723 3533
rect 2736 3527 2743 3573
rect 2753 3548 2767 3553
rect 2776 3547 2783 3693
rect 2796 3547 2803 3613
rect 2836 3607 2843 3713
rect 2876 3707 2883 3773
rect 2916 3687 2923 3783
rect 2956 3667 2963 3783
rect 2996 3707 3003 4073
rect 3036 4067 3043 4133
rect 3036 3947 3043 3993
rect 3056 3927 3063 4233
rect 3156 4147 3163 4393
rect 3196 4367 3203 4713
rect 3236 4683 3243 4793
rect 3256 4707 3263 4812
rect 3376 4803 3383 4812
rect 3356 4796 3383 4803
rect 3236 4676 3263 4683
rect 3236 4507 3243 4543
rect 3236 4307 3243 4453
rect 3256 4287 3263 4676
rect 3316 4543 3323 4733
rect 3336 4687 3343 4733
rect 3296 4536 3323 4543
rect 3336 4407 3343 4553
rect 3356 4467 3363 4796
rect 3396 4527 3403 4816
rect 3416 4547 3423 4733
rect 3536 4687 3543 4753
rect 3576 4747 3583 4852
rect 3596 4826 3603 4933
rect 3616 4867 3623 5232
rect 3656 5227 3663 5293
rect 3856 4987 3863 5312
rect 3876 5287 3883 5563
rect 3916 5560 3923 5563
rect 4036 5560 4043 5563
rect 3913 5547 3927 5560
rect 4033 5547 4047 5560
rect 3893 5388 3907 5393
rect 3876 5187 3883 5233
rect 3896 5167 3903 5193
rect 3936 5103 3943 5332
rect 3916 5096 3943 5103
rect 3676 4936 3713 4943
rect 3676 4907 3683 4936
rect 3696 4887 3703 4913
rect 3696 4856 3703 4873
rect 3616 4767 3623 4813
rect 3736 4767 3743 4853
rect 3836 4843 3843 4953
rect 3856 4868 3863 4973
rect 3836 4836 3863 4843
rect 3653 4687 3667 4693
rect 3396 4487 3403 4513
rect 3196 4083 3203 4273
rect 3276 4267 3283 4353
rect 3333 4340 3347 4353
rect 3376 4347 3383 4373
rect 3336 4336 3343 4340
rect 3296 4227 3303 4293
rect 3196 4076 3223 4083
rect 3216 4027 3223 4076
rect 3296 4023 3303 4173
rect 3356 4167 3363 4303
rect 3396 4068 3403 4413
rect 3416 4347 3423 4493
rect 3456 4336 3463 4393
rect 3496 4348 3503 4673
rect 3516 4607 3523 4633
rect 3556 4556 3563 4593
rect 3596 4507 3603 4553
rect 3536 4328 3543 4373
rect 3416 4087 3423 4293
rect 3436 4267 3443 4303
rect 3296 4016 3323 4023
rect 3296 3927 3303 4016
rect 3016 3727 3023 3793
rect 2836 3536 2843 3593
rect 2876 3567 2883 3633
rect 2793 3520 2807 3533
rect 2896 3527 2903 3613
rect 3016 3607 3023 3713
rect 3036 3627 3043 3873
rect 3096 3816 3103 3873
rect 3116 3807 3123 3913
rect 3156 3806 3163 3833
rect 3176 3796 3183 3913
rect 3416 3907 3423 4023
rect 3116 3756 3143 3763
rect 3116 3727 3123 3756
rect 3116 3687 3123 3713
rect 3136 3607 3143 3733
rect 3156 3647 3163 3713
rect 2796 3516 2803 3520
rect 2736 3367 2743 3473
rect 2776 3447 2783 3483
rect 2756 3303 2763 3413
rect 2736 3296 2763 3303
rect 2736 3107 2743 3296
rect 2816 3266 2823 3473
rect 2796 3260 2803 3263
rect 2793 3247 2807 3260
rect 2836 3187 2843 3393
rect 2856 3308 2863 3493
rect 2876 3107 2883 3503
rect 2996 3496 3003 3573
rect 3176 3567 3183 3733
rect 2896 3387 2903 3473
rect 3136 3407 3143 3533
rect 3196 3427 3203 3813
rect 3216 3547 3223 3573
rect 3236 3500 3243 3503
rect 3233 3487 3247 3500
rect 3216 3387 3223 3433
rect 2436 2327 2443 2353
rect 2416 2268 2423 2293
rect 2476 2287 2483 2593
rect 2433 2260 2447 2273
rect 2436 2256 2443 2260
rect 2416 2027 2423 2093
rect 2476 2047 2483 2223
rect 2496 2023 2503 2553
rect 2476 2016 2503 2023
rect 2236 1956 2243 1960
rect 2216 1827 2223 1923
rect 2076 1700 2083 1703
rect 2073 1687 2087 1700
rect 1987 1606 2000 1607
rect 1987 1593 1993 1606
rect 1956 1507 1963 1553
rect 1953 1448 1967 1453
rect 1996 1436 2003 1553
rect 2016 1483 2023 1593
rect 2036 1547 2043 1593
rect 2016 1476 2033 1483
rect 2036 1447 2043 1473
rect 1936 1307 1943 1393
rect 1836 1107 1843 1132
rect 1836 1027 1843 1093
rect 1856 1067 1863 1253
rect 1956 1227 1963 1373
rect 1976 1367 1983 1403
rect 1976 1356 1993 1367
rect 1980 1353 1993 1356
rect 1876 1123 1883 1153
rect 1896 1147 1903 1183
rect 1933 1147 1947 1151
rect 1976 1147 1983 1333
rect 1996 1227 2003 1313
rect 2016 1247 2023 1333
rect 2036 1267 2043 1393
rect 2056 1367 2063 1533
rect 2076 1403 2083 1613
rect 2116 1547 2123 1736
rect 2316 1736 2323 1954
rect 2336 1927 2343 1973
rect 2373 1960 2387 1973
rect 2376 1956 2383 1960
rect 2476 1927 2483 2016
rect 2516 2003 2523 2833
rect 2536 2788 2543 2933
rect 2556 2847 2563 2952
rect 2536 2607 2543 2653
rect 2536 2476 2543 2593
rect 2576 2587 2583 2743
rect 2616 2727 2623 2994
rect 2593 2480 2607 2493
rect 2596 2476 2603 2480
rect 2576 2440 2583 2443
rect 2573 2427 2587 2440
rect 2616 2403 2623 2713
rect 2636 2446 2643 2933
rect 2676 2927 2683 2963
rect 2676 2776 2683 2913
rect 2716 2807 2723 2953
rect 2736 2707 2743 3013
rect 2756 3007 2763 3033
rect 2776 3027 2783 3093
rect 2773 3000 2787 3013
rect 2813 3000 2827 3013
rect 2896 3008 2903 3263
rect 2956 3207 2963 3373
rect 2996 3107 3003 3373
rect 2776 2996 2783 3000
rect 2816 2996 2823 3000
rect 2793 2947 2807 2952
rect 2676 2483 2683 2693
rect 2656 2476 2683 2483
rect 2616 2396 2643 2403
rect 2496 1996 2523 2003
rect 2396 1787 2403 1923
rect 2176 1700 2183 1703
rect 2107 1536 2123 1547
rect 2107 1533 2120 1536
rect 2096 1427 2103 1453
rect 2116 1436 2123 1493
rect 2136 1463 2143 1693
rect 2173 1687 2187 1700
rect 2216 1687 2223 1703
rect 2216 1623 2223 1673
rect 2196 1616 2223 1623
rect 2156 1507 2163 1553
rect 2160 1483 2173 1487
rect 2156 1480 2173 1483
rect 2153 1473 2173 1480
rect 2153 1467 2167 1473
rect 2136 1456 2153 1463
rect 2076 1396 2103 1403
rect 2076 1227 2083 1373
rect 2016 1127 2023 1172
rect 1876 1116 1903 1123
rect 1896 1087 1903 1116
rect 2036 1087 2043 1153
rect 1853 947 1867 953
rect 1756 916 1763 920
rect 1796 916 1823 923
rect 1576 807 1583 883
rect 1816 883 1823 916
rect 1796 876 1823 883
rect 1556 796 1573 803
rect 1556 743 1563 796
rect 1596 787 1603 853
rect 1587 756 1613 763
rect 1636 743 1643 793
rect 1556 736 1643 743
rect 1476 607 1483 663
rect 1536 567 1543 713
rect 1376 456 1403 463
rect 1076 366 1083 392
rect 1213 383 1227 393
rect 1213 380 1243 383
rect 1216 376 1243 380
rect 956 327 963 363
rect 1116 307 1123 363
rect 1207 353 1213 367
rect 1236 347 1243 376
rect 1376 366 1383 456
rect 1296 360 1303 363
rect 676 107 683 133
rect 696 67 703 143
rect 816 107 823 233
rect 856 188 863 253
rect 916 176 963 183
rect 836 67 843 133
rect 916 87 923 176
rect 976 140 983 143
rect 973 127 987 140
rect 1056 127 1063 193
rect 1116 188 1123 213
rect 1136 207 1143 233
rect 1160 183 1173 187
rect 1156 176 1173 183
rect 1160 173 1173 176
rect 1196 147 1203 313
rect 1256 227 1263 353
rect 1293 347 1307 360
rect 1316 176 1323 273
rect 1336 207 1343 352
rect 1396 247 1403 433
rect 1416 407 1423 493
rect 1456 396 1463 433
rect 1616 407 1623 663
rect 1476 327 1483 363
rect 1456 247 1463 273
rect 1476 267 1483 313
rect 1536 187 1543 394
rect 1636 367 1643 593
rect 1656 447 1663 652
rect 1696 647 1703 753
rect 1736 703 1743 793
rect 1756 727 1763 773
rect 1776 767 1783 813
rect 1736 696 1763 703
rect 1796 696 1803 876
rect 1816 727 1823 833
rect 1836 707 1843 933
rect 1853 923 1867 933
rect 1853 920 1883 923
rect 1856 916 1883 920
rect 2056 916 2063 953
rect 2096 948 2103 1396
rect 2196 1387 2203 1616
rect 2236 1607 2243 1693
rect 2256 1567 2263 1734
rect 2276 1687 2283 1734
rect 2416 1727 2423 1893
rect 2436 1707 2443 1853
rect 2456 1747 2463 1873
rect 2476 1736 2483 1892
rect 2496 1867 2503 1996
rect 2536 1987 2543 2273
rect 2556 2256 2563 2313
rect 2596 2067 2603 2223
rect 2556 1956 2563 1993
rect 2516 1807 2523 1873
rect 2336 1700 2343 1703
rect 2333 1687 2347 1700
rect 2376 1696 2403 1703
rect 2216 1327 2223 1513
rect 2256 1448 2263 1513
rect 2296 1436 2303 1593
rect 2216 1227 2223 1253
rect 2236 1247 2243 1293
rect 2216 1226 2240 1227
rect 2216 1216 2233 1226
rect 2220 1213 2233 1216
rect 2116 1127 2123 1213
rect 2256 1187 2263 1373
rect 2136 1107 2143 1172
rect 2156 1087 2163 1183
rect 2196 1067 2203 1183
rect 1996 883 2003 913
rect 2136 887 2143 953
rect 2156 887 2163 1033
rect 2236 947 2243 1033
rect 2256 927 2263 1073
rect 2276 1047 2283 1353
rect 2296 1267 2303 1313
rect 2316 1243 2323 1393
rect 2336 1367 2343 1633
rect 2356 1447 2363 1473
rect 2376 1463 2383 1573
rect 2396 1567 2403 1696
rect 2516 1700 2523 1703
rect 2513 1687 2527 1700
rect 2396 1487 2403 1553
rect 2416 1507 2423 1553
rect 2376 1456 2403 1463
rect 2396 1436 2403 1456
rect 2436 1436 2443 1513
rect 2476 1407 2483 1673
rect 2536 1667 2543 1912
rect 2356 1347 2363 1393
rect 2376 1327 2383 1403
rect 2416 1327 2423 1403
rect 2496 1387 2503 1633
rect 2536 1547 2543 1593
rect 2536 1436 2543 1533
rect 2556 1467 2563 1893
rect 2596 1787 2603 1954
rect 2616 1907 2623 2373
rect 2636 2107 2643 2396
rect 2656 2327 2663 2476
rect 2756 2296 2763 2893
rect 2796 2776 2803 2833
rect 2836 2827 2843 2963
rect 2896 2743 2903 2994
rect 2916 2966 2923 3013
rect 2933 3007 2947 3013
rect 2813 2727 2827 2732
rect 2856 2707 2863 2743
rect 2876 2736 2903 2743
rect 2876 2607 2883 2736
rect 2836 2537 2873 2544
rect 2796 2387 2803 2533
rect 2836 2488 2843 2537
rect 2876 2476 2883 2512
rect 2896 2487 2903 2693
rect 2916 2527 2923 2853
rect 2936 2788 2943 2953
rect 2956 2887 2963 2952
rect 3016 2907 3023 3333
rect 3236 3327 3243 3353
rect 3256 3347 3263 3653
rect 3276 3547 3283 3593
rect 3296 3536 3303 3673
rect 3436 3667 3443 4013
rect 3456 3827 3463 4273
rect 3476 4167 3483 4303
rect 3513 4283 3527 4293
rect 3496 4280 3527 4283
rect 3496 4276 3523 4280
rect 3496 4067 3503 4276
rect 3576 4247 3583 4393
rect 3596 4316 3603 4493
rect 3756 4427 3763 4813
rect 3776 4447 3783 4513
rect 3796 4507 3803 4733
rect 3816 4556 3823 4593
rect 3856 4487 3863 4836
rect 3876 4707 3883 5063
rect 3876 4526 3883 4672
rect 3896 4607 3903 5053
rect 3956 4923 3963 5373
rect 3976 5267 3983 5353
rect 3996 5167 4003 5513
rect 4076 5507 4083 5593
rect 4107 5563 4120 5567
rect 4107 5556 4123 5563
rect 4156 5560 4163 5563
rect 4107 5553 4120 5556
rect 4153 5547 4167 5560
rect 4096 5388 4103 5413
rect 4116 5376 4163 5383
rect 4196 5376 4203 5473
rect 4016 5187 4023 5343
rect 3976 4987 3983 5113
rect 3996 5087 4003 5153
rect 4036 5076 4043 5113
rect 4053 5107 4067 5113
rect 3996 5036 4023 5043
rect 3996 4967 4003 5036
rect 4053 5023 4067 5033
rect 4036 5020 4067 5023
rect 4036 5016 4063 5020
rect 3956 4916 3983 4923
rect 3953 4860 3967 4873
rect 3976 4868 3983 4916
rect 3956 4856 3963 4860
rect 3916 4767 3923 4823
rect 3916 4647 3923 4753
rect 3976 4727 3983 4854
rect 4016 4667 4023 5013
rect 4007 4653 4023 4667
rect 4016 4567 4023 4653
rect 4036 4587 4043 5016
rect 4076 4967 4083 5293
rect 4096 5087 4103 5374
rect 4116 5127 4123 5376
rect 4176 5340 4183 5343
rect 4173 5327 4187 5340
rect 4153 5080 4167 5093
rect 4156 5076 4163 5080
rect 4093 5027 4107 5033
rect 4116 4887 4123 4933
rect 4136 4848 4143 4993
rect 4176 4983 4183 5043
rect 4156 4980 4183 4983
rect 4153 4976 4183 4980
rect 4153 4967 4167 4976
rect 4196 4963 4203 5033
rect 4176 4956 4203 4963
rect 4096 4707 4103 4823
rect 4176 4647 4183 4956
rect 4196 4836 4203 4933
rect 4216 4907 4223 5343
rect 4256 5307 4263 5593
rect 4353 5580 4367 5593
rect 4356 5576 4363 5580
rect 4496 5487 4503 5733
rect 4536 5487 4543 5583
rect 4396 5447 4403 5473
rect 4280 5383 4293 5387
rect 4276 5373 4293 5383
rect 4336 5376 4343 5413
rect 4373 5387 4387 5393
rect 4276 5107 4283 5373
rect 4396 5346 4403 5433
rect 4416 5387 4423 5413
rect 4496 5376 4503 5413
rect 4316 5340 4323 5343
rect 4313 5327 4327 5340
rect 4416 5267 4423 5333
rect 4436 5267 4443 5343
rect 4476 5307 4483 5343
rect 4296 5088 4303 5173
rect 4247 5083 4260 5087
rect 4247 5076 4263 5083
rect 4247 5073 4260 5076
rect 4236 5007 4243 5033
rect 4336 4947 4343 5133
rect 4356 5047 4363 5093
rect 4416 5076 4423 5173
rect 4453 5080 4467 5093
rect 4456 5076 4463 5080
rect 4396 4947 4403 5043
rect 4416 4967 4423 5013
rect 4436 5007 4443 5043
rect 4236 4747 4243 4933
rect 4476 4847 4483 4993
rect 4380 4843 4393 4847
rect 4376 4836 4393 4843
rect 4380 4833 4393 4836
rect 4496 4836 4503 5193
rect 4536 5087 4543 5313
rect 4556 5107 4563 5793
rect 4576 5627 4583 5833
rect 4596 5727 4603 5843
rect 4636 5807 4643 6113
rect 4896 6103 4903 6296
rect 5076 6267 5083 6303
rect 5036 6187 5043 6253
rect 4656 5908 4663 6092
rect 4716 6080 4723 6083
rect 4713 6067 4727 6080
rect 4636 5687 4643 5753
rect 4633 5627 4647 5633
rect 4656 5608 4663 5894
rect 4676 5667 4683 5993
rect 4736 5896 4743 5933
rect 4796 5866 4803 6013
rect 4856 6007 4863 6103
rect 4847 5996 4863 6007
rect 4876 6096 4903 6103
rect 5036 6096 5043 6152
rect 5056 6107 5063 6133
rect 4847 5993 4860 5996
rect 4856 5896 4863 5973
rect 4876 5927 4883 6096
rect 5136 6103 5143 6253
rect 5696 6207 5703 6303
rect 5836 6296 5863 6303
rect 5676 6196 5693 6203
rect 5196 6136 5243 6143
rect 5136 6096 5163 6103
rect 5136 6003 5143 6073
rect 5116 5996 5143 6003
rect 4896 5896 4903 5953
rect 4716 5807 4723 5863
rect 4956 5863 4963 5893
rect 4976 5866 4983 5953
rect 5076 5896 5083 5933
rect 4816 5856 4843 5863
rect 4796 5627 4803 5693
rect 4587 5583 4600 5587
rect 4587 5573 4603 5583
rect 4596 5523 4603 5573
rect 4616 5547 4623 5573
rect 4596 5516 4623 5523
rect 4616 5376 4623 5516
rect 4656 5327 4663 5594
rect 4676 5343 4683 5613
rect 4713 5600 4727 5613
rect 4716 5596 4723 5600
rect 4736 5388 4743 5413
rect 4676 5336 4703 5343
rect 4756 5327 4763 5473
rect 4576 5076 4583 5153
rect 3976 4527 3983 4554
rect 4056 4556 4063 4633
rect 4093 4560 4107 4573
rect 4096 4556 4103 4560
rect 3616 4327 3623 4353
rect 3636 4287 3643 4413
rect 3916 4327 3923 4473
rect 3616 4147 3623 4273
rect 3776 4247 3783 4323
rect 3876 4316 3903 4323
rect 3796 4267 3803 4313
rect 3876 4167 3883 4316
rect 3976 4287 3983 4492
rect 3996 4487 4003 4553
rect 4016 4463 4023 4513
rect 4036 4503 4043 4512
rect 4036 4496 4063 4503
rect 3996 4456 4023 4463
rect 3996 4327 4003 4456
rect 4016 4307 4023 4413
rect 4056 4336 4063 4496
rect 4076 4487 4083 4523
rect 4096 4447 4103 4473
rect 4136 4447 4143 4543
rect 4176 4427 4183 4573
rect 4196 4507 4203 4543
rect 4236 4387 4243 4693
rect 4376 4647 4383 4813
rect 4373 4540 4387 4553
rect 4376 4536 4383 4540
rect 4476 4507 4483 4733
rect 4536 4707 4543 4803
rect 4567 4753 4573 4767
rect 4596 4747 4603 5093
rect 4616 4967 4623 5213
rect 4656 5007 4663 5273
rect 4696 5147 4703 5313
rect 4796 5207 4803 5613
rect 4816 5387 4823 5856
rect 4876 5807 4883 5863
rect 4916 5856 4963 5863
rect 4847 5713 4853 5727
rect 4896 5687 4903 5833
rect 5016 5807 5023 5863
rect 5056 5787 5063 5863
rect 5116 5747 5123 5996
rect 5176 5896 5183 5933
rect 5236 5907 5243 6136
rect 5296 6116 5303 6153
rect 5336 6063 5343 6083
rect 5336 6056 5363 6063
rect 5256 5867 5263 5933
rect 5336 5896 5343 6033
rect 5356 6007 5363 6056
rect 5376 6043 5383 6113
rect 5396 6087 5403 6114
rect 5427 6123 5440 6127
rect 5427 6116 5443 6123
rect 5427 6113 5440 6116
rect 5376 6036 5403 6043
rect 4836 5467 4843 5653
rect 4856 5596 4863 5673
rect 5016 5596 5023 5693
rect 4836 5167 4843 5343
rect 4856 5187 4863 5513
rect 4896 5407 4903 5563
rect 4916 5507 4923 5573
rect 4936 5483 4943 5594
rect 5056 5547 5063 5733
rect 4916 5476 4943 5483
rect 4696 5076 4703 5133
rect 4776 5027 4783 5113
rect 4876 5087 4883 5374
rect 4916 5287 4923 5476
rect 4976 5343 4983 5453
rect 4956 5336 4983 5343
rect 5016 5327 5023 5533
rect 5076 5527 5083 5673
rect 5156 5596 5163 5693
rect 5196 5647 5203 5863
rect 5236 5827 5243 5853
rect 5236 5687 5243 5713
rect 5136 5527 5143 5563
rect 5136 5447 5143 5513
rect 5216 5507 5223 5583
rect 5256 5567 5263 5653
rect 5276 5467 5283 5583
rect 5316 5487 5323 5793
rect 5376 5767 5383 5894
rect 5396 5787 5403 6036
rect 5496 6007 5503 6083
rect 5476 5896 5483 5993
rect 5516 5896 5523 5933
rect 5533 5907 5547 5913
rect 5416 5807 5423 5853
rect 5496 5727 5503 5863
rect 5456 5576 5463 5673
rect 5556 5667 5563 6114
rect 5576 5967 5583 6073
rect 5676 6047 5683 6196
rect 5736 6116 5743 6193
rect 5773 6120 5787 6133
rect 5776 6116 5783 6120
rect 5756 6007 5763 6083
rect 5607 5996 5633 6003
rect 5816 5947 5823 6133
rect 5836 6127 5843 6296
rect 5867 6143 5880 6147
rect 5867 6133 5883 6143
rect 5876 6116 5883 6133
rect 5936 6086 5943 6133
rect 5996 6116 6003 6153
rect 6036 6128 6043 6193
rect 5976 6027 5983 6083
rect 6016 6047 6023 6083
rect 5627 5914 5633 5927
rect 5620 5913 5640 5914
rect 5576 5767 5583 5893
rect 5616 5628 5623 5813
rect 5696 5807 5703 5894
rect 5856 5867 5863 6013
rect 5913 5908 5927 5913
rect 5956 5896 5963 5933
rect 5053 5380 5067 5393
rect 5056 5376 5063 5380
rect 5116 5356 5123 5393
rect 5176 5356 5183 5453
rect 5556 5367 5563 5613
rect 5676 5566 5683 5673
rect 5736 5623 5743 5863
rect 5796 5827 5803 5863
rect 5936 5827 5943 5863
rect 5716 5616 5743 5623
rect 5716 5596 5723 5616
rect 5756 5596 5763 5653
rect 5816 5566 5823 5593
rect 5836 5566 5843 5713
rect 5896 5596 5903 5673
rect 5976 5627 5983 5863
rect 6016 5608 6023 5913
rect 6036 5667 6043 6033
rect 6076 5896 6083 6113
rect 6096 5927 6103 6133
rect 6156 6116 6163 6153
rect 6253 6120 6267 6133
rect 6256 6116 6263 6120
rect 6136 6047 6143 6083
rect 6107 5916 6123 5923
rect 6116 5896 6123 5916
rect 6033 5600 6047 5613
rect 6036 5596 6043 5600
rect 6096 5587 6103 5713
rect 6156 5687 6163 5893
rect 6156 5623 6163 5673
rect 6136 5616 6163 5623
rect 5876 5527 5883 5563
rect 5916 5487 5923 5563
rect 6136 5563 6143 5616
rect 6136 5556 6163 5563
rect 4936 5076 4943 5193
rect 4956 5187 4963 5213
rect 5056 5076 5063 5313
rect 5076 5167 5083 5343
rect 4996 5046 5003 5073
rect 5116 5047 5123 5253
rect 5356 5227 5363 5363
rect 5456 5356 5483 5363
rect 5456 5287 5463 5356
rect 5616 5356 5643 5363
rect 5220 5123 5233 5127
rect 5216 5120 5233 5123
rect 5213 5113 5233 5120
rect 5213 5108 5227 5113
rect 5293 5107 5307 5113
rect 4816 5007 4823 5043
rect 4656 4883 4663 4993
rect 4656 4876 4683 4883
rect 4676 4856 4683 4876
rect 4716 4856 4723 4933
rect 4893 4907 4907 4913
rect 4756 4826 4763 4893
rect 4853 4868 4867 4873
rect 4656 4820 4663 4823
rect 4653 4807 4667 4820
rect 4627 4753 4633 4767
rect 4536 4588 4543 4693
rect 4836 4687 4843 4823
rect 4916 4823 4923 4913
rect 4896 4816 4923 4823
rect 4093 4340 4107 4353
rect 4096 4336 4103 4340
rect 3996 4296 4013 4303
rect 3476 4020 3483 4023
rect 3473 4007 3487 4020
rect 3476 3803 3483 3993
rect 3496 3927 3503 4013
rect 3516 4007 3523 4073
rect 3656 4016 3663 4133
rect 3476 3796 3503 3803
rect 3536 3796 3563 3803
rect 3356 3506 3363 3613
rect 3296 3327 3303 3453
rect 3076 3227 3083 3263
rect 3076 3003 3083 3173
rect 3096 3067 3103 3153
rect 3116 3023 3123 3213
rect 3136 3067 3143 3133
rect 3116 3016 3143 3023
rect 3056 2996 3083 3003
rect 3136 2996 3143 3016
rect 3056 2923 3063 2996
rect 3156 2987 3163 3233
rect 3056 2916 3083 2923
rect 3056 2747 3063 2893
rect 3076 2867 3083 2916
rect 3096 2827 3103 2952
rect 3136 2907 3143 2933
rect 3136 2776 3143 2813
rect 3156 2807 3163 2952
rect 3176 2947 3183 3093
rect 3196 2987 3203 3263
rect 3216 3007 3223 3313
rect 3236 3127 3243 3313
rect 3316 3296 3323 3393
rect 3336 3303 3343 3503
rect 3456 3496 3463 3753
rect 3496 3687 3503 3796
rect 3556 3747 3563 3796
rect 3576 3787 3583 3813
rect 3596 3727 3603 3853
rect 3636 3816 3643 3913
rect 3736 3867 3743 3913
rect 3656 3780 3663 3783
rect 3653 3767 3667 3780
rect 3496 3627 3503 3673
rect 3596 3587 3603 3633
rect 3356 3327 3363 3413
rect 3336 3296 3363 3303
rect 3256 3067 3263 3253
rect 3296 3227 3303 3263
rect 3356 3127 3363 3296
rect 3436 3296 3443 3373
rect 3596 3367 3603 3552
rect 3656 3503 3663 3673
rect 3676 3547 3683 3573
rect 3636 3496 3663 3503
rect 3616 3467 3623 3492
rect 3376 3227 3383 3293
rect 3416 3260 3423 3263
rect 3413 3247 3427 3260
rect 3307 3113 3313 3127
rect 3256 3023 3263 3053
rect 3236 3016 3263 3023
rect 3236 2996 3243 3016
rect 3276 2996 3283 3113
rect 3396 3047 3403 3093
rect 3416 3087 3423 3233
rect 3436 3107 3443 3173
rect 3456 3167 3463 3252
rect 3476 3143 3483 3233
rect 3496 3207 3503 3293
rect 3516 3247 3523 3353
rect 3573 3300 3587 3313
rect 3576 3296 3583 3300
rect 3556 3260 3563 3263
rect 3553 3247 3567 3260
rect 3596 3207 3603 3263
rect 3636 3227 3643 3433
rect 3716 3427 3723 3653
rect 3736 3507 3743 3832
rect 3756 3786 3763 4113
rect 3776 3847 3783 3873
rect 3796 3847 3803 3993
rect 3856 3867 3863 4133
rect 3876 4007 3883 4073
rect 3896 4027 3903 4153
rect 3916 4147 3923 4213
rect 3936 4068 3943 4272
rect 3956 4036 3963 4193
rect 3976 4087 3983 4233
rect 3996 4127 4003 4296
rect 3993 4040 4007 4053
rect 4016 4047 4023 4272
rect 4036 4227 4043 4293
rect 4076 4267 4083 4292
rect 4156 4286 4163 4373
rect 4196 4267 4203 4303
rect 3996 4036 4003 4040
rect 3916 3947 3923 3993
rect 3936 3967 3943 4003
rect 3936 3828 3943 3853
rect 3736 3447 3743 3493
rect 3756 3423 3763 3673
rect 3796 3587 3803 3783
rect 3876 3767 3883 3793
rect 3796 3516 3803 3573
rect 3836 3516 3843 3553
rect 3876 3467 3883 3514
rect 3736 3416 3763 3423
rect 3696 3296 3703 3333
rect 3736 3307 3743 3416
rect 3607 3196 3623 3203
rect 3456 3136 3483 3143
rect 3436 3003 3443 3053
rect 3416 2996 3443 3003
rect 3176 2776 3183 2912
rect 3256 2907 3263 2963
rect 3236 2896 3253 2903
rect 3196 2787 3203 2873
rect 2956 2740 2963 2743
rect 2807 2256 2823 2263
rect 2816 2226 2823 2256
rect 2676 2216 2703 2223
rect 2676 1987 2683 2216
rect 2696 2007 2703 2153
rect 2696 1956 2703 1993
rect 2636 1787 2643 1833
rect 2596 1647 2603 1773
rect 2636 1736 2643 1773
rect 2616 1547 2623 1703
rect 2676 1700 2683 1703
rect 2673 1687 2687 1700
rect 2687 1676 2703 1683
rect 2573 1440 2587 1453
rect 2616 1447 2623 1512
rect 2576 1436 2583 1440
rect 2296 1240 2323 1243
rect 2293 1236 2323 1240
rect 2293 1227 2307 1236
rect 2336 1216 2343 1253
rect 2393 1247 2407 1253
rect 2416 1207 2423 1292
rect 1976 876 2003 883
rect 1896 787 1903 813
rect 1936 787 1943 843
rect 1927 760 1963 763
rect 1927 756 1967 760
rect 1953 747 1967 756
rect 1936 708 1943 733
rect 1976 696 1983 753
rect 1993 707 2007 713
rect 1716 627 1723 693
rect 1787 635 1813 642
rect 1856 607 1863 673
rect 1876 567 1883 693
rect 1956 660 1963 663
rect 1953 647 1967 660
rect 1993 647 2007 652
rect 1693 400 1707 413
rect 1696 396 1703 400
rect 1596 360 1603 363
rect 1593 347 1607 360
rect 1656 327 1663 393
rect 1716 267 1723 363
rect 1556 207 1563 233
rect 1096 47 1103 132
rect 1216 107 1223 174
rect 1353 167 1367 174
rect 1576 176 1583 213
rect 1233 127 1247 133
rect 1256 67 1263 143
rect 1356 47 1363 113
rect 1376 67 1383 133
rect 1396 47 1403 132
rect 1416 43 1423 113
rect 1436 107 1443 143
rect 1476 87 1483 113
rect 1496 83 1503 173
rect 1516 127 1523 173
rect 1656 147 1663 213
rect 1713 180 1727 193
rect 1733 187 1747 193
rect 1716 176 1723 180
rect 1596 140 1603 143
rect 1593 127 1607 140
rect 1593 107 1607 113
rect 1496 76 1523 83
rect 1467 56 1493 63
rect 1516 47 1523 76
rect 1587 76 1613 83
rect 1567 56 1633 63
rect 1756 47 1763 213
rect 1776 147 1783 353
rect 1796 187 1803 473
rect 2016 427 2023 773
rect 2036 627 2043 873
rect 2076 787 2083 883
rect 2187 883 2200 887
rect 2187 876 2203 883
rect 2236 880 2243 883
rect 2187 873 2200 876
rect 2233 867 2247 880
rect 2116 727 2123 773
rect 2136 767 2143 852
rect 2136 696 2143 753
rect 2176 707 2183 833
rect 1893 408 1907 413
rect 1933 407 1947 413
rect 1816 327 1823 394
rect 1836 267 1843 353
rect 1876 343 1883 363
rect 1876 340 1903 343
rect 1873 336 1903 340
rect 1873 327 1887 336
rect 1896 307 1903 336
rect 1916 327 1923 363
rect 1836 176 1843 213
rect 1876 176 1883 273
rect 1916 167 1923 213
rect 1956 207 1963 413
rect 1993 400 2007 413
rect 2033 400 2047 413
rect 2076 407 2083 663
rect 1996 396 2003 400
rect 2036 396 2043 400
rect 2056 356 2083 363
rect 1976 176 1983 213
rect 2016 176 2023 253
rect 2076 227 2083 356
rect 2096 327 2103 593
rect 2116 567 2123 663
rect 2156 627 2163 652
rect 2196 627 2203 793
rect 2236 767 2243 832
rect 2276 807 2283 993
rect 2296 867 2303 1173
rect 2316 1127 2323 1183
rect 2436 1186 2443 1253
rect 2456 1227 2463 1253
rect 2496 1216 2503 1313
rect 2556 1307 2563 1403
rect 2540 1223 2553 1227
rect 2536 1216 2553 1223
rect 2540 1213 2553 1216
rect 2393 1167 2407 1173
rect 2316 1047 2323 1113
rect 2416 1007 2423 1073
rect 2396 916 2403 993
rect 2336 880 2343 883
rect 2333 867 2347 880
rect 2256 708 2263 733
rect 2227 663 2240 667
rect 2296 666 2303 813
rect 2316 807 2323 833
rect 2376 807 2383 883
rect 2436 867 2443 914
rect 2456 847 2463 953
rect 2476 927 2483 1133
rect 2496 928 2503 1153
rect 2556 928 2563 1173
rect 2536 916 2553 923
rect 2473 867 2487 873
rect 2376 696 2383 753
rect 2416 727 2423 773
rect 2227 656 2243 663
rect 2227 653 2240 656
rect 2236 587 2243 613
rect 2116 347 2123 413
rect 2136 407 2143 513
rect 2213 447 2227 453
rect 2213 440 2233 447
rect 2216 436 2233 440
rect 2220 433 2233 436
rect 2173 408 2187 413
rect 2213 400 2227 413
rect 2216 396 2223 400
rect 2256 367 2263 613
rect 2396 587 2403 663
rect 2276 408 2283 453
rect 2316 396 2323 453
rect 2376 423 2383 453
rect 2436 423 2443 793
rect 2496 696 2503 853
rect 2516 723 2523 883
rect 2576 827 2583 1353
rect 2636 1287 2643 1453
rect 2656 1367 2663 1653
rect 2696 1547 2703 1676
rect 2716 1667 2723 1733
rect 2736 1687 2743 2173
rect 2756 1847 2763 2053
rect 2796 1956 2803 2073
rect 2836 2027 2843 2373
rect 2896 2256 2903 2433
rect 2916 2287 2923 2492
rect 2936 2447 2943 2733
rect 2953 2727 2967 2740
rect 2996 2707 3003 2743
rect 2956 2483 2963 2533
rect 2956 2476 2983 2483
rect 3056 2487 3063 2712
rect 3076 2667 3083 2773
rect 3116 2707 3123 2743
rect 3156 2740 3163 2743
rect 3153 2727 3167 2740
rect 3196 2707 3203 2733
rect 3140 2683 3153 2687
rect 3136 2680 3153 2683
rect 3133 2673 3153 2680
rect 3133 2667 3147 2673
rect 2996 2440 3003 2443
rect 2993 2427 3007 2440
rect 2956 2267 2963 2333
rect 2876 2167 2883 2223
rect 2956 2187 2963 2213
rect 2976 2167 2983 2313
rect 3016 2283 3023 2313
rect 3036 2307 3043 2443
rect 3076 2347 3083 2573
rect 3136 2563 3143 2593
rect 3216 2587 3223 2813
rect 3236 2787 3243 2896
rect 3273 2863 3287 2873
rect 3256 2860 3287 2863
rect 3256 2856 3283 2860
rect 3256 2787 3263 2856
rect 3316 2847 3323 2973
rect 3456 2963 3463 3136
rect 3516 3027 3523 3093
rect 3536 2996 3543 3093
rect 3576 3007 3583 3053
rect 3356 2887 3363 2963
rect 3396 2887 3403 2963
rect 3436 2956 3463 2963
rect 3276 2776 3283 2833
rect 3316 2776 3323 2812
rect 3376 2787 3383 2833
rect 3233 2746 3247 2752
rect 3136 2556 3193 2563
rect 3096 2427 3103 2493
rect 3136 2488 3143 2533
rect 3176 2476 3183 2533
rect 3216 2476 3223 2513
rect 3256 2447 3263 2693
rect 3276 2447 3283 2613
rect 3356 2507 3363 2553
rect 3376 2527 3383 2733
rect 3376 2487 3383 2513
rect 3396 2507 3403 2873
rect 3356 2476 3373 2483
rect 3416 2483 3423 2813
rect 3436 2787 3443 2956
rect 3476 2927 3483 2953
rect 3456 2776 3463 2893
rect 3556 2847 3563 2963
rect 3596 2887 3603 3093
rect 3616 2927 3623 3196
rect 3676 3087 3683 3263
rect 3716 3227 3723 3263
rect 3736 3167 3743 3253
rect 3653 3000 3667 3013
rect 3656 2996 3663 3000
rect 3696 2996 3703 3113
rect 3496 2788 3503 2813
rect 3553 2787 3567 2793
rect 3436 2667 3443 2733
rect 3476 2727 3483 2743
rect 3476 2716 3493 2727
rect 3480 2713 3493 2716
rect 3396 2476 3423 2483
rect 3456 2503 3463 2693
rect 3456 2496 3483 2503
rect 3433 2480 3447 2493
rect 3436 2476 3443 2480
rect 3476 2476 3483 2496
rect 3076 2336 3093 2347
rect 3080 2333 3093 2336
rect 3016 2276 3043 2283
rect 2996 2247 3003 2273
rect 3036 2256 3043 2276
rect 3096 2267 3103 2293
rect 3116 2283 3123 2433
rect 3156 2407 3163 2443
rect 3116 2276 3133 2283
rect 2993 2207 3007 2212
rect 2993 2167 3007 2172
rect 2876 2067 2883 2113
rect 2836 1956 2843 1992
rect 2776 1827 2783 1873
rect 2816 1743 2823 1923
rect 2876 1807 2883 2053
rect 2896 1867 2903 2013
rect 2936 1956 2943 2153
rect 2956 2067 2963 2152
rect 3016 2107 3023 2223
rect 3076 2147 3083 2223
rect 2976 2047 2983 2073
rect 3016 2063 3023 2093
rect 2996 2056 3023 2063
rect 2976 1956 2983 2033
rect 2996 2007 3003 2056
rect 2876 1748 2883 1793
rect 2956 1787 2963 1912
rect 2916 1748 2923 1773
rect 2816 1736 2843 1743
rect 2776 1667 2783 1703
rect 2616 1228 2623 1253
rect 2640 1186 2653 1187
rect 2647 1173 2653 1186
rect 2676 1167 2683 1473
rect 2696 1436 2703 1533
rect 2756 1436 2783 1443
rect 2696 1187 2703 1373
rect 2736 1367 2743 1392
rect 2716 1227 2723 1293
rect 2776 1247 2783 1436
rect 2796 1407 2803 1673
rect 2816 1627 2823 1693
rect 2836 1443 2843 1736
rect 2856 1687 2863 1713
rect 2876 1523 2883 1734
rect 2976 1706 2983 1853
rect 2896 1547 2903 1703
rect 2956 1696 2973 1703
rect 2876 1516 2903 1523
rect 2856 1487 2863 1513
rect 2816 1436 2843 1443
rect 2853 1440 2867 1452
rect 2896 1448 2903 1516
rect 2856 1436 2863 1440
rect 2796 1227 2803 1353
rect 2596 747 2603 1133
rect 2676 916 2703 923
rect 2516 716 2543 723
rect 2536 703 2543 716
rect 2536 696 2563 703
rect 2476 627 2483 652
rect 2516 607 2523 663
rect 2556 507 2563 696
rect 2616 696 2623 853
rect 2696 707 2703 916
rect 2576 607 2583 694
rect 2716 687 2723 1153
rect 2736 1027 2743 1183
rect 2776 1147 2783 1183
rect 2796 1107 2803 1173
rect 2816 1087 2823 1436
rect 2876 1400 2883 1403
rect 2836 1127 2843 1393
rect 2873 1387 2887 1400
rect 2853 1227 2867 1233
rect 2896 1216 2903 1293
rect 2936 1267 2943 1473
rect 2956 1243 2963 1533
rect 2976 1527 2983 1573
rect 2976 1436 2983 1513
rect 2996 1487 3003 1913
rect 3016 1667 3023 2033
rect 3096 1956 3103 2253
rect 3116 2187 3123 2252
rect 3136 1967 3143 2273
rect 3156 2267 3163 2393
rect 3196 2347 3203 2443
rect 3213 2407 3227 2413
rect 3173 2260 3187 2273
rect 3176 2256 3183 2260
rect 3216 2256 3223 2293
rect 3253 2267 3267 2273
rect 3196 2047 3203 2223
rect 3276 2187 3283 2293
rect 3296 2267 3303 2393
rect 3336 2256 3343 2333
rect 3356 2220 3363 2223
rect 3353 2207 3367 2220
rect 3296 2067 3303 2133
rect 3156 1926 3163 1953
rect 3076 1867 3083 1923
rect 3036 1767 3043 1793
rect 3056 1736 3063 1813
rect 3096 1736 3103 1773
rect 3056 1383 3063 1673
rect 3036 1376 3063 1383
rect 2936 1236 2963 1243
rect 2936 1216 2943 1236
rect 2876 1163 2883 1183
rect 2876 1156 2903 1163
rect 2816 967 2823 1073
rect 2776 916 2783 953
rect 2856 947 2863 1093
rect 2813 920 2827 932
rect 2816 916 2823 920
rect 2856 887 2863 933
rect 2756 807 2763 883
rect 2876 867 2883 1113
rect 2896 1047 2903 1156
rect 2916 987 2923 1183
rect 2976 1047 2983 1133
rect 2996 1107 3003 1373
rect 3036 1227 3043 1376
rect 3076 1307 3083 1703
rect 3136 1467 3143 1853
rect 3216 1847 3223 1912
rect 3256 1907 3263 1993
rect 3296 1968 3303 2053
rect 3316 2027 3323 2153
rect 3316 1987 3323 2013
rect 3376 1956 3383 2073
rect 3396 1963 3403 2476
rect 3416 2267 3423 2433
rect 3496 2256 3503 2393
rect 3516 2263 3523 2693
rect 3536 2687 3543 2774
rect 3633 2780 3647 2793
rect 3656 2787 3663 2913
rect 3716 2867 3723 2963
rect 3756 2907 3763 3393
rect 3776 3207 3783 3313
rect 3796 3263 3803 3333
rect 3836 3296 3843 3433
rect 3896 3267 3903 3713
rect 3936 3687 3943 3753
rect 3956 3747 3963 3783
rect 3936 3516 3943 3673
rect 3976 3567 3983 3773
rect 3996 3747 4003 3913
rect 3996 3523 4003 3673
rect 4016 3627 4023 3953
rect 4036 3707 4043 4093
rect 4056 3987 4063 4233
rect 4076 4047 4083 4213
rect 4113 4040 4127 4053
rect 4156 4047 4163 4213
rect 4216 4087 4223 4273
rect 4236 4187 4243 4303
rect 4276 4247 4283 4433
rect 4296 4227 4303 4353
rect 4356 4336 4363 4413
rect 4336 4247 4343 4303
rect 4116 4036 4123 4040
rect 4176 4003 4183 4053
rect 4233 4040 4247 4053
rect 4276 4048 4283 4193
rect 4236 4036 4243 4040
rect 4336 4007 4343 4034
rect 4076 3963 4083 3993
rect 4056 3956 4083 3963
rect 4056 3816 4063 3956
rect 4096 3927 4103 4003
rect 4136 3983 4143 4003
rect 4156 3996 4183 4003
rect 4156 3983 4163 3996
rect 4136 3976 4163 3983
rect 4096 3747 4103 3783
rect 4116 3667 4123 3973
rect 3987 3516 4003 3523
rect 3936 3407 3943 3453
rect 3956 3447 3963 3483
rect 3796 3256 3823 3263
rect 3876 3227 3883 3263
rect 3776 2966 3783 3073
rect 3796 3047 3803 3133
rect 3816 3008 3823 3213
rect 3856 2996 3863 3033
rect 3896 3007 3903 3153
rect 3916 3067 3923 3373
rect 4016 3367 4023 3613
rect 3956 3296 3963 3353
rect 4033 3307 4047 3313
rect 3896 2996 3913 3007
rect 3900 2993 3913 2996
rect 3876 2927 3883 2952
rect 3636 2776 3643 2780
rect 3676 2747 3683 2833
rect 3576 2740 3583 2743
rect 3556 2483 3563 2733
rect 3573 2727 3587 2740
rect 3696 2723 3703 2813
rect 3756 2776 3763 2872
rect 3727 2743 3740 2747
rect 3727 2736 3743 2743
rect 3776 2740 3783 2743
rect 3727 2733 3740 2736
rect 3773 2727 3787 2740
rect 3696 2716 3723 2723
rect 3536 2476 3563 2483
rect 3596 2476 3603 2613
rect 3656 2587 3663 2613
rect 3676 2567 3683 2712
rect 3636 2476 3643 2533
rect 3536 2287 3543 2476
rect 3696 2446 3703 2533
rect 3616 2367 3623 2443
rect 3636 2343 3643 2373
rect 3607 2336 3643 2343
rect 3516 2256 3543 2263
rect 3436 2220 3443 2223
rect 3476 2220 3483 2223
rect 3416 2007 3423 2213
rect 3433 2207 3447 2220
rect 3473 2207 3487 2220
rect 3476 2107 3483 2153
rect 3396 1956 3423 1963
rect 3476 1956 3483 2093
rect 3516 1956 3523 2073
rect 3536 2007 3543 2256
rect 3636 2256 3643 2313
rect 3656 2307 3663 2443
rect 3716 2347 3723 2716
rect 3816 2663 3823 2893
rect 3836 2787 3843 2913
rect 3876 2776 3883 2833
rect 3916 2807 3923 2953
rect 3856 2707 3863 2743
rect 3887 2725 3900 2727
rect 3887 2713 3893 2725
rect 3880 2683 3893 2687
rect 3876 2673 3893 2683
rect 3816 2656 3843 2663
rect 3736 2587 3743 2653
rect 3796 2487 3803 2573
rect 3816 2443 3823 2633
rect 3796 2436 3823 2443
rect 3656 2267 3663 2293
rect 3316 1920 3323 1923
rect 3313 1907 3327 1920
rect 3396 1827 3403 1913
rect 3193 1740 3207 1753
rect 3236 1748 3243 1773
rect 3196 1736 3203 1740
rect 3176 1587 3183 1703
rect 3156 1467 3163 1553
rect 3096 1267 3103 1453
rect 3176 1448 3183 1533
rect 3127 1443 3140 1447
rect 3127 1436 3143 1443
rect 3127 1433 3140 1436
rect 3196 1443 3203 1613
rect 3216 1527 3223 1703
rect 3296 1687 3303 1813
rect 3380 1703 3393 1707
rect 3196 1436 3223 1443
rect 3216 1406 3223 1436
rect 3296 1436 3303 1652
rect 3316 1627 3323 1693
rect 3336 1547 3343 1703
rect 3376 1696 3393 1703
rect 3380 1693 3393 1696
rect 3336 1487 3343 1533
rect 3116 1327 3123 1393
rect 3156 1367 3163 1403
rect 3056 1216 3063 1253
rect 3136 1227 3143 1253
rect 3016 1147 3023 1213
rect 3036 1127 3043 1173
rect 3076 1067 3083 1183
rect 3116 1180 3123 1183
rect 3113 1167 3127 1180
rect 3096 1007 3103 1053
rect 2893 927 2907 933
rect 2940 923 2953 927
rect 2936 916 2953 923
rect 2940 913 2953 916
rect 2996 916 3013 923
rect 2907 883 2920 887
rect 2996 886 3003 916
rect 3027 923 3040 927
rect 3027 916 3043 923
rect 3073 920 3087 933
rect 3116 927 3123 1113
rect 3136 927 3143 1173
rect 3156 1167 3163 1313
rect 3176 967 3183 1293
rect 3276 1243 3283 1403
rect 3256 1236 3283 1243
rect 3256 1216 3263 1236
rect 3296 1227 3303 1313
rect 3196 1007 3203 1173
rect 3236 1147 3243 1183
rect 3316 1186 3323 1253
rect 3336 1227 3343 1293
rect 3356 1247 3363 1673
rect 3376 1507 3383 1673
rect 3416 1587 3423 1956
rect 3436 1707 3443 1893
rect 3456 1867 3463 1923
rect 3556 1923 3563 2193
rect 3596 2127 3603 2193
rect 3616 2187 3623 2223
rect 3676 2167 3683 2333
rect 3736 2256 3743 2293
rect 3776 2267 3783 2313
rect 3796 2223 3803 2436
rect 3836 2427 3843 2656
rect 3876 2587 3883 2673
rect 3896 2547 3903 2613
rect 3916 2607 3923 2673
rect 3936 2647 3943 3253
rect 4016 3227 4023 3263
rect 4056 3163 4063 3393
rect 4076 3367 4083 3483
rect 4116 3327 4123 3653
rect 4136 3587 4143 3873
rect 4156 3787 4163 3976
rect 4176 3847 4183 3953
rect 4196 3887 4203 3993
rect 4216 3947 4223 4003
rect 4236 3923 4243 3973
rect 4216 3916 4243 3923
rect 4216 3828 4223 3916
rect 4296 3907 4303 4003
rect 4356 3967 4363 4173
rect 4376 4167 4383 4303
rect 4407 4273 4413 4287
rect 4436 4167 4443 4373
rect 4476 4363 4483 4472
rect 4496 4387 4503 4543
rect 4556 4447 4563 4533
rect 4516 4367 4523 4413
rect 4476 4356 4503 4363
rect 4496 4336 4503 4356
rect 4596 4347 4603 4473
rect 4636 4387 4643 4543
rect 4656 4487 4663 4633
rect 4756 4536 4763 4673
rect 4896 4447 4903 4816
rect 4936 4767 4943 4993
rect 4956 4887 4963 5032
rect 4987 4897 5013 4904
rect 5036 4887 5043 5032
rect 5156 4947 5163 5093
rect 5176 5003 5183 5033
rect 5176 4996 5223 5003
rect 4973 4860 4987 4872
rect 4976 4856 4983 4860
rect 4936 4507 4943 4543
rect 4476 4300 4483 4303
rect 4473 4287 4487 4300
rect 4376 4047 4383 4153
rect 4456 4143 4463 4253
rect 4473 4167 4487 4173
rect 4436 4136 4463 4143
rect 4436 4036 4443 4136
rect 4516 4087 4523 4292
rect 4556 4068 4563 4293
rect 4576 4267 4583 4333
rect 4656 4283 4663 4303
rect 4636 4276 4663 4283
rect 4636 4207 4643 4276
rect 4196 3516 4203 3772
rect 4256 3687 4263 3814
rect 4136 3323 4143 3514
rect 4276 3487 4283 3673
rect 4156 3343 4163 3433
rect 4176 3427 4183 3483
rect 4296 3483 4303 3613
rect 4316 3528 4323 3772
rect 4356 3767 4363 3953
rect 4376 3747 4383 3993
rect 4416 3967 4423 4003
rect 4476 3987 4483 4053
rect 4496 3967 4503 4033
rect 4636 4007 4643 4193
rect 4716 4167 4723 4433
rect 4736 4147 4743 4373
rect 4796 4336 4803 4433
rect 4956 4376 4963 4593
rect 5036 4546 5043 4873
rect 5056 4867 5063 4893
rect 5076 4856 5083 4913
rect 5216 4856 5223 4996
rect 5236 4927 5243 5043
rect 5267 5013 5273 5027
rect 5296 5007 5303 5072
rect 5316 5046 5323 5133
rect 5336 5083 5343 5153
rect 5373 5107 5387 5113
rect 5336 5076 5363 5083
rect 5396 5076 5403 5213
rect 5496 5207 5503 5273
rect 5636 5207 5643 5356
rect 5916 5356 5923 5433
rect 5976 5356 5983 5413
rect 6176 5383 6183 5413
rect 6176 5376 6203 5383
rect 5436 5167 5443 5193
rect 5416 5107 5423 5133
rect 5376 5040 5383 5043
rect 5373 5027 5387 5040
rect 5476 5027 5483 5074
rect 5373 5007 5387 5013
rect 5016 4343 5023 4413
rect 4996 4336 5023 4343
rect 4816 4267 4823 4303
rect 4876 4296 4903 4303
rect 4876 4207 4883 4296
rect 4776 4067 4783 4173
rect 4673 4040 4687 4053
rect 4676 4036 4683 4040
rect 4416 3816 4423 3893
rect 4456 3816 4463 3873
rect 4516 3786 4523 3833
rect 4536 3827 4543 4003
rect 4776 4003 4783 4053
rect 4776 3996 4803 4003
rect 4573 3820 4587 3833
rect 4576 3816 4583 3820
rect 4416 3527 4423 3753
rect 4556 3687 4563 3783
rect 4296 3476 4343 3483
rect 4196 3387 4203 3453
rect 4156 3336 4193 3343
rect 4136 3316 4203 3323
rect 4076 3187 4083 3313
rect 4136 3296 4143 3316
rect 4196 3303 4203 3316
rect 4196 3296 4223 3303
rect 4107 3263 4120 3267
rect 4107 3256 4123 3263
rect 4107 3253 4120 3256
rect 4156 3227 4163 3252
rect 4196 3207 4203 3253
rect 4216 3227 4223 3296
rect 4056 3156 4083 3163
rect 3967 3036 3993 3043
rect 3996 2960 4003 2963
rect 3993 2947 4007 2960
rect 3956 2727 3963 2913
rect 4036 2827 4043 2873
rect 4056 2867 4063 3093
rect 4076 2927 4083 3156
rect 4156 3056 4193 3063
rect 4136 2996 4143 3053
rect 4156 3027 4163 3056
rect 4176 3008 4183 3033
rect 4113 2947 4127 2952
rect 3876 2476 3883 2513
rect 3936 2488 3943 2533
rect 3816 2287 3823 2353
rect 3836 2288 3843 2392
rect 3856 2327 3863 2473
rect 3956 2467 3963 2713
rect 3976 2687 3983 2732
rect 3996 2727 4003 2743
rect 3896 2427 3903 2443
rect 3876 2307 3883 2353
rect 3896 2267 3903 2413
rect 3956 2383 3963 2453
rect 3976 2407 3983 2613
rect 3996 2547 4003 2713
rect 4036 2707 4043 2732
rect 4076 2667 4083 2793
rect 4096 2587 4103 2773
rect 4116 2740 4123 2743
rect 4113 2727 4127 2740
rect 4176 2707 4183 2743
rect 4073 2507 4087 2513
rect 4033 2480 4047 2493
rect 4036 2476 4043 2480
rect 4007 2443 4020 2447
rect 4007 2436 4023 2443
rect 4056 2440 4063 2443
rect 4007 2433 4020 2436
rect 4053 2427 4067 2440
rect 4096 2407 4103 2493
rect 4116 2427 4123 2692
rect 4156 2507 4163 2653
rect 4196 2627 4203 2931
rect 4236 2907 4243 3413
rect 4267 3323 4280 3327
rect 4267 3313 4283 3323
rect 4276 3296 4283 3313
rect 4256 3227 4263 3263
rect 4316 3187 4323 3263
rect 4256 2947 4263 3173
rect 4336 3107 4343 3476
rect 4356 3087 4363 3453
rect 4376 3443 4383 3483
rect 4376 3436 4403 3443
rect 4376 3187 4383 3413
rect 4396 3327 4403 3436
rect 4436 3407 4443 3573
rect 4500 3543 4513 3547
rect 4496 3533 4513 3543
rect 4496 3516 4503 3533
rect 4456 3323 4463 3473
rect 4476 3347 4483 3483
rect 4536 3427 4543 3514
rect 4556 3486 4563 3673
rect 4596 3667 4603 3783
rect 4636 3687 4643 3873
rect 4656 3823 4663 3953
rect 4716 3856 4723 3933
rect 4656 3816 4683 3823
rect 4796 3727 4803 3996
rect 4816 3947 4823 3992
rect 4593 3520 4607 3533
rect 4636 3528 4643 3652
rect 4596 3516 4603 3520
rect 4696 3483 4703 3653
rect 4656 3476 4703 3483
rect 4456 3316 4483 3323
rect 4433 3300 4447 3313
rect 4436 3296 4443 3300
rect 4456 3227 4463 3263
rect 4476 3207 4483 3316
rect 4516 3303 4523 3393
rect 4516 3296 4543 3303
rect 4576 3296 4583 3413
rect 4696 3387 4703 3453
rect 4716 3427 4723 3713
rect 4836 3627 4843 3953
rect 4876 3927 4883 4153
rect 4996 4007 5003 4233
rect 5056 4167 5063 4753
rect 5076 4427 5083 4573
rect 5096 4567 5103 4823
rect 5136 4820 5143 4823
rect 5133 4807 5147 4820
rect 5176 4727 5183 4854
rect 5376 4856 5383 4913
rect 5416 4867 5423 4893
rect 5276 4820 5283 4823
rect 5273 4807 5287 4820
rect 5227 4805 5240 4807
rect 5227 4793 5233 4805
rect 5136 4607 5143 4653
rect 5136 4556 5143 4593
rect 5176 4587 5183 4613
rect 5173 4560 5187 4573
rect 5176 4556 5183 4560
rect 5196 4447 5203 4512
rect 5216 4367 5223 4653
rect 5236 4507 5243 4713
rect 5336 4707 5343 4853
rect 5356 4763 5363 4793
rect 5373 4783 5387 4793
rect 5396 4787 5403 4823
rect 5436 4807 5443 5013
rect 5476 4887 5483 4933
rect 5496 4887 5503 5153
rect 5516 5087 5523 5173
rect 5516 5007 5523 5033
rect 5536 4983 5543 5043
rect 5516 4976 5543 4983
rect 5516 4907 5523 4976
rect 5576 4967 5583 5043
rect 5456 4856 5503 4863
rect 5536 4856 5543 4933
rect 5576 4867 5583 4913
rect 5373 4780 5393 4783
rect 5376 4776 5393 4780
rect 5356 4756 5383 4763
rect 5296 4556 5303 4613
rect 5336 4556 5343 4653
rect 5276 4520 5283 4523
rect 5273 4507 5287 4520
rect 5316 4447 5323 4512
rect 5376 4487 5383 4756
rect 5456 4747 5463 4856
rect 5476 4767 5483 4813
rect 5520 4805 5540 4807
rect 5527 4802 5540 4805
rect 5527 4793 5543 4802
rect 5536 4787 5543 4793
rect 5536 4776 5553 4787
rect 5540 4773 5553 4776
rect 5596 4747 5603 5013
rect 5636 5007 5643 5074
rect 5656 4967 5663 5173
rect 5736 5076 5743 5153
rect 5676 4927 5683 5033
rect 5716 5007 5723 5043
rect 5736 4967 5743 5013
rect 5756 4987 5763 5043
rect 5796 5027 5803 5113
rect 5876 5076 5883 5352
rect 5996 5303 6003 5374
rect 5976 5296 6003 5303
rect 5916 5107 5923 5133
rect 5936 5083 5943 5113
rect 5916 5076 5943 5083
rect 5856 5040 5863 5043
rect 5853 5027 5867 5040
rect 5673 4860 5687 4873
rect 5676 4856 5683 4860
rect 5616 4787 5623 4853
rect 5656 4787 5663 4823
rect 5696 4820 5703 4823
rect 5693 4807 5707 4820
rect 5196 4336 5223 4343
rect 5273 4340 5287 4353
rect 5276 4336 5283 4340
rect 5076 4296 5103 4303
rect 5076 4247 5083 4296
rect 5216 4187 5223 4336
rect 5356 4307 5363 4433
rect 5416 4336 5423 4473
rect 5456 4336 5463 4513
rect 5476 4447 5483 4693
rect 5300 4303 5313 4307
rect 5296 4296 5313 4303
rect 5300 4293 5313 4296
rect 5387 4303 5400 4307
rect 5387 4296 5403 4303
rect 5387 4293 5400 4296
rect 5056 4036 5063 4073
rect 5096 4007 5103 4093
rect 5176 4036 5183 4073
rect 4916 3967 4923 4003
rect 5036 3967 5043 4003
rect 5236 4003 5243 4053
rect 5196 3996 5243 4003
rect 5036 3816 5043 3953
rect 5073 3827 5087 3833
rect 5133 3820 5147 3833
rect 5136 3816 5143 3820
rect 4976 3786 4983 3813
rect 4876 3667 4883 3772
rect 4916 3687 4923 3783
rect 5056 3780 5063 3783
rect 5016 3727 5023 3772
rect 5053 3767 5067 3780
rect 5096 3767 5103 3793
rect 5216 3787 5223 3996
rect 4773 3520 4787 3533
rect 4776 3516 4783 3520
rect 4836 3527 4843 3613
rect 4756 3480 4763 3483
rect 4753 3467 4767 3480
rect 4833 3467 4847 3473
rect 4856 3407 4863 3533
rect 4953 3520 4967 3533
rect 4996 3527 5003 3693
rect 4956 3516 4963 3520
rect 4876 3467 4883 3514
rect 5053 3520 5067 3533
rect 5116 3528 5123 3653
rect 5056 3516 5063 3520
rect 4696 3296 4703 3373
rect 4496 3083 4503 3293
rect 4596 3187 4603 3263
rect 4496 3076 4523 3083
rect 4316 2996 4323 3073
rect 4216 2767 4223 2833
rect 4173 2480 4187 2493
rect 4176 2476 4183 2480
rect 4216 2476 4223 2753
rect 4236 2667 4243 2813
rect 4316 2807 4323 2933
rect 4336 2847 4343 2963
rect 4396 2947 4403 3053
rect 4496 2963 4503 3053
rect 4516 3007 4523 3076
rect 4476 2956 4503 2963
rect 4376 2743 4383 2833
rect 4476 2776 4483 2956
rect 4536 2907 4543 2963
rect 4356 2736 4383 2743
rect 4236 2487 4243 2593
rect 4256 2446 4263 2653
rect 4156 2407 4163 2443
rect 3956 2376 3983 2383
rect 3716 2167 3723 2223
rect 3536 1916 3563 1923
rect 3536 1767 3543 1916
rect 3520 1703 3533 1707
rect 3456 1696 3483 1703
rect 3516 1696 3533 1703
rect 3456 1663 3463 1696
rect 3520 1693 3533 1696
rect 3556 1687 3563 1833
rect 3576 1787 3583 1993
rect 3616 1956 3623 2073
rect 3636 1987 3643 2073
rect 3653 1960 3667 1973
rect 3696 1968 3703 2053
rect 3716 2007 3723 2093
rect 3656 1956 3663 1960
rect 3676 1920 3683 1923
rect 3673 1907 3687 1920
rect 3716 1847 3723 1913
rect 3736 1827 3743 2193
rect 3756 2107 3763 2223
rect 3776 2220 3803 2223
rect 3773 2216 3803 2220
rect 3773 2207 3787 2216
rect 3786 2200 3787 2207
rect 3756 1907 3763 2013
rect 3776 1967 3783 2153
rect 3796 2067 3803 2193
rect 3816 2127 3823 2213
rect 3836 2103 3843 2193
rect 3896 2167 3903 2193
rect 3916 2167 3923 2373
rect 3936 2287 3943 2353
rect 3956 2263 3963 2293
rect 3976 2287 3983 2376
rect 3956 2256 3983 2263
rect 3936 2227 3943 2252
rect 3816 2096 3843 2103
rect 3816 2047 3823 2096
rect 3836 1956 3843 2073
rect 3876 1923 3883 2113
rect 3976 2107 3983 2133
rect 3896 1963 3903 2013
rect 3996 1968 4003 2093
rect 4016 2087 4023 2173
rect 4036 2107 4043 2393
rect 4096 2256 4103 2313
rect 4116 2287 4123 2353
rect 4116 2167 4123 2223
rect 3896 1956 3923 1963
rect 3856 1916 3883 1923
rect 3436 1656 3463 1663
rect 3376 1447 3383 1472
rect 3416 1436 3423 1473
rect 3436 1447 3443 1656
rect 3456 1547 3463 1593
rect 3396 1307 3403 1392
rect 3433 1383 3447 1393
rect 3416 1380 3447 1383
rect 3416 1376 3443 1380
rect 3376 1216 3383 1253
rect 3416 1227 3423 1376
rect 3456 1367 3463 1434
rect 3173 948 3187 953
rect 3076 916 3083 920
rect 3027 913 3040 916
rect 3216 916 3223 1073
rect 3296 1027 3303 1173
rect 3396 1047 3403 1172
rect 3356 928 3363 953
rect 2907 876 2923 883
rect 2907 873 2920 876
rect 2916 767 2923 853
rect 2736 667 2743 694
rect 2636 660 2643 663
rect 2633 647 2647 660
rect 2876 666 2883 753
rect 2916 696 2923 732
rect 2953 700 2967 713
rect 2956 696 2963 700
rect 3056 703 3063 883
rect 3096 827 3103 883
rect 3136 847 3143 892
rect 3436 886 3443 1233
rect 3456 1147 3463 1353
rect 3476 1307 3483 1673
rect 3496 1447 3503 1673
rect 3576 1527 3583 1734
rect 3536 1436 3543 1513
rect 3496 1327 3503 1392
rect 3516 1263 3523 1403
rect 3556 1327 3563 1403
rect 3507 1256 3523 1263
rect 3496 1216 3503 1253
rect 3536 1223 3543 1293
rect 3616 1247 3623 1473
rect 3536 1216 3563 1223
rect 3533 1147 3547 1153
rect 3556 1107 3563 1216
rect 3576 1147 3583 1233
rect 3636 1216 3643 1703
rect 3653 1687 3667 1693
rect 3676 1667 3683 1813
rect 3696 1647 3703 1753
rect 3753 1740 3767 1753
rect 3816 1747 3823 1912
rect 3756 1736 3763 1740
rect 3813 1707 3827 1712
rect 3733 1687 3747 1692
rect 3776 1667 3783 1703
rect 3836 1687 3843 1853
rect 3856 1747 3863 1916
rect 3936 1887 3943 1923
rect 3876 1736 3883 1793
rect 3913 1748 3927 1753
rect 3676 1347 3683 1392
rect 3736 1363 3743 1433
rect 3756 1383 3763 1493
rect 3816 1400 3823 1403
rect 3813 1387 3827 1400
rect 3856 1387 3863 1473
rect 3756 1376 3783 1383
rect 3716 1356 3743 1363
rect 3716 1287 3723 1356
rect 3736 1307 3743 1333
rect 3656 1180 3663 1183
rect 3653 1167 3667 1180
rect 3533 920 3547 933
rect 3536 916 3543 920
rect 3036 696 3063 703
rect 3076 696 3083 813
rect 3113 708 3127 713
rect 3016 666 3023 693
rect 2536 496 2553 503
rect 2376 416 2403 423
rect 2416 420 2443 423
rect 2053 187 2067 193
rect 1793 122 1807 133
rect 1936 127 1943 173
rect 1996 127 2003 143
rect 1793 120 1853 122
rect 1796 115 1853 120
rect 1996 87 2003 113
rect 2076 107 2083 213
rect 2136 188 2143 353
rect 2156 227 2163 363
rect 2296 360 2303 363
rect 2096 107 2103 133
rect 2156 140 2163 143
rect 2153 127 2167 140
rect 2216 146 2223 253
rect 2276 203 2283 353
rect 2293 347 2307 360
rect 2276 196 2303 203
rect 2247 183 2260 187
rect 2247 176 2263 183
rect 2296 176 2303 196
rect 2336 183 2343 363
rect 2376 267 2383 353
rect 2396 327 2403 416
rect 2413 416 2443 420
rect 2413 407 2427 416
rect 2456 396 2463 433
rect 2436 307 2443 352
rect 2336 176 2363 183
rect 2247 173 2260 176
rect 2096 96 2113 107
rect 2100 93 2113 96
rect 2196 67 2203 133
rect 2316 140 2323 143
rect 2276 107 2283 132
rect 2313 127 2327 140
rect 2236 67 2243 93
rect 2356 87 2363 176
rect 2376 127 2383 213
rect 2396 187 2403 273
rect 2476 267 2483 363
rect 2516 303 2523 353
rect 2507 296 2523 303
rect 2416 176 2423 213
rect 2456 176 2463 213
rect 2496 187 2503 293
rect 2516 127 2523 213
rect 2440 125 2460 127
rect 2447 122 2460 125
rect 2447 113 2463 122
rect 2456 107 2463 113
rect 2536 107 2543 496
rect 2716 467 2723 652
rect 2753 647 2767 653
rect 2776 607 2783 663
rect 2816 567 2823 593
rect 2936 567 2943 663
rect 3036 547 3043 696
rect 3136 567 3143 663
rect 3176 587 3183 833
rect 3196 627 3203 793
rect 3216 703 3223 753
rect 3236 727 3243 883
rect 3376 847 3383 883
rect 3416 876 3433 883
rect 3416 827 3423 876
rect 3216 696 3243 703
rect 3276 696 3283 733
rect 3256 587 3263 663
rect 3296 656 3323 663
rect 2853 527 2867 533
rect 2847 520 2867 527
rect 2847 516 2863 520
rect 2847 513 2860 516
rect 2616 396 2623 433
rect 2756 396 2763 493
rect 2556 367 2563 394
rect 2696 367 2703 394
rect 2856 387 2863 493
rect 2896 407 2903 513
rect 2956 396 2963 453
rect 2993 408 3007 413
rect 3006 400 3007 408
rect 2596 327 2603 363
rect 2636 227 2643 352
rect 2696 267 2703 353
rect 2716 247 2723 373
rect 3016 367 3023 394
rect 2796 307 2803 333
rect 2816 327 2823 363
rect 2816 287 2823 313
rect 2836 267 2843 353
rect 2573 180 2587 193
rect 2576 176 2583 180
rect 2796 176 2803 253
rect 2676 147 2683 174
rect 2456 96 2473 107
rect 2460 93 2473 96
rect 2596 67 2603 143
rect 1987 56 2013 63
rect 2327 53 2333 67
rect 2387 53 2393 67
rect 2636 47 2643 143
rect 2696 47 2703 174
rect 2776 67 2783 143
rect 2856 107 2863 352
rect 2896 176 2903 353
rect 2976 227 2983 363
rect 3036 366 3043 453
rect 3127 414 3133 427
rect 3120 413 3140 414
rect 3176 366 3183 433
rect 3296 396 3303 613
rect 3316 407 3323 656
rect 3096 176 3103 293
rect 3116 247 3123 333
rect 3136 227 3143 363
rect 3176 227 3183 352
rect 3196 307 3203 394
rect 3236 287 3243 352
rect 3313 347 3327 353
rect 3113 207 3127 212
rect 3196 176 3203 253
rect 3236 176 3243 233
rect 3336 183 3343 793
rect 3516 747 3523 883
rect 3596 767 3603 993
rect 3653 920 3667 933
rect 3696 928 3703 1073
rect 3716 1007 3723 1213
rect 3736 967 3743 1233
rect 3756 1227 3763 1353
rect 3776 1347 3783 1376
rect 3776 1243 3783 1333
rect 3776 1236 3803 1243
rect 3796 1216 3803 1236
rect 3833 1220 3847 1233
rect 3856 1228 3863 1373
rect 3836 1216 3843 1220
rect 3876 1186 3883 1673
rect 3896 1547 3903 1703
rect 3956 1487 3963 1733
rect 3976 1627 3983 1893
rect 3996 1807 4003 1954
rect 4016 1748 4023 1973
rect 4036 1963 4043 1993
rect 4156 1987 4163 2213
rect 4176 2187 4183 2413
rect 4196 2087 4203 2333
rect 4256 2256 4263 2432
rect 4276 2407 4283 2613
rect 4316 2476 4323 2653
rect 4456 2627 4463 2743
rect 4496 2587 4503 2732
rect 4407 2476 4443 2483
rect 4336 2407 4343 2443
rect 4256 2107 4263 2133
rect 4036 1956 4063 1963
rect 4036 1927 4043 1956
rect 4276 1956 4283 2113
rect 4296 2047 4303 2273
rect 4356 2256 4363 2313
rect 4396 2267 4403 2474
rect 4456 2367 4463 2432
rect 4536 2307 4543 2853
rect 4576 2847 4583 2952
rect 4616 2867 4623 3193
rect 4676 2996 4683 3073
rect 4716 3047 4723 3263
rect 4756 3087 4763 3393
rect 4896 3363 4903 3473
rect 4936 3447 4943 3483
rect 4976 3463 4983 3483
rect 5016 3467 5023 3493
rect 5080 3483 5093 3487
rect 5076 3476 5093 3483
rect 5080 3473 5093 3476
rect 4956 3456 4983 3463
rect 4956 3407 4963 3456
rect 4896 3356 4923 3363
rect 4820 3323 4833 3327
rect 4816 3313 4833 3323
rect 4860 3323 4873 3327
rect 4856 3313 4873 3323
rect 4816 3296 4823 3313
rect 4856 3296 4863 3313
rect 4836 3247 4843 3263
rect 4833 3227 4847 3233
rect 4736 2966 4743 2993
rect 4696 2927 4703 2963
rect 4756 2867 4763 3073
rect 4840 3003 4853 3007
rect 4836 2996 4853 3003
rect 4840 2993 4853 2996
rect 4856 2927 4863 2953
rect 4876 2927 4883 3252
rect 4916 3203 4923 3356
rect 4933 3327 4947 3333
rect 4976 3327 4983 3433
rect 5036 3407 5043 3473
rect 5116 3467 5123 3514
rect 5136 3467 5143 3753
rect 5236 3627 5243 3973
rect 5256 3703 5263 4293
rect 5333 4040 5347 4053
rect 5336 4036 5343 4040
rect 5316 3967 5323 4003
rect 5396 3823 5403 4133
rect 5416 4007 5423 4253
rect 5496 4247 5503 4733
rect 5556 4556 5563 4593
rect 5636 4527 5643 4593
rect 5536 4303 5543 4523
rect 5656 4507 5663 4693
rect 5736 4556 5743 4813
rect 5756 4787 5763 4893
rect 5776 4887 5783 4953
rect 5836 4856 5843 5013
rect 5896 5007 5903 5043
rect 5876 4856 5883 4893
rect 5816 4767 5823 4823
rect 5856 4707 5863 4823
rect 5856 4556 5863 4613
rect 5916 4587 5923 5013
rect 5956 4927 5963 5273
rect 5976 5027 5983 5296
rect 6116 5287 6123 5343
rect 6176 5267 6183 5376
rect 6013 5080 6027 5093
rect 6016 5076 6023 5080
rect 6036 5007 6043 5043
rect 5956 4868 5963 4913
rect 6056 4827 6063 4873
rect 6076 4867 6083 5043
rect 6116 5007 6123 5193
rect 6136 5047 6143 5253
rect 6176 5076 6183 5113
rect 6236 5007 6243 5074
rect 6093 4860 6107 4873
rect 6096 4856 6103 4860
rect 6136 4856 6143 4913
rect 5616 4376 5623 4433
rect 5676 4387 5683 4513
rect 5676 4343 5683 4373
rect 5656 4336 5683 4343
rect 5536 4296 5563 4303
rect 5536 4267 5543 4296
rect 5456 4036 5463 4093
rect 5376 3816 5403 3823
rect 5436 3816 5443 3953
rect 5476 3887 5483 4003
rect 5536 3987 5543 4034
rect 5496 3863 5503 3973
rect 5556 3963 5563 4233
rect 5636 4036 5643 4093
rect 5616 4000 5623 4003
rect 5476 3856 5503 3863
rect 5536 3956 5563 3963
rect 5476 3816 5483 3856
rect 5276 3727 5283 3783
rect 5336 3767 5343 3783
rect 5376 3767 5383 3816
rect 5536 3827 5543 3956
rect 5516 3783 5523 3814
rect 5576 3816 5583 3993
rect 5613 3987 5627 4000
rect 5336 3756 5353 3767
rect 5340 3753 5353 3756
rect 5256 3696 5283 3703
rect 5276 3507 5283 3696
rect 5256 3476 5283 3483
rect 4976 3296 4983 3313
rect 4956 3260 4963 3263
rect 4953 3247 4967 3260
rect 4896 3196 4923 3203
rect 4896 2967 4903 3196
rect 4936 2996 4943 3033
rect 4976 2996 4983 3033
rect 4996 2927 5003 2963
rect 5036 2907 5043 2994
rect 4656 2747 4663 2813
rect 4616 2727 4623 2743
rect 4616 2716 4633 2727
rect 4620 2713 4633 2716
rect 4616 2647 4623 2673
rect 4636 2476 4643 2653
rect 4676 2563 4683 2833
rect 4736 2776 4743 2813
rect 4716 2740 4723 2743
rect 4713 2727 4727 2740
rect 4756 2707 4763 2743
rect 4816 2727 4823 2773
rect 4856 2607 4863 2743
rect 4896 2740 4903 2743
rect 4893 2727 4907 2740
rect 4907 2716 4923 2723
rect 4676 2556 4703 2563
rect 4616 2407 4623 2443
rect 4656 2407 4663 2443
rect 4416 2187 4423 2293
rect 4336 1968 4343 2173
rect 4376 1956 4383 1993
rect 4436 1956 4443 2212
rect 4456 2107 4463 2223
rect 4493 2207 4507 2212
rect 4536 2107 4543 2254
rect 4556 2226 4563 2353
rect 4656 2256 4663 2293
rect 4596 2220 4603 2223
rect 4593 2207 4607 2220
rect 4633 2207 4647 2212
rect 4596 2147 4603 2193
rect 4696 2107 4703 2556
rect 4816 2476 4823 2533
rect 4856 2446 4863 2593
rect 4916 2488 4923 2716
rect 4936 2667 4943 2773
rect 4956 2687 4963 2893
rect 5056 2788 5063 3333
rect 5076 3147 5083 3453
rect 5096 3307 5103 3452
rect 5216 3407 5223 3443
rect 5276 3427 5283 3476
rect 5296 3403 5303 3693
rect 5376 3647 5383 3753
rect 5376 3587 5383 3633
rect 5416 3627 5423 3783
rect 5456 3780 5463 3783
rect 5453 3767 5467 3780
rect 5516 3776 5563 3783
rect 5336 3516 5343 3573
rect 5536 3547 5543 3776
rect 5487 3516 5503 3523
rect 5556 3516 5563 3753
rect 5596 3707 5603 3772
rect 5636 3767 5643 3873
rect 5656 3707 5663 3953
rect 5673 3927 5687 3933
rect 5696 3907 5703 4493
rect 5776 4487 5783 4554
rect 5880 4523 5893 4527
rect 5836 4387 5843 4523
rect 5876 4516 5893 4523
rect 5880 4513 5893 4516
rect 5716 4287 5723 4373
rect 5796 4336 5803 4373
rect 5716 3947 5723 4233
rect 5796 4047 5803 4273
rect 5816 4247 5823 4303
rect 5856 4247 5863 4473
rect 5876 4287 5883 4493
rect 5916 4487 5923 4573
rect 5936 4547 5943 4793
rect 5976 4783 5983 4823
rect 6013 4807 6027 4812
rect 5956 4776 5983 4783
rect 5956 4687 5963 4776
rect 5956 4567 5963 4673
rect 6013 4560 6027 4573
rect 6036 4567 6043 4773
rect 6056 4627 6063 4693
rect 6016 4556 6023 4560
rect 5936 4447 5943 4533
rect 6056 4527 6063 4613
rect 6136 4556 6143 4773
rect 6176 4687 6183 4993
rect 6256 4856 6263 4953
rect 6196 4707 6203 4854
rect 6316 4567 6323 4812
rect 5936 4336 5943 4433
rect 5916 4207 5923 4303
rect 5956 4287 5963 4303
rect 6016 4283 6023 4493
rect 6116 4487 6123 4523
rect 6156 4503 6163 4512
rect 6136 4496 6163 4503
rect 6036 4303 6043 4473
rect 6036 4296 6063 4303
rect 6016 4276 6043 4283
rect 5747 4043 5760 4047
rect 5747 4036 5763 4043
rect 5747 4033 5760 4036
rect 5816 4027 5823 4193
rect 5916 4036 5923 4133
rect 5776 4000 5783 4003
rect 5736 3963 5743 3993
rect 5773 3987 5787 4000
rect 5836 3996 5863 4003
rect 5736 3956 5773 3963
rect 5736 3887 5743 3933
rect 5756 3816 5763 3913
rect 5776 3827 5783 3932
rect 5736 3780 5743 3783
rect 5733 3767 5747 3780
rect 5796 3747 5803 3993
rect 5836 3967 5843 3996
rect 5896 3907 5903 4003
rect 5856 3816 5863 3873
rect 5936 3847 5943 3992
rect 5956 3927 5963 4273
rect 6036 4036 6043 4276
rect 6056 4207 6063 4296
rect 6136 4267 6143 4496
rect 6216 4487 6223 4554
rect 6176 4336 6183 4413
rect 6196 4300 6203 4303
rect 6193 4287 6207 4300
rect 6236 4267 6243 4303
rect 6276 4283 6283 4473
rect 6267 4276 6283 4283
rect 5976 3887 5983 4034
rect 6016 3987 6023 4034
rect 5893 3820 5907 3833
rect 5896 3816 5903 3820
rect 5836 3780 5843 3783
rect 5816 3743 5823 3773
rect 5833 3767 5847 3780
rect 5936 3747 5943 3833
rect 6033 3820 6047 3833
rect 6036 3816 6043 3820
rect 5816 3736 5843 3743
rect 5396 3480 5403 3483
rect 5393 3467 5407 3480
rect 5276 3396 5303 3403
rect 5136 3296 5143 3333
rect 5116 3087 5123 3252
rect 5156 3167 5163 3263
rect 5076 3007 5083 3073
rect 5116 2996 5123 3033
rect 5076 2827 5083 2953
rect 5096 2867 5103 2963
rect 5076 2783 5083 2813
rect 5076 2776 5103 2783
rect 5156 2747 5163 3153
rect 5016 2740 5023 2743
rect 5013 2727 5027 2740
rect 4956 2476 4963 2593
rect 4976 2387 4983 2443
rect 5036 2407 5043 2653
rect 4976 2307 4983 2373
rect 5036 2323 5043 2393
rect 5016 2316 5043 2323
rect 4896 2256 4903 2293
rect 4996 2267 5003 2313
rect 5016 2256 5023 2316
rect 5056 2256 5063 2733
rect 5116 2727 5123 2743
rect 5176 2727 5183 3093
rect 5196 3007 5203 3233
rect 5216 3107 5223 3333
rect 5276 3308 5283 3396
rect 5313 3300 5327 3313
rect 5316 3296 5323 3300
rect 5256 3067 5263 3263
rect 5296 3260 5303 3263
rect 5293 3247 5307 3260
rect 5276 2996 5283 3153
rect 5356 3127 5363 3413
rect 5476 3367 5483 3514
rect 5536 3467 5543 3483
rect 5547 3460 5563 3463
rect 5547 3456 5567 3460
rect 5553 3447 5567 3456
rect 5576 3323 5583 3533
rect 5636 3516 5643 3653
rect 5736 3487 5743 3732
rect 5616 3427 5623 3473
rect 5656 3387 5663 3483
rect 5756 3447 5763 3693
rect 5836 3516 5843 3736
rect 5956 3707 5963 3814
rect 5873 3520 5887 3533
rect 5876 3516 5883 3520
rect 5567 3316 5583 3323
rect 5296 3047 5303 3093
rect 5376 3067 5383 3293
rect 5496 3266 5503 3313
rect 5553 3300 5567 3313
rect 5556 3296 5563 3300
rect 5416 3227 5423 3263
rect 5536 3260 5543 3263
rect 5533 3247 5547 3260
rect 5576 3243 5583 3263
rect 5576 3236 5603 3243
rect 5473 3227 5487 3233
rect 5196 2927 5203 2953
rect 5216 2788 5223 2963
rect 5256 2943 5263 2963
rect 5256 2936 5283 2943
rect 5256 2776 5263 2913
rect 5276 2887 5283 2936
rect 5296 2783 5303 2953
rect 5316 2807 5323 3053
rect 5296 2776 5323 2783
rect 5236 2740 5243 2743
rect 5233 2727 5247 2740
rect 5116 2713 5133 2727
rect 5116 2687 5123 2713
rect 5136 2476 5143 2533
rect 5196 2443 5203 2474
rect 5076 2327 5083 2433
rect 5116 2387 5123 2443
rect 5156 2263 5163 2443
rect 5176 2436 5203 2443
rect 5176 2268 5183 2436
rect 5216 2427 5223 2513
rect 5256 2476 5263 2533
rect 5316 2507 5323 2776
rect 5336 2743 5343 3013
rect 5376 2996 5383 3032
rect 5413 3000 5427 3013
rect 5456 3007 5463 3153
rect 5416 2996 5423 3000
rect 5440 2963 5453 2967
rect 5396 2827 5403 2963
rect 5436 2956 5453 2963
rect 5440 2953 5453 2956
rect 5476 2947 5483 3213
rect 5553 3000 5567 3013
rect 5596 3007 5603 3236
rect 5616 3207 5623 3253
rect 5556 2996 5563 3000
rect 5616 2963 5623 2994
rect 5373 2780 5387 2793
rect 5376 2776 5383 2780
rect 5436 2747 5443 2933
rect 5536 2887 5543 2963
rect 5576 2960 5583 2963
rect 5573 2947 5587 2960
rect 5596 2956 5623 2963
rect 5596 2907 5603 2956
rect 5636 2947 5643 3353
rect 5716 3327 5723 3433
rect 5713 3300 5727 3313
rect 5736 3307 5743 3413
rect 5716 3296 5723 3300
rect 5656 3007 5663 3253
rect 5736 3163 5743 3253
rect 5756 3187 5763 3433
rect 5776 3307 5783 3472
rect 5816 3447 5823 3483
rect 5816 3296 5823 3433
rect 5916 3387 5923 3533
rect 5936 3528 5943 3553
rect 5987 3543 6000 3547
rect 5987 3533 6003 3543
rect 5996 3516 6003 3533
rect 5896 3267 5903 3293
rect 5796 3260 5803 3263
rect 5836 3260 5843 3263
rect 5773 3247 5787 3253
rect 5793 3247 5807 3260
rect 5833 3247 5847 3260
rect 5736 3156 5763 3163
rect 5696 3008 5703 3033
rect 5756 3007 5763 3156
rect 5667 2956 5683 2963
rect 5716 2960 5723 2963
rect 5536 2776 5543 2833
rect 5336 2736 5353 2743
rect 5356 2443 5363 2732
rect 5376 2487 5383 2593
rect 5476 2547 5483 2733
rect 5516 2723 5523 2743
rect 5496 2716 5523 2723
rect 5416 2476 5423 2513
rect 5136 2256 5163 2263
rect 4756 2147 4763 2223
rect 4796 2220 4803 2223
rect 4793 2207 4807 2220
rect 4956 2187 4963 2253
rect 5116 2223 5123 2254
rect 5096 2216 5123 2223
rect 5036 2202 5043 2212
rect 5036 2195 5073 2202
rect 5096 2187 5103 2216
rect 5136 2187 5143 2256
rect 5216 2256 5223 2293
rect 5256 2267 5263 2393
rect 5276 2367 5283 2443
rect 5316 2436 5363 2443
rect 5196 2220 5203 2223
rect 5193 2207 5207 2220
rect 5276 2226 5283 2293
rect 5296 2267 5303 2413
rect 5333 2260 5347 2273
rect 5336 2256 5343 2260
rect 5376 2256 5383 2333
rect 5396 2327 5403 2432
rect 4536 2007 4543 2093
rect 4616 2047 4623 2093
rect 4156 1916 4183 1923
rect 4256 1920 4263 1923
rect 4176 1887 4183 1916
rect 4253 1907 4267 1920
rect 4116 1827 4123 1883
rect 3916 1347 3923 1403
rect 3896 1227 3903 1253
rect 3913 1228 3927 1233
rect 3956 1216 3963 1253
rect 3976 1243 3983 1533
rect 4036 1507 4043 1703
rect 4076 1700 4083 1703
rect 4073 1687 4087 1700
rect 4116 1607 4123 1792
rect 4136 1687 4143 1733
rect 4156 1703 4163 1753
rect 4296 1743 4303 1853
rect 4276 1736 4303 1743
rect 4156 1696 4183 1703
rect 4076 1436 4083 1533
rect 3996 1387 4003 1433
rect 4056 1400 4063 1403
rect 4053 1387 4067 1400
rect 4007 1376 4023 1383
rect 3993 1243 4007 1253
rect 3976 1236 4007 1243
rect 3993 1227 4007 1236
rect 4016 1186 4023 1376
rect 4067 1376 4083 1383
rect 4036 1227 4043 1373
rect 4076 1216 4083 1376
rect 4096 1367 4103 1403
rect 4136 1307 4143 1553
rect 4176 1447 4183 1593
rect 4296 1567 4303 1713
rect 4316 1706 4323 1813
rect 4336 1747 4343 1954
rect 4396 1867 4403 1923
rect 4576 1920 4583 1923
rect 4573 1907 4587 1920
rect 4616 1907 4623 2033
rect 4676 2027 4683 2053
rect 4676 1956 4683 2013
rect 4713 1960 4727 1973
rect 4716 1956 4723 1960
rect 4756 1926 4763 1973
rect 4876 1963 4883 2013
rect 4796 1956 4823 1963
rect 4876 1956 4903 1963
rect 4976 1956 4983 2073
rect 5036 1987 5043 2073
rect 4433 1767 4447 1773
rect 4616 1767 4623 1893
rect 4396 1700 4403 1703
rect 4247 1460 4263 1463
rect 4247 1456 4267 1460
rect 4156 1367 4163 1434
rect 4233 1440 4247 1453
rect 4253 1447 4267 1456
rect 4236 1436 4243 1440
rect 4173 1387 4187 1393
rect 4176 1227 4183 1253
rect 4116 1216 4163 1223
rect 3656 916 3663 920
rect 3896 927 3903 1173
rect 4096 1180 4103 1183
rect 4093 1167 4107 1180
rect 3876 916 3893 923
rect 3676 847 3683 883
rect 3506 733 3507 740
rect 3493 723 3507 733
rect 3493 720 3523 723
rect 3496 716 3523 720
rect 3516 696 3523 716
rect 3396 527 3403 652
rect 3436 627 3443 663
rect 3476 643 3483 694
rect 3713 700 3727 713
rect 3716 696 3723 700
rect 3476 636 3503 643
rect 3476 367 3483 553
rect 3496 507 3503 636
rect 3536 623 3543 652
rect 3536 616 3563 623
rect 3376 287 3383 363
rect 3496 347 3503 493
rect 3536 408 3543 593
rect 3556 507 3563 616
rect 3576 607 3583 663
rect 3636 563 3643 693
rect 3776 666 3783 733
rect 3796 666 3803 853
rect 3816 727 3823 883
rect 3916 886 3923 953
rect 3896 827 3903 873
rect 3853 700 3867 713
rect 3936 708 3943 993
rect 3976 916 3983 953
rect 4156 947 4163 1216
rect 4193 1220 4207 1233
rect 4233 1220 4247 1233
rect 4276 1227 4283 1493
rect 4316 1467 4323 1692
rect 4393 1687 4407 1700
rect 4436 1507 4443 1732
rect 4456 1687 4463 1753
rect 4493 1748 4507 1753
rect 4533 1740 4547 1753
rect 4536 1736 4543 1740
rect 4516 1700 4523 1703
rect 4476 1436 4483 1693
rect 4513 1687 4527 1700
rect 4576 1687 4583 1753
rect 4696 1748 4703 1923
rect 4796 1847 4803 1956
rect 4616 1700 4623 1703
rect 4613 1687 4627 1700
rect 4293 1387 4307 1392
rect 4316 1367 4323 1403
rect 4396 1327 4403 1433
rect 4196 1216 4203 1220
rect 4236 1216 4243 1220
rect 4296 1007 4303 1233
rect 4316 1127 4323 1313
rect 4356 1216 4363 1273
rect 4416 1223 4423 1333
rect 4516 1247 4523 1613
rect 4556 1447 4563 1493
rect 4696 1467 4703 1734
rect 4536 1407 4543 1434
rect 4613 1440 4627 1453
rect 4653 1447 4667 1453
rect 4616 1436 4623 1440
rect 4596 1400 4603 1403
rect 4593 1387 4607 1400
rect 4396 1216 4423 1223
rect 4456 1187 4463 1214
rect 4476 1007 4483 1233
rect 4496 1087 4503 1183
rect 4556 1127 4563 1172
rect 4576 1047 4583 1333
rect 4636 1287 4643 1403
rect 4676 1347 4683 1433
rect 4696 1406 4703 1453
rect 4716 1447 4723 1753
rect 4796 1736 4803 1793
rect 4836 1767 4843 1912
rect 4820 1703 4833 1707
rect 4776 1700 4783 1703
rect 4773 1687 4787 1700
rect 4816 1696 4833 1703
rect 4820 1693 4833 1696
rect 4836 1667 4843 1693
rect 4736 1436 4743 1493
rect 4836 1467 4843 1653
rect 4773 1440 4787 1453
rect 4856 1448 4863 1833
rect 4896 1767 4903 1956
rect 5056 1927 5063 2033
rect 4913 1740 4927 1753
rect 4916 1736 4923 1740
rect 4936 1467 4943 1703
rect 4976 1607 4983 1703
rect 5016 1687 5023 1793
rect 5076 1767 5083 1993
rect 5256 1963 5263 2213
rect 5416 2223 5423 2413
rect 5436 2367 5443 2443
rect 5456 2327 5463 2393
rect 5496 2347 5503 2716
rect 5556 2707 5563 2743
rect 5596 2647 5603 2893
rect 5616 2847 5623 2933
rect 5656 2776 5663 2953
rect 5713 2947 5727 2960
rect 5616 2736 5643 2743
rect 5616 2667 5623 2736
rect 5556 2476 5563 2513
rect 5593 2480 5607 2493
rect 5616 2487 5623 2653
rect 5596 2476 5603 2480
rect 5536 2407 5543 2443
rect 5576 2403 5583 2443
rect 5576 2396 5603 2403
rect 5476 2316 5523 2323
rect 5476 2287 5483 2316
rect 5407 2216 5423 2223
rect 5393 2207 5407 2212
rect 5236 1956 5263 1963
rect 5276 1956 5283 2033
rect 5156 1880 5163 1883
rect 5153 1867 5167 1880
rect 5216 1867 5223 1954
rect 5236 1787 5243 1956
rect 5296 1847 5303 1923
rect 5336 1887 5343 1912
rect 5076 1736 5083 1753
rect 4776 1436 4783 1440
rect 4873 1440 4887 1453
rect 4876 1436 4883 1440
rect 4976 1406 4983 1593
rect 5056 1587 5063 1703
rect 5096 1700 5103 1703
rect 5093 1687 5107 1700
rect 5096 1627 5103 1673
rect 5156 1507 5163 1753
rect 5213 1740 5227 1753
rect 5216 1736 5223 1740
rect 5196 1587 5203 1703
rect 5236 1627 5243 1703
rect 4596 1147 4603 1233
rect 4616 1187 4623 1253
rect 4676 1243 4683 1333
rect 4796 1307 4803 1403
rect 4896 1387 4903 1403
rect 4896 1376 4913 1387
rect 4900 1373 4913 1376
rect 4676 1236 4703 1243
rect 4653 1220 4667 1233
rect 4656 1216 4663 1220
rect 4696 1216 4703 1236
rect 4013 920 4027 933
rect 4016 916 4023 920
rect 4176 916 4183 993
rect 3956 747 3963 873
rect 3976 723 3983 753
rect 3956 716 3983 723
rect 4036 723 4043 883
rect 4096 847 4103 914
rect 4256 886 4263 933
rect 4296 916 4303 993
rect 4576 923 4583 1033
rect 4556 916 4583 923
rect 4596 916 4603 973
rect 4636 928 4643 1133
rect 4676 1067 4683 1183
rect 4756 1007 4763 1293
rect 4936 1267 4943 1403
rect 4996 1327 5003 1453
rect 5073 1440 5087 1453
rect 5076 1436 5083 1440
rect 5096 1367 5103 1403
rect 4796 1228 4803 1253
rect 4940 1243 4953 1247
rect 4833 1220 4847 1233
rect 4936 1233 4953 1243
rect 4836 1216 4843 1220
rect 4936 1216 4943 1233
rect 4876 1186 4883 1213
rect 4816 1167 4823 1183
rect 4996 1186 5003 1233
rect 5016 1187 5023 1233
rect 5036 1187 5043 1273
rect 4816 1156 4833 1167
rect 4820 1153 4833 1156
rect 4876 1147 4883 1172
rect 4913 1143 4927 1151
rect 4913 1140 4953 1143
rect 4916 1136 4953 1140
rect 4196 867 4203 883
rect 4196 856 4213 867
rect 4200 853 4213 856
rect 4036 716 4063 723
rect 3856 696 3863 700
rect 3786 652 3787 660
rect 3876 660 3883 663
rect 3773 647 3787 652
rect 3873 647 3887 660
rect 3956 663 3963 716
rect 3956 656 3983 663
rect 3636 556 3663 563
rect 3576 396 3583 433
rect 3636 367 3643 533
rect 3600 363 3613 367
rect 3556 360 3563 363
rect 3456 247 3463 273
rect 3316 176 3343 183
rect 1416 36 1473 43
rect 2876 23 2883 132
rect 2916 127 2923 143
rect 2896 116 2913 123
rect 2896 87 2903 116
rect 2916 47 2923 92
rect 2996 67 3003 174
rect 3136 146 3143 174
rect 3036 67 3043 143
rect 3076 140 3083 143
rect 3073 127 3087 140
rect 3136 107 3143 132
rect 3156 127 3163 174
rect 3316 146 3323 176
rect 3356 140 3363 143
rect 3396 140 3403 143
rect 3313 127 3327 132
rect 3353 127 3367 140
rect 3393 127 3407 140
rect 3456 127 3463 233
rect 3516 227 3523 353
rect 3553 347 3567 360
rect 3596 356 3613 363
rect 3600 353 3613 356
rect 3656 327 3663 556
rect 3676 527 3683 613
rect 3916 587 3923 653
rect 4036 647 4043 663
rect 3676 407 3683 473
rect 3716 427 3723 573
rect 3720 363 3733 367
rect 3716 356 3733 363
rect 3720 353 3733 356
rect 3736 267 3743 293
rect 3756 287 3763 394
rect 3776 367 3783 513
rect 3876 396 3883 493
rect 3936 367 3943 453
rect 3956 408 3963 533
rect 4036 507 4043 633
rect 4056 587 4063 716
rect 4076 627 4083 753
rect 4156 627 4163 663
rect 4196 647 4203 833
rect 4256 696 4263 793
rect 4296 696 4303 733
rect 4356 723 4363 883
rect 4373 867 4387 873
rect 4396 847 4403 914
rect 4416 767 4423 893
rect 4556 886 4563 916
rect 4476 863 4483 883
rect 4476 856 4503 863
rect 4453 847 4467 853
rect 4347 716 4363 723
rect 4336 687 4343 713
rect 4376 703 4383 733
rect 4356 696 4383 703
rect 4227 663 4240 667
rect 4227 653 4243 663
rect 4236 642 4243 653
rect 4236 635 4273 642
rect 3996 396 4003 493
rect 4033 400 4047 413
rect 4056 403 4063 573
rect 4076 427 4083 513
rect 4136 408 4143 473
rect 4036 396 4043 400
rect 4056 396 4083 403
rect 4076 366 4083 396
rect 4173 400 4187 413
rect 4176 396 4183 400
rect 4216 366 4223 413
rect 4276 396 4283 473
rect 4316 427 4323 653
rect 4356 647 4363 696
rect 4456 696 4463 753
rect 4396 627 4403 663
rect 4476 447 4483 653
rect 4496 587 4503 856
rect 4516 827 4523 883
rect 4347 436 4363 443
rect 4336 403 4343 433
rect 4316 396 4343 403
rect 3976 307 3983 363
rect 3787 293 3793 307
rect 4116 267 4123 363
rect 4156 327 4163 363
rect 3553 180 3567 193
rect 3556 176 3563 180
rect 3693 180 3707 193
rect 3756 188 3763 233
rect 3696 176 3703 180
rect 3476 107 3483 173
rect 3533 127 3547 132
rect 3287 93 3293 107
rect 3360 106 3380 107
rect 3056 47 3063 93
rect 3367 93 3373 106
rect 2907 36 2923 47
rect 2907 33 2920 36
rect 3387 36 3413 43
rect 3616 27 3623 173
rect 3776 146 3783 233
rect 3836 176 3843 253
rect 3676 140 3683 143
rect 3673 127 3687 140
rect 3716 107 3723 143
rect 3916 47 3923 253
rect 3936 127 3943 213
rect 3996 176 4003 253
rect 4056 187 4063 253
rect 4116 207 4123 253
rect 4076 146 4083 193
rect 4196 183 4203 213
rect 4256 207 4263 363
rect 4356 327 4363 436
rect 4516 407 4523 753
rect 4596 708 4603 833
rect 4616 723 4623 883
rect 4616 720 4643 723
rect 4616 716 4647 720
rect 4633 707 4647 716
rect 4576 587 4583 663
rect 4656 666 4663 733
rect 4696 703 4703 993
rect 4716 807 4723 973
rect 4676 696 4703 703
rect 4716 696 4723 733
rect 4756 696 4763 833
rect 4796 703 4803 883
rect 4856 847 4863 973
rect 4896 847 4903 883
rect 4896 807 4903 833
rect 4936 807 4943 873
rect 4956 787 4963 1053
rect 4976 1047 4983 1173
rect 5056 1180 5063 1183
rect 5053 1167 5067 1180
rect 5013 1147 5027 1152
rect 5040 1146 5060 1147
rect 5047 1133 5053 1146
rect 5016 916 5023 1073
rect 5096 1067 5103 1153
rect 5096 886 5103 1053
rect 5136 1027 5143 1253
rect 5156 987 5163 1453
rect 5196 1448 5203 1573
rect 5296 1523 5303 1773
rect 5356 1736 5363 1913
rect 5376 1847 5383 2073
rect 5396 1927 5403 2193
rect 5436 2187 5443 2273
rect 5496 2268 5503 2293
rect 5516 2287 5523 2316
rect 5536 2256 5543 2293
rect 5476 2187 5483 2223
rect 5516 2220 5523 2223
rect 5513 2207 5527 2220
rect 5576 2183 5583 2373
rect 5596 2347 5603 2396
rect 5616 2263 5623 2433
rect 5636 2427 5643 2693
rect 5716 2687 5723 2833
rect 5736 2707 5743 2813
rect 5756 2788 5763 2953
rect 5776 2887 5783 3233
rect 5796 2827 5803 3013
rect 5816 3007 5823 3113
rect 5916 3087 5923 3333
rect 5936 3307 5943 3514
rect 5976 3427 5983 3483
rect 6016 3407 6023 3483
rect 5976 3296 5983 3373
rect 6056 3347 6063 3733
rect 6020 3303 6033 3307
rect 6016 3296 6033 3303
rect 6020 3293 6033 3296
rect 5947 3263 5960 3267
rect 5947 3256 5963 3263
rect 5947 3253 5960 3256
rect 5833 3000 5847 3013
rect 5836 2996 5843 3000
rect 5876 2996 5883 3053
rect 5936 2967 5943 3232
rect 5956 3007 5963 3153
rect 5996 3027 6003 3263
rect 6056 3247 6063 3293
rect 6076 3263 6083 3971
rect 6096 3827 6103 3853
rect 6116 3816 6123 3873
rect 6136 3867 6143 4003
rect 6236 3987 6243 4253
rect 6153 3828 6167 3833
rect 6176 3776 6203 3783
rect 6136 3763 6143 3772
rect 6116 3756 6143 3763
rect 6116 3516 6123 3756
rect 6196 3707 6203 3776
rect 6176 3487 6183 3653
rect 6136 3480 6143 3483
rect 6096 3407 6103 3473
rect 6133 3467 6147 3480
rect 6096 3307 6103 3393
rect 6136 3296 6143 3413
rect 6176 3307 6183 3452
rect 6076 3256 6103 3263
rect 6016 3067 6023 3233
rect 5993 3000 6007 3013
rect 5996 2996 6003 3000
rect 6036 2996 6043 3173
rect 6056 3007 6063 3073
rect 5816 2847 5823 2953
rect 5836 2807 5843 2893
rect 5756 2746 5763 2774
rect 5636 2307 5643 2413
rect 5656 2387 5663 2493
rect 5696 2476 5703 2533
rect 5716 2436 5733 2443
rect 5640 2286 5660 2287
rect 5647 2283 5660 2286
rect 5647 2273 5663 2283
rect 5596 2256 5623 2263
rect 5656 2256 5663 2273
rect 5696 2256 5703 2393
rect 5596 2223 5603 2256
rect 5596 2216 5623 2223
rect 5576 2176 5593 2183
rect 5416 1956 5433 1963
rect 5416 1867 5423 1956
rect 5496 1767 5503 1883
rect 5596 1867 5603 2173
rect 5393 1740 5407 1753
rect 5396 1736 5403 1740
rect 5427 1733 5433 1747
rect 5456 1706 5463 1753
rect 5487 1743 5500 1747
rect 5487 1736 5503 1743
rect 5487 1733 5500 1736
rect 5276 1516 5303 1523
rect 5236 1436 5243 1493
rect 5216 1307 5223 1403
rect 5236 1216 5243 1253
rect 5276 1227 5283 1516
rect 5296 1406 5303 1493
rect 5336 1487 5343 1692
rect 5516 1683 5523 1703
rect 5567 1696 5583 1703
rect 5496 1676 5523 1683
rect 5496 1587 5503 1676
rect 5496 1436 5503 1573
rect 5396 1363 5403 1403
rect 5436 1367 5443 1434
rect 5556 1407 5563 1671
rect 5396 1356 5423 1363
rect 5396 1216 5403 1333
rect 5416 1247 5423 1356
rect 5456 1327 5463 1373
rect 5476 1367 5483 1403
rect 5487 1356 5503 1363
rect 5256 1107 5263 1183
rect 5296 1147 5303 1193
rect 5316 1107 5323 1214
rect 5333 1167 5347 1173
rect 5376 1147 5383 1183
rect 5176 927 5183 1093
rect 4996 863 5003 883
rect 4996 856 5023 863
rect 4796 696 4823 703
rect 4876 696 4883 753
rect 4913 700 4927 713
rect 4916 696 4923 700
rect 4213 183 4227 193
rect 4196 180 4227 183
rect 4196 176 4223 180
rect 3976 140 3983 143
rect 3973 127 3987 140
rect 3933 107 3947 113
rect 4096 67 4103 173
rect 4136 140 4143 143
rect 4133 127 4147 140
rect 4236 107 4243 173
rect 4256 146 4263 193
rect 4276 187 4283 253
rect 4416 227 4423 363
rect 4316 176 4323 213
rect 4476 207 4483 393
rect 4496 307 4503 394
rect 4556 396 4563 433
rect 4636 366 4643 653
rect 4676 587 4683 696
rect 4816 666 4823 696
rect 4696 627 4703 653
rect 4776 627 4783 663
rect 4676 408 4683 573
rect 4696 527 4703 613
rect 4716 396 4723 433
rect 4696 327 4703 363
rect 4347 193 4353 207
rect 4356 176 4403 183
rect 4396 107 4403 176
rect 4436 123 4443 143
rect 4436 116 4463 123
rect 4427 93 4433 107
rect 4456 87 4463 116
rect 4516 87 4523 193
rect 4536 146 4543 313
rect 4686 293 4687 300
rect 4673 283 4687 293
rect 4716 283 4723 313
rect 4673 280 4723 283
rect 4676 276 4723 280
rect 4596 176 4603 273
rect 4796 227 4803 513
rect 4816 366 4823 613
rect 4896 423 4903 652
rect 4936 587 4943 663
rect 4976 627 4983 713
rect 4996 707 5003 833
rect 5016 767 5023 856
rect 5076 707 5083 793
rect 5096 666 5103 773
rect 5216 707 5223 973
rect 5233 967 5247 973
rect 5236 927 5243 953
rect 5256 916 5263 993
rect 5336 927 5343 1013
rect 5236 708 5243 873
rect 5276 747 5283 883
rect 5316 787 5323 883
rect 5336 827 5343 873
rect 5356 727 5363 1033
rect 5376 967 5383 1073
rect 5416 1067 5423 1183
rect 5436 1027 5443 1173
rect 5456 1147 5463 1233
rect 5476 1027 5483 1253
rect 5496 1227 5503 1356
rect 5516 1307 5523 1403
rect 5516 1247 5523 1293
rect 5536 1216 5543 1273
rect 5576 1227 5583 1696
rect 5596 1647 5603 1733
rect 5616 1687 5623 2216
rect 5676 2187 5683 2223
rect 5736 2087 5743 2433
rect 5756 2223 5763 2732
rect 5776 2667 5783 2743
rect 5856 2707 5863 2963
rect 5876 2747 5883 2933
rect 5896 2743 5903 2893
rect 5956 2776 5963 2953
rect 5976 2807 5983 2963
rect 6076 2847 6083 3133
rect 6096 3127 6103 3256
rect 6116 3227 6123 3263
rect 6116 3147 6123 3173
rect 6116 3027 6123 3133
rect 6136 3027 6143 3233
rect 6156 3207 6163 3263
rect 6176 3023 6183 3253
rect 6196 3167 6203 3693
rect 6216 3667 6223 3853
rect 6256 3827 6263 4273
rect 6236 3787 6243 3814
rect 6296 3816 6303 3853
rect 6236 3516 6243 3553
rect 6256 3327 6263 3483
rect 6296 3443 6303 3473
rect 6287 3436 6303 3443
rect 6216 3267 6223 3313
rect 6276 3296 6283 3433
rect 6316 3387 6323 3773
rect 6253 3247 6267 3252
rect 6176 3020 6203 3023
rect 6176 3016 6207 3020
rect 6133 3000 6147 3013
rect 6136 2996 6143 3000
rect 6193 3007 6207 3016
rect 6216 2963 6223 3232
rect 6296 3207 6303 3263
rect 6233 3007 6247 3013
rect 6256 2996 6263 3133
rect 6196 2956 6223 2963
rect 6136 2776 6143 2933
rect 6156 2787 6163 2833
rect 5896 2736 5923 2743
rect 5776 2407 5783 2474
rect 5807 2483 5820 2487
rect 5807 2476 5823 2483
rect 5853 2480 5867 2493
rect 5856 2476 5863 2480
rect 5807 2473 5820 2476
rect 5836 2440 5843 2443
rect 5876 2440 5883 2443
rect 5833 2427 5847 2440
rect 5873 2427 5887 2440
rect 5916 2407 5923 2736
rect 5976 2727 5983 2743
rect 6036 2727 6043 2774
rect 6067 2743 6080 2747
rect 6067 2736 6083 2743
rect 6067 2733 6080 2736
rect 5956 2716 5973 2723
rect 5856 2256 5863 2393
rect 5936 2347 5943 2493
rect 5956 2487 5963 2716
rect 5976 2476 5983 2533
rect 6056 2487 6063 2673
rect 5956 2307 5963 2433
rect 5996 2367 6003 2443
rect 6036 2387 6043 2443
rect 6076 2427 6083 2693
rect 6156 2527 6163 2733
rect 6176 2727 6183 2913
rect 6196 2703 6203 2956
rect 6216 2787 6223 2933
rect 6256 2788 6263 2933
rect 6276 2907 6283 2963
rect 6316 2927 6323 3113
rect 6236 2723 6243 2743
rect 6236 2716 6263 2723
rect 6196 2696 6213 2703
rect 5756 2216 5803 2223
rect 5656 1736 5663 1853
rect 5676 1767 5683 1883
rect 5693 1740 5707 1753
rect 5696 1736 5703 1740
rect 5720 1703 5733 1707
rect 5616 1436 5623 1473
rect 5656 1448 5663 1653
rect 5676 1587 5683 1703
rect 5716 1696 5733 1703
rect 5720 1693 5733 1696
rect 5596 1183 5603 1393
rect 5613 1227 5627 1233
rect 5636 1216 5643 1353
rect 5676 1307 5683 1403
rect 5716 1283 5723 1673
rect 5736 1667 5743 1693
rect 5756 1643 5763 1753
rect 5776 1687 5783 2216
rect 5836 2103 5843 2223
rect 5896 2207 5903 2253
rect 5916 2127 5923 2293
rect 6076 2267 6083 2413
rect 6096 2387 6103 2493
rect 6153 2480 6167 2492
rect 6193 2480 6207 2493
rect 6216 2487 6223 2693
rect 6156 2476 6163 2480
rect 6196 2476 6203 2480
rect 6096 2287 6103 2373
rect 5816 2096 5843 2103
rect 5796 1867 5803 2033
rect 5816 1967 5823 2096
rect 5976 1987 5983 2223
rect 6016 2216 6033 2223
rect 6007 2193 6013 2207
rect 5853 1960 5867 1973
rect 5856 1956 5863 1960
rect 5936 1923 5943 1973
rect 5996 1956 6003 2113
rect 6036 1967 6043 2213
rect 5833 1907 5847 1912
rect 5876 1903 5883 1923
rect 5936 1916 5963 1923
rect 5976 1920 5983 1923
rect 5876 1896 5903 1903
rect 5876 1736 5883 1853
rect 5896 1807 5903 1896
rect 5816 1647 5823 1703
rect 5856 1683 5863 1703
rect 5836 1676 5863 1683
rect 5736 1636 5763 1643
rect 5736 1447 5743 1636
rect 5836 1623 5843 1676
rect 5816 1620 5843 1623
rect 5816 1616 5847 1620
rect 5796 1436 5803 1473
rect 5816 1467 5823 1616
rect 5833 1607 5847 1616
rect 5836 1447 5843 1553
rect 5856 1407 5863 1653
rect 5733 1387 5747 1393
rect 5876 1403 5883 1673
rect 5916 1667 5923 1734
rect 5896 1567 5903 1653
rect 5896 1447 5903 1513
rect 5916 1436 5923 1632
rect 5936 1467 5943 1853
rect 5956 1747 5963 1916
rect 5973 1907 5987 1920
rect 6016 1867 6023 1923
rect 6036 1767 6043 1913
rect 6056 1807 6063 2254
rect 6116 2256 6123 2433
rect 6176 2440 6183 2443
rect 6173 2427 6187 2440
rect 6186 2420 6187 2427
rect 6096 2220 6103 2223
rect 6076 2067 6083 2213
rect 6093 2207 6107 2220
rect 6076 1967 6083 1993
rect 6096 1987 6103 2073
rect 6116 2007 6123 2193
rect 6136 1988 6143 2223
rect 6153 2207 6167 2213
rect 6156 1987 6163 2033
rect 6093 1960 6107 1973
rect 6176 1968 6183 2273
rect 6096 1956 6103 1960
rect 6036 1736 6043 1753
rect 6076 1747 6083 1913
rect 5956 1647 5963 1693
rect 5976 1667 5983 1703
rect 6016 1683 6023 1703
rect 5996 1676 6023 1683
rect 5996 1607 6003 1676
rect 6027 1663 6040 1667
rect 6027 1653 6043 1663
rect 6016 1563 6023 1632
rect 6036 1587 6043 1653
rect 6016 1556 6043 1563
rect 5980 1543 5993 1547
rect 5976 1540 5993 1543
rect 5973 1533 5993 1540
rect 5973 1527 5987 1533
rect 5996 1447 6003 1493
rect 5876 1396 5903 1403
rect 5716 1276 5743 1283
rect 5676 1216 5683 1253
rect 5596 1176 5623 1183
rect 5556 1127 5563 1172
rect 5576 1147 5583 1173
rect 5396 916 5403 993
rect 5436 916 5443 973
rect 5496 887 5503 933
rect 5416 827 5423 872
rect 5376 747 5383 813
rect 5096 587 5103 652
rect 5116 627 5123 693
rect 5147 663 5160 667
rect 5147 656 5163 663
rect 5147 653 5160 656
rect 4947 576 4963 583
rect 4876 416 4903 423
rect 4876 396 4883 416
rect 4956 366 4963 576
rect 5136 447 5143 632
rect 5196 587 5203 663
rect 5256 587 5263 693
rect 5316 567 5323 652
rect 5136 396 5143 433
rect 5273 400 5287 413
rect 5276 396 5283 400
rect 4856 327 4863 363
rect 5056 307 5063 394
rect 5336 366 5343 633
rect 5356 587 5363 663
rect 5396 423 5403 773
rect 5476 727 5483 833
rect 5416 427 5423 713
rect 5473 700 5487 713
rect 5516 708 5523 1013
rect 5536 927 5543 1013
rect 5556 916 5563 993
rect 5596 916 5603 973
rect 5616 967 5623 1176
rect 5656 1047 5663 1183
rect 5696 1176 5723 1183
rect 5620 883 5633 887
rect 5576 827 5583 883
rect 5616 876 5633 883
rect 5620 873 5633 876
rect 5476 696 5483 700
rect 5536 666 5543 753
rect 5556 707 5563 773
rect 5616 747 5623 853
rect 5636 696 5643 813
rect 5656 787 5663 953
rect 5676 707 5683 933
rect 5696 927 5703 1153
rect 5716 1127 5723 1176
rect 5736 1167 5743 1276
rect 5756 1087 5763 1333
rect 5776 1287 5783 1392
rect 5816 1287 5823 1392
rect 5836 1327 5843 1393
rect 5853 1347 5867 1353
rect 5787 1223 5800 1227
rect 5787 1216 5803 1223
rect 5836 1216 5843 1253
rect 5787 1213 5800 1216
rect 5776 1127 5783 1173
rect 5896 1167 5903 1396
rect 5916 1227 5923 1373
rect 5936 1287 5943 1403
rect 5956 1267 5963 1373
rect 5976 1367 5983 1403
rect 5976 1243 5983 1313
rect 5956 1236 5983 1243
rect 5956 1216 5963 1236
rect 5996 1228 6003 1293
rect 6016 1223 6023 1453
rect 6036 1447 6043 1556
rect 6056 1507 6063 1693
rect 6076 1667 6083 1712
rect 6076 1436 6083 1573
rect 6096 1467 6103 1753
rect 6116 1747 6123 1853
rect 6176 1827 6183 1913
rect 6196 1867 6203 2413
rect 6236 2343 6243 2493
rect 6256 2407 6263 2716
rect 6276 2707 6283 2743
rect 6216 2336 6243 2343
rect 6216 2267 6223 2336
rect 6276 2287 6283 2513
rect 6296 2427 6303 2713
rect 6296 2256 6303 2392
rect 6316 2267 6323 2773
rect 6236 2087 6243 2223
rect 6276 2203 6283 2223
rect 6276 2196 6303 2203
rect 6256 1987 6263 2193
rect 6276 1956 6283 2053
rect 6296 1967 6303 2196
rect 6136 1736 6143 1793
rect 6216 1747 6223 1912
rect 6113 1687 6127 1693
rect 6116 1436 6123 1533
rect 6156 1487 6163 1703
rect 6156 1406 6163 1452
rect 6036 1247 6043 1393
rect 6120 1384 6133 1387
rect 6116 1373 6133 1384
rect 6056 1327 6063 1353
rect 6116 1327 6123 1373
rect 6056 1316 6073 1327
rect 6060 1313 6073 1316
rect 6116 1287 6123 1313
rect 6136 1263 6143 1352
rect 6156 1347 6163 1392
rect 6176 1323 6183 1673
rect 6196 1447 6203 1653
rect 6216 1436 6223 1693
rect 6236 1647 6243 1813
rect 6256 1747 6263 1773
rect 6296 1767 6303 1893
rect 6316 1787 6323 2213
rect 6300 1743 6313 1747
rect 6296 1736 6313 1743
rect 6300 1733 6313 1736
rect 6236 1463 6243 1573
rect 6256 1487 6263 1693
rect 6296 1547 6303 1653
rect 6236 1456 6263 1463
rect 6256 1436 6263 1456
rect 6296 1447 6303 1473
rect 6196 1367 6203 1393
rect 6236 1347 6243 1403
rect 6116 1256 6143 1263
rect 6156 1316 6183 1323
rect 6016 1216 6043 1223
rect 5733 920 5747 933
rect 5773 920 5787 933
rect 5736 916 5743 920
rect 5776 916 5783 920
rect 5496 656 5533 663
rect 5553 647 5567 653
rect 5376 416 5403 423
rect 5376 408 5383 416
rect 5416 396 5423 413
rect 5476 367 5483 633
rect 5616 527 5623 663
rect 5656 660 5663 663
rect 5653 647 5667 660
rect 5696 647 5703 873
rect 5716 847 5723 883
rect 5756 880 5763 883
rect 5753 867 5767 880
rect 5816 863 5823 1151
rect 5836 883 5843 1053
rect 5856 927 5863 953
rect 5896 916 5903 1033
rect 5916 967 5923 1173
rect 5936 1167 5943 1183
rect 5936 963 5943 1153
rect 5976 1127 5983 1183
rect 6036 1167 6043 1216
rect 6116 1216 6123 1256
rect 6156 1227 6163 1316
rect 5936 956 5963 963
rect 5956 927 5963 956
rect 5836 876 5883 883
rect 5816 856 5843 863
rect 5716 647 5723 693
rect 5733 663 5747 673
rect 5733 660 5763 663
rect 5736 656 5763 660
rect 5836 643 5843 856
rect 5856 767 5863 876
rect 5916 827 5923 883
rect 5876 707 5883 813
rect 5956 807 5963 873
rect 5976 867 5983 914
rect 5976 783 5983 832
rect 5996 827 6003 1013
rect 6056 1007 6063 1173
rect 6076 916 6083 1153
rect 6096 1127 6103 1183
rect 6136 967 6143 1183
rect 6113 920 6127 933
rect 6116 916 6123 920
rect 5956 776 5983 783
rect 5893 727 5907 733
rect 5927 714 5933 727
rect 5920 713 5933 714
rect 5816 636 5843 643
rect 5856 696 5873 703
rect 5516 396 5523 493
rect 5696 396 5703 473
rect 5716 427 5723 633
rect 5756 407 5763 453
rect 5116 327 5123 363
rect 4636 176 4643 213
rect 4716 176 4723 213
rect 4576 107 4583 132
rect 4616 107 4623 143
rect 4736 107 4743 143
rect 4776 140 4783 143
rect 4773 127 4787 140
rect 4816 107 4823 253
rect 4916 176 4923 233
rect 5036 176 5043 233
rect 5076 176 5083 293
rect 5176 176 5183 233
rect 5216 207 5223 363
rect 5316 360 5333 363
rect 5313 356 5333 360
rect 5313 347 5327 356
rect 5396 360 5403 363
rect 5393 347 5407 360
rect 5216 176 5263 183
rect 4836 47 4843 173
rect 5056 140 5063 143
rect 5053 127 5067 140
rect 5116 87 5123 173
rect 5196 140 5203 143
rect 5193 127 5207 140
rect 5256 127 5263 176
rect 5376 176 5383 333
rect 5276 47 5283 174
rect 5356 140 5363 143
rect 5316 87 5323 132
rect 5353 127 5367 140
rect 5333 103 5347 113
rect 5333 100 5393 103
rect 5336 96 5393 100
rect 5416 67 5423 293
rect 5436 267 5443 363
rect 5536 176 5543 293
rect 5576 267 5583 363
rect 5636 307 5643 394
rect 5776 387 5783 633
rect 5760 366 5780 367
rect 5767 353 5773 366
rect 5796 327 5803 413
rect 5816 407 5823 636
rect 5856 428 5863 696
rect 5956 696 5963 776
rect 5896 443 5903 652
rect 5936 627 5943 663
rect 5896 436 5923 443
rect 5893 400 5907 413
rect 5916 407 5923 436
rect 5896 396 5903 400
rect 5656 176 5663 313
rect 5816 303 5823 353
rect 5796 296 5823 303
rect 5676 267 5683 293
rect 5716 176 5763 183
rect 5796 176 5803 296
rect 5836 247 5843 363
rect 5876 327 5883 363
rect 5936 203 5943 493
rect 6016 467 6023 872
rect 6156 867 6163 1173
rect 6176 1147 6183 1253
rect 6016 427 6023 453
rect 6036 403 6043 853
rect 6176 847 6183 933
rect 6196 927 6203 1253
rect 6216 1227 6223 1273
rect 6256 1243 6263 1353
rect 6276 1287 6283 1403
rect 6296 1267 6303 1393
rect 6256 1236 6283 1243
rect 6276 1216 6283 1236
rect 6316 1227 6323 1693
rect 6216 928 6223 1173
rect 6236 947 6243 1153
rect 6256 1147 6263 1183
rect 6296 1087 6303 1183
rect 6316 1023 6323 1153
rect 6296 1016 6323 1023
rect 6256 916 6263 1013
rect 6296 927 6303 1016
rect 6316 887 6323 993
rect 6076 696 6083 753
rect 6136 696 6143 773
rect 6116 587 6123 663
rect 6176 627 6183 663
rect 6196 507 6203 873
rect 6053 403 6067 413
rect 6036 400 6067 403
rect 6036 396 6063 400
rect 6076 367 6083 413
rect 6133 400 6147 413
rect 6136 396 6143 400
rect 5976 307 5983 363
rect 6016 287 6023 363
rect 5916 196 5943 203
rect 5916 176 5923 196
rect 5953 180 5967 193
rect 5956 176 5963 180
rect 5476 140 5483 143
rect 5516 140 5523 143
rect 5453 127 5467 133
rect 5473 127 5487 140
rect 5513 127 5527 140
rect 5596 107 5603 153
rect 5636 140 5643 143
rect 5633 127 5647 140
rect 5716 127 5723 176
rect 6036 146 6043 333
rect 6096 176 6103 273
rect 6136 176 6143 313
rect 6156 287 6163 363
rect 6216 227 6223 853
rect 6236 847 6243 883
rect 6236 188 6243 413
rect 6256 327 6263 813
rect 5500 106 5520 107
rect 5507 93 5513 106
rect 5816 67 5823 143
rect 5936 47 5943 143
rect 5976 107 5983 143
rect 6176 67 6183 174
rect 6276 47 6283 713
rect 6296 107 6303 853
rect 2876 16 2913 23
rect 3407 16 3433 23
<< m3contact >>
rect 1693 6253 1707 6267
rect 1793 6253 1807 6267
rect 1633 6213 1647 6227
rect 1473 6193 1487 6207
rect 113 6173 127 6187
rect 713 6173 727 6187
rect 373 6153 387 6167
rect 653 6153 667 6167
rect 353 6114 367 6128
rect 93 5933 107 5947
rect 133 5894 147 5908
rect 173 5894 187 5908
rect 273 6033 287 6047
rect 253 5894 267 5908
rect 153 5853 167 5867
rect 233 5852 247 5866
rect 273 5813 287 5827
rect 153 5793 167 5807
rect 313 5852 327 5866
rect 293 5773 307 5787
rect 113 5594 127 5608
rect 193 5594 207 5608
rect 133 5552 147 5566
rect 273 5594 287 5608
rect 313 5593 327 5607
rect 153 5533 167 5547
rect 213 5533 227 5547
rect 93 5513 107 5527
rect 193 5512 207 5526
rect 113 5433 127 5447
rect 153 5433 167 5447
rect 13 5374 27 5388
rect 153 5374 167 5388
rect 93 5313 107 5327
rect 193 5332 207 5346
rect 33 5074 47 5088
rect 93 5074 107 5088
rect 133 5074 147 5088
rect 53 5032 67 5046
rect 33 4993 47 5007
rect 33 4933 47 4947
rect 13 4753 27 4767
rect 13 4653 27 4667
rect 113 5032 127 5046
rect 153 5033 167 5047
rect 113 4993 127 5007
rect 153 4854 167 4868
rect 313 5553 327 5567
rect 293 5533 307 5547
rect 413 6114 427 6128
rect 453 6114 467 6128
rect 513 6114 527 6128
rect 553 6114 567 6128
rect 373 6033 387 6047
rect 353 6013 367 6027
rect 452 6013 466 6027
rect 473 6013 487 6027
rect 433 5933 447 5947
rect 373 5894 387 5908
rect 353 5853 367 5867
rect 393 5852 407 5866
rect 433 5813 447 5827
rect 353 5793 367 5807
rect 673 6133 687 6147
rect 653 6093 667 6107
rect 573 6072 587 6086
rect 593 6053 607 6067
rect 593 6013 607 6027
rect 813 6153 827 6167
rect 1233 6153 1247 6167
rect 753 6133 767 6147
rect 713 6114 727 6128
rect 913 6114 927 6128
rect 953 6114 967 6128
rect 993 6114 1007 6128
rect 1053 6114 1067 6128
rect 1093 6114 1107 6128
rect 1133 6114 1147 6128
rect 1353 6133 1367 6147
rect 1433 6133 1447 6147
rect 1273 6114 1287 6128
rect 813 6093 827 6107
rect 733 6033 747 6047
rect 633 5993 647 6007
rect 673 5993 687 6007
rect 713 5993 727 6007
rect 613 5953 627 5967
rect 573 5933 587 5947
rect 673 5894 687 5908
rect 533 5852 547 5866
rect 573 5853 587 5867
rect 493 5813 507 5827
rect 493 5773 507 5787
rect 693 5853 707 5867
rect 933 6072 947 6086
rect 973 6072 987 6086
rect 913 6053 927 6067
rect 873 6033 887 6047
rect 933 6032 947 6046
rect 1113 6072 1127 6086
rect 1293 6072 1307 6086
rect 1253 6053 1267 6067
rect 1053 6033 1067 6047
rect 1013 6013 1027 6027
rect 1393 6114 1407 6128
rect 1513 6114 1527 6128
rect 1553 6114 1567 6128
rect 1613 6114 1627 6128
rect 1373 6072 1387 6086
rect 1413 6072 1427 6086
rect 1473 6073 1487 6087
rect 1353 6013 1367 6027
rect 1713 6193 1727 6207
rect 1673 6153 1687 6167
rect 1613 6053 1627 6067
rect 1533 6013 1547 6027
rect 1613 6013 1627 6027
rect 933 5993 947 6007
rect 1333 5993 1347 6007
rect 1373 5993 1387 6007
rect 1593 5993 1607 6007
rect 853 5973 867 5987
rect 893 5973 907 5987
rect 773 5894 787 5908
rect 833 5893 847 5907
rect 993 5953 1007 5967
rect 1313 5953 1327 5967
rect 1453 5953 1467 5967
rect 1493 5953 1507 5967
rect 653 5733 667 5747
rect 393 5713 407 5727
rect 453 5713 467 5727
rect 613 5713 627 5727
rect 353 5673 367 5687
rect 733 5813 747 5827
rect 493 5673 507 5687
rect 693 5673 707 5687
rect 433 5633 447 5647
rect 593 5633 607 5647
rect 513 5594 527 5608
rect 553 5594 567 5608
rect 593 5594 607 5608
rect 653 5594 667 5608
rect 793 5793 807 5807
rect 1113 5933 1127 5947
rect 1033 5913 1047 5927
rect 1073 5913 1087 5927
rect 1053 5894 1067 5908
rect 1173 5894 1187 5908
rect 1253 5893 1267 5907
rect 1473 5933 1487 5947
rect 1533 5933 1547 5947
rect 1373 5893 1387 5907
rect 1433 5894 1447 5908
rect 873 5852 887 5866
rect 993 5852 1007 5866
rect 1033 5852 1047 5866
rect 1073 5852 1087 5866
rect 1113 5852 1127 5866
rect 833 5833 847 5847
rect 913 5833 927 5847
rect 1053 5833 1067 5847
rect 1033 5813 1047 5827
rect 733 5594 747 5608
rect 773 5594 787 5608
rect 1193 5852 1207 5866
rect 1253 5852 1267 5866
rect 1293 5852 1307 5866
rect 1333 5852 1347 5866
rect 1733 6072 1747 6086
rect 1713 5953 1727 5967
rect 1753 5953 1767 5967
rect 1733 5933 1747 5947
rect 1733 5894 1747 5908
rect 1153 5813 1167 5827
rect 1053 5773 1067 5787
rect 1033 5733 1047 5747
rect 493 5573 507 5587
rect 413 5552 427 5566
rect 353 5533 367 5547
rect 253 5493 267 5507
rect 313 5493 327 5507
rect 313 5413 327 5427
rect 273 5393 287 5407
rect 273 5374 287 5388
rect 253 5332 267 5346
rect 453 5513 467 5527
rect 573 5533 587 5547
rect 533 5513 547 5527
rect 473 5453 487 5467
rect 373 5413 387 5427
rect 393 5374 407 5388
rect 513 5374 527 5388
rect 373 5332 387 5346
rect 313 5313 327 5327
rect 353 5313 367 5327
rect 233 5273 247 5287
rect 293 5273 307 5287
rect 253 4953 267 4967
rect 233 4893 247 4907
rect 213 4854 227 4868
rect 53 4793 67 4807
rect 133 4793 147 4807
rect 93 4773 107 4787
rect 53 4713 67 4727
rect 33 4493 47 4507
rect 13 4333 27 4347
rect 73 4613 87 4627
rect 93 4593 107 4607
rect 73 4554 87 4568
rect 113 4512 127 4526
rect 73 4493 87 4507
rect 13 3853 27 3867
rect 53 4034 67 4048
rect 153 4593 167 4607
rect 153 4513 167 4527
rect 133 4413 147 4427
rect 93 4334 107 4348
rect 133 4213 147 4227
rect 133 4173 147 4187
rect 213 4813 227 4827
rect 413 5332 427 5346
rect 393 5273 407 5287
rect 333 5133 347 5147
rect 553 5473 567 5487
rect 593 5393 607 5407
rect 713 5552 727 5566
rect 653 5473 667 5487
rect 753 5453 767 5467
rect 813 5594 827 5608
rect 853 5594 867 5608
rect 993 5594 1007 5608
rect 833 5552 847 5566
rect 1373 5833 1387 5847
rect 1533 5852 1547 5866
rect 1573 5852 1587 5866
rect 1453 5833 1467 5847
rect 1473 5813 1487 5827
rect 1473 5773 1487 5787
rect 1713 5813 1727 5827
rect 1833 6213 1847 6227
rect 1913 6173 1927 6187
rect 1873 6114 1887 6128
rect 1973 6114 1987 6128
rect 1853 6072 1867 6086
rect 1913 6072 1927 6086
rect 1993 6013 2007 6027
rect 1973 5953 1987 5967
rect 2013 5953 2027 5967
rect 1853 5894 1867 5908
rect 1613 5753 1627 5767
rect 1753 5753 1767 5767
rect 1793 5753 1807 5767
rect 1333 5673 1347 5687
rect 1313 5633 1327 5647
rect 1053 5593 1067 5607
rect 1273 5594 1287 5608
rect 793 5513 807 5527
rect 873 5513 887 5527
rect 973 5513 987 5527
rect 633 5413 647 5427
rect 773 5413 787 5427
rect 713 5374 727 5388
rect 753 5374 767 5388
rect 853 5413 867 5427
rect 913 5393 927 5407
rect 973 5374 987 5388
rect 813 5332 827 5346
rect 853 5332 867 5346
rect 1193 5553 1207 5567
rect 1113 5513 1127 5527
rect 1173 5433 1187 5447
rect 1053 5413 1067 5427
rect 1113 5413 1127 5427
rect 1073 5374 1087 5388
rect 553 5273 567 5287
rect 613 5273 627 5287
rect 533 5113 547 5127
rect 593 5113 607 5127
rect 333 5074 347 5088
rect 373 5074 387 5088
rect 413 5074 427 5088
rect 453 5074 467 5088
rect 513 5074 527 5088
rect 553 5074 567 5088
rect 293 4873 307 4887
rect 253 4812 267 4826
rect 233 4773 247 4787
rect 393 5032 407 5046
rect 353 4993 367 5007
rect 373 4973 387 4987
rect 433 4893 447 4907
rect 573 5033 587 5047
rect 513 5013 527 5027
rect 553 5013 567 5027
rect 493 4953 507 4967
rect 393 4854 407 4868
rect 473 4854 487 4868
rect 513 4854 527 4868
rect 593 5013 607 5027
rect 573 4973 587 4987
rect 653 5313 667 5327
rect 713 5313 727 5327
rect 753 5313 767 5327
rect 633 5253 647 5267
rect 733 5253 747 5267
rect 633 5153 647 5167
rect 693 5113 707 5127
rect 653 5074 667 5088
rect 733 5073 747 5087
rect 713 5032 727 5046
rect 613 4953 627 4967
rect 593 4854 607 4868
rect 533 4812 547 4826
rect 433 4773 447 4787
rect 473 4773 487 4787
rect 413 4753 427 4767
rect 353 4713 367 4727
rect 313 4653 327 4667
rect 213 4593 227 4607
rect 293 4593 307 4607
rect 193 4513 207 4527
rect 233 4512 247 4526
rect 333 4512 347 4526
rect 373 4473 387 4487
rect 393 4453 407 4467
rect 273 4393 287 4407
rect 193 4253 207 4267
rect 213 4113 227 4127
rect 173 4073 187 4087
rect 93 4034 107 4048
rect 153 4033 167 4047
rect 113 3992 127 4006
rect 73 3933 87 3947
rect 153 3933 167 3947
rect 53 3814 67 3828
rect 113 3814 127 3828
rect 33 3772 47 3786
rect 33 3633 47 3647
rect 13 3553 27 3567
rect 13 3333 27 3347
rect 13 3252 27 3266
rect 293 4273 307 4287
rect 333 4413 347 4427
rect 513 4753 527 4767
rect 573 4753 587 4767
rect 473 4733 487 4747
rect 493 4673 507 4687
rect 473 4593 487 4607
rect 1013 5333 1027 5347
rect 1193 5393 1207 5407
rect 1233 5393 1247 5407
rect 1093 5332 1107 5346
rect 1133 5332 1147 5346
rect 1173 5332 1187 5346
rect 1053 5313 1067 5327
rect 773 5293 787 5307
rect 893 5293 907 5307
rect 1053 5273 1067 5287
rect 913 5193 927 5207
rect 893 5173 907 5187
rect 833 5153 847 5167
rect 773 5113 787 5127
rect 793 5093 807 5107
rect 793 5074 807 5088
rect 893 5133 907 5147
rect 813 5032 827 5046
rect 853 5032 867 5046
rect 773 5013 787 5027
rect 733 4933 747 4947
rect 713 4854 727 4868
rect 753 4854 767 4868
rect 793 4953 807 4967
rect 873 4933 887 4947
rect 953 5113 967 5127
rect 1033 5113 1047 5127
rect 993 5074 1007 5088
rect 933 5032 947 5046
rect 973 5032 987 5046
rect 793 4893 807 4907
rect 833 4893 847 4907
rect 893 4893 907 4907
rect 2073 6114 2087 6128
rect 2353 6193 2367 6207
rect 2273 6114 2287 6128
rect 2333 6093 2347 6107
rect 2553 6094 2567 6108
rect 2713 6134 2727 6148
rect 2753 6134 2767 6148
rect 2153 6072 2167 6086
rect 2253 6072 2267 6086
rect 2313 6073 2327 6087
rect 2073 5953 2087 5967
rect 2193 5953 2207 5967
rect 2053 5933 2067 5947
rect 2073 5894 2087 5908
rect 2113 5894 2127 5908
rect 2153 5894 2167 5908
rect 1993 5852 2007 5866
rect 2073 5853 2087 5867
rect 1933 5813 1947 5827
rect 1433 5633 1447 5647
rect 1813 5633 1827 5647
rect 1873 5633 1887 5647
rect 1973 5633 1987 5647
rect 2133 5633 2147 5647
rect 1393 5594 1407 5608
rect 1553 5594 1567 5608
rect 1633 5593 1647 5607
rect 1753 5594 1767 5608
rect 1813 5594 1827 5608
rect 1873 5594 1887 5608
rect 1373 5552 1387 5566
rect 1413 5552 1427 5566
rect 1333 5513 1347 5527
rect 1633 5552 1647 5566
rect 1693 5513 1707 5527
rect 1773 5513 1787 5527
rect 1953 5593 1967 5607
rect 1893 5533 1907 5547
rect 2013 5552 2027 5566
rect 1973 5533 1987 5547
rect 1853 5513 1867 5527
rect 1953 5513 1967 5527
rect 1573 5433 1587 5447
rect 1813 5433 1827 5447
rect 1273 5374 1287 5388
rect 1333 5374 1347 5388
rect 1373 5374 1387 5388
rect 1413 5374 1427 5388
rect 1533 5374 1547 5388
rect 1633 5374 1647 5388
rect 1673 5374 1687 5388
rect 1853 5374 1867 5388
rect 2133 5594 2147 5608
rect 2172 5594 2186 5608
rect 2253 5933 2267 5947
rect 2293 5894 2307 5908
rect 2233 5852 2247 5866
rect 2273 5852 2287 5866
rect 2653 6073 2667 6087
rect 2453 5993 2467 6007
rect 2413 5894 2427 5908
rect 2593 5973 2607 5987
rect 2533 5913 2547 5927
rect 2513 5894 2527 5908
rect 2353 5852 2367 5866
rect 2393 5852 2407 5866
rect 2433 5852 2447 5866
rect 2253 5813 2267 5827
rect 2333 5813 2347 5827
rect 2233 5773 2247 5787
rect 2213 5753 2227 5767
rect 2253 5753 2267 5767
rect 2213 5693 2227 5707
rect 2193 5593 2207 5607
rect 2053 5513 2067 5527
rect 2153 5473 2167 5487
rect 2153 5413 2167 5427
rect 2093 5374 2107 5388
rect 1293 5332 1307 5346
rect 1333 5333 1347 5347
rect 1253 5273 1267 5287
rect 1433 5332 1447 5346
rect 1533 5293 1547 5307
rect 1393 5273 1407 5287
rect 1293 5133 1307 5147
rect 1353 5133 1367 5147
rect 1113 5074 1127 5088
rect 1153 5074 1167 5088
rect 1193 5074 1207 5088
rect 1173 5033 1187 5047
rect 1033 5013 1047 5027
rect 1093 5013 1107 5027
rect 1133 5013 1147 5027
rect 1073 4953 1087 4967
rect 793 4853 807 4867
rect 833 4854 847 4868
rect 873 4854 887 4868
rect 933 4854 947 4868
rect 673 4813 687 4827
rect 573 4713 587 4727
rect 653 4713 667 4727
rect 533 4613 547 4627
rect 553 4554 567 4568
rect 613 4633 627 4647
rect 633 4573 647 4587
rect 733 4812 747 4826
rect 693 4773 707 4787
rect 693 4673 707 4687
rect 433 4513 447 4527
rect 573 4513 587 4527
rect 553 4433 567 4447
rect 493 4413 507 4427
rect 413 4373 427 4387
rect 453 4373 467 4387
rect 333 4193 347 4207
rect 533 4413 547 4427
rect 693 4553 707 4567
rect 653 4512 667 4526
rect 773 4773 787 4787
rect 753 4733 767 4747
rect 733 4693 747 4707
rect 613 4473 627 4487
rect 593 4433 607 4447
rect 593 4393 607 4407
rect 573 4373 587 4387
rect 593 4333 607 4347
rect 493 4292 507 4306
rect 432 4253 446 4267
rect 453 4253 467 4267
rect 393 4213 407 4227
rect 313 4173 327 4187
rect 373 4173 387 4187
rect 473 4233 487 4247
rect 593 4293 607 4307
rect 533 4213 547 4227
rect 493 4193 507 4207
rect 533 4173 547 4187
rect 493 4133 507 4147
rect 412 4113 426 4127
rect 433 4113 447 4127
rect 393 4073 407 4087
rect 253 4033 267 4047
rect 313 4013 327 4027
rect 233 3992 247 4006
rect 273 3953 287 3967
rect 173 3853 187 3867
rect 213 3814 227 3828
rect 313 3953 327 3967
rect 293 3933 307 3947
rect 473 4073 487 4087
rect 453 3993 467 4007
rect 413 3933 427 3947
rect 373 3913 387 3927
rect 433 3893 447 3907
rect 393 3853 407 3867
rect 353 3833 367 3847
rect 93 3772 107 3786
rect 153 3773 167 3787
rect 193 3772 207 3786
rect 133 3533 147 3547
rect 53 3513 67 3527
rect 93 3514 107 3528
rect 53 3373 67 3387
rect 153 3433 167 3447
rect 252 3773 266 3787
rect 273 3773 287 3787
rect 233 3753 247 3767
rect 633 4453 647 4467
rect 753 4613 767 4627
rect 853 4812 867 4826
rect 913 4812 927 4826
rect 953 4812 967 4826
rect 933 4793 947 4807
rect 893 4773 907 4787
rect 893 4713 907 4727
rect 833 4693 847 4707
rect 793 4673 807 4687
rect 993 4793 1007 4807
rect 973 4673 987 4687
rect 873 4633 887 4647
rect 913 4633 927 4647
rect 953 4633 967 4647
rect 853 4593 867 4607
rect 793 4573 807 4587
rect 853 4553 867 4567
rect 733 4413 747 4427
rect 833 4512 847 4526
rect 813 4373 827 4387
rect 893 4553 907 4567
rect 873 4473 887 4487
rect 853 4353 867 4367
rect 633 4292 647 4306
rect 673 4292 687 4306
rect 773 4292 787 4306
rect 713 4213 727 4227
rect 773 4213 787 4227
rect 1273 5093 1287 5107
rect 1273 5074 1287 5088
rect 1313 5074 1327 5088
rect 1213 5032 1227 5046
rect 1253 5032 1267 5046
rect 1233 4973 1247 4987
rect 1293 4973 1307 4987
rect 1193 4953 1207 4967
rect 1153 4893 1167 4907
rect 1193 4854 1207 4868
rect 1173 4812 1187 4826
rect 1093 4753 1107 4767
rect 1153 4753 1167 4767
rect 1013 4653 1027 4667
rect 1053 4653 1067 4667
rect 993 4633 1007 4647
rect 973 4573 987 4587
rect 933 4554 947 4568
rect 953 4433 967 4447
rect 993 4393 1007 4407
rect 933 4353 947 4367
rect 993 4353 1007 4367
rect 913 4313 927 4327
rect 833 4292 847 4306
rect 873 4292 887 4306
rect 853 4253 867 4267
rect 613 4173 627 4187
rect 713 4113 727 4127
rect 633 4073 647 4087
rect 553 4053 567 4067
rect 533 4034 547 4048
rect 593 4032 607 4046
rect 673 4034 687 4048
rect 833 4173 847 4187
rect 813 4153 827 4167
rect 813 4113 827 4127
rect 773 4053 787 4067
rect 793 4034 807 4048
rect 553 3973 567 3987
rect 513 3913 527 3927
rect 613 3973 627 3987
rect 592 3893 606 3907
rect 613 3893 627 3907
rect 673 3973 687 3987
rect 573 3873 587 3887
rect 653 3873 667 3887
rect 553 3853 567 3867
rect 513 3833 527 3847
rect 432 3813 446 3827
rect 373 3772 387 3786
rect 413 3772 427 3786
rect 293 3753 307 3767
rect 413 3713 427 3727
rect 433 3633 447 3647
rect 313 3613 327 3627
rect 213 3513 227 3527
rect 253 3514 267 3528
rect 273 3453 287 3467
rect 213 3433 227 3447
rect 193 3373 207 3387
rect 133 3333 147 3347
rect 333 3593 347 3607
rect 313 3413 327 3427
rect 253 3353 267 3367
rect 213 3314 227 3328
rect 173 3293 187 3307
rect 213 3293 227 3307
rect 313 3313 327 3327
rect 113 3193 127 3207
rect 53 3113 67 3127
rect 33 3093 47 3107
rect 133 3093 147 3107
rect 33 3053 47 3067
rect 13 3033 27 3047
rect 13 2953 27 2967
rect 13 2913 27 2927
rect 13 2773 27 2787
rect 93 3013 107 3027
rect 233 3233 247 3247
rect 313 3233 327 3247
rect 313 3212 327 3226
rect 273 3053 287 3067
rect 173 3013 187 3027
rect 273 3013 287 3027
rect 133 2994 147 3008
rect 193 2994 207 3008
rect 233 2994 247 3008
rect 473 3814 487 3828
rect 553 3832 567 3846
rect 593 3853 607 3867
rect 493 3753 507 3767
rect 573 3772 587 3786
rect 533 3693 547 3707
rect 493 3633 507 3647
rect 453 3573 467 3587
rect 433 3533 447 3547
rect 373 3514 387 3528
rect 353 3473 367 3487
rect 393 3453 407 3467
rect 413 3433 427 3447
rect 393 3294 407 3308
rect 533 3573 547 3587
rect 493 3533 507 3547
rect 633 3814 647 3828
rect 693 3953 707 3967
rect 713 3913 727 3927
rect 713 3853 727 3867
rect 593 3713 607 3727
rect 653 3772 667 3786
rect 753 3973 767 3987
rect 1053 4613 1067 4627
rect 1033 4573 1047 4587
rect 953 4292 967 4306
rect 933 4213 947 4227
rect 913 4153 927 4167
rect 993 4253 1007 4267
rect 973 4073 987 4087
rect 893 4034 907 4048
rect 913 3992 927 4006
rect 953 3992 967 4006
rect 853 3973 867 3987
rect 773 3953 787 3967
rect 833 3953 847 3967
rect 773 3873 787 3887
rect 753 3813 767 3827
rect 833 3814 847 3828
rect 753 3773 767 3787
rect 733 3753 747 3767
rect 713 3673 727 3687
rect 693 3633 707 3647
rect 673 3613 687 3627
rect 613 3553 627 3567
rect 553 3472 567 3486
rect 513 3433 527 3447
rect 453 3373 467 3387
rect 373 3252 387 3266
rect 413 3213 427 3227
rect 533 3353 547 3367
rect 553 3313 567 3327
rect 573 3294 587 3308
rect 633 3514 647 3528
rect 713 3573 727 3587
rect 713 3552 727 3566
rect 693 3453 707 3467
rect 673 3413 687 3427
rect 673 3373 687 3387
rect 633 3353 647 3367
rect 453 3193 467 3207
rect 493 3253 507 3267
rect 493 3193 507 3207
rect 473 3173 487 3187
rect 453 3153 467 3167
rect 433 3133 447 3147
rect 373 3053 387 3067
rect 333 3013 347 3027
rect 573 3233 587 3247
rect 513 3073 527 3087
rect 513 3052 527 3066
rect 493 3033 507 3047
rect 393 2994 407 3008
rect 73 2952 87 2966
rect 113 2952 127 2966
rect 193 2953 207 2967
rect 173 2913 187 2927
rect 113 2774 127 2788
rect 313 2953 327 2967
rect 373 2952 387 2966
rect 333 2893 347 2907
rect 393 2893 407 2907
rect 253 2873 267 2887
rect 273 2813 287 2827
rect 213 2774 227 2788
rect 153 2732 167 2746
rect 313 2773 327 2787
rect 453 2994 467 3008
rect 633 3293 647 3307
rect 932 3814 946 3828
rect 1053 4553 1067 4567
rect 1093 4554 1107 4568
rect 1133 4554 1147 4568
rect 1053 4513 1067 4527
rect 1033 4233 1047 4247
rect 1113 4513 1127 4527
rect 1073 4473 1087 4487
rect 1093 4433 1107 4447
rect 1133 4493 1147 4507
rect 1133 4393 1147 4407
rect 1213 4733 1227 4747
rect 1193 4713 1207 4727
rect 1173 4673 1187 4687
rect 1193 4653 1207 4667
rect 1273 4953 1287 4967
rect 1313 4854 1327 4868
rect 1433 5093 1447 5107
rect 1373 5074 1387 5088
rect 1473 5074 1487 5088
rect 1513 5074 1527 5088
rect 1373 5033 1387 5047
rect 1413 5032 1427 5046
rect 1393 4933 1407 4947
rect 1373 4893 1387 4907
rect 1353 4853 1367 4867
rect 1353 4813 1367 4827
rect 1333 4773 1347 4787
rect 1253 4753 1267 4767
rect 1233 4693 1247 4707
rect 1333 4713 1347 4727
rect 1253 4653 1267 4667
rect 1313 4653 1327 4667
rect 1253 4632 1267 4646
rect 1213 4613 1227 4627
rect 1193 4593 1207 4607
rect 1313 4612 1327 4626
rect 1273 4593 1287 4607
rect 1193 4493 1207 4507
rect 1173 4453 1187 4467
rect 1113 4373 1127 4387
rect 1073 4333 1087 4347
rect 1193 4413 1207 4427
rect 1213 4373 1227 4387
rect 1253 4373 1267 4387
rect 1233 4333 1247 4347
rect 1053 4153 1067 4167
rect 1013 4073 1027 4087
rect 1013 4033 1027 4047
rect 1233 4312 1247 4326
rect 1093 4233 1107 4247
rect 1153 4292 1167 4306
rect 1453 4993 1467 5007
rect 1513 4973 1527 4987
rect 1593 5332 1607 5346
rect 1553 5153 1567 5167
rect 1693 5332 1707 5346
rect 1793 5332 1807 5346
rect 1753 5273 1767 5287
rect 1673 5253 1687 5267
rect 1633 5113 1647 5127
rect 1573 5074 1587 5088
rect 1613 5074 1627 5088
rect 1593 5032 1607 5046
rect 1633 4993 1647 5007
rect 1633 4953 1647 4967
rect 1533 4933 1547 4947
rect 1413 4873 1427 4887
rect 1493 4893 1507 4907
rect 1593 4893 1607 4907
rect 1473 4873 1487 4887
rect 1533 4854 1547 4868
rect 1633 4854 1647 4868
rect 1333 4554 1347 4568
rect 1373 4554 1387 4568
rect 1413 4554 1427 4568
rect 1513 4812 1527 4826
rect 1453 4593 1467 4607
rect 1453 4554 1467 4568
rect 1273 4333 1287 4347
rect 1393 4453 1407 4467
rect 1353 4433 1367 4447
rect 1353 4334 1367 4348
rect 1333 4292 1347 4306
rect 1253 4273 1267 4287
rect 1293 4273 1307 4287
rect 1113 4213 1127 4227
rect 1333 4173 1347 4187
rect 1373 4173 1387 4187
rect 1253 4153 1267 4167
rect 1233 4133 1247 4147
rect 1133 4053 1147 4067
rect 1073 4034 1087 4048
rect 1113 4034 1127 4048
rect 1193 4053 1207 4067
rect 1153 4034 1167 4048
rect 1053 3992 1067 4006
rect 1112 3993 1126 4007
rect 1133 3993 1147 4007
rect 1053 3953 1067 3967
rect 1093 3953 1107 3967
rect 953 3813 967 3827
rect 1013 3913 1027 3927
rect 1033 3893 1047 3907
rect 1013 3873 1027 3887
rect 993 3853 1007 3867
rect 853 3772 867 3786
rect 833 3753 847 3767
rect 773 3713 787 3727
rect 753 3593 767 3607
rect 1013 3833 1027 3847
rect 1093 3814 1107 3828
rect 993 3772 1007 3786
rect 913 3733 927 3747
rect 933 3713 947 3727
rect 913 3693 927 3707
rect 833 3673 847 3687
rect 873 3673 887 3687
rect 793 3633 807 3647
rect 773 3553 787 3567
rect 833 3593 847 3607
rect 853 3514 867 3528
rect 913 3593 927 3607
rect 993 3593 1007 3607
rect 973 3553 987 3567
rect 733 3353 747 3367
rect 713 3294 727 3308
rect 833 3472 847 3486
rect 913 3514 927 3528
rect 953 3514 967 3528
rect 853 3453 867 3467
rect 773 3413 787 3427
rect 893 3472 907 3486
rect 873 3433 887 3447
rect 913 3433 927 3447
rect 793 3353 807 3367
rect 853 3353 867 3367
rect 653 3252 667 3266
rect 613 3153 627 3167
rect 633 3073 647 3087
rect 573 2993 587 3007
rect 453 2953 467 2967
rect 493 2952 507 2966
rect 533 2952 547 2966
rect 573 2953 587 2967
rect 573 2873 587 2887
rect 733 3133 747 3147
rect 713 3113 727 3127
rect 713 3073 727 3087
rect 693 3053 707 3067
rect 673 3013 687 3027
rect 653 2952 667 2966
rect 693 2933 707 2947
rect 693 2893 707 2907
rect 633 2873 647 2887
rect 593 2853 607 2867
rect 433 2773 447 2787
rect 513 2774 527 2788
rect 573 2773 587 2787
rect 633 2774 647 2788
rect 213 2713 227 2727
rect 253 2713 267 2727
rect 33 2593 47 2607
rect 193 2573 207 2587
rect 33 2513 47 2527
rect 113 2432 127 2446
rect 73 2393 87 2407
rect 133 2313 147 2327
rect 373 2732 387 2746
rect 413 2732 427 2746
rect 973 3472 987 3486
rect 933 3413 947 3427
rect 933 3392 947 3406
rect 893 3313 907 3327
rect 853 3294 867 3308
rect 833 3252 847 3266
rect 913 3253 927 3267
rect 793 3233 807 3247
rect 833 3213 847 3227
rect 793 3193 807 3207
rect 913 3213 927 3227
rect 873 3173 887 3187
rect 913 3153 927 3167
rect 773 3093 787 3107
rect 873 3093 887 3107
rect 793 3013 807 3027
rect 793 2994 807 3008
rect 833 2994 847 3008
rect 913 3053 927 3067
rect 913 2994 927 3008
rect 753 2973 767 2987
rect 853 2952 867 2966
rect 813 2873 827 2887
rect 853 2853 867 2867
rect 733 2833 747 2847
rect 713 2774 727 2788
rect 773 2774 787 2788
rect 813 2774 827 2788
rect 613 2732 627 2746
rect 493 2693 507 2707
rect 353 2613 367 2627
rect 313 2513 327 2527
rect 253 2474 267 2488
rect 413 2573 427 2587
rect 353 2474 367 2488
rect 453 2474 467 2488
rect 193 2453 207 2467
rect 273 2353 287 2367
rect 273 2293 287 2307
rect 313 2293 327 2307
rect 133 2254 147 2268
rect 173 2254 187 2268
rect 153 2193 167 2207
rect 93 1993 107 2007
rect 113 1954 127 1968
rect 153 1913 167 1927
rect 133 1893 147 1907
rect 93 1873 107 1887
rect 273 2254 287 2268
rect 193 2212 207 2226
rect 253 2212 267 2226
rect 293 2212 307 2226
rect 253 2191 267 2205
rect 193 1993 207 2007
rect 173 1893 187 1907
rect 293 2113 307 2127
rect 473 2433 487 2447
rect 433 2413 447 2427
rect 393 2393 407 2407
rect 373 2293 387 2307
rect 453 2293 467 2307
rect 372 2253 386 2267
rect 393 2254 407 2268
rect 413 2212 427 2226
rect 353 2033 367 2047
rect 693 2732 707 2746
rect 713 2653 727 2667
rect 773 2653 787 2667
rect 653 2613 667 2627
rect 653 2513 667 2527
rect 593 2474 607 2488
rect 513 2413 527 2427
rect 553 2353 567 2367
rect 533 2313 547 2327
rect 513 2273 527 2287
rect 493 2253 507 2267
rect 593 2273 607 2287
rect 473 2213 487 2227
rect 753 2613 767 2627
rect 713 2474 727 2488
rect 993 3413 1007 3427
rect 1033 3772 1047 3786
rect 1113 3773 1127 3787
rect 1073 3713 1087 3727
rect 1073 3573 1087 3587
rect 1033 3553 1047 3567
rect 1173 3992 1187 4006
rect 1213 3953 1227 3967
rect 1213 3913 1227 3927
rect 1153 3853 1167 3867
rect 1133 3673 1147 3687
rect 1133 3533 1147 3547
rect 1113 3513 1127 3527
rect 1013 3393 1027 3407
rect 973 3373 987 3387
rect 972 3293 986 3307
rect 993 3294 1007 3308
rect 1053 3472 1067 3486
rect 1073 3433 1087 3447
rect 1053 3413 1067 3427
rect 1033 3293 1047 3307
rect 1033 3253 1047 3267
rect 1013 3233 1027 3247
rect 973 3173 987 3187
rect 1033 3093 1047 3107
rect 1013 3013 1027 3027
rect 973 2994 987 3008
rect 1113 3473 1127 3487
rect 1093 3353 1107 3367
rect 1093 3313 1107 3327
rect 1213 3833 1227 3847
rect 1273 4034 1287 4048
rect 1393 4153 1407 4167
rect 1573 4812 1587 4826
rect 1573 4773 1587 4787
rect 1512 4753 1526 4767
rect 1533 4753 1547 4767
rect 1553 4733 1567 4747
rect 1533 4613 1547 4627
rect 1513 4554 1527 4568
rect 1573 4693 1587 4707
rect 1473 4513 1487 4527
rect 1533 4512 1547 4526
rect 1453 4473 1467 4487
rect 1613 4613 1627 4627
rect 1693 5233 1707 5247
rect 1693 5193 1707 5207
rect 1833 5193 1847 5207
rect 1873 5193 1887 5207
rect 1953 5193 1967 5207
rect 1753 5173 1767 5187
rect 1853 5153 1867 5167
rect 1713 5113 1727 5127
rect 1693 5074 1707 5088
rect 1733 5074 1747 5088
rect 1713 5033 1727 5047
rect 1832 5032 1846 5046
rect 1853 5033 1867 5047
rect 1933 5113 1947 5127
rect 1973 5074 1987 5088
rect 2113 5332 2127 5346
rect 2233 5633 2247 5647
rect 2293 5594 2307 5608
rect 2253 5533 2267 5547
rect 2233 5453 2247 5467
rect 2233 5432 2247 5446
rect 2233 5393 2247 5407
rect 2173 5374 2187 5388
rect 2213 5374 2227 5388
rect 2312 5552 2326 5566
rect 2333 5553 2347 5567
rect 2273 5513 2287 5527
rect 2273 5473 2287 5487
rect 2253 5373 2267 5387
rect 2173 5333 2187 5347
rect 2473 5833 2487 5847
rect 2493 5773 2507 5787
rect 2453 5713 2467 5727
rect 2373 5594 2387 5608
rect 2413 5594 2427 5608
rect 2493 5593 2507 5607
rect 2373 5553 2387 5567
rect 2373 5493 2387 5507
rect 2353 5473 2367 5487
rect 2373 5374 2387 5388
rect 2413 5374 2427 5388
rect 2153 5293 2167 5307
rect 2013 5173 2027 5187
rect 1913 5032 1927 5046
rect 1793 4993 1807 5007
rect 1873 4993 1887 5007
rect 1833 4953 1847 4967
rect 1893 4953 1907 4967
rect 1773 4913 1787 4927
rect 1993 5013 2007 5027
rect 1973 4993 1987 5007
rect 1953 4913 1967 4927
rect 1873 4893 1887 4907
rect 1853 4873 1867 4887
rect 1833 4833 1847 4847
rect 1673 4733 1687 4747
rect 1633 4593 1647 4607
rect 1613 4554 1627 4568
rect 1673 4554 1687 4568
rect 1733 4733 1747 4747
rect 1633 4493 1647 4507
rect 1533 4453 1547 4467
rect 1593 4453 1607 4467
rect 1473 4353 1487 4367
rect 1433 4293 1447 4307
rect 1673 4493 1687 4507
rect 1653 4473 1667 4487
rect 1593 4334 1607 4348
rect 1633 4334 1647 4348
rect 1453 4273 1467 4287
rect 1533 4292 1547 4306
rect 1573 4292 1587 4306
rect 1653 4293 1667 4307
rect 1433 4233 1447 4247
rect 1413 4133 1427 4147
rect 1393 4113 1407 4127
rect 1472 4253 1486 4267
rect 1493 4253 1507 4267
rect 1613 4253 1627 4267
rect 1453 4193 1467 4207
rect 1473 4173 1487 4187
rect 1553 4133 1567 4147
rect 1373 4052 1387 4066
rect 1373 4034 1387 4048
rect 1273 3993 1287 4007
rect 1353 3992 1367 4006
rect 1473 4073 1487 4087
rect 1513 4073 1527 4087
rect 1433 4034 1447 4048
rect 1473 4034 1487 4048
rect 1573 4053 1587 4067
rect 1613 4053 1627 4067
rect 1313 3973 1327 3987
rect 1293 3953 1307 3967
rect 1273 3833 1287 3847
rect 1433 3993 1447 4007
rect 1333 3953 1347 3967
rect 1393 3953 1407 3967
rect 1453 3953 1467 3967
rect 1313 3812 1327 3826
rect 1413 3913 1427 3927
rect 1413 3873 1427 3887
rect 1373 3814 1387 3828
rect 1533 3992 1547 4006
rect 1753 4653 1767 4667
rect 1773 4593 1787 4607
rect 1753 4553 1767 4567
rect 1893 4872 1907 4886
rect 1873 4853 1887 4867
rect 1953 4853 1967 4867
rect 1853 4673 1867 4687
rect 1833 4553 1847 4567
rect 1733 4493 1747 4507
rect 1713 4473 1727 4487
rect 1713 4413 1727 4427
rect 1733 4393 1747 4407
rect 1873 4532 1887 4546
rect 1793 4512 1807 4526
rect 1853 4513 1867 4527
rect 1813 4493 1827 4507
rect 1793 4433 1807 4447
rect 1753 4373 1767 4387
rect 1793 4373 1807 4387
rect 1693 4293 1707 4307
rect 1753 4273 1767 4287
rect 1713 4253 1727 4267
rect 1733 4073 1747 4087
rect 1673 4053 1687 4067
rect 1693 4034 1707 4048
rect 1733 4034 1747 4048
rect 1513 3873 1527 3887
rect 1493 3813 1507 3827
rect 1573 3992 1587 4006
rect 1693 3973 1707 3987
rect 1633 3953 1647 3967
rect 1673 3933 1687 3947
rect 1573 3893 1587 3907
rect 1593 3873 1607 3887
rect 1552 3853 1566 3867
rect 1573 3853 1587 3867
rect 1273 3772 1287 3786
rect 1312 3772 1326 3786
rect 1333 3773 1347 3787
rect 1293 3753 1307 3767
rect 1193 3713 1207 3727
rect 1252 3713 1266 3727
rect 1273 3713 1287 3727
rect 1193 3613 1207 3627
rect 1233 3593 1247 3607
rect 1193 3533 1207 3547
rect 1153 3513 1167 3527
rect 1293 3693 1307 3707
rect 1393 3772 1407 3786
rect 1473 3772 1487 3786
rect 1533 3772 1547 3786
rect 1353 3613 1367 3627
rect 1313 3593 1327 3607
rect 1353 3573 1367 3587
rect 1433 3733 1447 3747
rect 1493 3733 1507 3747
rect 1473 3713 1487 3727
rect 1533 3713 1547 3727
rect 1493 3692 1507 3706
rect 1413 3673 1427 3687
rect 1393 3633 1407 3647
rect 1373 3553 1387 3567
rect 1553 3673 1567 3687
rect 1493 3533 1507 3547
rect 1533 3533 1547 3547
rect 1393 3513 1407 3527
rect 1213 3472 1227 3486
rect 1273 3473 1287 3487
rect 1193 3453 1207 3467
rect 1173 3373 1187 3387
rect 1133 3353 1147 3367
rect 1133 3294 1147 3308
rect 1173 3293 1187 3307
rect 1233 3433 1247 3447
rect 1373 3472 1387 3486
rect 1513 3513 1527 3527
rect 1473 3472 1487 3486
rect 1513 3473 1527 3487
rect 1333 3433 1347 3447
rect 1413 3433 1427 3447
rect 1253 3413 1267 3427
rect 1273 3393 1287 3407
rect 1413 3393 1427 3407
rect 1213 3353 1227 3367
rect 1413 3353 1427 3367
rect 1273 3333 1287 3347
rect 1353 3333 1367 3347
rect 1213 3313 1227 3327
rect 1073 3253 1087 3267
rect 1053 2973 1067 2987
rect 993 2952 1007 2966
rect 933 2933 947 2947
rect 973 2933 987 2947
rect 893 2813 907 2827
rect 953 2793 967 2807
rect 1192 3253 1206 3267
rect 1313 3294 1327 3308
rect 1213 3252 1227 3266
rect 1253 3252 1267 3266
rect 1173 3213 1187 3227
rect 1153 3173 1167 3187
rect 1173 3153 1187 3167
rect 1253 3153 1267 3167
rect 1193 3113 1207 3127
rect 1113 3033 1127 3047
rect 1113 2994 1127 3008
rect 1173 2993 1187 3007
rect 1133 2952 1147 2966
rect 1173 2952 1187 2966
rect 1433 3333 1447 3347
rect 1453 3294 1467 3308
rect 1673 3773 1687 3787
rect 1653 3633 1667 3647
rect 1573 3613 1587 3627
rect 1573 3513 1587 3527
rect 1613 3514 1627 3528
rect 1593 3472 1607 3486
rect 1533 3313 1547 3327
rect 1473 3252 1487 3266
rect 1513 3253 1527 3267
rect 1433 3193 1447 3207
rect 1673 3473 1687 3487
rect 1673 3413 1687 3427
rect 1633 3353 1647 3367
rect 1673 3353 1687 3367
rect 1573 3294 1587 3308
rect 1633 3294 1647 3308
rect 1673 3273 1687 3287
rect 1593 3252 1607 3266
rect 1653 3213 1667 3227
rect 1553 3173 1567 3187
rect 1373 3133 1387 3147
rect 1513 3133 1527 3147
rect 1613 3133 1627 3147
rect 1313 3113 1327 3127
rect 1353 3113 1367 3127
rect 1593 3113 1607 3127
rect 1492 3093 1506 3107
rect 1513 3093 1527 3107
rect 1372 3053 1386 3067
rect 1393 3053 1407 3067
rect 1313 3033 1327 3047
rect 1353 2994 1367 3008
rect 1513 3033 1527 3047
rect 1433 2994 1447 3008
rect 1472 2994 1486 3008
rect 1493 2994 1507 3008
rect 1533 2994 1547 3008
rect 1573 2994 1587 3008
rect 1613 3093 1627 3107
rect 1613 2994 1627 3008
rect 1233 2952 1247 2966
rect 1313 2952 1327 2966
rect 1373 2952 1387 2966
rect 1473 2953 1487 2967
rect 1513 2952 1527 2966
rect 1553 2952 1567 2966
rect 1593 2952 1607 2966
rect 1433 2933 1447 2947
rect 1193 2913 1207 2927
rect 1413 2913 1427 2927
rect 1173 2893 1187 2907
rect 1073 2873 1087 2887
rect 1213 2873 1227 2887
rect 1293 2873 1307 2887
rect 1053 2813 1067 2827
rect 1173 2813 1187 2827
rect 1033 2793 1047 2807
rect 1093 2793 1107 2807
rect 1013 2773 1027 2787
rect 853 2673 867 2687
rect 793 2613 807 2627
rect 773 2473 787 2487
rect 733 2432 747 2446
rect 773 2432 787 2446
rect 833 2432 847 2446
rect 973 2713 987 2727
rect 1033 2713 1047 2727
rect 933 2474 947 2488
rect 693 2393 707 2407
rect 693 2313 707 2327
rect 513 2212 527 2226
rect 593 2212 607 2226
rect 633 2173 647 2187
rect 553 2053 567 2067
rect 513 2013 527 2027
rect 833 2393 847 2407
rect 813 2254 827 2268
rect 853 2254 867 2268
rect 753 2212 767 2226
rect 953 2432 967 2446
rect 1073 2693 1087 2707
rect 1253 2733 1267 2747
rect 1233 2713 1247 2727
rect 1193 2673 1207 2687
rect 1093 2653 1107 2667
rect 1073 2474 1087 2488
rect 1033 2433 1047 2447
rect 1093 2432 1107 2446
rect 933 2393 947 2407
rect 1013 2393 1027 2407
rect 993 2313 1007 2327
rect 1253 2573 1267 2587
rect 1213 2474 1227 2488
rect 1413 2833 1427 2847
rect 1333 2774 1347 2788
rect 1413 2774 1427 2788
rect 1392 2733 1406 2747
rect 1413 2733 1427 2747
rect 1393 2693 1407 2707
rect 1373 2653 1387 2667
rect 1353 2613 1367 2627
rect 1333 2593 1347 2607
rect 1373 2593 1387 2607
rect 1353 2553 1367 2567
rect 1333 2533 1347 2547
rect 1313 2513 1327 2527
rect 1293 2333 1307 2347
rect 1193 2313 1207 2327
rect 1253 2313 1267 2327
rect 1113 2273 1127 2287
rect 1153 2273 1167 2287
rect 1013 2254 1027 2268
rect 1073 2254 1087 2268
rect 1293 2273 1307 2287
rect 853 2193 867 2207
rect 793 2173 807 2187
rect 833 2113 847 2127
rect 773 2013 787 2027
rect 693 1993 707 2007
rect 753 1993 767 2007
rect 293 1954 307 1968
rect 333 1954 347 1968
rect 373 1954 387 1968
rect 413 1954 427 1968
rect 473 1954 487 1968
rect 213 1913 227 1927
rect 193 1873 207 1887
rect 153 1853 167 1867
rect 153 1753 167 1767
rect 193 1753 207 1767
rect 53 1734 67 1748
rect 113 1734 127 1748
rect 193 1732 207 1746
rect 393 1912 407 1926
rect 533 1954 547 1968
rect 633 1954 647 1968
rect 713 1954 727 1968
rect 373 1893 387 1907
rect 233 1853 247 1867
rect 273 1853 287 1867
rect 333 1853 347 1867
rect 333 1773 347 1787
rect 233 1734 247 1748
rect 273 1734 287 1748
rect 53 1653 67 1667
rect 133 1692 147 1706
rect 73 1633 87 1647
rect 33 1593 47 1607
rect 433 1813 447 1827
rect 373 1753 387 1767
rect 353 1733 367 1747
rect 413 1734 427 1748
rect 493 1912 507 1926
rect 513 1893 527 1907
rect 493 1773 507 1787
rect 253 1692 267 1706
rect 293 1692 307 1706
rect 333 1692 347 1706
rect 193 1613 207 1627
rect 273 1613 287 1627
rect 233 1573 247 1587
rect 193 1533 207 1547
rect 93 1392 107 1406
rect 233 1434 247 1448
rect 333 1493 347 1507
rect 373 1693 387 1707
rect 433 1692 447 1706
rect 493 1693 507 1707
rect 393 1653 407 1667
rect 433 1653 447 1667
rect 373 1633 387 1647
rect 433 1613 447 1627
rect 353 1473 367 1487
rect 413 1473 427 1487
rect 373 1434 387 1448
rect 213 1392 227 1406
rect 273 1393 287 1407
rect 153 1233 167 1247
rect 213 1233 227 1247
rect 33 1214 47 1228
rect 113 1214 127 1228
rect 173 1213 187 1227
rect 93 1113 107 1127
rect 133 1073 147 1087
rect 53 914 67 928
rect 93 914 107 928
rect 133 914 147 928
rect 113 872 127 886
rect 53 813 67 827
rect 313 1214 327 1228
rect 473 1593 487 1607
rect 433 1433 447 1447
rect 553 1853 567 1867
rect 593 1853 607 1867
rect 633 1912 647 1926
rect 613 1773 627 1787
rect 573 1753 587 1767
rect 533 1692 547 1706
rect 593 1692 607 1706
rect 593 1573 607 1587
rect 513 1493 527 1507
rect 593 1473 607 1487
rect 653 1893 667 1907
rect 793 1954 807 1968
rect 993 2212 1007 2226
rect 1153 2252 1167 2266
rect 1193 2254 1207 2268
rect 1233 2254 1247 2268
rect 973 2193 987 2207
rect 913 2153 927 2167
rect 973 2113 987 2127
rect 913 2093 927 2107
rect 893 2053 907 2067
rect 873 2013 887 2027
rect 993 2033 1007 2047
rect 993 1953 1007 1967
rect 693 1873 707 1887
rect 753 1873 767 1887
rect 653 1833 667 1847
rect 753 1833 767 1847
rect 713 1793 727 1807
rect 653 1753 667 1767
rect 693 1753 707 1767
rect 813 1912 827 1926
rect 913 1913 927 1927
rect 853 1873 867 1887
rect 793 1793 807 1807
rect 752 1734 766 1748
rect 773 1734 787 1748
rect 653 1692 667 1706
rect 693 1692 707 1706
rect 813 1733 827 1747
rect 872 1734 886 1748
rect 953 1912 967 1926
rect 1053 2212 1067 2226
rect 1033 2153 1047 2167
rect 1093 1954 1107 1968
rect 1033 1913 1047 1927
rect 1013 1893 1027 1907
rect 933 1873 947 1887
rect 913 1753 927 1767
rect 893 1733 907 1747
rect 793 1653 807 1667
rect 733 1573 747 1587
rect 633 1533 647 1547
rect 673 1533 687 1547
rect 513 1434 527 1448
rect 553 1434 567 1448
rect 633 1434 647 1448
rect 453 1392 467 1406
rect 453 1253 467 1267
rect 413 1233 427 1247
rect 353 1214 367 1228
rect 253 1172 267 1186
rect 293 1172 307 1186
rect 353 1173 367 1187
rect 273 1053 287 1067
rect 253 1033 267 1047
rect 233 973 247 987
rect 213 914 227 928
rect 253 914 267 928
rect 353 1113 367 1127
rect 333 913 347 927
rect 373 1073 387 1087
rect 273 872 287 886
rect 313 853 327 867
rect 193 813 207 827
rect 253 733 267 747
rect 133 694 147 708
rect 173 693 187 707
rect 273 694 287 708
rect 33 653 47 667
rect 73 652 87 666
rect 353 873 367 887
rect 333 753 347 767
rect 393 1053 407 1067
rect 553 1393 567 1407
rect 613 1392 627 1406
rect 593 1333 607 1347
rect 513 1214 527 1228
rect 553 1214 567 1228
rect 733 1473 747 1487
rect 833 1693 847 1707
rect 893 1693 907 1707
rect 833 1613 847 1627
rect 813 1453 827 1467
rect 1113 1893 1127 1907
rect 1073 1853 1087 1867
rect 973 1813 987 1827
rect 1033 1793 1047 1807
rect 993 1692 1007 1706
rect 1253 2212 1267 2226
rect 1293 2212 1307 2226
rect 1213 2153 1227 2167
rect 1293 2153 1307 2167
rect 1153 2013 1167 2027
rect 1133 1793 1147 1807
rect 1213 1954 1227 1968
rect 1253 1954 1267 1968
rect 1193 1912 1207 1926
rect 1273 1913 1287 1927
rect 1253 1853 1267 1867
rect 1193 1813 1207 1827
rect 1233 1813 1247 1827
rect 1293 1892 1307 1906
rect 1273 1793 1287 1807
rect 1232 1753 1246 1767
rect 1253 1753 1267 1767
rect 1093 1692 1107 1706
rect 993 1653 1007 1667
rect 1033 1653 1047 1667
rect 1133 1653 1147 1667
rect 933 1573 947 1587
rect 773 1434 787 1448
rect 833 1434 847 1448
rect 873 1434 887 1448
rect 913 1434 927 1448
rect 673 1373 687 1387
rect 973 1433 987 1447
rect 833 1333 847 1347
rect 753 1313 767 1327
rect 813 1313 827 1327
rect 693 1273 707 1287
rect 653 1253 667 1267
rect 613 1233 627 1247
rect 493 1113 507 1127
rect 433 1033 447 1047
rect 573 1172 587 1186
rect 633 1173 647 1187
rect 733 1253 747 1267
rect 793 1253 807 1267
rect 693 1214 707 1228
rect 613 1153 627 1167
rect 653 1153 667 1167
rect 573 1113 587 1127
rect 533 1073 547 1087
rect 513 973 527 987
rect 753 1153 767 1167
rect 713 1113 727 1127
rect 613 993 627 1007
rect 653 993 667 1007
rect 473 914 487 928
rect 633 933 647 947
rect 333 713 347 727
rect 373 713 387 727
rect 213 652 227 666
rect 313 652 327 666
rect 253 613 267 627
rect 113 553 127 567
rect 273 473 287 487
rect 153 394 167 408
rect 113 333 127 347
rect 213 333 227 347
rect 293 353 307 367
rect 253 313 267 327
rect 153 253 167 267
rect 113 174 127 188
rect 193 174 207 188
rect 253 174 267 188
rect 453 872 467 886
rect 413 813 427 827
rect 593 813 607 827
rect 453 733 467 747
rect 533 733 547 747
rect 593 733 607 747
rect 433 694 447 708
rect 473 694 487 708
rect 373 652 387 666
rect 593 693 607 707
rect 473 613 487 627
rect 453 573 467 587
rect 413 553 427 567
rect 333 473 347 487
rect 393 433 407 447
rect 353 394 367 408
rect 393 394 407 408
rect 313 333 327 347
rect 333 313 347 327
rect 413 352 427 366
rect 433 313 447 327
rect 373 293 387 307
rect 393 273 407 287
rect 353 173 367 187
rect 613 653 627 667
rect 593 593 607 607
rect 513 553 527 567
rect 513 493 527 507
rect 473 473 487 487
rect 613 533 627 547
rect 513 394 527 408
rect 553 394 567 408
rect 713 973 727 987
rect 933 1392 947 1406
rect 953 1333 967 1347
rect 913 1313 927 1327
rect 893 1233 907 1247
rect 873 1214 887 1228
rect 1153 1613 1167 1627
rect 1073 1533 1087 1547
rect 1033 1453 1047 1467
rect 1113 1473 1127 1487
rect 993 1393 1007 1407
rect 1013 1273 1027 1287
rect 973 1214 987 1228
rect 1193 1733 1207 1747
rect 1273 1734 1287 1748
rect 1213 1692 1227 1706
rect 1253 1692 1267 1706
rect 1293 1693 1307 1707
rect 1233 1653 1247 1667
rect 1173 1593 1187 1607
rect 1213 1593 1227 1607
rect 1133 1373 1147 1387
rect 1113 1333 1127 1347
rect 1073 1253 1087 1267
rect 1053 1233 1067 1247
rect 1093 1233 1107 1247
rect 853 1172 867 1186
rect 893 1172 907 1186
rect 953 1172 967 1186
rect 993 1153 1007 1167
rect 1053 1153 1067 1167
rect 853 1133 867 1147
rect 933 1133 947 1147
rect 1033 1133 1047 1147
rect 813 1073 827 1087
rect 793 1013 807 1027
rect 833 973 847 987
rect 753 953 767 967
rect 793 953 807 967
rect 753 914 767 928
rect 733 872 747 886
rect 713 813 727 827
rect 693 773 707 787
rect 653 693 667 707
rect 733 753 747 767
rect 773 694 787 708
rect 873 953 887 967
rect 833 914 847 928
rect 953 1073 967 1087
rect 853 872 867 886
rect 893 872 907 886
rect 933 873 947 887
rect 933 753 947 767
rect 753 633 767 647
rect 693 613 707 627
rect 833 694 847 708
rect 813 652 827 666
rect 773 593 787 607
rect 893 633 907 647
rect 773 553 787 567
rect 813 553 827 567
rect 873 553 887 567
rect 693 433 707 447
rect 633 394 647 408
rect 733 394 747 408
rect 493 353 507 367
rect 573 352 587 366
rect 613 353 627 367
rect 493 313 507 327
rect 473 293 487 307
rect 453 273 467 287
rect 513 253 527 267
rect 433 174 447 188
rect 93 113 107 127
rect 193 133 207 147
rect 233 132 247 146
rect 273 132 287 146
rect 333 133 347 147
rect 173 113 187 127
rect 233 93 247 107
rect 453 132 467 146
rect 613 233 627 247
rect 573 174 587 188
rect 873 493 887 507
rect 853 473 867 487
rect 832 433 846 447
rect 853 433 867 447
rect 713 352 727 366
rect 773 353 787 367
rect 793 333 807 347
rect 633 174 647 188
rect 673 293 687 307
rect 753 193 767 207
rect 713 174 727 188
rect 853 352 867 366
rect 813 293 827 307
rect 1013 1053 1027 1067
rect 973 933 987 947
rect 1013 933 1027 947
rect 1033 914 1047 928
rect 993 872 1007 886
rect 1053 873 1067 887
rect 1173 1313 1187 1327
rect 1173 1253 1187 1267
rect 1133 1213 1147 1227
rect 1173 1214 1187 1228
rect 1153 1153 1167 1167
rect 1213 1173 1227 1187
rect 1173 1053 1187 1067
rect 1153 933 1167 947
rect 1113 914 1127 928
rect 1293 1653 1307 1667
rect 1353 2474 1367 2488
rect 1393 2474 1407 2488
rect 1513 2913 1527 2927
rect 1453 2893 1467 2907
rect 1473 2774 1487 2788
rect 1533 2873 1547 2887
rect 1533 2833 1547 2847
rect 1773 4233 1787 4247
rect 1813 4173 1827 4187
rect 1873 4493 1887 4507
rect 1873 4453 1887 4467
rect 1913 4733 1927 4747
rect 1933 4673 1947 4687
rect 2032 5074 2046 5088
rect 2273 5332 2287 5346
rect 2313 5332 2327 5346
rect 2353 5253 2367 5267
rect 2393 5173 2407 5187
rect 2293 5133 2307 5147
rect 2373 5133 2387 5147
rect 2053 5073 2067 5087
rect 2133 5074 2147 5088
rect 2173 5074 2187 5088
rect 2253 5074 2267 5088
rect 2033 5033 2047 5047
rect 2073 5032 2087 5046
rect 2173 5033 2187 5047
rect 2233 5032 2247 5046
rect 2153 4993 2167 5007
rect 2113 4953 2127 4967
rect 2153 4953 2167 4967
rect 2133 4933 2147 4947
rect 2053 4913 2067 4927
rect 2113 4913 2127 4927
rect 2013 4893 2027 4907
rect 1973 4773 1987 4787
rect 1953 4593 1967 4607
rect 2093 4853 2107 4867
rect 2013 4813 2027 4827
rect 1993 4453 2007 4467
rect 1973 4433 1987 4447
rect 1913 4373 1927 4387
rect 1913 4334 1927 4348
rect 1853 4273 1867 4287
rect 1893 4273 1907 4287
rect 1833 4133 1847 4147
rect 1793 4034 1807 4048
rect 1773 3993 1787 4007
rect 1753 3973 1767 3987
rect 1733 3933 1747 3947
rect 1733 3893 1747 3907
rect 1833 3972 1847 3986
rect 1913 4253 1927 4267
rect 1873 4213 1887 4227
rect 1873 4173 1887 4187
rect 1873 4133 1887 4147
rect 1953 4293 1967 4307
rect 1933 4233 1947 4247
rect 1933 4034 1947 4048
rect 1993 4373 2007 4387
rect 1973 4113 1987 4127
rect 2033 4673 2047 4687
rect 2053 4593 2067 4607
rect 2033 4573 2047 4587
rect 2093 4753 2107 4767
rect 2193 4893 2207 4907
rect 2133 4873 2147 4887
rect 2333 5032 2347 5046
rect 2393 5032 2407 5046
rect 2313 4973 2327 4987
rect 2253 4913 2267 4927
rect 2293 4913 2307 4927
rect 2133 4813 2147 4827
rect 2173 4812 2187 4826
rect 2213 4812 2227 4826
rect 2273 4893 2287 4907
rect 2273 4853 2287 4867
rect 2353 4913 2367 4927
rect 2353 4873 2367 4887
rect 2193 4773 2207 4787
rect 2253 4773 2267 4787
rect 2193 4752 2207 4766
rect 2293 4812 2307 4826
rect 2113 4733 2127 4747
rect 2093 4673 2107 4687
rect 2033 4512 2047 4526
rect 2073 4512 2087 4526
rect 2113 4512 2127 4526
rect 2093 4473 2107 4487
rect 2133 4453 2147 4467
rect 2193 4533 2207 4547
rect 2153 4433 2167 4447
rect 2333 4753 2347 4767
rect 2533 5853 2547 5867
rect 2713 6013 2727 6027
rect 3333 6253 3347 6267
rect 3673 6253 3687 6267
rect 2953 6193 2967 6207
rect 2893 6093 2907 6107
rect 2753 5993 2767 6007
rect 2853 6013 2867 6027
rect 2833 5973 2847 5987
rect 2753 5894 2767 5908
rect 2813 5894 2827 5908
rect 2933 6093 2947 6107
rect 2913 5973 2927 5987
rect 2853 5893 2867 5907
rect 2573 5833 2587 5847
rect 2653 5833 2667 5847
rect 2733 5833 2747 5847
rect 2693 5813 2707 5827
rect 2733 5793 2747 5807
rect 2733 5753 2747 5767
rect 2633 5653 2647 5667
rect 2713 5653 2727 5667
rect 2573 5594 2587 5608
rect 2653 5613 2667 5627
rect 2633 5573 2647 5587
rect 2553 5552 2567 5566
rect 2473 5533 2487 5547
rect 2513 5533 2527 5547
rect 2493 5453 2507 5467
rect 2533 5453 2547 5467
rect 2453 5293 2467 5307
rect 2553 5333 2567 5347
rect 2533 5313 2547 5327
rect 2513 5233 2527 5247
rect 2473 5113 2487 5127
rect 2473 5074 2487 5088
rect 2413 4913 2427 4927
rect 2493 5032 2507 5046
rect 2653 5512 2667 5526
rect 2593 5493 2607 5507
rect 2633 5493 2647 5507
rect 2653 5413 2667 5427
rect 2633 5393 2647 5407
rect 2733 5552 2747 5566
rect 2893 5833 2907 5847
rect 2893 5753 2907 5767
rect 2873 5733 2887 5747
rect 2853 5713 2867 5727
rect 2953 5693 2967 5707
rect 2933 5673 2947 5687
rect 2893 5613 2907 5627
rect 2913 5594 2927 5608
rect 2733 5513 2747 5527
rect 2713 5433 2727 5447
rect 2693 5373 2707 5387
rect 2593 5173 2607 5187
rect 2773 5374 2787 5388
rect 2853 5552 2867 5566
rect 2893 5552 2907 5566
rect 2933 5553 2947 5567
rect 2713 5313 2727 5327
rect 2793 5253 2807 5267
rect 2753 5193 2767 5207
rect 2693 5133 2707 5147
rect 2553 5073 2567 5087
rect 2593 5074 2607 5088
rect 2653 5072 2667 5086
rect 2813 5233 2827 5247
rect 2933 5393 2947 5407
rect 2873 5373 2887 5387
rect 2993 6094 3007 6108
rect 3153 6094 3167 6108
rect 3313 6134 3327 6148
rect 3373 6134 3387 6148
rect 3293 6093 3307 6107
rect 3533 6094 3547 6108
rect 3273 6073 3287 6087
rect 3033 5993 3047 6007
rect 2993 5933 3007 5947
rect 3873 6133 3887 6147
rect 3713 6073 3727 6087
rect 3833 6094 3847 6108
rect 3393 6053 3407 6067
rect 3673 6053 3687 6067
rect 3773 6053 3787 6067
rect 3293 5993 3307 6007
rect 3213 5973 3227 5987
rect 3273 5973 3287 5987
rect 3093 5933 3107 5947
rect 3133 5894 3147 5908
rect 3173 5894 3187 5908
rect 3113 5833 3127 5847
rect 3333 5953 3347 5967
rect 3313 5933 3327 5947
rect 3313 5894 3327 5908
rect 3373 5894 3387 5908
rect 3133 5813 3147 5827
rect 3073 5793 3087 5807
rect 2973 5633 2987 5647
rect 3033 5594 3047 5608
rect 2973 5552 2987 5566
rect 3013 5552 3027 5566
rect 3053 5513 3067 5527
rect 3033 5493 3047 5507
rect 2973 5473 2987 5487
rect 3013 5473 3027 5487
rect 2973 5413 2987 5427
rect 2973 5354 2987 5368
rect 2873 5293 2887 5307
rect 2933 5313 2947 5327
rect 2913 5253 2927 5267
rect 2953 5253 2967 5267
rect 2933 5233 2947 5247
rect 2853 5173 2867 5187
rect 2873 5153 2887 5167
rect 2813 5133 2827 5147
rect 2773 5093 2787 5107
rect 2533 5013 2547 5027
rect 2453 4933 2467 4947
rect 2493 4913 2507 4927
rect 2533 4893 2547 4907
rect 2413 4853 2427 4867
rect 2493 4873 2507 4887
rect 2473 4854 2487 4868
rect 2453 4812 2467 4826
rect 2493 4812 2507 4826
rect 2633 5012 2647 5026
rect 2593 4913 2607 4927
rect 2552 4853 2566 4867
rect 2573 4853 2587 4867
rect 2713 5032 2727 5046
rect 2833 5074 2847 5088
rect 2912 5073 2926 5087
rect 2933 5074 2947 5088
rect 3133 5773 3147 5787
rect 3093 5753 3107 5767
rect 3093 5693 3107 5707
rect 3233 5852 3247 5866
rect 3293 5852 3307 5866
rect 3353 5833 3367 5847
rect 3313 5813 3327 5827
rect 3193 5733 3207 5747
rect 3253 5633 3267 5647
rect 3193 5594 3207 5608
rect 3093 5552 3107 5566
rect 3153 5552 3167 5566
rect 3193 5553 3207 5567
rect 3173 5533 3187 5547
rect 3073 5473 3087 5487
rect 3273 5533 3287 5547
rect 3253 5493 3267 5507
rect 3273 5473 3287 5487
rect 3053 5453 3067 5467
rect 3093 5453 3107 5467
rect 3173 5453 3187 5467
rect 3253 5453 3267 5467
rect 3073 5393 3087 5407
rect 3073 5354 3087 5368
rect 3053 5273 3067 5287
rect 3013 5213 3027 5227
rect 2793 5033 2807 5047
rect 2853 5013 2867 5027
rect 2713 4973 2727 4987
rect 2773 4973 2787 4987
rect 2873 4973 2887 4987
rect 2693 4913 2707 4927
rect 2653 4812 2667 4826
rect 2553 4793 2567 4807
rect 2612 4793 2626 4807
rect 2633 4793 2647 4807
rect 2613 4753 2627 4767
rect 2453 4733 2467 4747
rect 2533 4733 2547 4747
rect 2393 4633 2407 4647
rect 2493 4633 2507 4647
rect 2393 4553 2407 4567
rect 2253 4433 2267 4447
rect 2293 4433 2307 4447
rect 2473 4433 2487 4447
rect 2213 4413 2227 4427
rect 2433 4413 2447 4427
rect 2013 4353 2027 4367
rect 2093 4353 2107 4367
rect 2133 4353 2147 4367
rect 2033 4334 2047 4348
rect 2013 4292 2027 4306
rect 2052 4292 2066 4306
rect 2073 4293 2087 4307
rect 2073 4233 2087 4247
rect 2153 4334 2167 4348
rect 2133 4253 2147 4267
rect 2053 4153 2067 4167
rect 2093 4153 2107 4167
rect 2093 4113 2107 4127
rect 1873 3993 1887 4007
rect 1953 3993 1967 4007
rect 1913 3973 1927 3987
rect 1893 3933 1907 3947
rect 1853 3893 1867 3907
rect 1833 3853 1847 3867
rect 1813 3813 1827 3827
rect 1713 3773 1727 3787
rect 1753 3693 1767 3707
rect 1833 3772 1847 3786
rect 1793 3593 1807 3607
rect 1713 3513 1727 3527
rect 1753 3514 1767 3528
rect 1813 3533 1827 3547
rect 1713 3433 1727 3447
rect 1753 3453 1767 3467
rect 1753 3393 1767 3407
rect 1733 3353 1747 3367
rect 1753 3313 1767 3327
rect 1793 3453 1807 3467
rect 1733 3252 1747 3266
rect 1713 3233 1727 3247
rect 1693 3213 1707 3227
rect 1673 3093 1687 3107
rect 1673 3053 1687 3067
rect 1673 3013 1687 3027
rect 1653 2993 1667 3007
rect 1733 2994 1747 3008
rect 1773 2994 1787 3008
rect 1673 2952 1687 2966
rect 1713 2952 1727 2966
rect 1773 2933 1787 2947
rect 1653 2913 1667 2927
rect 1713 2913 1727 2927
rect 1593 2773 1607 2787
rect 1453 2733 1467 2747
rect 1493 2732 1507 2746
rect 1633 2732 1647 2746
rect 1693 2733 1707 2747
rect 1493 2553 1507 2567
rect 1893 3833 1907 3847
rect 1993 3973 2007 3987
rect 1973 3873 1987 3887
rect 2153 4093 2167 4107
rect 2113 4053 2127 4067
rect 2193 4293 2207 4307
rect 2393 4314 2407 4328
rect 2233 4253 2247 4267
rect 2193 4233 2207 4247
rect 2193 4173 2207 4187
rect 2173 4073 2187 4087
rect 2253 4113 2267 4127
rect 2233 4093 2247 4107
rect 2113 3933 2127 3947
rect 2093 3913 2107 3927
rect 1853 3653 1867 3667
rect 1893 3772 1907 3786
rect 1913 3713 1927 3727
rect 2033 3853 2047 3867
rect 2073 3853 2087 3867
rect 1993 3814 2007 3828
rect 2033 3814 2047 3828
rect 2073 3813 2087 3827
rect 2093 3794 2107 3808
rect 2173 3992 2187 4006
rect 2153 3973 2167 3987
rect 2213 3973 2227 3987
rect 2153 3933 2167 3947
rect 1993 3733 2007 3747
rect 1973 3713 1987 3727
rect 1933 3693 1947 3707
rect 2073 3773 2087 3787
rect 1913 3673 1927 3687
rect 1953 3673 1967 3687
rect 2053 3673 2067 3687
rect 1873 3633 1887 3647
rect 1973 3653 1987 3667
rect 1953 3613 1967 3627
rect 1933 3593 1947 3607
rect 1893 3514 1907 3528
rect 1873 3472 1887 3486
rect 1893 3453 1907 3467
rect 1853 3433 1867 3447
rect 1833 3373 1847 3387
rect 1853 3353 1867 3367
rect 1813 3313 1827 3327
rect 1853 3294 1867 3308
rect 2013 3514 2027 3528
rect 2053 3514 2067 3528
rect 2113 3753 2127 3767
rect 2113 3713 2127 3727
rect 1913 3413 1927 3427
rect 1973 3413 1987 3427
rect 1993 3393 2007 3407
rect 2093 3473 2107 3487
rect 2033 3373 2047 3387
rect 2033 3352 2047 3366
rect 1933 3333 1947 3347
rect 1973 3333 1987 3347
rect 1953 3273 1967 3287
rect 1813 3252 1827 3266
rect 1873 3252 1887 3266
rect 1933 3253 1947 3267
rect 1913 3233 1927 3247
rect 1913 3212 1927 3226
rect 1873 3173 1887 3187
rect 1813 3093 1827 3107
rect 1833 3053 1847 3067
rect 1813 2993 1827 3007
rect 1893 2953 1907 2967
rect 1853 2933 1867 2947
rect 2113 3353 2127 3367
rect 2073 3333 2087 3347
rect 2073 3294 2087 3308
rect 2113 3294 2127 3308
rect 2153 3772 2167 3786
rect 2153 3751 2167 3765
rect 2313 4093 2327 4107
rect 2393 4233 2407 4247
rect 2373 4193 2387 4207
rect 2353 4073 2367 4087
rect 2273 4034 2287 4048
rect 2313 4034 2327 4048
rect 2313 3973 2327 3987
rect 2293 3953 2307 3967
rect 2233 3853 2247 3867
rect 2273 3853 2287 3867
rect 2233 3794 2247 3808
rect 2473 4313 2487 4327
rect 2473 4273 2487 4287
rect 2433 4193 2447 4207
rect 2393 4073 2407 4087
rect 2553 4613 2567 4627
rect 2513 4473 2527 4487
rect 2593 4473 2607 4487
rect 2853 4893 2867 4907
rect 2813 4873 2827 4887
rect 2773 4854 2787 4868
rect 2792 4793 2806 4807
rect 2813 4793 2827 4807
rect 2692 4773 2706 4787
rect 2713 4773 2727 4787
rect 2733 4753 2747 4767
rect 2673 4713 2687 4727
rect 2793 4713 2807 4727
rect 2693 4693 2707 4707
rect 2673 4673 2687 4687
rect 2673 4593 2687 4607
rect 2733 4613 2747 4627
rect 2793 4612 2807 4626
rect 2733 4554 2747 4568
rect 2773 4553 2787 4567
rect 2833 4713 2847 4727
rect 2833 4692 2847 4706
rect 2893 4913 2907 4927
rect 2873 4793 2887 4807
rect 2873 4733 2887 4747
rect 2853 4673 2867 4687
rect 2833 4613 2847 4627
rect 2853 4593 2867 4607
rect 2973 5074 2987 5088
rect 3213 5352 3227 5366
rect 3353 5713 3367 5727
rect 3353 5413 3367 5427
rect 3413 6013 3427 6027
rect 3773 6013 3787 6027
rect 3453 5953 3467 5967
rect 3413 5893 3427 5907
rect 3573 5913 3587 5927
rect 3713 5913 3727 5927
rect 3493 5894 3507 5908
rect 3573 5894 3587 5908
rect 3613 5894 3627 5908
rect 3653 5894 3667 5908
rect 3973 6134 3987 6148
rect 4393 6173 4407 6187
rect 4133 6094 4147 6108
rect 4293 6073 4307 6087
rect 3893 6053 3907 6067
rect 3993 5993 4007 6007
rect 3873 5933 3887 5947
rect 3933 5933 3947 5947
rect 3873 5894 3887 5908
rect 3913 5893 3927 5907
rect 3433 5852 3447 5866
rect 3473 5852 3487 5866
rect 3653 5853 3667 5867
rect 3653 5813 3667 5827
rect 3593 5793 3607 5807
rect 3653 5733 3667 5747
rect 3413 5713 3427 5727
rect 3693 5693 3707 5707
rect 3393 5594 3407 5608
rect 3433 5594 3447 5608
rect 3533 5594 3547 5608
rect 3572 5593 3586 5607
rect 3593 5593 3607 5607
rect 3653 5594 3667 5608
rect 3793 5594 3807 5608
rect 3913 5852 3927 5866
rect 3853 5793 3867 5807
rect 4113 5973 4127 5987
rect 4053 5913 4067 5927
rect 4153 5894 4167 5908
rect 4193 5874 4207 5888
rect 3973 5852 3987 5866
rect 4053 5852 4067 5866
rect 4133 5852 4147 5866
rect 4013 5813 4027 5827
rect 4093 5813 4107 5827
rect 3933 5653 3947 5667
rect 3853 5633 3867 5647
rect 3513 5552 3527 5566
rect 3393 5513 3407 5527
rect 3433 5513 3447 5527
rect 3373 5393 3387 5407
rect 3533 5473 3547 5487
rect 3573 5473 3587 5487
rect 3433 5413 3447 5427
rect 3353 5353 3367 5367
rect 3393 5353 3407 5367
rect 3413 5333 3427 5347
rect 3213 5313 3227 5327
rect 3313 5313 3327 5327
rect 3073 5193 3087 5207
rect 3373 5312 3387 5326
rect 3373 5273 3387 5287
rect 3453 5373 3467 5387
rect 3573 5452 3587 5466
rect 3613 5552 3627 5566
rect 3773 5552 3787 5566
rect 3773 5493 3787 5507
rect 3713 5433 3727 5447
rect 3653 5413 3667 5427
rect 3453 5312 3467 5326
rect 3513 5332 3527 5346
rect 3492 5293 3506 5307
rect 3513 5293 3527 5307
rect 3473 5253 3487 5267
rect 3233 5193 3247 5207
rect 3433 5193 3447 5207
rect 3233 5153 3247 5167
rect 3473 5153 3487 5167
rect 3213 5133 3227 5147
rect 3053 5094 3067 5108
rect 3413 5113 3427 5127
rect 3113 5093 3127 5107
rect 3213 5093 3227 5107
rect 3093 5052 3107 5066
rect 2953 5033 2967 5047
rect 2953 4993 2967 5007
rect 2973 4953 2987 4967
rect 2933 4873 2947 4887
rect 2913 4854 2927 4868
rect 2953 4713 2967 4727
rect 2953 4692 2967 4706
rect 2913 4673 2927 4687
rect 2913 4593 2927 4607
rect 2673 4512 2687 4526
rect 2913 4533 2927 4547
rect 2713 4473 2727 4487
rect 2773 4473 2787 4487
rect 2633 4453 2647 4467
rect 2833 4512 2847 4526
rect 2833 4453 2847 4467
rect 2873 4453 2887 4467
rect 2613 4413 2627 4427
rect 2793 4413 2807 4427
rect 2733 4393 2747 4407
rect 2493 4113 2507 4127
rect 2452 4053 2466 4067
rect 2473 4053 2487 4067
rect 2413 4034 2427 4048
rect 2453 4034 2467 4048
rect 2373 3973 2387 3987
rect 2333 3933 2347 3947
rect 2333 3912 2347 3926
rect 2273 3773 2287 3787
rect 2253 3733 2267 3747
rect 2213 3573 2227 3587
rect 2253 3533 2267 3547
rect 2153 3514 2167 3528
rect 2213 3513 2227 3527
rect 2193 3472 2207 3486
rect 2232 3492 2246 3506
rect 2253 3493 2267 3507
rect 1973 3252 1987 3266
rect 2013 3252 2027 3266
rect 1953 3213 1967 3227
rect 1973 3133 1987 3147
rect 1933 3093 1947 3107
rect 1973 3093 1987 3107
rect 1913 2913 1927 2927
rect 1893 2893 1907 2907
rect 1793 2873 1807 2887
rect 1833 2793 1847 2807
rect 1773 2774 1787 2788
rect 1813 2774 1827 2788
rect 1753 2732 1767 2746
rect 1813 2733 1827 2747
rect 1793 2713 1807 2727
rect 1793 2653 1807 2667
rect 1713 2593 1727 2607
rect 1513 2533 1527 2547
rect 1653 2533 1667 2547
rect 1733 2533 1747 2547
rect 1533 2513 1547 2527
rect 1613 2493 1627 2507
rect 1553 2432 1567 2446
rect 1513 2413 1527 2427
rect 1433 2393 1447 2407
rect 1373 2353 1387 2367
rect 1413 2333 1427 2347
rect 1433 2313 1447 2327
rect 1433 2273 1447 2287
rect 1473 2273 1487 2287
rect 1373 2213 1387 2227
rect 1393 2193 1407 2207
rect 1433 2193 1447 2207
rect 1373 2173 1387 2187
rect 1413 2113 1427 2127
rect 1373 2053 1387 2067
rect 1373 1973 1387 1987
rect 1313 1633 1327 1647
rect 1353 1873 1367 1887
rect 1553 2411 1567 2425
rect 1513 2333 1527 2347
rect 1533 2293 1547 2307
rect 1513 2153 1527 2167
rect 1493 2093 1507 2107
rect 1593 2393 1607 2407
rect 1553 2253 1567 2267
rect 1633 2373 1647 2387
rect 1633 2313 1647 2327
rect 1613 2293 1627 2307
rect 1553 2213 1567 2227
rect 1613 2212 1627 2226
rect 1573 2173 1587 2187
rect 1553 2133 1567 2147
rect 1773 2473 1787 2487
rect 1693 2432 1707 2446
rect 2093 3053 2107 3067
rect 2213 3293 2227 3307
rect 2153 3252 2167 3266
rect 2213 3173 2227 3187
rect 2193 3113 2207 3127
rect 2153 2994 2167 3008
rect 2013 2952 2027 2966
rect 2093 2953 2107 2967
rect 2173 2952 2187 2966
rect 1953 2933 1967 2947
rect 2013 2931 2027 2945
rect 2133 2933 2147 2947
rect 1953 2873 1967 2887
rect 1933 2833 1947 2847
rect 1873 2732 1887 2746
rect 1833 2693 1847 2707
rect 1813 2633 1827 2647
rect 1913 2713 1927 2727
rect 1873 2553 1887 2567
rect 1813 2474 1827 2488
rect 1893 2453 1907 2467
rect 1793 2432 1807 2446
rect 1673 2313 1687 2327
rect 1613 2073 1627 2087
rect 1653 2073 1667 2087
rect 1533 2033 1547 2047
rect 1493 1954 1507 1968
rect 1453 1893 1467 1907
rect 1413 1833 1427 1847
rect 1373 1793 1387 1807
rect 1433 1734 1447 1748
rect 1393 1692 1407 1706
rect 1393 1633 1407 1647
rect 1333 1613 1347 1627
rect 1373 1613 1387 1627
rect 1293 1553 1307 1567
rect 1273 1533 1287 1547
rect 1313 1533 1327 1547
rect 1293 1392 1307 1406
rect 1293 1353 1307 1367
rect 1253 1214 1267 1228
rect 1333 1333 1347 1347
rect 1333 1214 1347 1228
rect 1233 1133 1247 1147
rect 1473 1853 1487 1867
rect 1573 1954 1587 1968
rect 1593 1912 1607 1926
rect 1633 1893 1647 1907
rect 1533 1853 1547 1867
rect 1573 1833 1587 1847
rect 1613 1833 1627 1847
rect 1513 1773 1527 1787
rect 1513 1734 1527 1748
rect 1553 1613 1567 1627
rect 1453 1593 1467 1607
rect 1533 1593 1547 1607
rect 1433 1553 1447 1567
rect 1513 1553 1527 1567
rect 1433 1513 1447 1527
rect 1413 1493 1427 1507
rect 1473 1434 1487 1448
rect 1533 1453 1547 1467
rect 1513 1433 1527 1447
rect 1453 1392 1467 1406
rect 1493 1373 1507 1387
rect 1413 1333 1427 1347
rect 1473 1333 1487 1347
rect 1493 1273 1507 1287
rect 1493 1233 1507 1247
rect 1593 1793 1607 1807
rect 1593 1733 1607 1747
rect 1713 2273 1727 2287
rect 1773 2353 1787 2367
rect 1753 2253 1767 2267
rect 1732 2212 1746 2226
rect 1753 2213 1767 2227
rect 1693 2133 1707 2147
rect 1873 2333 1887 2347
rect 1853 2313 1867 2327
rect 1793 2293 1807 2307
rect 1773 2153 1787 2167
rect 1693 1953 1707 1967
rect 1713 1873 1727 1887
rect 1633 1692 1647 1706
rect 1653 1673 1667 1687
rect 1633 1653 1647 1667
rect 1573 1453 1587 1467
rect 1593 1434 1607 1448
rect 1573 1392 1587 1406
rect 1973 2853 1987 2867
rect 2253 3393 2267 3407
rect 2593 4053 2607 4067
rect 2553 4034 2567 4048
rect 2753 4314 2767 4328
rect 2772 4273 2786 4287
rect 2793 4272 2807 4286
rect 2813 4213 2827 4227
rect 2673 4153 2687 4167
rect 2733 4153 2747 4167
rect 2793 4153 2807 4167
rect 2513 3973 2527 3987
rect 2433 3893 2447 3907
rect 2473 3792 2487 3806
rect 2613 3992 2627 4006
rect 2593 3973 2607 3987
rect 2773 4132 2787 4146
rect 2693 4033 2707 4047
rect 2673 3993 2687 4007
rect 2653 3953 2667 3967
rect 2673 3893 2687 3907
rect 2613 3833 2627 3847
rect 2613 3793 2627 3807
rect 2673 3773 2687 3787
rect 2653 3753 2667 3767
rect 2573 3633 2587 3647
rect 2573 3612 2587 3626
rect 2333 3573 2347 3587
rect 2313 3533 2327 3547
rect 2473 3494 2487 3508
rect 2653 3673 2667 3687
rect 2713 3992 2727 4006
rect 2853 4413 2867 4427
rect 2853 4133 2867 4147
rect 2833 4093 2847 4107
rect 2933 4513 2947 4527
rect 2933 4373 2947 4387
rect 2913 4353 2927 4367
rect 3073 4973 3087 4987
rect 3353 5073 3367 5087
rect 3213 5054 3227 5068
rect 3413 5013 3427 5027
rect 3453 5013 3467 5027
rect 3213 4953 3227 4967
rect 3353 4953 3367 4967
rect 3113 4933 3127 4947
rect 3113 4912 3127 4926
rect 3113 4873 3127 4887
rect 3353 4932 3367 4946
rect 3213 4854 3227 4868
rect 2993 4812 3007 4826
rect 3053 4812 3067 4826
rect 3253 4812 3267 4826
rect 3333 4812 3347 4826
rect 3373 4812 3387 4826
rect 3433 4973 3447 4987
rect 3473 4953 3487 4967
rect 3533 5253 3547 5267
rect 3593 5333 3607 5347
rect 3813 5493 3827 5507
rect 3893 5594 3907 5608
rect 4093 5693 4107 5707
rect 4493 6114 4507 6128
rect 4633 6113 4647 6127
rect 4393 6073 4407 6087
rect 4473 6072 4487 6086
rect 4373 6053 4387 6067
rect 4373 5993 4387 6007
rect 4573 5933 4587 5947
rect 4433 5872 4447 5886
rect 4573 5873 4587 5887
rect 4613 5873 4627 5887
rect 4533 5833 4547 5847
rect 4573 5833 4587 5847
rect 4553 5793 4567 5807
rect 4253 5733 4267 5747
rect 4293 5733 4307 5747
rect 4493 5733 4507 5747
rect 4253 5673 4267 5687
rect 4193 5653 4207 5667
rect 4233 5653 4247 5667
rect 4073 5593 4087 5607
rect 4133 5594 4147 5608
rect 4253 5593 4267 5607
rect 4353 5593 4367 5607
rect 3973 5573 3987 5587
rect 3853 5373 3867 5387
rect 3573 5293 3587 5307
rect 3553 5193 3567 5207
rect 3533 5153 3547 5167
rect 3573 5153 3587 5167
rect 3673 5332 3687 5346
rect 3713 5332 3727 5346
rect 3753 5332 3767 5346
rect 3793 5332 3807 5346
rect 3832 5333 3846 5347
rect 3853 5333 3867 5347
rect 3653 5293 3667 5307
rect 3613 5253 3627 5267
rect 3613 5232 3627 5246
rect 3553 5113 3567 5127
rect 3593 5113 3607 5127
rect 3533 5053 3547 5067
rect 3593 5033 3607 5047
rect 3573 5013 3587 5027
rect 3533 4893 3547 4907
rect 3513 4873 3527 4887
rect 3593 4973 3607 4987
rect 3593 4933 3607 4947
rect 3552 4853 3566 4867
rect 3573 4852 3587 4866
rect 3093 4793 3107 4807
rect 3233 4793 3247 4807
rect 3053 4713 3067 4727
rect 3193 4713 3207 4727
rect 2973 4673 2987 4687
rect 3033 4573 3047 4587
rect 3053 4553 3067 4567
rect 3093 4433 3107 4447
rect 2993 4373 3007 4387
rect 2973 4333 2987 4347
rect 2953 4292 2967 4306
rect 2933 4273 2947 4287
rect 2913 4233 2927 4247
rect 2913 4173 2927 4187
rect 2913 4133 2927 4147
rect 2893 4113 2907 4127
rect 2893 4053 2907 4067
rect 2873 4033 2887 4047
rect 3013 4353 3027 4367
rect 3073 4353 3087 4367
rect 2993 4133 3007 4147
rect 3153 4393 3167 4407
rect 3093 4313 3107 4327
rect 3033 4272 3047 4286
rect 3053 4233 3067 4247
rect 3033 4193 3047 4207
rect 3033 4133 3047 4147
rect 3013 4113 3027 4127
rect 2993 4073 3007 4087
rect 2933 4033 2947 4047
rect 2813 3993 2827 4007
rect 2793 3913 2807 3927
rect 2713 3853 2727 3867
rect 2813 3853 2827 3867
rect 2773 3833 2787 3847
rect 2853 3953 2867 3967
rect 2893 3933 2907 3947
rect 2853 3913 2867 3927
rect 2833 3813 2847 3827
rect 2753 3772 2767 3786
rect 2973 4013 2987 4027
rect 2953 3893 2967 3907
rect 2893 3853 2907 3867
rect 2933 3833 2947 3847
rect 2873 3773 2887 3787
rect 2713 3752 2727 3766
rect 2793 3753 2807 3767
rect 2853 3753 2867 3767
rect 2713 3713 2727 3727
rect 2833 3713 2847 3727
rect 2773 3693 2787 3707
rect 2713 3673 2727 3687
rect 2693 3653 2707 3667
rect 2673 3633 2687 3647
rect 2653 3533 2667 3547
rect 2313 3473 2327 3487
rect 2573 3473 2587 3487
rect 2293 3453 2307 3467
rect 2293 3313 2307 3327
rect 2273 3293 2287 3307
rect 2573 3413 2587 3427
rect 2493 3393 2507 3407
rect 2413 3313 2427 3327
rect 2373 3293 2387 3307
rect 2253 3252 2267 3266
rect 2293 3252 2307 3266
rect 2333 3252 2347 3266
rect 2373 3253 2387 3267
rect 2273 3193 2287 3207
rect 2073 2893 2087 2907
rect 2233 2893 2247 2907
rect 2013 2813 2027 2827
rect 1973 2773 1987 2787
rect 2113 2793 2127 2807
rect 2173 2793 2187 2807
rect 1993 2732 2007 2746
rect 2033 2732 2047 2746
rect 2073 2732 2087 2746
rect 1953 2713 1967 2727
rect 2013 2713 2027 2727
rect 1933 2593 1947 2607
rect 1993 2673 2007 2687
rect 1953 2573 1967 2587
rect 1953 2493 1967 2507
rect 2013 2633 2027 2647
rect 2133 2693 2147 2707
rect 2053 2633 2067 2647
rect 2033 2533 2047 2547
rect 1993 2474 2007 2488
rect 1953 2432 1967 2446
rect 2013 2432 2027 2446
rect 1933 2393 1947 2407
rect 1913 2373 1927 2387
rect 2013 2393 2027 2407
rect 1953 2333 1967 2347
rect 1993 2333 2007 2347
rect 1893 2293 1907 2307
rect 1853 2254 1867 2268
rect 1933 2273 1947 2287
rect 1993 2273 2007 2287
rect 2033 2273 2047 2287
rect 2013 2254 2027 2268
rect 2113 2613 2127 2627
rect 2193 2774 2207 2788
rect 2233 2774 2247 2788
rect 2353 3173 2367 3187
rect 2333 2873 2347 2887
rect 2453 3294 2467 3308
rect 2553 3373 2567 3387
rect 2513 3252 2527 3266
rect 2473 3233 2487 3247
rect 2413 3213 2427 3227
rect 2473 3212 2487 3226
rect 2393 3153 2407 3167
rect 2433 3133 2447 3147
rect 2433 3093 2447 3107
rect 2493 3093 2507 3107
rect 2453 3073 2467 3087
rect 2393 3033 2407 3047
rect 2373 2953 2387 2967
rect 2413 2952 2427 2966
rect 2353 2793 2367 2807
rect 2333 2774 2347 2788
rect 2373 2774 2387 2788
rect 2453 2833 2467 2847
rect 2473 2793 2487 2807
rect 2233 2693 2247 2707
rect 2293 2713 2307 2727
rect 2313 2693 2327 2707
rect 2253 2613 2267 2627
rect 2173 2453 2187 2467
rect 2093 2432 2107 2446
rect 2133 2413 2147 2427
rect 2173 2413 2187 2427
rect 2253 2413 2267 2427
rect 2093 2333 2107 2347
rect 2113 2253 2127 2267
rect 1873 2212 1887 2226
rect 1933 2212 1947 2226
rect 2033 2212 2047 2226
rect 2093 2212 2107 2226
rect 1993 2193 2007 2207
rect 2053 2193 2067 2207
rect 1833 2173 1847 2187
rect 1993 2152 2007 2166
rect 1853 2113 1867 2127
rect 1973 2113 1987 2127
rect 1873 2093 1887 2107
rect 1853 1953 1867 1967
rect 1933 2053 1947 2067
rect 1973 2013 1987 2027
rect 1953 1993 1967 2007
rect 1853 1913 1867 1927
rect 1893 1912 1907 1926
rect 1893 1873 1907 1887
rect 1813 1833 1827 1847
rect 1853 1833 1867 1847
rect 1793 1813 1807 1827
rect 1813 1793 1827 1807
rect 1773 1734 1787 1748
rect 1833 1734 1847 1748
rect 1692 1653 1706 1667
rect 1713 1653 1727 1667
rect 1713 1613 1727 1627
rect 1753 1692 1767 1706
rect 1813 1653 1827 1667
rect 1793 1633 1807 1647
rect 1753 1613 1767 1627
rect 1733 1553 1747 1567
rect 1673 1493 1687 1507
rect 1713 1493 1727 1507
rect 1653 1473 1667 1487
rect 1793 1513 1807 1527
rect 1773 1493 1787 1507
rect 1813 1493 1827 1507
rect 1773 1452 1787 1466
rect 1753 1433 1767 1447
rect 1533 1353 1547 1367
rect 1533 1313 1547 1327
rect 1553 1293 1567 1307
rect 1533 1213 1547 1227
rect 1253 1113 1267 1127
rect 1332 1153 1346 1167
rect 1353 1153 1367 1167
rect 1313 1133 1327 1147
rect 1333 1073 1347 1087
rect 1293 1033 1307 1047
rect 1333 1033 1347 1047
rect 1233 1013 1247 1027
rect 1093 813 1107 827
rect 1033 793 1047 807
rect 993 694 1007 708
rect 1073 773 1087 787
rect 1213 873 1227 887
rect 1253 973 1267 987
rect 1313 973 1327 987
rect 1273 872 1287 886
rect 1353 993 1367 1007
rect 1353 933 1367 947
rect 1353 893 1367 907
rect 1093 733 1107 747
rect 1153 733 1167 747
rect 1193 733 1207 747
rect 1013 652 1027 666
rect 1073 652 1087 666
rect 973 593 987 607
rect 1153 694 1167 708
rect 1233 694 1247 708
rect 1173 652 1187 666
rect 1333 853 1347 867
rect 1353 793 1367 807
rect 1353 772 1367 786
rect 1393 973 1407 987
rect 1493 1172 1507 1186
rect 1613 1233 1627 1247
rect 1693 1392 1707 1406
rect 1713 1373 1727 1387
rect 1693 1233 1707 1247
rect 1593 1172 1607 1186
rect 1553 1153 1567 1167
rect 1453 1113 1467 1127
rect 1493 1113 1507 1127
rect 1473 1093 1487 1107
rect 1453 1073 1467 1087
rect 1553 1073 1567 1087
rect 1493 993 1507 1007
rect 1533 953 1547 967
rect 1413 933 1427 947
rect 1453 914 1467 928
rect 1513 893 1527 907
rect 1413 853 1427 867
rect 1393 793 1407 807
rect 1333 753 1347 767
rect 1313 694 1327 708
rect 1393 673 1407 687
rect 1273 653 1287 667
rect 1313 633 1327 647
rect 1173 613 1187 627
rect 1233 613 1247 627
rect 1293 613 1307 627
rect 1133 573 1147 587
rect 1093 553 1107 567
rect 973 513 987 527
rect 1133 513 1147 527
rect 933 473 947 487
rect 933 393 947 407
rect 1093 453 1107 467
rect 1033 433 1047 447
rect 1073 432 1087 446
rect 1073 392 1087 406
rect 1353 593 1367 607
rect 1313 573 1327 587
rect 1193 493 1207 507
rect 1173 473 1187 487
rect 1193 433 1207 447
rect 1173 394 1187 408
rect 1213 393 1227 407
rect 1273 394 1287 408
rect 1313 394 1327 408
rect 1473 872 1487 886
rect 1493 833 1507 847
rect 1433 733 1447 747
rect 1453 713 1467 727
rect 1653 1153 1667 1167
rect 1633 993 1647 1007
rect 1633 953 1647 967
rect 1793 1433 1807 1447
rect 1873 1793 1887 1807
rect 1973 1873 1987 1887
rect 1953 1853 1967 1867
rect 2013 2113 2027 2127
rect 2013 1973 2027 1987
rect 2073 1973 2087 1987
rect 2053 1954 2067 1968
rect 2353 2733 2367 2747
rect 2333 2633 2347 2647
rect 2433 2713 2447 2727
rect 2393 2693 2407 2707
rect 2393 2633 2407 2647
rect 2353 2593 2367 2607
rect 2393 2573 2407 2587
rect 2433 2533 2447 2547
rect 2433 2474 2447 2488
rect 2373 2413 2387 2427
rect 2353 2333 2367 2347
rect 2353 2293 2367 2307
rect 2313 2253 2327 2267
rect 2373 2253 2387 2267
rect 2253 2212 2267 2226
rect 2293 2212 2307 2226
rect 2173 2093 2187 2107
rect 2153 1973 2167 1987
rect 2133 1953 2147 1967
rect 2013 1912 2027 1926
rect 2073 1912 2087 1926
rect 1993 1793 2007 1807
rect 1893 1773 1907 1787
rect 1973 1773 1987 1787
rect 1913 1734 1927 1748
rect 1873 1653 1887 1667
rect 1913 1673 1927 1687
rect 1893 1633 1907 1647
rect 1853 1613 1867 1627
rect 1833 1453 1847 1467
rect 1833 1392 1847 1406
rect 1773 1353 1787 1367
rect 1833 1353 1847 1367
rect 1793 1293 1807 1307
rect 1733 1233 1747 1247
rect 1713 1213 1727 1227
rect 1753 1214 1767 1228
rect 1793 1214 1807 1228
rect 1712 1173 1726 1187
rect 1693 1073 1707 1087
rect 1693 1033 1707 1047
rect 1553 913 1567 927
rect 1593 914 1607 928
rect 1673 933 1687 947
rect 1653 913 1667 927
rect 1733 1172 1747 1186
rect 1813 1173 1827 1187
rect 1733 1053 1747 1067
rect 1793 993 1807 1007
rect 1713 933 1727 947
rect 1913 1573 1927 1587
rect 1893 1333 1907 1347
rect 1973 1693 1987 1707
rect 2113 1893 2127 1907
rect 2053 1833 2067 1847
rect 2193 2013 2207 2027
rect 2233 1973 2247 1987
rect 2473 2713 2487 2727
rect 2533 3053 2547 3067
rect 2573 3353 2587 3367
rect 2613 3493 2627 3507
rect 2673 3493 2687 3507
rect 2753 3613 2767 3627
rect 2733 3573 2747 3587
rect 2713 3533 2727 3547
rect 2693 3433 2707 3447
rect 2673 3393 2687 3407
rect 2613 3373 2627 3387
rect 2693 3353 2707 3367
rect 2593 3313 2607 3327
rect 2573 3293 2587 3307
rect 2633 3294 2647 3308
rect 2573 3252 2587 3266
rect 2653 3252 2667 3266
rect 2633 3233 2647 3247
rect 2613 3193 2627 3207
rect 2573 3073 2587 3087
rect 2552 3033 2566 3047
rect 2573 3033 2587 3047
rect 2533 2993 2547 3007
rect 2753 3553 2767 3567
rect 2793 3613 2807 3627
rect 2873 3693 2887 3707
rect 2913 3673 2927 3687
rect 3033 4053 3047 4067
rect 3013 4012 3027 4026
rect 3033 3993 3047 4007
rect 3033 3933 3047 3947
rect 3312 4733 3326 4747
rect 3333 4733 3347 4747
rect 3253 4693 3267 4707
rect 3233 4493 3247 4507
rect 3233 4453 3247 4467
rect 3193 4353 3207 4367
rect 3213 4334 3227 4348
rect 3173 4292 3187 4306
rect 3333 4553 3347 4567
rect 3433 4812 3447 4826
rect 3473 4812 3487 4826
rect 3513 4812 3527 4826
rect 3533 4753 3547 4767
rect 3413 4733 3427 4747
rect 3653 5213 3667 5227
rect 3753 5054 3767 5068
rect 3913 5533 3927 5547
rect 4033 5533 4047 5547
rect 3993 5513 4007 5527
rect 3893 5393 3907 5407
rect 3893 5374 3907 5388
rect 3953 5373 3967 5387
rect 3933 5332 3947 5346
rect 3873 5273 3887 5287
rect 3873 5233 3887 5247
rect 3893 5193 3907 5207
rect 3873 5173 3887 5187
rect 3893 5153 3907 5167
rect 3853 4973 3867 4987
rect 3833 4953 3847 4967
rect 3713 4933 3727 4947
rect 3693 4913 3707 4927
rect 3673 4893 3687 4907
rect 3693 4873 3707 4887
rect 3613 4853 3627 4867
rect 3653 4854 3667 4868
rect 3733 4853 3747 4867
rect 3773 4854 3787 4868
rect 3593 4812 3607 4826
rect 3633 4812 3647 4826
rect 3673 4812 3687 4826
rect 3853 4854 3867 4868
rect 3753 4813 3767 4827
rect 3613 4753 3627 4767
rect 3733 4753 3747 4767
rect 3573 4733 3587 4747
rect 3653 4693 3667 4707
rect 3493 4673 3507 4687
rect 3533 4673 3547 4687
rect 3433 4554 3447 4568
rect 3413 4533 3427 4547
rect 3393 4513 3407 4527
rect 3413 4493 3427 4507
rect 3393 4473 3407 4487
rect 3353 4453 3367 4467
rect 3393 4413 3407 4427
rect 3333 4393 3347 4407
rect 3373 4373 3387 4387
rect 3273 4353 3287 4367
rect 3333 4353 3347 4367
rect 3193 4273 3207 4287
rect 3253 4273 3267 4287
rect 3153 4133 3167 4147
rect 3373 4333 3387 4347
rect 3273 4253 3287 4267
rect 3313 4292 3327 4306
rect 3293 4213 3307 4227
rect 3192 4014 3206 4028
rect 3213 4013 3227 4027
rect 3353 4153 3367 4167
rect 3453 4393 3467 4407
rect 3413 4333 3427 4347
rect 3513 4633 3527 4647
rect 3513 4593 3527 4607
rect 3553 4593 3567 4607
rect 3593 4553 3607 4567
rect 3693 4554 3707 4568
rect 3593 4493 3607 4507
rect 3573 4393 3587 4407
rect 3533 4373 3547 4387
rect 3493 4334 3507 4348
rect 3533 4314 3547 4328
rect 3413 4293 3427 4307
rect 3453 4273 3467 4287
rect 3433 4253 3447 4267
rect 3413 4073 3427 4087
rect 3353 4054 3367 4068
rect 3393 4054 3407 4068
rect 3053 3913 3067 3927
rect 3113 3913 3127 3927
rect 3173 3913 3187 3927
rect 3293 3913 3307 3927
rect 3033 3873 3047 3887
rect 3093 3873 3107 3887
rect 3013 3713 3027 3727
rect 2993 3693 3007 3707
rect 2953 3653 2967 3667
rect 2873 3633 2887 3647
rect 2833 3593 2847 3607
rect 2772 3533 2786 3547
rect 2793 3533 2807 3547
rect 2893 3613 2907 3627
rect 2873 3553 2887 3567
rect 2753 3513 2767 3527
rect 3153 3833 3167 3847
rect 3113 3793 3127 3807
rect 3153 3792 3167 3806
rect 3433 4013 3447 4027
rect 3413 3893 3427 3907
rect 3193 3813 3207 3827
rect 3053 3772 3067 3786
rect 3133 3733 3147 3747
rect 3173 3733 3187 3747
rect 3113 3713 3127 3727
rect 3113 3673 3127 3687
rect 3033 3613 3047 3627
rect 3153 3713 3167 3727
rect 3153 3633 3167 3647
rect 3013 3593 3027 3607
rect 3133 3593 3147 3607
rect 2993 3573 3007 3587
rect 2893 3513 2907 3527
rect 2853 3493 2867 3507
rect 2733 3473 2747 3487
rect 2813 3473 2827 3487
rect 2773 3433 2787 3447
rect 2753 3413 2767 3427
rect 2733 3353 2747 3367
rect 2713 3213 2727 3227
rect 2833 3393 2847 3407
rect 2813 3252 2827 3266
rect 2793 3233 2807 3247
rect 2853 3294 2867 3308
rect 2833 3173 2847 3187
rect 3173 3553 3187 3567
rect 3133 3533 3147 3547
rect 2893 3473 2907 3487
rect 3173 3492 3187 3506
rect 3293 3792 3307 3806
rect 3293 3673 3307 3687
rect 3253 3653 3267 3667
rect 3213 3573 3227 3587
rect 3213 3533 3227 3547
rect 3233 3473 3247 3487
rect 3213 3433 3227 3447
rect 3193 3413 3207 3427
rect 3133 3393 3147 3407
rect 2893 3373 2907 3387
rect 2953 3373 2967 3387
rect 2993 3373 3007 3387
rect 3213 3373 3227 3387
rect 2933 3294 2947 3308
rect 2733 3093 2747 3107
rect 2773 3093 2787 3107
rect 2753 3033 2767 3047
rect 2613 2994 2627 3008
rect 2653 2994 2667 3008
rect 2693 2994 2707 3008
rect 2553 2952 2567 2966
rect 2533 2933 2547 2947
rect 2513 2873 2527 2887
rect 2513 2833 2527 2847
rect 2493 2673 2507 2687
rect 2473 2593 2487 2607
rect 2453 2373 2467 2387
rect 2433 2353 2447 2367
rect 2433 2313 2447 2327
rect 2413 2293 2427 2307
rect 2493 2553 2507 2567
rect 2433 2273 2447 2287
rect 2473 2273 2487 2287
rect 2413 2254 2427 2268
rect 2393 2113 2407 2127
rect 2413 2093 2427 2107
rect 2333 2053 2347 2067
rect 2473 2033 2487 2047
rect 2413 2013 2427 2027
rect 2273 1954 2287 1968
rect 2313 1954 2327 1968
rect 2173 1893 2187 1907
rect 2253 1912 2267 1926
rect 2213 1813 2227 1827
rect 2013 1673 2027 1687
rect 2073 1673 2087 1687
rect 1993 1613 2007 1627
rect 2073 1613 2087 1627
rect 1973 1593 1987 1607
rect 2013 1593 2027 1607
rect 1953 1553 1967 1567
rect 1993 1553 2007 1567
rect 1953 1493 1967 1507
rect 1953 1434 1967 1448
rect 2053 1533 2067 1547
rect 2033 1473 2047 1487
rect 1933 1393 1947 1407
rect 1953 1373 1967 1387
rect 1933 1293 1947 1307
rect 1853 1253 1867 1267
rect 1913 1253 1927 1267
rect 1833 1153 1847 1167
rect 1833 1093 1847 1107
rect 1913 1214 1927 1228
rect 2013 1392 2027 1406
rect 1993 1353 2007 1367
rect 1973 1333 1987 1347
rect 2013 1333 2027 1347
rect 1933 1172 1947 1186
rect 1993 1313 2007 1327
rect 2193 1734 2207 1748
rect 2252 1734 2266 1748
rect 2273 1734 2287 1748
rect 2413 1954 2427 1968
rect 2553 2833 2567 2847
rect 2533 2774 2547 2788
rect 2533 2653 2547 2667
rect 2533 2593 2547 2607
rect 2633 2933 2647 2947
rect 2613 2713 2627 2727
rect 2573 2573 2587 2587
rect 2593 2493 2607 2507
rect 2573 2413 2587 2427
rect 2713 2953 2727 2967
rect 2673 2913 2687 2927
rect 2713 2793 2727 2807
rect 2693 2732 2707 2746
rect 2753 2993 2767 3007
rect 2813 3013 2827 3027
rect 2953 3193 2967 3207
rect 3233 3353 3247 3367
rect 3013 3333 3027 3347
rect 2993 3093 3007 3107
rect 2913 3013 2927 3027
rect 2853 2994 2867 3008
rect 2893 2994 2907 3008
rect 2793 2952 2807 2966
rect 2793 2933 2807 2947
rect 2753 2893 2767 2907
rect 2673 2693 2687 2707
rect 2733 2693 2747 2707
rect 2633 2432 2647 2446
rect 2613 2373 2627 2387
rect 2553 2313 2567 2327
rect 2533 2273 2547 2287
rect 2333 1913 2347 1927
rect 2433 1912 2447 1926
rect 2473 1913 2487 1927
rect 2413 1893 2427 1907
rect 2393 1773 2407 1787
rect 2353 1734 2367 1748
rect 2133 1693 2147 1707
rect 2113 1493 2127 1507
rect 2093 1453 2107 1467
rect 2233 1693 2247 1707
rect 2173 1673 2187 1687
rect 2213 1673 2227 1687
rect 2153 1553 2167 1567
rect 2153 1493 2167 1507
rect 2173 1473 2187 1487
rect 2153 1453 2167 1467
rect 2173 1434 2187 1448
rect 2093 1413 2107 1427
rect 2073 1373 2087 1387
rect 2053 1353 2067 1367
rect 2033 1253 2047 1267
rect 2013 1233 2027 1247
rect 1993 1213 2007 1227
rect 2033 1214 2047 1228
rect 2073 1213 2087 1227
rect 2013 1172 2027 1186
rect 2053 1172 2067 1186
rect 1933 1133 1947 1147
rect 1973 1133 1987 1147
rect 2033 1153 2047 1167
rect 2013 1113 2027 1127
rect 1893 1073 1907 1087
rect 2033 1073 2047 1087
rect 1853 1053 1867 1067
rect 1833 1013 1847 1027
rect 1853 953 1867 967
rect 2053 953 2067 967
rect 1833 933 1847 947
rect 1533 813 1547 827
rect 1613 872 1627 886
rect 1673 872 1687 886
rect 1733 872 1747 886
rect 1773 872 1787 886
rect 1593 853 1607 867
rect 1573 793 1587 807
rect 1773 813 1787 827
rect 1633 793 1647 807
rect 1733 793 1747 807
rect 1593 773 1607 787
rect 1613 753 1627 767
rect 1693 753 1707 767
rect 1533 713 1547 727
rect 1413 653 1427 667
rect 1473 593 1487 607
rect 1593 694 1607 708
rect 1633 694 1647 708
rect 1533 553 1547 567
rect 1413 493 1427 507
rect 1353 393 1367 407
rect 993 352 1007 366
rect 1073 352 1087 366
rect 953 313 967 327
rect 1153 352 1167 366
rect 1193 353 1207 367
rect 1253 353 1267 367
rect 1393 433 1407 447
rect 1233 333 1247 347
rect 1193 313 1207 327
rect 1113 293 1127 307
rect 853 253 867 267
rect 913 253 927 267
rect 813 233 827 247
rect 653 153 667 167
rect 793 153 807 167
rect 513 133 527 147
rect 553 132 567 146
rect 593 132 607 146
rect 673 133 687 147
rect 673 93 687 107
rect 353 73 367 87
rect 733 132 747 146
rect 1133 233 1147 247
rect 1113 213 1127 227
rect 853 174 867 188
rect 833 133 847 147
rect 813 93 827 107
rect 873 132 887 146
rect 993 174 1007 188
rect 1013 132 1027 146
rect 1113 174 1127 188
rect 1333 352 1347 366
rect 1373 352 1387 366
rect 1293 333 1307 347
rect 1313 273 1327 287
rect 1253 213 1267 227
rect 1213 174 1227 188
rect 1273 174 1287 188
rect 1453 433 1467 447
rect 1413 393 1427 407
rect 1493 394 1507 408
rect 1533 394 1547 408
rect 1573 394 1587 408
rect 1653 652 1667 666
rect 1633 593 1647 607
rect 1433 352 1447 366
rect 1473 313 1487 327
rect 1453 273 1467 287
rect 1473 253 1487 267
rect 1393 233 1407 247
rect 1453 233 1467 247
rect 1333 193 1347 207
rect 1353 174 1367 188
rect 1413 174 1427 188
rect 1453 174 1467 188
rect 1613 393 1627 407
rect 1713 693 1727 707
rect 1753 773 1767 787
rect 1773 753 1787 767
rect 1753 713 1767 727
rect 1813 833 1827 847
rect 1813 713 1827 727
rect 1993 913 2007 927
rect 2153 1392 2167 1406
rect 2233 1593 2247 1607
rect 2453 1873 2467 1887
rect 2433 1853 2447 1867
rect 2413 1713 2427 1727
rect 2453 1733 2467 1747
rect 2593 2053 2607 2067
rect 2553 1993 2567 2007
rect 2593 1954 2607 1968
rect 2533 1912 2547 1926
rect 2513 1873 2527 1887
rect 2493 1853 2507 1867
rect 2513 1793 2527 1807
rect 2333 1673 2347 1687
rect 2333 1633 2347 1647
rect 2293 1593 2307 1607
rect 2253 1553 2267 1567
rect 2213 1513 2227 1527
rect 2253 1513 2267 1527
rect 2193 1373 2207 1387
rect 2253 1434 2267 1448
rect 2273 1392 2287 1406
rect 2313 1393 2327 1407
rect 2253 1373 2267 1387
rect 2213 1313 2227 1327
rect 2233 1293 2247 1307
rect 2213 1253 2227 1267
rect 2113 1213 2127 1227
rect 2173 1214 2187 1228
rect 2233 1233 2247 1247
rect 2273 1353 2287 1367
rect 2133 1172 2147 1186
rect 2113 1113 2127 1127
rect 2133 1093 2147 1107
rect 2153 1073 2167 1087
rect 2253 1173 2267 1187
rect 2253 1073 2267 1087
rect 2193 1053 2207 1067
rect 2153 1033 2167 1047
rect 2233 1033 2247 1047
rect 2133 953 2147 967
rect 2093 934 2107 948
rect 2093 913 2107 927
rect 2213 914 2227 928
rect 2293 1313 2307 1327
rect 2373 1573 2387 1587
rect 2353 1473 2367 1487
rect 2433 1693 2447 1707
rect 2473 1673 2487 1687
rect 2513 1673 2527 1687
rect 2392 1553 2406 1567
rect 2413 1553 2427 1567
rect 2433 1513 2447 1527
rect 2413 1493 2427 1507
rect 2393 1473 2407 1487
rect 2353 1433 2367 1447
rect 2553 1893 2567 1907
rect 2533 1653 2547 1667
rect 2493 1633 2507 1647
rect 2353 1393 2367 1407
rect 2333 1353 2347 1367
rect 2353 1333 2367 1347
rect 2473 1393 2487 1407
rect 2533 1593 2547 1607
rect 2533 1533 2547 1547
rect 2733 2474 2747 2488
rect 2713 2432 2727 2446
rect 2653 2313 2667 2327
rect 2793 2833 2807 2847
rect 2833 2813 2847 2827
rect 2833 2774 2847 2788
rect 2813 2732 2827 2746
rect 2933 2993 2947 3007
rect 2973 2994 2987 3008
rect 2913 2952 2927 2966
rect 2913 2853 2927 2867
rect 2853 2693 2867 2707
rect 2893 2693 2907 2707
rect 2873 2593 2887 2607
rect 2793 2533 2807 2547
rect 2833 2474 2847 2488
rect 2953 2952 2967 2966
rect 3273 3593 3287 3607
rect 3273 3533 3287 3547
rect 3513 4293 3527 4307
rect 3473 4153 3487 4167
rect 3813 4812 3827 4826
rect 3793 4733 3807 4747
rect 3773 4513 3787 4527
rect 3813 4593 3827 4607
rect 3793 4493 3807 4507
rect 3893 5053 3907 5067
rect 3873 4693 3887 4707
rect 3873 4672 3887 4686
rect 3973 5353 3987 5367
rect 3973 5253 3987 5267
rect 4233 5572 4247 5586
rect 4153 5533 4167 5547
rect 4073 5493 4087 5507
rect 4193 5473 4207 5487
rect 4093 5413 4107 5427
rect 4053 5374 4067 5388
rect 4093 5374 4107 5388
rect 4073 5293 4087 5307
rect 4013 5173 4027 5187
rect 3993 5153 4007 5167
rect 3973 5113 3987 5127
rect 4033 5113 4047 5127
rect 3993 5073 4007 5087
rect 4053 5093 4067 5107
rect 3973 4973 3987 4987
rect 4053 5033 4067 5047
rect 4013 5013 4027 5027
rect 3993 4953 4007 4967
rect 3953 4873 3967 4887
rect 3973 4854 3987 4868
rect 3913 4753 3927 4767
rect 3973 4713 3987 4727
rect 3993 4653 4007 4667
rect 3913 4633 3927 4647
rect 3893 4593 3907 4607
rect 3933 4554 3947 4568
rect 3972 4554 3986 4568
rect 4173 5313 4187 5327
rect 4113 5113 4127 5127
rect 4153 5093 4167 5107
rect 4113 5074 4127 5088
rect 4133 5032 4147 5046
rect 4093 5013 4107 5027
rect 4133 4993 4147 5007
rect 4073 4953 4087 4967
rect 4113 4933 4127 4947
rect 4113 4873 4127 4887
rect 4053 4854 4067 4868
rect 4193 5033 4207 5047
rect 4153 4953 4167 4967
rect 4133 4834 4147 4848
rect 4093 4693 4107 4707
rect 4193 4933 4207 4947
rect 4393 5473 4407 5487
rect 4493 5473 4507 5487
rect 4533 5473 4547 5487
rect 4393 5433 4407 5447
rect 4333 5413 4347 5427
rect 4293 5373 4307 5387
rect 4373 5373 4387 5387
rect 4253 5293 4267 5307
rect 4413 5413 4427 5427
rect 4493 5413 4507 5427
rect 4453 5374 4467 5388
rect 4353 5332 4367 5346
rect 4392 5332 4406 5346
rect 4413 5333 4427 5347
rect 4313 5313 4327 5327
rect 4513 5332 4527 5346
rect 4533 5313 4547 5327
rect 4473 5293 4487 5307
rect 4412 5253 4426 5267
rect 4433 5253 4447 5267
rect 4293 5173 4307 5187
rect 4413 5173 4427 5187
rect 4273 5093 4287 5107
rect 4333 5133 4347 5147
rect 4293 5074 4307 5088
rect 4273 5032 4287 5046
rect 4233 4993 4247 5007
rect 4353 5093 4367 5107
rect 4453 5093 4467 5107
rect 4353 5033 4367 5047
rect 4413 5013 4427 5027
rect 4433 4993 4447 5007
rect 4473 4993 4487 5007
rect 4413 4953 4427 4967
rect 4233 4933 4247 4947
rect 4333 4933 4347 4947
rect 4393 4933 4407 4947
rect 4213 4893 4227 4907
rect 4393 4833 4407 4847
rect 4473 4833 4487 4847
rect 4653 6092 4667 6106
rect 4793 6092 4807 6106
rect 5033 6253 5047 6267
rect 5073 6253 5087 6267
rect 5033 6173 5047 6187
rect 5033 6152 5047 6166
rect 4713 6053 4727 6067
rect 4793 6013 4807 6027
rect 4673 5993 4687 6007
rect 4653 5894 4667 5908
rect 4633 5793 4647 5807
rect 4633 5753 4647 5767
rect 4593 5713 4607 5727
rect 4633 5673 4647 5687
rect 4633 5633 4647 5647
rect 4573 5613 4587 5627
rect 4733 5933 4747 5947
rect 4833 5993 4847 6007
rect 5053 6133 5067 6147
rect 4853 5973 4867 5987
rect 5053 6093 5067 6107
rect 5293 6153 5307 6167
rect 5133 6073 5147 6087
rect 4893 5953 4907 5967
rect 4973 5953 4987 5967
rect 4873 5913 4887 5927
rect 4953 5893 4967 5907
rect 4753 5852 4767 5866
rect 4793 5852 4807 5866
rect 5073 5933 5087 5947
rect 5033 5894 5047 5908
rect 4713 5793 4727 5807
rect 4793 5693 4807 5707
rect 4673 5653 4687 5667
rect 4793 5613 4807 5627
rect 4653 5594 4667 5608
rect 4573 5573 4587 5587
rect 4613 5573 4627 5587
rect 4613 5533 4627 5547
rect 4593 5332 4607 5346
rect 4753 5594 4767 5608
rect 4733 5552 4747 5566
rect 4753 5473 4767 5487
rect 4733 5413 4747 5427
rect 4733 5374 4747 5388
rect 4653 5313 4667 5327
rect 4693 5313 4707 5327
rect 4753 5313 4767 5327
rect 4653 5273 4667 5287
rect 4613 5213 4627 5227
rect 4573 5153 4587 5167
rect 4553 5093 4567 5107
rect 4533 5073 4547 5087
rect 4593 5093 4607 5107
rect 4373 4813 4387 4827
rect 4233 4733 4247 4747
rect 4233 4693 4247 4707
rect 4053 4633 4067 4647
rect 4173 4633 4187 4647
rect 3993 4553 4007 4567
rect 4093 4573 4107 4587
rect 4173 4573 4187 4587
rect 3873 4512 3887 4526
rect 3913 4512 3927 4526
rect 3973 4513 3987 4527
rect 3773 4433 3787 4447
rect 3633 4413 3647 4427
rect 3753 4413 3767 4427
rect 3613 4353 3627 4367
rect 3612 4313 3626 4327
rect 3612 4273 3626 4287
rect 3633 4273 3647 4287
rect 3573 4233 3587 4247
rect 3793 4313 3807 4327
rect 3793 4253 3807 4267
rect 3773 4233 3787 4247
rect 3913 4313 3927 4327
rect 3993 4473 4007 4487
rect 4033 4512 4047 4526
rect 4013 4413 4027 4427
rect 4072 4473 4086 4487
rect 4093 4473 4107 4487
rect 4093 4433 4107 4447
rect 4133 4433 4147 4447
rect 4193 4493 4207 4507
rect 4173 4413 4187 4427
rect 4473 4733 4487 4747
rect 4373 4633 4387 4647
rect 4373 4553 4387 4567
rect 4553 4753 4567 4767
rect 4973 5852 4987 5866
rect 4893 5833 4907 5847
rect 4873 5793 4887 5807
rect 4853 5713 4867 5727
rect 5013 5793 5027 5807
rect 5053 5773 5067 5787
rect 5173 5933 5187 5947
rect 5213 5894 5227 5908
rect 5353 6114 5367 6128
rect 5393 6114 5407 6128
rect 5333 6033 5347 6047
rect 5253 5933 5267 5947
rect 5473 6114 5487 6128
rect 5553 6114 5567 6128
rect 5593 6114 5607 6128
rect 5393 6073 5407 6087
rect 5453 6072 5467 6086
rect 5353 5993 5367 6007
rect 5373 5894 5387 5908
rect 5153 5852 5167 5866
rect 5053 5733 5067 5747
rect 5113 5733 5127 5747
rect 5013 5693 5027 5707
rect 4853 5673 4867 5687
rect 4893 5673 4907 5687
rect 4833 5653 4847 5667
rect 4933 5594 4947 5608
rect 4913 5573 4927 5587
rect 4853 5513 4867 5527
rect 4833 5453 4847 5467
rect 4813 5373 4827 5387
rect 4793 5193 4807 5207
rect 4913 5493 4927 5507
rect 4993 5552 5007 5566
rect 5153 5693 5167 5707
rect 5073 5673 5087 5687
rect 5013 5533 5027 5547
rect 5053 5533 5067 5547
rect 4893 5393 4907 5407
rect 4873 5374 4887 5388
rect 4853 5173 4867 5187
rect 4833 5153 4847 5167
rect 4693 5133 4707 5147
rect 4773 5113 4787 5127
rect 4833 5074 4847 5088
rect 4973 5453 4987 5467
rect 5113 5594 5127 5608
rect 5253 5853 5267 5867
rect 5313 5852 5327 5866
rect 5233 5813 5247 5827
rect 5313 5793 5327 5807
rect 5233 5713 5247 5727
rect 5233 5673 5247 5687
rect 5253 5653 5267 5667
rect 5193 5633 5207 5647
rect 5173 5552 5187 5566
rect 5073 5513 5087 5527
rect 5133 5513 5147 5527
rect 5253 5553 5267 5567
rect 5213 5493 5227 5507
rect 5472 5993 5486 6007
rect 5493 5993 5507 6007
rect 5433 5894 5447 5908
rect 5513 5933 5527 5947
rect 5533 5893 5547 5907
rect 5413 5853 5427 5867
rect 5453 5852 5467 5866
rect 5413 5793 5427 5807
rect 5393 5773 5407 5787
rect 5373 5753 5387 5767
rect 5493 5713 5507 5727
rect 5453 5673 5467 5687
rect 5573 6073 5587 6087
rect 5613 6072 5627 6086
rect 5693 6193 5707 6207
rect 5733 6193 5747 6207
rect 5773 6133 5787 6147
rect 5713 6072 5727 6086
rect 5673 6033 5687 6047
rect 5593 5993 5607 6007
rect 5633 5993 5647 6007
rect 5753 5993 5767 6007
rect 5573 5953 5587 5967
rect 6033 6193 6047 6207
rect 5993 6153 6007 6167
rect 5933 6133 5947 6147
rect 5833 6113 5847 6127
rect 6153 6153 6167 6167
rect 6093 6133 6107 6147
rect 6033 6114 6047 6128
rect 6073 6113 6087 6127
rect 5853 6072 5867 6086
rect 5893 6072 5907 6086
rect 5933 6072 5947 6086
rect 6012 6033 6026 6047
rect 6033 6033 6047 6047
rect 5853 6013 5867 6027
rect 5973 6013 5987 6027
rect 5813 5933 5827 5947
rect 5633 5914 5647 5928
rect 5573 5893 5587 5907
rect 5613 5893 5627 5907
rect 5693 5894 5707 5908
rect 5753 5894 5767 5908
rect 5633 5852 5647 5866
rect 5613 5813 5627 5827
rect 5573 5753 5587 5767
rect 5553 5653 5567 5667
rect 5953 5933 5967 5947
rect 5913 5913 5927 5927
rect 5913 5894 5927 5908
rect 6013 5913 6027 5927
rect 5693 5793 5707 5807
rect 5673 5673 5687 5687
rect 5553 5613 5567 5627
rect 5613 5614 5627 5628
rect 5313 5473 5327 5487
rect 5173 5453 5187 5467
rect 5273 5453 5287 5467
rect 5133 5433 5147 5447
rect 5053 5393 5067 5407
rect 5113 5393 5127 5407
rect 5573 5572 5587 5586
rect 5853 5853 5867 5867
rect 5893 5852 5907 5866
rect 5793 5813 5807 5827
rect 5933 5813 5947 5827
rect 5833 5713 5847 5727
rect 5753 5653 5767 5667
rect 5813 5593 5827 5607
rect 5893 5673 5907 5687
rect 5973 5613 5987 5627
rect 6253 6133 6267 6147
rect 6173 6072 6187 6086
rect 6273 6072 6287 6086
rect 6133 6033 6147 6047
rect 6093 5913 6107 5927
rect 6153 5893 6167 5907
rect 6193 5894 6207 5908
rect 6093 5852 6107 5866
rect 6033 5653 6047 5667
rect 6033 5613 6047 5627
rect 5933 5594 5947 5608
rect 6013 5594 6027 5608
rect 6233 5852 6247 5866
rect 6153 5673 6167 5687
rect 6093 5573 6107 5587
rect 5673 5552 5687 5566
rect 5733 5552 5747 5566
rect 5773 5552 5787 5566
rect 5812 5552 5826 5566
rect 5833 5552 5847 5566
rect 5873 5513 5887 5527
rect 6053 5552 6067 5566
rect 6193 5594 6207 5608
rect 5913 5473 5927 5487
rect 5913 5433 5927 5447
rect 5013 5313 5027 5327
rect 5053 5313 5067 5327
rect 4913 5273 4927 5287
rect 4953 5213 4967 5227
rect 4933 5193 4947 5207
rect 4873 5073 4887 5087
rect 4953 5173 4967 5187
rect 4993 5073 5007 5087
rect 5113 5253 5127 5267
rect 5073 5153 5087 5167
rect 5553 5353 5567 5367
rect 5513 5312 5527 5326
rect 5573 5312 5587 5326
rect 5453 5273 5467 5287
rect 5493 5273 5507 5287
rect 5353 5213 5367 5227
rect 5393 5213 5407 5227
rect 5333 5153 5347 5167
rect 5313 5133 5327 5147
rect 5233 5113 5247 5127
rect 5293 5113 5307 5127
rect 4773 5013 4787 5027
rect 4913 5032 4927 5046
rect 4953 5032 4967 5046
rect 4993 5032 5007 5046
rect 5033 5032 5047 5046
rect 5093 5032 5107 5046
rect 4653 4993 4667 5007
rect 4813 4993 4827 5007
rect 4933 4993 4947 5007
rect 4613 4953 4627 4967
rect 4713 4933 4727 4947
rect 4913 4913 4927 4927
rect 4753 4893 4767 4907
rect 4893 4893 4907 4907
rect 4813 4854 4827 4868
rect 4853 4854 4867 4868
rect 4693 4812 4707 4826
rect 4753 4812 4767 4826
rect 4793 4812 4807 4826
rect 4653 4793 4667 4807
rect 4633 4753 4647 4767
rect 4593 4733 4607 4747
rect 4533 4693 4547 4707
rect 4873 4812 4887 4826
rect 4753 4673 4767 4687
rect 4833 4673 4847 4687
rect 4653 4633 4667 4647
rect 4533 4574 4547 4588
rect 4593 4574 4607 4588
rect 4473 4493 4487 4507
rect 4473 4472 4487 4486
rect 4273 4433 4287 4447
rect 4153 4373 4167 4387
rect 4233 4373 4247 4387
rect 4093 4353 4107 4367
rect 3933 4272 3947 4286
rect 3913 4213 3927 4227
rect 3613 4133 3627 4147
rect 3653 4133 3667 4147
rect 3513 4073 3527 4087
rect 3493 4053 3507 4067
rect 3493 4013 3507 4027
rect 3473 3993 3487 4007
rect 3453 3813 3467 3827
rect 3753 4113 3767 4127
rect 3513 3993 3527 4007
rect 3493 3913 3507 3927
rect 3633 3913 3647 3927
rect 3733 3913 3747 3927
rect 3593 3853 3607 3867
rect 3573 3813 3587 3827
rect 3453 3753 3467 3767
rect 3433 3653 3447 3667
rect 3353 3613 3367 3627
rect 3293 3453 3307 3467
rect 3253 3333 3267 3347
rect 3313 3393 3327 3407
rect 3233 3313 3247 3327
rect 3033 3294 3047 3308
rect 3153 3294 3167 3308
rect 3153 3233 3167 3247
rect 3073 3213 3087 3227
rect 3113 3213 3127 3227
rect 3073 3173 3087 3187
rect 3093 3153 3107 3167
rect 3093 3053 3107 3067
rect 3133 3133 3147 3147
rect 3133 3053 3147 3067
rect 3173 3093 3187 3107
rect 3153 2973 3167 2987
rect 3093 2952 3107 2966
rect 3013 2893 3027 2907
rect 3053 2893 3067 2907
rect 2953 2873 2967 2887
rect 2933 2774 2947 2788
rect 2973 2774 2987 2788
rect 3013 2774 3027 2788
rect 3073 2853 3087 2867
rect 3133 2933 3147 2947
rect 3133 2893 3147 2907
rect 3093 2813 3107 2827
rect 3133 2813 3147 2827
rect 3073 2773 3087 2787
rect 3353 3492 3367 3506
rect 3573 3773 3587 3787
rect 3553 3733 3567 3747
rect 3733 3853 3747 3867
rect 3673 3814 3687 3828
rect 3693 3772 3707 3786
rect 3653 3753 3667 3767
rect 3593 3713 3607 3727
rect 3493 3673 3507 3687
rect 3653 3673 3667 3687
rect 3593 3633 3607 3647
rect 3493 3613 3507 3627
rect 3593 3573 3607 3587
rect 3593 3552 3607 3566
rect 3353 3413 3367 3427
rect 3433 3373 3447 3387
rect 3353 3313 3367 3327
rect 3253 3253 3267 3267
rect 3233 3113 3247 3127
rect 3293 3213 3307 3227
rect 3373 3293 3387 3307
rect 3613 3492 3627 3506
rect 3713 3653 3727 3667
rect 3673 3573 3687 3587
rect 3673 3533 3687 3547
rect 3693 3492 3707 3506
rect 3613 3453 3627 3467
rect 3633 3433 3647 3447
rect 3513 3353 3527 3367
rect 3593 3353 3607 3367
rect 3493 3293 3507 3307
rect 3453 3252 3467 3266
rect 3413 3233 3427 3247
rect 3373 3213 3387 3227
rect 3273 3113 3287 3127
rect 3313 3113 3327 3127
rect 3353 3113 3367 3127
rect 3253 3053 3267 3067
rect 3393 3093 3407 3107
rect 3433 3173 3447 3187
rect 3473 3233 3487 3247
rect 3453 3153 3467 3167
rect 3573 3313 3587 3327
rect 3513 3233 3527 3247
rect 3553 3233 3567 3247
rect 3813 4054 3827 4068
rect 3773 4012 3787 4026
rect 3793 3993 3807 4007
rect 3773 3873 3787 3887
rect 3873 4073 3887 4087
rect 3973 4233 3987 4247
rect 3953 4193 3967 4207
rect 3933 4054 3947 4068
rect 4013 4293 4027 4307
rect 3993 4113 4007 4127
rect 3973 4073 3987 4087
rect 3993 4053 4007 4067
rect 4073 4292 4087 4306
rect 4113 4292 4127 4306
rect 4213 4334 4227 4348
rect 4153 4272 4167 4286
rect 4213 4273 4227 4287
rect 4073 4253 4087 4267
rect 4193 4253 4207 4267
rect 4053 4233 4067 4247
rect 4033 4213 4047 4227
rect 4033 4093 4047 4107
rect 4013 4033 4027 4047
rect 3893 4013 3907 4027
rect 3873 3993 3887 4007
rect 3913 3993 3927 4007
rect 3973 3992 3987 4006
rect 3933 3953 3947 3967
rect 4013 3953 4027 3967
rect 3913 3933 3927 3947
rect 3993 3913 4007 3927
rect 3773 3833 3787 3847
rect 3813 3814 3827 3828
rect 3933 3814 3947 3828
rect 3873 3793 3887 3807
rect 3753 3772 3767 3786
rect 3753 3673 3767 3687
rect 3733 3493 3747 3507
rect 3733 3433 3747 3447
rect 3713 3413 3727 3427
rect 3833 3772 3847 3786
rect 3893 3713 3907 3727
rect 3793 3573 3807 3587
rect 3833 3553 3847 3567
rect 3873 3514 3887 3528
rect 3813 3472 3827 3486
rect 3873 3453 3887 3467
rect 3833 3433 3847 3447
rect 3693 3333 3707 3347
rect 3753 3393 3767 3407
rect 3733 3293 3747 3307
rect 3633 3213 3647 3227
rect 3493 3193 3507 3207
rect 3593 3193 3607 3207
rect 3433 3093 3447 3107
rect 3413 3073 3427 3087
rect 3433 3053 3447 3067
rect 3393 3033 3407 3047
rect 3373 2994 3387 3008
rect 3193 2973 3207 2987
rect 3313 2973 3327 2987
rect 3173 2933 3187 2947
rect 3173 2912 3187 2926
rect 3153 2793 3167 2807
rect 3193 2873 3207 2887
rect 3213 2813 3227 2827
rect 2933 2733 2947 2747
rect 2913 2492 2927 2506
rect 2893 2473 2907 2487
rect 2853 2432 2867 2446
rect 2893 2433 2907 2447
rect 2793 2373 2807 2387
rect 2833 2373 2847 2387
rect 2793 2254 2807 2268
rect 2633 2093 2647 2107
rect 2813 2212 2827 2226
rect 2733 2173 2747 2187
rect 2693 2153 2707 2167
rect 2693 1993 2707 2007
rect 2673 1973 2687 1987
rect 2653 1954 2667 1968
rect 2673 1912 2687 1926
rect 2613 1893 2627 1907
rect 2633 1833 2647 1847
rect 2593 1773 2607 1787
rect 2633 1773 2647 1787
rect 2713 1733 2727 1747
rect 2593 1633 2607 1647
rect 2673 1673 2687 1687
rect 2653 1653 2667 1667
rect 2613 1533 2627 1547
rect 2613 1512 2627 1526
rect 2553 1453 2567 1467
rect 2613 1433 2627 1447
rect 2493 1373 2507 1387
rect 2373 1313 2387 1327
rect 2413 1313 2427 1327
rect 2493 1313 2507 1327
rect 2413 1292 2427 1306
rect 2333 1253 2347 1267
rect 2393 1253 2407 1267
rect 2293 1213 2307 1227
rect 2373 1214 2387 1228
rect 2433 1253 2447 1267
rect 2413 1193 2427 1207
rect 2293 1173 2307 1187
rect 2273 1033 2287 1047
rect 2273 993 2287 1007
rect 2253 913 2267 927
rect 2033 873 2047 887
rect 1893 813 1907 827
rect 1893 773 1907 787
rect 1933 773 1947 787
rect 2013 773 2027 787
rect 1913 753 1927 767
rect 1973 753 1987 767
rect 1932 733 1946 747
rect 1953 733 1967 747
rect 1933 694 1947 708
rect 1993 713 2007 727
rect 1853 673 1867 687
rect 1773 652 1787 666
rect 1813 652 1827 666
rect 1713 613 1727 627
rect 1853 593 1867 607
rect 1913 652 1927 666
rect 1993 652 2007 666
rect 1873 553 1887 567
rect 1793 473 1807 487
rect 1653 433 1667 447
rect 1693 413 1707 427
rect 1653 393 1667 407
rect 1733 394 1747 408
rect 1633 353 1647 367
rect 1593 333 1607 347
rect 1653 313 1667 327
rect 1753 352 1767 366
rect 1713 253 1727 267
rect 1553 233 1567 247
rect 1573 213 1587 227
rect 1653 213 1667 227
rect 1753 213 1767 227
rect 1553 193 1567 207
rect 1093 132 1107 146
rect 1133 132 1147 146
rect 1193 133 1207 147
rect 913 73 927 87
rect 693 53 707 67
rect 833 53 847 67
rect 1513 173 1527 187
rect 1613 174 1627 188
rect 1233 113 1247 127
rect 1213 93 1227 107
rect 1293 132 1307 146
rect 1253 53 1267 67
rect 1393 132 1407 146
rect 1373 53 1387 67
rect 1093 33 1107 47
rect 1353 33 1367 47
rect 1393 33 1407 47
rect 1473 113 1487 127
rect 1433 93 1447 107
rect 1473 73 1487 87
rect 1713 193 1727 207
rect 1733 173 1747 187
rect 1553 132 1567 146
rect 1653 133 1667 147
rect 1693 132 1707 146
rect 1593 93 1607 107
rect 1453 53 1467 67
rect 1493 53 1507 67
rect 1573 73 1587 87
rect 1613 73 1627 87
rect 1553 53 1567 67
rect 1633 53 1647 67
rect 2133 873 2147 887
rect 2173 873 2187 887
rect 2073 773 2087 787
rect 2113 773 2127 787
rect 2173 833 2187 847
rect 2133 753 2147 767
rect 2113 713 2127 727
rect 2093 694 2107 708
rect 2193 793 2207 807
rect 2173 693 2187 707
rect 2033 613 2047 627
rect 1813 394 1827 408
rect 1853 394 1867 408
rect 1893 394 1907 408
rect 1953 413 1967 427
rect 2013 413 2027 427
rect 1933 393 1947 407
rect 1833 353 1847 367
rect 1813 313 1827 327
rect 1873 313 1887 327
rect 1913 313 1927 327
rect 1893 293 1907 307
rect 1873 273 1887 287
rect 1833 253 1847 267
rect 1833 213 1847 227
rect 1793 173 1807 187
rect 1913 213 1927 227
rect 2093 593 2107 607
rect 2073 393 2087 407
rect 2013 352 2027 366
rect 2013 253 2027 267
rect 1973 213 1987 227
rect 1953 193 1967 207
rect 1933 173 1947 187
rect 2153 652 2167 666
rect 2353 1172 2367 1186
rect 2393 1173 2407 1187
rect 2453 1213 2467 1227
rect 2593 1392 2607 1406
rect 2573 1353 2587 1367
rect 2553 1293 2567 1307
rect 2433 1172 2447 1186
rect 2473 1172 2487 1186
rect 2513 1172 2527 1186
rect 2473 1133 2487 1147
rect 2313 1113 2327 1127
rect 2413 1073 2427 1087
rect 2313 1033 2327 1047
rect 2392 993 2406 1007
rect 2413 993 2427 1007
rect 2353 914 2367 928
rect 2453 953 2467 967
rect 2433 914 2447 928
rect 2293 853 2307 867
rect 2333 853 2347 867
rect 2293 813 2307 827
rect 2273 793 2287 807
rect 2233 753 2247 767
rect 2253 733 2267 747
rect 2253 694 2267 708
rect 2213 653 2227 667
rect 2493 914 2507 928
rect 2553 914 2567 928
rect 2473 853 2487 867
rect 2453 833 2467 847
rect 2313 793 2327 807
rect 2373 793 2387 807
rect 2433 793 2447 807
rect 2413 773 2427 787
rect 2373 753 2387 767
rect 2333 694 2347 708
rect 2413 713 2427 727
rect 2293 652 2307 666
rect 2353 652 2367 666
rect 2153 613 2167 627
rect 2193 613 2207 627
rect 2232 613 2246 627
rect 2253 613 2267 627
rect 2233 573 2247 587
rect 2113 553 2127 567
rect 2133 513 2147 527
rect 2113 413 2127 427
rect 2213 453 2227 467
rect 2233 433 2247 447
rect 2133 393 2147 407
rect 2173 394 2187 408
rect 2213 413 2227 427
rect 2393 573 2407 587
rect 2273 453 2287 467
rect 2313 453 2327 467
rect 2373 453 2387 467
rect 2273 394 2287 408
rect 2793 2073 2807 2087
rect 2753 2053 2767 2067
rect 3053 2733 3067 2747
rect 3053 2712 3067 2726
rect 2993 2693 3007 2707
rect 3013 2474 3027 2488
rect 3193 2733 3207 2747
rect 3113 2693 3127 2707
rect 3193 2693 3207 2707
rect 3153 2673 3167 2687
rect 3073 2653 3087 2667
rect 3133 2653 3147 2667
rect 3133 2593 3147 2607
rect 3073 2573 3087 2587
rect 3053 2473 3067 2487
rect 2933 2433 2947 2447
rect 2993 2413 3007 2427
rect 2953 2333 2967 2347
rect 2913 2273 2927 2287
rect 2933 2254 2947 2268
rect 2973 2313 2987 2327
rect 3013 2313 3027 2327
rect 2913 2212 2927 2226
rect 2953 2213 2967 2227
rect 2953 2173 2967 2187
rect 2993 2273 3007 2287
rect 3253 2893 3267 2907
rect 3273 2873 3287 2887
rect 3512 3093 3526 3107
rect 3533 3093 3547 3107
rect 3593 3093 3607 3107
rect 3513 3013 3527 3027
rect 3493 2994 3507 3008
rect 3573 3053 3587 3067
rect 3573 2993 3587 3007
rect 3353 2873 3367 2887
rect 3393 2873 3407 2887
rect 3273 2833 3287 2847
rect 3313 2833 3327 2847
rect 3373 2833 3387 2847
rect 3233 2773 3247 2787
rect 3313 2812 3327 2826
rect 3353 2774 3367 2788
rect 3233 2732 3247 2746
rect 3293 2732 3307 2746
rect 3333 2732 3347 2746
rect 3253 2693 3267 2707
rect 3213 2573 3227 2587
rect 3193 2553 3207 2567
rect 3133 2533 3147 2547
rect 3173 2533 3187 2547
rect 3093 2493 3107 2507
rect 3133 2474 3147 2488
rect 3213 2513 3227 2527
rect 3273 2613 3287 2627
rect 3353 2553 3367 2567
rect 3373 2513 3387 2527
rect 3313 2474 3327 2488
rect 3413 2813 3427 2827
rect 3393 2493 3407 2507
rect 3473 2953 3487 2967
rect 3513 2952 3527 2966
rect 3473 2913 3487 2927
rect 3453 2893 3467 2907
rect 3733 3253 3747 3267
rect 3713 3213 3727 3227
rect 3733 3153 3747 3167
rect 3693 3113 3707 3127
rect 3673 3073 3687 3087
rect 3653 3013 3667 3027
rect 3673 2952 3687 2966
rect 3613 2913 3627 2927
rect 3653 2913 3667 2927
rect 3593 2873 3607 2887
rect 3553 2833 3567 2847
rect 3493 2813 3507 2827
rect 3553 2793 3567 2807
rect 3493 2774 3507 2788
rect 3533 2774 3547 2788
rect 3633 2793 3647 2807
rect 3453 2693 3467 2707
rect 3513 2693 3527 2707
rect 3433 2653 3447 2667
rect 3113 2433 3127 2447
rect 3093 2413 3107 2427
rect 3093 2333 3107 2347
rect 3033 2293 3047 2307
rect 3093 2293 3107 2307
rect 3153 2393 3167 2407
rect 3133 2273 3147 2287
rect 3093 2253 3107 2267
rect 2993 2233 3007 2247
rect 2993 2193 3007 2207
rect 2993 2172 3007 2186
rect 2873 2153 2887 2167
rect 2933 2153 2947 2167
rect 2873 2113 2887 2127
rect 2873 2053 2887 2067
rect 2833 1992 2847 2006
rect 2773 1873 2787 1887
rect 2753 1833 2767 1847
rect 2773 1813 2787 1827
rect 2793 1734 2807 1748
rect 2973 2153 2987 2167
rect 3073 2133 3087 2147
rect 3013 2093 3027 2107
rect 2973 2073 2987 2087
rect 2953 2053 2967 2067
rect 2973 2033 2987 2047
rect 3013 2033 3027 2047
rect 2993 1993 3007 2007
rect 2953 1912 2967 1926
rect 2993 1913 3007 1927
rect 2893 1853 2907 1867
rect 2873 1793 2887 1807
rect 2973 1853 2987 1867
rect 2913 1773 2927 1787
rect 2953 1773 2967 1787
rect 2733 1673 2747 1687
rect 2813 1693 2827 1707
rect 2793 1673 2807 1687
rect 2713 1653 2727 1667
rect 2773 1653 2787 1667
rect 2693 1533 2707 1547
rect 2673 1473 2687 1487
rect 2653 1353 2667 1367
rect 2633 1273 2647 1287
rect 2613 1253 2627 1267
rect 2613 1214 2627 1228
rect 2633 1172 2647 1186
rect 2733 1392 2747 1406
rect 2693 1373 2707 1387
rect 2733 1353 2747 1367
rect 2713 1293 2727 1307
rect 2813 1613 2827 1627
rect 2873 1734 2887 1748
rect 2913 1734 2927 1748
rect 2853 1713 2867 1727
rect 2853 1673 2867 1687
rect 2853 1513 2867 1527
rect 2973 1692 2987 1706
rect 2973 1573 2987 1587
rect 2893 1533 2907 1547
rect 2953 1533 2967 1547
rect 2853 1473 2867 1487
rect 2853 1452 2867 1466
rect 2933 1473 2947 1487
rect 2793 1393 2807 1407
rect 2793 1353 2807 1367
rect 2773 1233 2787 1247
rect 2753 1214 2767 1228
rect 2793 1213 2807 1227
rect 2693 1173 2707 1187
rect 2593 1133 2607 1147
rect 2573 813 2587 827
rect 2613 914 2627 928
rect 2653 872 2667 886
rect 2613 853 2627 867
rect 2593 733 2607 747
rect 2473 652 2487 666
rect 2473 613 2487 627
rect 2513 593 2527 607
rect 2573 694 2587 708
rect 2653 694 2667 708
rect 2793 1173 2807 1187
rect 2773 1133 2787 1147
rect 2793 1093 2807 1107
rect 2893 1434 2907 1448
rect 2833 1393 2847 1407
rect 2873 1373 2887 1387
rect 2893 1293 2907 1307
rect 2853 1213 2867 1227
rect 2933 1253 2947 1267
rect 2973 1513 2987 1527
rect 3053 1954 3067 1968
rect 3113 2173 3127 2187
rect 3273 2433 3287 2447
rect 3333 2432 3347 2446
rect 3213 2393 3227 2407
rect 3293 2393 3307 2407
rect 3193 2333 3207 2347
rect 3213 2293 3227 2307
rect 3273 2293 3287 2307
rect 3173 2273 3187 2287
rect 3253 2253 3267 2267
rect 3233 2212 3247 2226
rect 3333 2333 3347 2347
rect 3313 2212 3327 2226
rect 3353 2193 3367 2207
rect 3273 2173 3287 2187
rect 3313 2153 3327 2167
rect 3293 2133 3307 2147
rect 3293 2053 3307 2067
rect 3193 2033 3207 2047
rect 3253 1993 3267 2007
rect 3132 1953 3146 1967
rect 3153 1953 3167 1967
rect 3193 1954 3207 1968
rect 3113 1912 3127 1926
rect 3153 1912 3167 1926
rect 3213 1912 3227 1926
rect 3073 1853 3087 1867
rect 3133 1853 3147 1867
rect 3053 1813 3067 1827
rect 3033 1793 3047 1807
rect 3033 1753 3047 1767
rect 3093 1773 3107 1787
rect 3053 1673 3067 1687
rect 3013 1653 3027 1667
rect 2993 1473 3007 1487
rect 3033 1434 3047 1448
rect 3013 1392 3027 1406
rect 2993 1373 3007 1387
rect 2833 1113 2847 1127
rect 2873 1113 2887 1127
rect 2853 1093 2867 1107
rect 2813 1073 2827 1087
rect 2733 1013 2747 1027
rect 2773 953 2787 967
rect 2813 953 2827 967
rect 2853 933 2867 947
rect 2793 872 2807 886
rect 2853 873 2867 886
rect 2853 872 2867 873
rect 2893 1033 2907 1047
rect 2953 1172 2967 1186
rect 2973 1133 2987 1147
rect 3373 2073 3387 2087
rect 3313 2013 3327 2027
rect 3313 1973 3327 1987
rect 3293 1954 3307 1968
rect 3333 1954 3347 1968
rect 3453 2432 3467 2446
rect 3493 2393 3507 2407
rect 3413 2253 3427 2267
rect 3453 2254 3467 2268
rect 3593 2774 3607 2788
rect 3793 3333 3807 3347
rect 3773 3313 3787 3327
rect 3973 3773 3987 3787
rect 3953 3733 3967 3747
rect 3933 3673 3947 3687
rect 3993 3733 4007 3747
rect 3993 3673 4007 3687
rect 3973 3553 3987 3567
rect 3973 3514 3987 3528
rect 4073 4213 4087 4227
rect 4153 4213 4167 4227
rect 4113 4053 4127 4067
rect 4353 4413 4367 4427
rect 4293 4353 4307 4367
rect 4273 4233 4287 4247
rect 4433 4373 4447 4387
rect 4333 4233 4347 4247
rect 4293 4213 4307 4227
rect 4273 4193 4287 4207
rect 4233 4173 4247 4187
rect 4213 4073 4227 4087
rect 4153 4033 4167 4047
rect 4353 4173 4367 4187
rect 4273 4034 4287 4048
rect 4333 4034 4347 4048
rect 4053 3973 4067 3987
rect 4113 3973 4127 3987
rect 4193 3993 4207 4007
rect 4093 3913 4107 3927
rect 4093 3733 4107 3747
rect 4033 3693 4047 3707
rect 4133 3873 4147 3887
rect 4113 3653 4127 3667
rect 4013 3613 4027 3627
rect 3933 3453 3947 3467
rect 3953 3433 3967 3447
rect 3933 3393 3947 3407
rect 3913 3373 3927 3387
rect 3893 3253 3907 3267
rect 3813 3213 3827 3227
rect 3873 3213 3887 3227
rect 3773 3193 3787 3207
rect 3793 3133 3807 3147
rect 3773 3073 3787 3087
rect 3793 3033 3807 3047
rect 3893 3153 3907 3167
rect 3853 3033 3867 3047
rect 3813 2994 3827 3008
rect 4053 3514 4067 3528
rect 4053 3393 4067 3407
rect 3953 3353 3967 3367
rect 4013 3353 4027 3367
rect 4033 3313 4047 3327
rect 3993 3294 4007 3308
rect 3933 3253 3947 3267
rect 3913 3053 3927 3067
rect 3773 2952 3787 2966
rect 3833 2952 3847 2966
rect 3873 2952 3887 2966
rect 3833 2913 3847 2927
rect 3873 2913 3887 2927
rect 3753 2893 3767 2907
rect 3813 2893 3827 2907
rect 3753 2872 3767 2886
rect 3713 2853 3727 2867
rect 3673 2833 3687 2847
rect 3693 2813 3707 2827
rect 3533 2673 3547 2687
rect 3613 2732 3627 2746
rect 3673 2733 3687 2747
rect 3673 2712 3687 2726
rect 3593 2613 3607 2627
rect 3653 2613 3667 2627
rect 3653 2573 3667 2587
rect 3673 2553 3687 2567
rect 3633 2533 3647 2547
rect 3693 2533 3707 2547
rect 3573 2432 3587 2446
rect 3633 2373 3647 2387
rect 3613 2353 3627 2367
rect 3593 2333 3607 2347
rect 3633 2313 3647 2327
rect 3413 2213 3427 2227
rect 3473 2193 3487 2207
rect 3473 2153 3487 2167
rect 3473 2093 3487 2107
rect 3413 1993 3427 2007
rect 3513 2073 3527 2087
rect 3593 2254 3607 2268
rect 3693 2432 3707 2446
rect 3773 2713 3787 2727
rect 3733 2653 3747 2667
rect 3873 2833 3887 2847
rect 3833 2773 3847 2787
rect 3913 2793 3927 2807
rect 3893 2732 3907 2746
rect 3873 2713 3887 2727
rect 3853 2693 3867 2707
rect 3913 2673 3927 2687
rect 3813 2633 3827 2647
rect 3733 2573 3747 2587
rect 3793 2573 3807 2587
rect 3773 2474 3787 2488
rect 3753 2432 3767 2446
rect 3673 2333 3687 2347
rect 3713 2333 3727 2347
rect 3653 2293 3667 2307
rect 3653 2253 3667 2267
rect 3573 2212 3587 2226
rect 3553 2193 3567 2207
rect 3533 1993 3547 2007
rect 3353 1912 3367 1926
rect 3393 1913 3407 1927
rect 3253 1893 3267 1907
rect 3313 1893 3327 1907
rect 3213 1833 3227 1847
rect 3293 1813 3307 1827
rect 3393 1813 3407 1827
rect 3233 1773 3247 1787
rect 3193 1753 3207 1767
rect 3233 1734 3247 1748
rect 3193 1613 3207 1627
rect 3173 1573 3187 1587
rect 3153 1553 3167 1567
rect 3173 1533 3187 1547
rect 3093 1453 3107 1467
rect 3132 1453 3146 1467
rect 3153 1453 3167 1467
rect 3073 1293 3087 1307
rect 3113 1433 3127 1447
rect 3173 1434 3187 1448
rect 3253 1692 3267 1706
rect 3353 1734 3367 1748
rect 3313 1693 3327 1707
rect 3293 1673 3307 1687
rect 3293 1652 3307 1666
rect 3213 1513 3227 1527
rect 3113 1393 3127 1407
rect 3253 1434 3267 1448
rect 3313 1613 3327 1627
rect 3393 1693 3407 1707
rect 3352 1673 3366 1687
rect 3373 1673 3387 1687
rect 3333 1533 3347 1547
rect 3333 1473 3347 1487
rect 3213 1392 3227 1406
rect 3153 1353 3167 1367
rect 3113 1313 3127 1327
rect 3153 1313 3167 1327
rect 3053 1253 3067 1267
rect 3093 1253 3107 1267
rect 3133 1253 3147 1267
rect 3013 1213 3027 1227
rect 3093 1214 3107 1228
rect 3133 1213 3147 1227
rect 3013 1133 3027 1147
rect 3033 1113 3047 1127
rect 2993 1093 3007 1107
rect 3133 1173 3147 1187
rect 3113 1113 3127 1127
rect 3072 1053 3086 1067
rect 3093 1053 3107 1067
rect 2973 1033 2987 1047
rect 3093 993 3107 1007
rect 2913 973 2927 987
rect 2893 913 2907 927
rect 3173 1293 3187 1307
rect 3313 1392 3327 1406
rect 3293 1313 3307 1327
rect 3213 1214 3227 1228
rect 3333 1293 3347 1307
rect 3313 1253 3327 1267
rect 3293 1213 3307 1227
rect 3193 1173 3207 1187
rect 3273 1172 3287 1186
rect 3433 1893 3447 1907
rect 3493 1912 3507 1926
rect 3613 2173 3627 2187
rect 3773 2313 3787 2327
rect 3733 2293 3747 2307
rect 3773 2253 3787 2267
rect 3893 2613 3907 2627
rect 3873 2573 3887 2587
rect 3973 3252 3987 3266
rect 4013 3213 4027 3227
rect 4073 3353 4087 3367
rect 4173 3953 4187 3967
rect 4253 3992 4267 4006
rect 4233 3973 4247 3987
rect 4213 3933 4227 3947
rect 4193 3873 4207 3887
rect 4173 3833 4187 3847
rect 4333 3993 4347 4007
rect 4393 4273 4407 4287
rect 4553 4533 4567 4547
rect 4593 4473 4607 4487
rect 4553 4433 4567 4447
rect 4513 4413 4527 4427
rect 4493 4373 4507 4387
rect 4513 4353 4527 4367
rect 4533 4334 4547 4348
rect 4653 4473 4667 4487
rect 5213 5073 5227 5087
rect 5253 5074 5267 5088
rect 5293 5072 5307 5086
rect 5193 5032 5207 5046
rect 5153 4933 5167 4947
rect 5073 4913 5087 4927
rect 4973 4872 4987 4886
rect 5033 4873 5047 4887
rect 4993 4812 5007 4826
rect 4933 4753 4947 4767
rect 4953 4593 4967 4607
rect 4933 4493 4947 4507
rect 4713 4433 4727 4447
rect 4793 4433 4807 4447
rect 4893 4433 4907 4447
rect 4633 4373 4647 4387
rect 4573 4333 4587 4347
rect 4633 4334 4647 4348
rect 4673 4334 4687 4348
rect 4513 4292 4527 4306
rect 4453 4253 4467 4267
rect 4373 4153 4387 4167
rect 4433 4153 4447 4167
rect 4473 4173 4487 4187
rect 4393 4034 4407 4048
rect 4513 4073 4527 4087
rect 4613 4292 4627 4306
rect 4573 4253 4587 4267
rect 4633 4193 4647 4207
rect 4353 3953 4367 3967
rect 4293 3893 4307 3907
rect 4213 3814 4227 3828
rect 4253 3814 4267 3828
rect 4293 3814 4307 3828
rect 4153 3773 4167 3787
rect 4193 3772 4207 3786
rect 4133 3573 4147 3587
rect 4133 3514 4147 3528
rect 4313 3772 4327 3786
rect 4252 3673 4266 3687
rect 4273 3673 4287 3687
rect 4233 3514 4247 3528
rect 4073 3313 4087 3327
rect 4113 3313 4127 3327
rect 4293 3613 4307 3627
rect 4153 3433 4167 3447
rect 4213 3472 4227 3486
rect 4273 3473 4287 3487
rect 4493 4033 4507 4047
rect 4553 4033 4567 4047
rect 4593 4034 4607 4048
rect 4473 3973 4487 3987
rect 4733 4373 4747 4387
rect 4713 4153 4727 4167
rect 5053 4853 5067 4867
rect 5113 4854 5127 4868
rect 5173 4854 5187 4868
rect 5253 5013 5267 5027
rect 5373 5113 5387 5127
rect 5733 5352 5747 5366
rect 5873 5352 5887 5366
rect 5973 5413 5987 5427
rect 6173 5413 6187 5427
rect 5993 5374 6007 5388
rect 6093 5374 6107 5388
rect 5433 5193 5447 5207
rect 5513 5173 5527 5187
rect 5653 5173 5667 5187
rect 5433 5153 5447 5167
rect 5493 5153 5507 5167
rect 5413 5133 5427 5147
rect 5413 5093 5427 5107
rect 5433 5074 5447 5088
rect 5473 5074 5487 5088
rect 5313 5032 5327 5046
rect 5413 5032 5427 5046
rect 5433 5013 5447 5027
rect 5473 5013 5487 5027
rect 5293 4993 5307 5007
rect 5373 4993 5387 5007
rect 5233 4913 5247 4927
rect 5373 4913 5387 4927
rect 5253 4854 5267 4868
rect 5053 4753 5067 4767
rect 4993 4532 5007 4546
rect 5033 4532 5047 4546
rect 5013 4413 5027 4427
rect 4773 4292 4787 4306
rect 4813 4253 4827 4267
rect 4993 4233 5007 4247
rect 4873 4193 4887 4207
rect 4773 4173 4787 4187
rect 4873 4153 4887 4167
rect 4673 4053 4687 4067
rect 4773 4053 4787 4067
rect 4713 4034 4727 4048
rect 4413 3953 4427 3967
rect 4493 3953 4507 3967
rect 4413 3893 4427 3907
rect 4453 3873 4467 3887
rect 4513 3833 4527 3847
rect 4573 3992 4587 4006
rect 4633 3993 4647 4007
rect 4693 3992 4707 4006
rect 4833 4034 4847 4048
rect 4653 3953 4667 3967
rect 4633 3873 4647 3887
rect 4573 3833 4587 3847
rect 4533 3813 4547 3827
rect 4433 3772 4447 3786
rect 4473 3772 4487 3786
rect 4513 3772 4527 3786
rect 4373 3733 4387 3747
rect 4313 3514 4327 3528
rect 4353 3514 4367 3528
rect 4393 3514 4407 3528
rect 4553 3673 4567 3687
rect 4433 3573 4447 3587
rect 4193 3453 4207 3467
rect 4173 3413 4187 3427
rect 4233 3413 4247 3427
rect 4193 3373 4207 3387
rect 4193 3333 4207 3347
rect 4173 3294 4187 3308
rect 4153 3252 4167 3266
rect 4153 3213 4167 3227
rect 4213 3213 4227 3227
rect 4193 3193 4207 3207
rect 4073 3173 4087 3187
rect 4053 3093 4067 3107
rect 3953 3033 3967 3047
rect 3993 3033 4007 3047
rect 3973 2994 3987 3008
rect 4013 2994 4027 3008
rect 3993 2933 4007 2947
rect 3953 2913 3967 2927
rect 4033 2873 4047 2887
rect 4133 3053 4147 3067
rect 4193 3053 4207 3067
rect 4173 3033 4187 3047
rect 4153 3013 4167 3027
rect 4173 2994 4187 3008
rect 4113 2952 4127 2966
rect 4153 2952 4167 2966
rect 4193 2952 4207 2966
rect 4113 2933 4127 2947
rect 4073 2913 4087 2927
rect 4053 2853 4067 2867
rect 4033 2813 4047 2827
rect 4073 2793 4087 2807
rect 4013 2774 4027 2788
rect 3973 2732 3987 2746
rect 3933 2633 3947 2647
rect 3913 2593 3927 2607
rect 3893 2533 3907 2547
rect 3933 2533 3947 2547
rect 3873 2513 3887 2527
rect 3853 2473 3867 2487
rect 3933 2474 3947 2488
rect 3833 2413 3847 2427
rect 3813 2353 3827 2367
rect 4033 2732 4047 2746
rect 3993 2713 4007 2727
rect 3973 2613 3987 2627
rect 3953 2453 3967 2467
rect 3893 2413 3907 2427
rect 3873 2353 3887 2367
rect 3853 2313 3867 2327
rect 3813 2273 3827 2287
rect 3833 2253 3847 2267
rect 3872 2254 3886 2268
rect 3913 2373 3927 2387
rect 4033 2693 4047 2707
rect 4093 2773 4107 2787
rect 4133 2774 4147 2788
rect 4073 2653 4087 2667
rect 4113 2713 4127 2727
rect 4113 2692 4127 2706
rect 4173 2693 4187 2707
rect 4093 2573 4107 2587
rect 3993 2533 4007 2547
rect 4073 2513 4087 2527
rect 4033 2493 4047 2507
rect 4093 2493 4107 2507
rect 3993 2433 4007 2447
rect 4053 2413 4067 2427
rect 4153 2653 4167 2667
rect 4253 3213 4267 3227
rect 4253 3173 4267 3187
rect 4313 3173 4327 3187
rect 4353 3453 4367 3467
rect 4333 3093 4347 3107
rect 4373 3413 4387 3427
rect 4533 3514 4547 3528
rect 4433 3393 4447 3407
rect 4393 3313 4407 3327
rect 4433 3313 4447 3327
rect 4713 3933 4727 3947
rect 4773 3772 4787 3786
rect 4813 3992 4827 4006
rect 4833 3953 4847 3967
rect 4813 3933 4827 3947
rect 4713 3713 4727 3727
rect 4793 3713 4807 3727
rect 4633 3673 4647 3687
rect 4593 3653 4607 3667
rect 4633 3652 4647 3666
rect 4693 3653 4707 3667
rect 4633 3514 4647 3528
rect 4553 3472 4567 3486
rect 4613 3472 4627 3486
rect 4693 3453 4707 3467
rect 4533 3413 4547 3427
rect 4573 3413 4587 3427
rect 4513 3393 4527 3407
rect 4473 3333 4487 3347
rect 4393 3252 4407 3266
rect 4453 3213 4467 3227
rect 4493 3293 4507 3307
rect 4933 4034 4947 4048
rect 5073 4573 5087 4587
rect 5133 4793 5147 4807
rect 5333 4853 5347 4867
rect 5413 4893 5427 4907
rect 5413 4853 5427 4867
rect 5233 4812 5247 4826
rect 5213 4793 5227 4807
rect 5173 4713 5187 4727
rect 5233 4713 5247 4727
rect 5133 4653 5147 4667
rect 5213 4653 5227 4667
rect 5173 4613 5187 4627
rect 5133 4593 5147 4607
rect 5093 4553 5107 4567
rect 5173 4573 5187 4587
rect 5113 4512 5127 4526
rect 5153 4512 5167 4526
rect 5193 4512 5207 4526
rect 5193 4433 5207 4447
rect 5073 4413 5087 4427
rect 5153 4373 5167 4387
rect 5353 4793 5367 4807
rect 5473 4933 5487 4947
rect 5513 5073 5527 5087
rect 5553 5074 5567 5088
rect 5593 5074 5607 5088
rect 5633 5074 5647 5088
rect 5513 5033 5527 5047
rect 5513 4993 5527 5007
rect 5593 5013 5607 5027
rect 5573 4953 5587 4967
rect 5533 4933 5547 4947
rect 5513 4893 5527 4907
rect 5472 4873 5486 4887
rect 5493 4873 5507 4887
rect 5573 4913 5587 4927
rect 5393 4773 5407 4787
rect 5333 4693 5347 4707
rect 5333 4653 5347 4667
rect 5293 4613 5307 4627
rect 5313 4512 5327 4526
rect 5233 4493 5247 4507
rect 5273 4493 5287 4507
rect 5573 4853 5587 4867
rect 5473 4813 5487 4827
rect 5513 4812 5527 4826
rect 5553 4812 5567 4826
rect 5473 4753 5487 4767
rect 5633 4993 5647 5007
rect 5733 5153 5747 5167
rect 5693 5074 5707 5088
rect 5793 5113 5807 5127
rect 5673 5033 5687 5047
rect 5653 4953 5667 4967
rect 5733 5013 5747 5027
rect 5713 4993 5727 5007
rect 5833 5074 5847 5088
rect 5953 5273 5967 5287
rect 5913 5133 5927 5147
rect 5933 5113 5947 5127
rect 5833 5013 5847 5027
rect 5753 4973 5767 4987
rect 5733 4953 5747 4967
rect 5773 4953 5787 4967
rect 5673 4913 5687 4927
rect 5753 4893 5767 4907
rect 5673 4873 5687 4887
rect 5613 4853 5627 4867
rect 5713 4854 5727 4868
rect 5733 4813 5747 4827
rect 5693 4793 5707 4807
rect 5653 4773 5667 4787
rect 5453 4733 5467 4747
rect 5493 4733 5507 4747
rect 5593 4733 5607 4747
rect 5473 4693 5487 4707
rect 5413 4554 5427 4568
rect 5433 4512 5447 4526
rect 5453 4513 5467 4527
rect 5373 4473 5387 4487
rect 5413 4473 5427 4487
rect 5313 4433 5327 4447
rect 5353 4433 5367 4447
rect 5213 4353 5227 4367
rect 5273 4353 5287 4367
rect 5073 4233 5087 4247
rect 5473 4433 5487 4447
rect 5253 4293 5267 4307
rect 5353 4293 5367 4307
rect 5213 4173 5227 4187
rect 5053 4153 5067 4167
rect 5093 4093 5107 4107
rect 5053 4073 5067 4087
rect 5173 4073 5187 4087
rect 5133 4034 5147 4048
rect 4993 3993 5007 4007
rect 5093 3993 5107 4007
rect 5153 3992 5167 4006
rect 4913 3953 4927 3967
rect 5033 3953 5047 3967
rect 4873 3913 4887 3927
rect 4893 3814 4907 3828
rect 4973 3813 4987 3827
rect 5073 3813 5087 3827
rect 5173 3814 5187 3828
rect 5093 3793 5107 3807
rect 4873 3772 4887 3786
rect 4973 3772 4987 3786
rect 5013 3772 5027 3786
rect 5233 3973 5247 3987
rect 5153 3772 5167 3786
rect 5213 3773 5227 3787
rect 5053 3753 5067 3767
rect 5093 3753 5107 3767
rect 5133 3753 5147 3767
rect 5013 3713 5027 3727
rect 4993 3693 5007 3707
rect 4913 3673 4927 3687
rect 4873 3653 4887 3667
rect 4833 3613 4847 3627
rect 4773 3533 4787 3547
rect 4813 3514 4827 3528
rect 4853 3533 4867 3547
rect 4953 3533 4967 3547
rect 4793 3472 4807 3486
rect 4833 3473 4847 3487
rect 4753 3453 4767 3467
rect 4713 3413 4727 3427
rect 4873 3514 4887 3528
rect 4913 3514 4927 3528
rect 5113 3653 5127 3667
rect 5053 3533 5067 3547
rect 5113 3514 5127 3528
rect 5013 3493 5027 3507
rect 4893 3473 4907 3487
rect 4872 3453 4886 3467
rect 4753 3393 4767 3407
rect 4853 3393 4867 3407
rect 4693 3373 4707 3387
rect 4473 3193 4487 3207
rect 4373 3173 4387 3187
rect 4313 3073 4327 3087
rect 4353 3073 4367 3087
rect 4553 3252 4567 3266
rect 4613 3193 4627 3207
rect 4593 3173 4607 3187
rect 4393 3053 4407 3067
rect 4493 3053 4507 3067
rect 4353 2994 4367 3008
rect 4293 2952 4307 2966
rect 4313 2933 4327 2947
rect 4233 2893 4247 2907
rect 4213 2833 4227 2847
rect 4233 2813 4247 2827
rect 4293 2813 4307 2827
rect 4213 2753 4227 2767
rect 4193 2613 4207 2627
rect 4153 2493 4167 2507
rect 4453 2994 4467 3008
rect 4433 2952 4447 2966
rect 4513 2993 4527 3007
rect 4553 2994 4567 3008
rect 4393 2933 4407 2947
rect 4333 2833 4347 2847
rect 4373 2833 4387 2847
rect 4313 2793 4327 2807
rect 4253 2774 4267 2788
rect 4433 2774 4447 2788
rect 4573 2952 4587 2966
rect 4533 2893 4547 2907
rect 4533 2853 4547 2867
rect 4233 2653 4247 2667
rect 4253 2653 4267 2667
rect 4313 2653 4327 2667
rect 4233 2593 4247 2607
rect 4233 2473 4247 2487
rect 4273 2613 4287 2627
rect 4113 2413 4127 2427
rect 4193 2432 4207 2446
rect 4253 2432 4267 2446
rect 4173 2413 4187 2427
rect 3973 2393 3987 2407
rect 4033 2393 4047 2407
rect 4093 2393 4107 2407
rect 4153 2393 4167 2407
rect 3893 2253 3907 2267
rect 3733 2193 3747 2207
rect 3673 2153 3687 2167
rect 3713 2153 3727 2167
rect 3593 2113 3607 2127
rect 3713 2093 3727 2107
rect 3612 2073 3626 2087
rect 3633 2073 3647 2087
rect 3573 1993 3587 2007
rect 3453 1853 3467 1867
rect 3553 1833 3567 1847
rect 3533 1753 3547 1767
rect 3493 1734 3507 1748
rect 3433 1693 3447 1707
rect 3533 1693 3547 1707
rect 3693 2053 3707 2067
rect 3632 1973 3646 1987
rect 3653 1973 3667 1987
rect 3713 1993 3727 2007
rect 3693 1954 3707 1968
rect 3633 1912 3647 1926
rect 3673 1893 3687 1907
rect 3713 1833 3727 1847
rect 3772 2193 3786 2207
rect 3793 2193 3807 2207
rect 3773 2153 3787 2167
rect 3753 2093 3767 2107
rect 3753 2013 3767 2027
rect 3853 2212 3867 2226
rect 3833 2193 3847 2207
rect 3893 2193 3907 2207
rect 3813 2113 3827 2127
rect 3933 2353 3947 2367
rect 3933 2273 3947 2287
rect 3933 2252 3947 2266
rect 3973 2273 3987 2287
rect 3933 2213 3947 2227
rect 3993 2212 4007 2226
rect 4013 2173 4027 2187
rect 3892 2153 3906 2167
rect 3913 2153 3927 2167
rect 3973 2133 3987 2147
rect 3873 2113 3887 2127
rect 3793 2053 3807 2067
rect 3833 2073 3847 2087
rect 3813 2033 3827 2047
rect 3793 1954 3807 1968
rect 3813 1912 3827 1926
rect 3972 2093 3986 2107
rect 3993 2093 4007 2107
rect 3893 2013 3907 2027
rect 4113 2353 4127 2367
rect 4093 2313 4107 2327
rect 4113 2273 4127 2287
rect 4133 2254 4147 2268
rect 4073 2212 4087 2226
rect 4153 2213 4167 2227
rect 4113 2153 4127 2167
rect 4033 2093 4047 2107
rect 4013 2073 4027 2087
rect 4033 1993 4047 2007
rect 4013 1973 4027 1987
rect 3953 1954 3967 1968
rect 3993 1954 4007 1968
rect 3753 1893 3767 1907
rect 3673 1813 3687 1827
rect 3733 1813 3747 1827
rect 3573 1773 3587 1787
rect 3573 1734 3587 1748
rect 3613 1734 3627 1748
rect 3472 1673 3486 1687
rect 3493 1673 3507 1687
rect 3553 1673 3567 1687
rect 3413 1573 3427 1587
rect 3373 1493 3387 1507
rect 3373 1472 3387 1486
rect 3413 1473 3427 1487
rect 3373 1433 3387 1447
rect 3453 1593 3467 1607
rect 3453 1533 3467 1547
rect 3432 1433 3446 1447
rect 3453 1434 3467 1448
rect 3393 1392 3407 1406
rect 3393 1293 3407 1307
rect 3373 1253 3387 1267
rect 3353 1233 3367 1247
rect 3453 1353 3467 1367
rect 3433 1233 3447 1247
rect 3413 1213 3427 1227
rect 3233 1133 3247 1147
rect 3213 1073 3227 1087
rect 3193 993 3207 1007
rect 3173 953 3187 967
rect 3133 913 3147 927
rect 3173 913 3187 927
rect 3313 1172 3327 1186
rect 3353 1172 3367 1186
rect 3393 1172 3407 1186
rect 3393 1033 3407 1047
rect 3293 1013 3307 1027
rect 3353 953 3367 967
rect 3313 914 3327 928
rect 3353 914 3367 928
rect 2993 872 3007 886
rect 2873 853 2887 867
rect 2913 853 2927 867
rect 2753 793 2767 807
rect 2873 753 2887 767
rect 2913 753 2927 767
rect 2733 694 2747 708
rect 2793 694 2807 708
rect 2833 694 2847 708
rect 2713 673 2727 687
rect 2673 652 2687 666
rect 2732 653 2746 667
rect 2753 653 2767 667
rect 2913 732 2927 746
rect 2953 713 2967 727
rect 3013 693 3027 707
rect 3533 1513 3547 1527
rect 3573 1513 3587 1527
rect 3613 1473 3627 1487
rect 3573 1434 3587 1448
rect 3493 1392 3507 1406
rect 3493 1313 3507 1327
rect 3473 1293 3487 1307
rect 3493 1253 3507 1267
rect 3553 1313 3567 1327
rect 3533 1293 3547 1307
rect 3573 1233 3587 1247
rect 3613 1233 3627 1247
rect 3513 1172 3527 1186
rect 3453 1133 3467 1147
rect 3533 1133 3547 1147
rect 3653 1693 3667 1707
rect 3693 1753 3707 1767
rect 3753 1753 3767 1767
rect 3673 1653 3687 1667
rect 3833 1853 3847 1867
rect 3813 1733 3827 1747
rect 3733 1692 3747 1706
rect 3813 1693 3827 1707
rect 3973 1893 3987 1907
rect 3933 1873 3947 1887
rect 3873 1793 3887 1807
rect 3913 1753 3927 1767
rect 3913 1734 3927 1748
rect 3953 1733 3967 1747
rect 3833 1673 3847 1687
rect 3873 1673 3887 1687
rect 3773 1653 3787 1667
rect 3693 1633 3707 1647
rect 3753 1493 3767 1507
rect 3693 1434 3707 1448
rect 3733 1433 3747 1447
rect 3673 1392 3687 1406
rect 3853 1473 3867 1487
rect 3793 1434 3807 1448
rect 3673 1333 3687 1347
rect 3753 1353 3767 1367
rect 3733 1333 3747 1347
rect 3733 1293 3747 1307
rect 3713 1273 3727 1287
rect 3733 1233 3747 1247
rect 3673 1214 3687 1228
rect 3713 1213 3727 1227
rect 3613 1172 3627 1186
rect 3573 1133 3587 1147
rect 3553 1093 3567 1107
rect 3693 1073 3707 1087
rect 3593 993 3607 1007
rect 3533 933 3547 947
rect 3493 914 3507 928
rect 3193 872 3207 886
rect 3133 833 3147 847
rect 3173 833 3187 847
rect 3072 813 3086 827
rect 3093 813 3107 827
rect 3113 713 3127 727
rect 2573 593 2587 607
rect 2453 433 2467 447
rect 2353 394 2367 408
rect 2133 353 2147 367
rect 2113 333 2127 347
rect 2093 313 2107 327
rect 2073 213 2087 227
rect 2053 193 2067 207
rect 1913 153 1927 167
rect 1773 133 1787 147
rect 1813 132 1827 146
rect 1853 132 1867 146
rect 2033 132 2047 146
rect 2193 352 2207 366
rect 2252 353 2266 367
rect 2273 353 2287 367
rect 2213 253 2227 267
rect 2153 213 2167 227
rect 2133 174 2147 188
rect 2173 174 2187 188
rect 2113 132 2127 146
rect 2293 333 2307 347
rect 2493 394 2507 408
rect 2433 352 2447 366
rect 2393 313 2407 327
rect 2433 293 2447 307
rect 2393 273 2407 287
rect 2373 253 2387 267
rect 2373 213 2387 227
rect 2073 93 2087 107
rect 2113 93 2127 107
rect 1993 73 2007 87
rect 2213 132 2227 146
rect 2273 132 2287 146
rect 2233 93 2247 107
rect 2273 93 2287 107
rect 2513 353 2527 367
rect 2493 293 2507 307
rect 2473 253 2487 267
rect 2413 213 2427 227
rect 2453 213 2467 227
rect 2393 173 2407 187
rect 2513 213 2527 227
rect 2493 173 2507 187
rect 2433 132 2447 146
rect 2473 132 2487 146
rect 2513 113 2527 127
rect 2553 493 2567 507
rect 2813 652 2827 666
rect 2873 652 2887 666
rect 2773 593 2787 607
rect 2813 593 2827 607
rect 2973 652 2987 666
rect 3013 652 3027 666
rect 2813 553 2827 567
rect 2933 553 2947 567
rect 3113 694 3127 708
rect 3093 652 3107 666
rect 3193 793 3207 807
rect 3213 753 3227 767
rect 3333 872 3347 886
rect 3373 833 3387 847
rect 3433 872 3447 886
rect 3473 872 3487 886
rect 3413 813 3427 827
rect 3333 793 3347 807
rect 3273 733 3287 747
rect 3233 713 3247 727
rect 3193 613 3207 627
rect 3293 613 3307 627
rect 3173 573 3187 587
rect 3253 573 3267 587
rect 3133 553 3147 567
rect 2853 533 2867 547
rect 3033 533 3047 547
rect 2833 513 2847 527
rect 2893 513 2907 527
rect 2753 493 2767 507
rect 2853 493 2867 507
rect 2713 453 2727 467
rect 2613 433 2627 447
rect 2553 394 2567 408
rect 2653 394 2667 408
rect 2693 394 2707 408
rect 2793 394 2807 408
rect 2953 453 2967 467
rect 3033 453 3047 467
rect 2913 394 2927 408
rect 2992 394 3006 408
rect 3013 394 3027 408
rect 2713 373 2727 387
rect 2553 353 2567 367
rect 2633 352 2647 366
rect 2693 353 2707 367
rect 2593 313 2607 327
rect 2693 253 2707 267
rect 2773 352 2787 366
rect 2793 333 2807 347
rect 2813 313 2827 327
rect 2793 293 2807 307
rect 2813 273 2827 287
rect 2853 352 2867 366
rect 2793 253 2807 267
rect 2833 253 2847 267
rect 2713 233 2727 247
rect 2633 213 2647 227
rect 2573 193 2587 207
rect 2613 174 2627 188
rect 2672 174 2686 188
rect 2693 174 2707 188
rect 2753 174 2767 188
rect 2353 73 2367 87
rect 1973 53 1987 67
rect 2013 53 2027 67
rect 2193 53 2207 67
rect 2233 53 2247 67
rect 2313 53 2327 67
rect 2393 53 2407 67
rect 2593 53 2607 67
rect 2673 133 2687 147
rect 2733 132 2747 146
rect 2933 352 2947 366
rect 3012 353 3026 367
rect 3173 433 3187 447
rect 3133 414 3147 428
rect 3073 394 3087 408
rect 3113 393 3127 407
rect 3193 394 3207 408
rect 3253 394 3267 408
rect 3033 352 3047 366
rect 3093 352 3107 366
rect 3113 333 3127 347
rect 3093 293 3107 307
rect 2973 213 2987 227
rect 2933 174 2947 188
rect 2993 174 3007 188
rect 3053 174 3067 188
rect 3113 233 3127 247
rect 3173 352 3187 366
rect 3233 352 3247 366
rect 3273 352 3287 366
rect 3193 293 3207 307
rect 3313 333 3327 347
rect 3233 273 3247 287
rect 3193 253 3207 267
rect 3133 213 3147 227
rect 3113 193 3127 207
rect 3132 174 3146 188
rect 3153 174 3167 188
rect 3233 233 3247 247
rect 3653 933 3667 947
rect 3713 993 3727 1007
rect 3773 1333 3787 1347
rect 3753 1213 3767 1227
rect 3833 1233 3847 1247
rect 3853 1214 3867 1228
rect 3893 1533 3907 1547
rect 3993 1793 4007 1807
rect 4193 2333 4207 2347
rect 4173 2173 4187 2187
rect 4493 2732 4507 2746
rect 4453 2613 4467 2627
rect 4493 2573 4507 2587
rect 4353 2474 4367 2488
rect 4393 2474 4407 2488
rect 4493 2474 4507 2488
rect 4273 2393 4287 2407
rect 4333 2393 4347 2407
rect 4353 2313 4367 2327
rect 4293 2273 4307 2287
rect 4233 2212 4247 2226
rect 4253 2133 4267 2147
rect 4273 2113 4287 2127
rect 4253 2093 4267 2107
rect 4193 2073 4207 2087
rect 4153 1973 4167 1987
rect 4233 1954 4247 1968
rect 4453 2432 4467 2446
rect 4453 2353 4467 2367
rect 4673 3073 4687 3087
rect 5093 3473 5107 3487
rect 4933 3433 4947 3447
rect 5013 3453 5027 3467
rect 4973 3433 4987 3447
rect 4953 3393 4967 3407
rect 4873 3313 4887 3327
rect 4873 3252 4887 3266
rect 4833 3213 4847 3227
rect 4753 3073 4767 3087
rect 4713 3033 4727 3047
rect 4733 2993 4747 3007
rect 4653 2952 4667 2966
rect 4733 2952 4747 2966
rect 4693 2913 4707 2927
rect 4793 2994 4807 3008
rect 4813 2952 4827 2966
rect 4933 3333 4947 3347
rect 5433 4292 5447 4306
rect 5413 4253 5427 4267
rect 5393 4133 5407 4147
rect 5293 4034 5307 4048
rect 5353 3992 5367 4006
rect 5313 3953 5327 3967
rect 5293 3814 5307 3828
rect 5653 4693 5667 4707
rect 5553 4593 5567 4607
rect 5633 4593 5647 4607
rect 5593 4554 5607 4568
rect 5573 4512 5587 4526
rect 5693 4554 5707 4568
rect 5773 4873 5787 4887
rect 5913 5013 5927 5027
rect 5893 4993 5907 5007
rect 5873 4893 5887 4907
rect 5753 4773 5767 4787
rect 5813 4753 5827 4767
rect 5853 4693 5867 4707
rect 5853 4613 5867 4627
rect 5773 4554 5787 4568
rect 5813 4554 5827 4568
rect 6113 5273 6127 5287
rect 6233 5332 6247 5346
rect 6133 5253 6147 5267
rect 6173 5253 6187 5267
rect 6113 5193 6127 5207
rect 6053 5074 6067 5088
rect 5973 5013 5987 5027
rect 6033 4993 6047 5007
rect 5953 4913 5967 4927
rect 5953 4854 5967 4868
rect 5993 4854 6007 4868
rect 6173 5113 6187 5127
rect 6233 5074 6247 5088
rect 6133 5033 6147 5047
rect 6193 5032 6207 5046
rect 6113 4993 6127 5007
rect 6173 4993 6187 5007
rect 6233 4993 6247 5007
rect 6133 4913 6147 4927
rect 6073 4853 6087 4867
rect 5933 4793 5947 4807
rect 5913 4573 5927 4587
rect 5653 4493 5667 4507
rect 5613 4433 5627 4447
rect 5713 4512 5727 4526
rect 5693 4493 5707 4507
rect 5673 4373 5687 4387
rect 5533 4253 5547 4267
rect 5493 4233 5507 4247
rect 5553 4233 5567 4247
rect 5453 4093 5467 4107
rect 5493 4034 5507 4048
rect 5533 4034 5547 4048
rect 5413 3993 5427 4007
rect 5433 3953 5447 3967
rect 5493 3973 5507 3987
rect 5533 3973 5547 3987
rect 5473 3873 5487 3887
rect 5633 4093 5647 4107
rect 5593 4034 5607 4048
rect 5573 3993 5587 4007
rect 5513 3814 5527 3828
rect 5653 3992 5667 4006
rect 5613 3973 5627 3987
rect 5653 3953 5667 3967
rect 5633 3873 5647 3887
rect 5373 3753 5387 3767
rect 5273 3713 5287 3727
rect 5233 3613 5247 3627
rect 5153 3514 5167 3528
rect 5293 3693 5307 3707
rect 5273 3493 5287 3507
rect 5073 3453 5087 3467
rect 5033 3393 5047 3407
rect 5053 3333 5067 3347
rect 4973 3313 4987 3327
rect 5013 3294 5027 3308
rect 4993 3252 5007 3266
rect 4933 3033 4947 3047
rect 4973 3033 4987 3047
rect 5033 2994 5047 3008
rect 4893 2953 4907 2967
rect 4953 2952 4967 2966
rect 4852 2913 4866 2927
rect 4873 2913 4887 2927
rect 4993 2913 5007 2927
rect 4953 2893 4967 2907
rect 5033 2893 5047 2907
rect 4613 2853 4627 2867
rect 4753 2853 4767 2867
rect 4573 2833 4587 2847
rect 4673 2833 4687 2847
rect 4653 2813 4667 2827
rect 4593 2774 4607 2788
rect 4653 2733 4667 2747
rect 4613 2673 4627 2687
rect 4633 2653 4647 2667
rect 4613 2633 4627 2647
rect 4593 2474 4607 2488
rect 4733 2813 4747 2827
rect 4773 2774 4787 2788
rect 4813 2773 4827 2787
rect 4873 2774 4887 2788
rect 4933 2773 4947 2787
rect 4813 2713 4827 2727
rect 4753 2693 4767 2707
rect 4893 2713 4907 2727
rect 4853 2593 4867 2607
rect 4613 2393 4627 2407
rect 4653 2393 4667 2407
rect 4553 2353 4567 2367
rect 4413 2293 4427 2307
rect 4533 2293 4547 2307
rect 4393 2253 4407 2267
rect 4333 2212 4347 2226
rect 4373 2212 4387 2226
rect 4473 2254 4487 2268
rect 4533 2254 4547 2268
rect 4433 2212 4447 2226
rect 4333 2173 4347 2187
rect 4413 2173 4427 2187
rect 4293 2033 4307 2047
rect 4373 1993 4387 2007
rect 4333 1954 4347 1968
rect 4493 2212 4507 2226
rect 4653 2293 4667 2307
rect 4613 2254 4627 2268
rect 4553 2212 4567 2226
rect 4633 2212 4647 2226
rect 4633 2193 4647 2207
rect 4593 2133 4607 2147
rect 4813 2533 4827 2547
rect 4753 2474 4767 2488
rect 5113 3453 5127 3467
rect 5273 3413 5287 3427
rect 5213 3393 5227 3407
rect 5373 3633 5387 3647
rect 5413 3613 5427 3627
rect 5333 3573 5347 3587
rect 5373 3573 5387 3587
rect 5593 3772 5607 3786
rect 5533 3533 5547 3547
rect 5373 3514 5387 3528
rect 5473 3514 5487 3528
rect 5673 3913 5687 3927
rect 5773 4473 5787 4487
rect 5873 4493 5887 4507
rect 5853 4473 5867 4487
rect 5713 4373 5727 4387
rect 5793 4373 5807 4387
rect 5833 4373 5847 4387
rect 5753 4334 5767 4348
rect 5773 4292 5787 4306
rect 5713 4273 5727 4287
rect 5793 4273 5807 4287
rect 5713 4233 5727 4247
rect 6013 4812 6027 4826
rect 6053 4813 6067 4827
rect 6113 4812 6127 4826
rect 6013 4793 6027 4807
rect 6033 4773 6047 4787
rect 6133 4773 6147 4787
rect 5953 4673 5967 4687
rect 6013 4573 6027 4587
rect 5973 4554 5987 4568
rect 6053 4693 6067 4707
rect 6053 4613 6067 4627
rect 5933 4533 5947 4547
rect 5913 4473 5927 4487
rect 6093 4554 6107 4568
rect 6253 4953 6267 4967
rect 6193 4854 6207 4868
rect 6293 4854 6307 4868
rect 6233 4812 6247 4826
rect 6273 4812 6287 4826
rect 6313 4812 6327 4826
rect 6193 4693 6207 4707
rect 6173 4673 6187 4687
rect 6173 4554 6187 4568
rect 6213 4554 6227 4568
rect 6253 4554 6267 4568
rect 6292 4554 6306 4568
rect 5993 4512 6007 4526
rect 6053 4513 6067 4527
rect 5933 4433 5947 4447
rect 5973 4334 5987 4348
rect 5813 4233 5827 4247
rect 5853 4233 5867 4247
rect 6153 4512 6167 4526
rect 6033 4473 6047 4487
rect 6113 4473 6127 4487
rect 6073 4334 6087 4348
rect 5813 4193 5827 4207
rect 5913 4193 5927 4207
rect 5913 4133 5927 4147
rect 5873 4034 5887 4048
rect 5813 4013 5827 4027
rect 5773 3973 5787 3987
rect 5713 3933 5727 3947
rect 5693 3893 5707 3907
rect 5773 3932 5787 3946
rect 5753 3913 5767 3927
rect 5733 3873 5747 3887
rect 5713 3814 5727 3828
rect 5773 3813 5787 3827
rect 5693 3772 5707 3786
rect 5933 3992 5947 4006
rect 5893 3893 5907 3907
rect 5853 3873 5867 3887
rect 5973 4034 5987 4048
rect 6013 4034 6027 4048
rect 6093 4292 6107 4306
rect 6313 4553 6327 4567
rect 6273 4512 6287 4526
rect 6213 4473 6227 4487
rect 6273 4473 6287 4487
rect 6173 4413 6187 4427
rect 6213 4334 6227 4348
rect 6133 4253 6147 4267
rect 6233 4253 6247 4267
rect 6053 4193 6067 4207
rect 6093 4034 6107 4048
rect 5953 3913 5967 3927
rect 6073 3992 6087 4006
rect 6013 3973 6027 3987
rect 5973 3873 5987 3887
rect 5893 3833 5907 3847
rect 5933 3833 5947 3847
rect 6033 3833 6047 3847
rect 5813 3773 5827 3787
rect 5733 3732 5747 3746
rect 5793 3733 5807 3747
rect 5873 3772 5887 3786
rect 5833 3753 5847 3767
rect 5953 3814 5967 3828
rect 5993 3814 6007 3828
rect 5593 3693 5607 3707
rect 5653 3693 5667 3707
rect 5633 3653 5647 3667
rect 5573 3533 5587 3547
rect 5353 3472 5367 3486
rect 5393 3453 5407 3467
rect 5353 3413 5367 3427
rect 5133 3333 5147 3347
rect 5213 3333 5227 3347
rect 5093 3293 5107 3307
rect 5173 3294 5187 3308
rect 5113 3252 5127 3266
rect 5073 3133 5087 3147
rect 5193 3233 5207 3247
rect 5153 3153 5167 3167
rect 5073 3073 5087 3087
rect 5113 3073 5127 3087
rect 5113 3033 5127 3047
rect 5093 2853 5107 2867
rect 5073 2813 5087 2827
rect 4993 2774 5007 2788
rect 5053 2774 5067 2788
rect 5173 3093 5187 3107
rect 5053 2733 5067 2747
rect 5013 2713 5027 2727
rect 4953 2673 4967 2687
rect 4933 2653 4947 2667
rect 5033 2653 5047 2667
rect 4953 2593 4967 2607
rect 4913 2474 4927 2488
rect 4993 2474 5007 2488
rect 4793 2432 4807 2446
rect 4853 2432 4867 2446
rect 4933 2432 4947 2446
rect 5033 2393 5047 2407
rect 4973 2373 4987 2387
rect 4993 2313 5007 2327
rect 4893 2293 4907 2307
rect 4973 2293 4987 2307
rect 4773 2254 4787 2268
rect 4813 2254 4827 2268
rect 4953 2253 4967 2267
rect 4993 2253 5007 2267
rect 5153 2733 5167 2747
rect 5313 3313 5327 3327
rect 5273 3294 5287 3308
rect 5213 3093 5227 3107
rect 5293 3233 5307 3247
rect 5273 3153 5287 3167
rect 5253 3053 5267 3067
rect 5233 2994 5247 3008
rect 5533 3453 5547 3467
rect 5553 3433 5567 3447
rect 5473 3353 5487 3367
rect 5493 3313 5507 3327
rect 5553 3313 5567 3327
rect 5673 3514 5687 3528
rect 5753 3693 5767 3707
rect 5613 3473 5627 3487
rect 5613 3413 5627 3427
rect 5693 3472 5707 3486
rect 5733 3473 5747 3487
rect 5793 3514 5807 3528
rect 5933 3733 5947 3747
rect 6013 3772 6027 3786
rect 6053 3733 6067 3747
rect 5953 3693 5967 3707
rect 5933 3553 5947 3567
rect 5773 3472 5787 3486
rect 5713 3433 5727 3447
rect 5753 3433 5767 3447
rect 5653 3373 5667 3387
rect 5633 3353 5647 3367
rect 5373 3293 5387 3307
rect 5433 3294 5447 3308
rect 5353 3113 5367 3127
rect 5293 3093 5307 3107
rect 5593 3294 5607 3308
rect 5453 3252 5467 3266
rect 5493 3252 5507 3266
rect 5613 3253 5627 3267
rect 5413 3213 5427 3227
rect 5473 3213 5487 3227
rect 5453 3153 5467 3167
rect 5313 3053 5327 3067
rect 5373 3053 5387 3067
rect 5193 2913 5207 2927
rect 5293 2953 5307 2967
rect 5253 2913 5267 2927
rect 5213 2774 5227 2788
rect 5273 2873 5287 2887
rect 5313 2793 5327 2807
rect 5273 2732 5287 2746
rect 5173 2713 5187 2727
rect 5113 2673 5127 2687
rect 5133 2533 5147 2547
rect 5253 2533 5267 2547
rect 5093 2474 5107 2488
rect 5213 2513 5227 2527
rect 5193 2474 5207 2488
rect 5073 2433 5087 2447
rect 5113 2373 5127 2387
rect 5073 2313 5087 2327
rect 5113 2254 5127 2268
rect 5453 2993 5467 3007
rect 5513 2994 5527 3008
rect 5613 3193 5627 3207
rect 5613 2994 5627 3008
rect 5433 2933 5447 2947
rect 5473 2933 5487 2947
rect 5393 2813 5407 2827
rect 5373 2793 5387 2807
rect 5573 2933 5587 2947
rect 5733 3413 5747 3427
rect 5673 3294 5687 3308
rect 5733 3293 5747 3307
rect 5653 3253 5667 3267
rect 5693 3252 5707 3266
rect 5853 3472 5867 3486
rect 5813 3433 5827 3447
rect 5773 3293 5787 3307
rect 5933 3514 5947 3528
rect 5913 3373 5927 3387
rect 5913 3333 5927 3347
rect 5853 3294 5867 3308
rect 5893 3293 5907 3307
rect 5773 3253 5787 3267
rect 5793 3233 5807 3247
rect 5753 3173 5767 3187
rect 5693 3033 5707 3047
rect 5693 2994 5707 3008
rect 5733 2994 5747 3008
rect 5633 2933 5647 2947
rect 5593 2893 5607 2907
rect 5533 2873 5547 2887
rect 5533 2833 5547 2847
rect 5493 2774 5507 2788
rect 5353 2732 5367 2746
rect 5393 2732 5407 2746
rect 5433 2733 5447 2747
rect 5473 2733 5487 2747
rect 5313 2493 5327 2507
rect 5293 2474 5307 2488
rect 5373 2593 5387 2607
rect 5473 2533 5487 2547
rect 5413 2513 5427 2527
rect 5373 2473 5387 2487
rect 5453 2474 5467 2488
rect 5213 2413 5227 2427
rect 5253 2393 5267 2407
rect 5213 2293 5227 2307
rect 4913 2212 4927 2226
rect 4793 2193 4807 2207
rect 5033 2212 5047 2226
rect 5073 2212 5087 2226
rect 5173 2254 5187 2268
rect 5393 2432 5407 2446
rect 5293 2413 5307 2427
rect 5273 2353 5287 2367
rect 5273 2293 5287 2307
rect 5253 2253 5267 2267
rect 5233 2212 5247 2226
rect 5373 2333 5387 2347
rect 5333 2273 5347 2287
rect 5413 2413 5427 2427
rect 5393 2313 5407 2327
rect 4953 2173 4967 2187
rect 5093 2173 5107 2187
rect 5133 2173 5147 2187
rect 4753 2133 4767 2147
rect 4453 2093 4467 2107
rect 4533 2093 4547 2107
rect 4613 2093 4627 2107
rect 4693 2093 4707 2107
rect 4973 2073 4987 2087
rect 5033 2073 5047 2087
rect 4673 2053 4687 2067
rect 4613 2033 4627 2047
rect 4533 1993 4547 2007
rect 4553 1954 4567 1968
rect 4033 1913 4047 1927
rect 4253 1893 4267 1907
rect 4173 1873 4187 1887
rect 4293 1853 4307 1867
rect 4113 1813 4127 1827
rect 4113 1792 4127 1806
rect 4013 1734 4027 1748
rect 4053 1734 4067 1748
rect 3973 1613 3987 1627
rect 3973 1533 3987 1547
rect 3953 1473 3967 1487
rect 3933 1434 3947 1448
rect 3913 1333 3927 1347
rect 3893 1253 3907 1267
rect 3953 1253 3967 1267
rect 3913 1233 3927 1247
rect 3913 1214 3927 1228
rect 4073 1673 4087 1687
rect 4233 1773 4247 1787
rect 4153 1753 4167 1767
rect 4133 1733 4147 1747
rect 4313 1813 4327 1827
rect 4293 1713 4307 1727
rect 4133 1673 4147 1687
rect 4113 1593 4127 1607
rect 4173 1593 4187 1607
rect 4133 1553 4147 1567
rect 4073 1533 4087 1547
rect 4033 1493 4047 1507
rect 3993 1433 4007 1447
rect 4033 1434 4047 1448
rect 3993 1253 4007 1267
rect 3993 1213 4007 1227
rect 3773 1172 3787 1186
rect 3813 1172 3827 1186
rect 3873 1172 3887 1186
rect 4033 1373 4047 1387
rect 4033 1213 4047 1227
rect 4093 1353 4107 1367
rect 4153 1434 4167 1448
rect 4533 1912 4547 1926
rect 4673 2013 4687 2027
rect 4873 2013 4887 2027
rect 4713 1973 4727 1987
rect 4753 1973 4767 1987
rect 5053 2033 5067 2047
rect 5033 1973 5047 1987
rect 4393 1853 4407 1867
rect 4433 1773 4447 1787
rect 4453 1753 4467 1767
rect 4333 1733 4347 1747
rect 4373 1734 4387 1748
rect 4433 1732 4447 1746
rect 4313 1692 4327 1706
rect 4353 1692 4367 1706
rect 4293 1553 4307 1567
rect 4273 1493 4287 1507
rect 4233 1453 4247 1467
rect 4193 1434 4207 1448
rect 4213 1392 4227 1406
rect 4173 1373 4187 1387
rect 4153 1353 4167 1367
rect 4133 1293 4147 1307
rect 4173 1253 4187 1267
rect 4193 1233 4207 1247
rect 3733 953 3747 967
rect 3693 914 3707 928
rect 3793 914 3807 928
rect 3833 914 3847 928
rect 3933 1172 3947 1186
rect 3973 1172 3987 1186
rect 4013 1172 4027 1186
rect 4053 1172 4067 1186
rect 4093 1153 4107 1167
rect 3933 993 3947 1007
rect 3913 953 3927 967
rect 3893 913 3907 927
rect 3633 872 3647 886
rect 3793 853 3807 867
rect 3673 833 3687 847
rect 3593 753 3607 767
rect 3492 733 3506 747
rect 3513 733 3527 747
rect 3773 733 3787 747
rect 3373 694 3387 708
rect 3413 694 3427 708
rect 3473 694 3487 708
rect 3713 713 3727 727
rect 3553 694 3567 708
rect 3393 652 3407 666
rect 3633 693 3647 707
rect 3673 694 3687 708
rect 3533 652 3547 666
rect 3433 613 3447 627
rect 3473 553 3487 567
rect 3393 513 3407 527
rect 3393 394 3407 408
rect 3433 394 3447 408
rect 3533 593 3547 607
rect 3493 493 3507 507
rect 3413 352 3427 366
rect 3473 353 3487 367
rect 3573 593 3587 607
rect 3853 872 3867 886
rect 3913 872 3927 886
rect 3893 813 3907 827
rect 3813 713 3827 727
rect 3853 713 3867 727
rect 3973 953 3987 967
rect 4173 1213 4187 1227
rect 4233 1233 4247 1247
rect 4393 1673 4407 1687
rect 4493 1734 4507 1748
rect 4533 1753 4547 1767
rect 4573 1753 4587 1767
rect 4613 1753 4627 1767
rect 4473 1693 4487 1707
rect 4453 1673 4467 1687
rect 4433 1493 4447 1507
rect 4313 1453 4327 1467
rect 4333 1434 4347 1448
rect 4393 1433 4407 1447
rect 4433 1434 4447 1448
rect 4753 1912 4767 1926
rect 4833 1912 4847 1926
rect 4793 1833 4807 1847
rect 4793 1793 4807 1807
rect 4713 1753 4727 1767
rect 4633 1734 4647 1748
rect 4693 1734 4707 1748
rect 4653 1692 4667 1706
rect 4513 1673 4527 1687
rect 4513 1613 4527 1627
rect 4293 1392 4307 1406
rect 4353 1392 4367 1406
rect 4313 1353 4327 1367
rect 4453 1392 4467 1406
rect 4413 1333 4427 1347
rect 4313 1313 4327 1327
rect 4393 1313 4407 1327
rect 4293 1233 4307 1247
rect 4273 1213 4287 1227
rect 4213 1172 4227 1186
rect 4253 1172 4267 1186
rect 4353 1273 4367 1287
rect 4553 1493 4567 1507
rect 4533 1434 4547 1448
rect 4613 1453 4627 1467
rect 4573 1434 4587 1448
rect 4693 1453 4707 1467
rect 4653 1433 4667 1447
rect 4533 1393 4547 1407
rect 4573 1333 4587 1347
rect 4473 1233 4487 1247
rect 4513 1233 4527 1247
rect 4453 1214 4467 1228
rect 4373 1172 4387 1186
rect 4453 1173 4467 1187
rect 4313 1113 4327 1127
rect 4533 1214 4547 1228
rect 4553 1172 4567 1186
rect 4553 1113 4567 1127
rect 4493 1073 4507 1087
rect 4753 1734 4767 1748
rect 4853 1833 4867 1847
rect 4833 1693 4847 1707
rect 4773 1673 4787 1687
rect 4833 1653 4847 1667
rect 4733 1493 4747 1507
rect 5013 1954 5027 1968
rect 5073 1993 5087 2007
rect 4993 1912 5007 1926
rect 5053 1913 5067 1927
rect 5013 1793 5027 1807
rect 4893 1753 4907 1767
rect 4953 1734 4967 1748
rect 4893 1692 4907 1706
rect 5093 1954 5107 1968
rect 5213 1954 5227 1968
rect 5273 2212 5287 2226
rect 5313 2212 5327 2226
rect 5353 2212 5367 2226
rect 5393 2212 5407 2226
rect 5453 2393 5467 2407
rect 5433 2353 5447 2367
rect 5613 2833 5627 2847
rect 5753 2953 5767 2967
rect 5713 2933 5727 2947
rect 5713 2833 5727 2847
rect 5673 2732 5687 2746
rect 5633 2693 5647 2707
rect 5613 2653 5627 2667
rect 5593 2633 5607 2647
rect 5553 2513 5567 2527
rect 5613 2473 5627 2487
rect 5533 2393 5547 2407
rect 5613 2433 5627 2447
rect 5573 2373 5587 2387
rect 5493 2333 5507 2347
rect 5453 2313 5467 2327
rect 5493 2293 5507 2307
rect 5433 2273 5447 2287
rect 5473 2273 5487 2287
rect 5373 2073 5387 2087
rect 5273 2033 5287 2047
rect 5193 1912 5207 1926
rect 5153 1853 5167 1867
rect 5213 1853 5227 1867
rect 5313 1954 5327 1968
rect 5333 1912 5347 1926
rect 5333 1873 5347 1887
rect 5293 1833 5307 1847
rect 5233 1773 5247 1787
rect 5293 1773 5307 1787
rect 5073 1753 5087 1767
rect 5153 1753 5167 1767
rect 5213 1753 5227 1767
rect 5113 1734 5127 1748
rect 5013 1673 5027 1687
rect 4973 1593 4987 1607
rect 4933 1453 4947 1467
rect 4853 1434 4867 1448
rect 4913 1434 4927 1448
rect 5093 1673 5107 1687
rect 5093 1613 5107 1627
rect 5053 1573 5067 1587
rect 5253 1734 5267 1748
rect 5233 1613 5247 1627
rect 5193 1573 5207 1587
rect 5153 1493 5167 1507
rect 5153 1453 5167 1467
rect 4693 1392 4707 1406
rect 4753 1392 4767 1406
rect 4673 1333 4687 1347
rect 4633 1273 4647 1287
rect 4613 1253 4627 1267
rect 4913 1373 4927 1387
rect 4753 1293 4767 1307
rect 4793 1293 4807 1307
rect 4613 1173 4627 1187
rect 4593 1133 4607 1147
rect 4633 1133 4647 1147
rect 4573 1033 4587 1047
rect 4173 993 4187 1007
rect 4293 993 4307 1007
rect 4473 993 4487 1007
rect 4153 933 4167 947
rect 4093 914 4107 928
rect 4133 914 4147 928
rect 4253 933 4267 947
rect 3953 873 3967 887
rect 3993 872 4007 886
rect 3973 753 3987 767
rect 3953 733 3967 747
rect 4333 914 4347 928
rect 4393 914 4407 928
rect 4453 914 4467 928
rect 4493 914 4507 928
rect 4593 973 4607 987
rect 4673 1053 4687 1067
rect 4973 1392 4987 1406
rect 5033 1434 5047 1448
rect 5053 1392 5067 1406
rect 5093 1353 5107 1367
rect 4993 1313 5007 1327
rect 5033 1273 5047 1287
rect 4793 1253 4807 1267
rect 4933 1253 4947 1267
rect 4833 1233 4847 1247
rect 4793 1214 4807 1228
rect 4993 1233 5007 1247
rect 4873 1213 4887 1227
rect 4873 1172 4887 1186
rect 4913 1172 4927 1186
rect 4953 1172 4967 1186
rect 5133 1253 5147 1267
rect 5093 1214 5107 1228
rect 4873 1133 4887 1147
rect 4953 1053 4967 1067
rect 4693 993 4707 1007
rect 4753 993 4767 1007
rect 4153 872 4167 886
rect 4253 872 4267 886
rect 4313 872 4327 886
rect 4213 853 4227 867
rect 4093 833 4107 847
rect 4193 833 4207 847
rect 4073 753 4087 767
rect 3893 694 3907 708
rect 3933 694 3947 708
rect 3693 652 3707 666
rect 3733 652 3747 666
rect 3772 652 3786 666
rect 3793 652 3807 666
rect 3833 652 3847 666
rect 3913 653 3927 667
rect 4013 694 4027 708
rect 3673 613 3687 627
rect 3633 533 3647 547
rect 3553 493 3567 507
rect 3573 433 3587 447
rect 3533 394 3547 408
rect 3513 353 3527 367
rect 3493 333 3507 347
rect 3373 273 3387 287
rect 3453 273 3467 287
rect 3453 233 3467 247
rect 2873 132 2887 146
rect 2853 93 2867 107
rect 2773 53 2787 67
rect 1753 33 1767 47
rect 2633 33 2647 47
rect 2693 33 2707 47
rect 2953 132 2967 146
rect 2913 92 2927 106
rect 2893 73 2907 87
rect 3133 132 3147 146
rect 3373 174 3387 188
rect 3413 174 3427 188
rect 3213 132 3227 146
rect 3253 132 3267 146
rect 3313 132 3327 146
rect 3153 113 3167 127
rect 3353 113 3367 127
rect 3633 353 3647 367
rect 3553 333 3567 347
rect 4033 633 4047 647
rect 3713 573 3727 587
rect 3913 573 3927 587
rect 3673 513 3687 527
rect 3673 473 3687 487
rect 3953 533 3967 547
rect 3773 513 3787 527
rect 3713 413 3727 427
rect 3693 394 3707 408
rect 3753 394 3767 408
rect 3653 313 3667 327
rect 3873 493 3887 507
rect 3833 394 3847 408
rect 3933 453 3947 467
rect 4133 694 4147 708
rect 4113 652 4127 666
rect 4253 793 4267 807
rect 4293 733 4307 747
rect 4333 713 4347 727
rect 4373 873 4387 887
rect 4413 893 4427 907
rect 4393 833 4407 847
rect 4633 914 4647 928
rect 4453 833 4467 847
rect 4413 753 4427 767
rect 4453 753 4467 767
rect 4373 733 4387 747
rect 4333 673 4347 687
rect 4213 653 4227 667
rect 4193 633 4207 647
rect 4273 652 4287 666
rect 4313 653 4327 667
rect 4073 613 4087 627
rect 4153 613 4167 627
rect 4053 573 4067 587
rect 3993 493 4007 507
rect 4033 493 4047 507
rect 3953 394 3967 408
rect 4073 513 4087 527
rect 4133 473 4147 487
rect 4273 473 4287 487
rect 4173 413 4187 427
rect 4213 413 4227 427
rect 3773 353 3787 366
rect 3773 352 3787 353
rect 3813 352 3827 366
rect 3853 352 3867 366
rect 3933 353 3947 367
rect 4133 394 4147 408
rect 4413 694 4427 708
rect 4433 652 4447 666
rect 4473 653 4487 667
rect 4393 613 4407 627
rect 4553 872 4567 886
rect 4593 833 4607 847
rect 4513 813 4527 827
rect 4513 753 4527 767
rect 4493 573 4507 587
rect 4333 433 4347 447
rect 4313 413 4327 427
rect 4013 352 4027 366
rect 4073 352 4087 366
rect 3793 293 3807 307
rect 3973 293 3987 307
rect 3753 273 3767 287
rect 4213 352 4227 366
rect 4153 313 4167 327
rect 3733 253 3747 267
rect 3833 253 3847 267
rect 3913 253 3927 267
rect 3993 253 4007 267
rect 4053 253 4067 267
rect 4113 253 4127 267
rect 3752 233 3766 247
rect 3773 233 3787 247
rect 3513 213 3527 227
rect 3553 193 3567 207
rect 3473 173 3487 187
rect 3513 174 3527 188
rect 3693 193 3707 207
rect 3613 173 3627 187
rect 3653 174 3667 188
rect 3753 174 3767 188
rect 3453 113 3467 127
rect 3533 132 3547 146
rect 3573 132 3587 146
rect 3533 113 3547 127
rect 3053 93 3067 107
rect 3133 93 3147 107
rect 3273 93 3287 107
rect 2993 53 3007 67
rect 3033 53 3047 67
rect 3373 92 3387 106
rect 3473 93 3487 107
rect 2893 33 2907 47
rect 3053 33 3067 47
rect 3373 33 3387 47
rect 3413 33 3427 47
rect 3873 174 3887 188
rect 3673 113 3687 127
rect 3773 132 3787 146
rect 3813 132 3827 146
rect 3853 132 3867 146
rect 3713 93 3727 107
rect 3933 213 3947 227
rect 4033 174 4047 188
rect 4193 213 4207 227
rect 4153 174 4167 188
rect 4293 352 4307 366
rect 4473 433 4487 447
rect 4393 394 4407 408
rect 4433 394 4447 408
rect 4493 394 4507 408
rect 4653 872 4667 886
rect 4653 733 4667 747
rect 4553 694 4567 708
rect 4593 694 4607 708
rect 4613 652 4627 666
rect 4713 973 4727 987
rect 4853 973 4867 987
rect 4773 914 4787 928
rect 4813 914 4827 928
rect 4753 872 4767 886
rect 4753 833 4767 847
rect 4713 793 4727 807
rect 4713 733 4727 747
rect 4913 914 4927 928
rect 4933 873 4947 887
rect 4853 833 4867 847
rect 4893 833 4907 847
rect 4893 793 4907 807
rect 4933 793 4947 807
rect 4992 1172 5006 1186
rect 5013 1173 5027 1187
rect 5113 1172 5127 1186
rect 5093 1153 5107 1167
rect 5013 1133 5027 1147
rect 5053 1132 5067 1146
rect 5013 1073 5027 1087
rect 4973 1033 4987 1047
rect 5093 1053 5107 1067
rect 5053 914 5067 928
rect 5133 1013 5147 1027
rect 5533 2293 5547 2307
rect 5513 2273 5527 2287
rect 5493 2254 5507 2268
rect 5433 2173 5447 2187
rect 5473 2173 5487 2187
rect 5593 2333 5607 2347
rect 5733 2813 5747 2827
rect 5813 3113 5827 3127
rect 5773 2873 5787 2887
rect 5973 3413 5987 3427
rect 6013 3393 6027 3407
rect 5973 3373 5987 3387
rect 5933 3293 5947 3307
rect 6053 3333 6067 3347
rect 6053 3293 6067 3307
rect 5933 3232 5947 3246
rect 5913 3073 5927 3087
rect 5873 3053 5887 3067
rect 5813 2993 5827 3007
rect 5953 3153 5967 3167
rect 6113 3873 6127 3887
rect 6093 3853 6107 3867
rect 6093 3813 6107 3827
rect 6133 3853 6147 3867
rect 6213 3853 6227 3867
rect 6153 3833 6167 3847
rect 6153 3814 6167 3828
rect 6133 3772 6147 3786
rect 6193 3693 6207 3707
rect 6173 3653 6187 3667
rect 6093 3473 6107 3487
rect 6173 3473 6187 3487
rect 6133 3413 6147 3427
rect 6093 3393 6107 3407
rect 6093 3293 6107 3307
rect 6173 3293 6187 3307
rect 6053 3233 6067 3247
rect 6033 3173 6047 3187
rect 6013 3053 6027 3067
rect 5953 2993 5967 3007
rect 6073 3133 6087 3147
rect 6053 3073 6067 3087
rect 6053 2993 6067 3007
rect 5833 2893 5847 2907
rect 5813 2833 5827 2847
rect 5793 2813 5807 2827
rect 5833 2793 5847 2807
rect 5753 2774 5767 2788
rect 5813 2774 5827 2788
rect 5753 2732 5767 2746
rect 5733 2693 5747 2707
rect 5713 2673 5727 2687
rect 5693 2533 5707 2547
rect 5633 2413 5647 2427
rect 5693 2393 5707 2407
rect 5653 2373 5667 2387
rect 5633 2293 5647 2307
rect 5633 2272 5647 2286
rect 5433 1954 5447 1968
rect 5533 1912 5547 1926
rect 5413 1853 5427 1867
rect 5373 1833 5387 1847
rect 5593 1853 5607 1867
rect 5393 1753 5407 1767
rect 5453 1753 5467 1767
rect 5493 1753 5507 1767
rect 5413 1733 5427 1747
rect 5533 1734 5547 1748
rect 5593 1733 5607 1747
rect 5333 1692 5347 1706
rect 5373 1692 5387 1706
rect 5453 1692 5467 1706
rect 5233 1493 5247 1507
rect 5193 1434 5207 1448
rect 5213 1293 5227 1307
rect 5233 1253 5247 1267
rect 5193 1214 5207 1228
rect 5293 1493 5307 1507
rect 5553 1692 5567 1706
rect 5493 1573 5507 1587
rect 5333 1473 5347 1487
rect 5333 1434 5347 1448
rect 5373 1434 5387 1448
rect 5433 1434 5447 1448
rect 5293 1392 5307 1406
rect 5353 1392 5367 1406
rect 5453 1373 5467 1387
rect 5393 1333 5407 1347
rect 5313 1214 5327 1228
rect 5353 1214 5367 1228
rect 5433 1353 5447 1367
rect 5473 1353 5487 1367
rect 5453 1313 5467 1327
rect 5473 1253 5487 1267
rect 5413 1233 5427 1247
rect 5453 1233 5467 1247
rect 5293 1193 5307 1207
rect 5213 1172 5227 1186
rect 5293 1133 5307 1147
rect 5333 1173 5347 1187
rect 5373 1133 5387 1147
rect 5173 1093 5187 1107
rect 5253 1093 5267 1107
rect 5313 1093 5327 1107
rect 5133 914 5147 928
rect 5373 1073 5387 1087
rect 5353 1033 5367 1047
rect 5333 1013 5347 1027
rect 5253 993 5267 1007
rect 5213 973 5227 987
rect 5173 913 5187 927
rect 5033 872 5047 886
rect 5093 872 5107 886
rect 5153 872 5167 886
rect 4993 833 5007 847
rect 4953 773 4967 787
rect 4873 753 4887 767
rect 4913 713 4927 727
rect 4973 713 4987 727
rect 4573 573 4587 587
rect 4553 433 4567 447
rect 4353 313 4367 327
rect 4273 253 4287 267
rect 4253 193 4267 207
rect 4233 173 4247 187
rect 4013 132 4027 146
rect 4073 132 4087 146
rect 3933 93 3947 107
rect 4173 132 4187 146
rect 4133 113 4147 127
rect 4313 213 4327 227
rect 4413 213 4427 227
rect 4273 173 4287 187
rect 4593 394 4607 408
rect 4653 652 4667 666
rect 4693 653 4707 667
rect 4733 652 4747 666
rect 4813 652 4827 666
rect 4893 652 4907 666
rect 4693 613 4707 627
rect 4773 613 4787 627
rect 4813 613 4827 627
rect 4673 573 4687 587
rect 4693 513 4707 527
rect 4793 513 4807 527
rect 4713 433 4727 447
rect 4673 394 4687 408
rect 4753 394 4767 408
rect 4533 352 4547 366
rect 4573 352 4587 366
rect 4633 352 4647 366
rect 4733 352 4747 366
rect 4533 313 4547 327
rect 4692 313 4706 327
rect 4713 313 4727 327
rect 4493 293 4507 307
rect 4353 193 4367 207
rect 4473 193 4487 207
rect 4513 193 4527 207
rect 4253 132 4267 146
rect 4293 132 4307 146
rect 4333 132 4347 146
rect 4453 174 4467 188
rect 4473 132 4487 146
rect 4233 93 4247 107
rect 4433 93 4447 107
rect 4672 293 4686 307
rect 4593 273 4607 287
rect 5073 793 5087 807
rect 5013 753 5027 767
rect 4993 693 5007 707
rect 5033 694 5047 708
rect 5093 773 5107 787
rect 5113 693 5127 707
rect 5173 694 5187 708
rect 5233 953 5247 967
rect 5233 913 5247 927
rect 5293 914 5307 928
rect 5333 913 5347 927
rect 5233 873 5247 887
rect 5333 873 5347 887
rect 5333 813 5347 827
rect 5313 773 5327 787
rect 5273 733 5287 747
rect 5433 1173 5447 1187
rect 5413 1053 5427 1067
rect 5453 1133 5467 1147
rect 5553 1393 5567 1407
rect 5513 1293 5527 1307
rect 5533 1273 5547 1287
rect 5513 1233 5527 1247
rect 5493 1213 5507 1227
rect 5633 2212 5647 2226
rect 5833 2732 5847 2746
rect 5893 2952 5907 2966
rect 5933 2953 5947 2967
rect 5873 2933 5887 2947
rect 5893 2893 5907 2907
rect 5873 2733 5887 2747
rect 6013 2952 6027 2966
rect 6133 3233 6147 3247
rect 6113 3213 6127 3227
rect 6113 3173 6127 3187
rect 6113 3133 6127 3147
rect 6093 3113 6107 3127
rect 6153 3193 6167 3207
rect 6113 3013 6127 3027
rect 6232 3814 6246 3828
rect 6293 3853 6307 3867
rect 6253 3813 6267 3827
rect 6233 3773 6247 3787
rect 6273 3772 6287 3786
rect 6313 3773 6327 3787
rect 6213 3653 6227 3667
rect 6233 3553 6247 3567
rect 6273 3514 6287 3528
rect 6293 3473 6307 3487
rect 6273 3433 6287 3447
rect 6213 3313 6227 3327
rect 6253 3313 6267 3327
rect 6313 3373 6327 3387
rect 6253 3252 6267 3266
rect 6193 3153 6207 3167
rect 6173 2994 6187 3008
rect 6113 2952 6127 2966
rect 6153 2952 6167 2966
rect 6293 3193 6307 3207
rect 6253 3133 6267 3147
rect 6233 2993 6247 3007
rect 6313 3113 6327 3127
rect 6133 2933 6147 2947
rect 6073 2833 6087 2847
rect 5973 2793 5987 2807
rect 6033 2774 6047 2788
rect 6093 2774 6107 2788
rect 6173 2913 6187 2927
rect 6153 2833 6167 2847
rect 5853 2693 5867 2707
rect 5773 2653 5787 2667
rect 5853 2493 5867 2507
rect 5773 2474 5787 2488
rect 5833 2413 5847 2427
rect 5873 2413 5887 2427
rect 5933 2732 5947 2746
rect 6153 2773 6167 2787
rect 6053 2733 6067 2747
rect 6113 2732 6127 2746
rect 5933 2493 5947 2507
rect 5773 2393 5787 2407
rect 5853 2393 5867 2407
rect 5913 2393 5927 2407
rect 5813 2254 5827 2268
rect 6073 2693 6087 2707
rect 6053 2673 6067 2687
rect 5973 2533 5987 2547
rect 6013 2474 6027 2488
rect 5933 2333 5947 2347
rect 6173 2713 6187 2727
rect 6253 2933 6267 2947
rect 6313 2913 6327 2927
rect 6273 2893 6287 2907
rect 6253 2774 6267 2788
rect 6313 2773 6327 2787
rect 6213 2693 6227 2707
rect 6153 2513 6167 2527
rect 6093 2493 6107 2507
rect 6073 2413 6087 2427
rect 6033 2373 6047 2387
rect 5993 2353 6007 2367
rect 5913 2293 5927 2307
rect 5953 2293 5967 2307
rect 5893 2253 5907 2267
rect 5733 2073 5747 2087
rect 5733 1954 5747 1968
rect 5633 1912 5647 1926
rect 5653 1853 5667 1867
rect 5673 1753 5687 1767
rect 5653 1653 5667 1667
rect 5593 1633 5607 1647
rect 5613 1473 5627 1487
rect 5733 1693 5747 1707
rect 5713 1673 5727 1687
rect 5673 1573 5687 1587
rect 5653 1434 5667 1448
rect 5593 1393 5607 1407
rect 5573 1213 5587 1227
rect 5513 1172 5527 1186
rect 5553 1172 5567 1186
rect 5633 1392 5647 1406
rect 5633 1353 5647 1367
rect 5613 1233 5627 1247
rect 5673 1293 5687 1307
rect 5733 1653 5747 1667
rect 5893 2193 5907 2207
rect 5953 2254 5967 2268
rect 5993 2254 6007 2268
rect 6053 2254 6067 2268
rect 6193 2493 6207 2507
rect 6213 2473 6227 2487
rect 6093 2373 6107 2387
rect 6093 2273 6107 2287
rect 5913 2113 5927 2127
rect 5793 2033 5807 2047
rect 6033 2213 6047 2227
rect 5993 2193 6007 2207
rect 5993 2113 6007 2127
rect 5813 1953 5827 1967
rect 5893 1954 5907 1968
rect 5833 1912 5847 1926
rect 6033 1953 6047 1967
rect 5833 1893 5847 1907
rect 5793 1853 5807 1867
rect 5873 1853 5887 1867
rect 5833 1734 5847 1748
rect 5933 1853 5947 1867
rect 5893 1793 5907 1807
rect 5913 1734 5927 1748
rect 5773 1673 5787 1687
rect 5813 1633 5827 1647
rect 5873 1673 5887 1687
rect 5853 1653 5867 1667
rect 5793 1473 5807 1487
rect 5753 1434 5767 1448
rect 5833 1593 5847 1607
rect 5833 1553 5847 1567
rect 5813 1453 5827 1467
rect 5773 1392 5787 1406
rect 5813 1392 5827 1406
rect 5853 1393 5867 1407
rect 5913 1653 5927 1667
rect 5913 1632 5927 1646
rect 5893 1553 5907 1567
rect 5893 1513 5907 1527
rect 5973 1893 5987 1907
rect 6013 1853 6027 1867
rect 6133 2432 6147 2446
rect 6172 2413 6186 2427
rect 6193 2413 6207 2427
rect 6173 2273 6187 2287
rect 6113 2193 6127 2207
rect 6093 2073 6107 2087
rect 6073 2053 6087 2067
rect 6073 1993 6087 2007
rect 6113 1993 6127 2007
rect 6153 2193 6167 2207
rect 6153 2033 6167 2047
rect 6153 1973 6167 1987
rect 6073 1953 6087 1967
rect 6133 1953 6147 1967
rect 6173 1954 6187 1968
rect 6073 1913 6087 1927
rect 6053 1793 6067 1807
rect 6033 1753 6047 1767
rect 5953 1733 5967 1747
rect 5993 1734 6007 1748
rect 6113 1912 6127 1926
rect 6153 1912 6167 1926
rect 6113 1853 6127 1867
rect 6093 1753 6107 1767
rect 6073 1712 6087 1726
rect 5953 1693 5967 1707
rect 5973 1653 5987 1667
rect 5953 1633 5967 1647
rect 6013 1632 6027 1646
rect 5993 1593 6007 1607
rect 6033 1573 6047 1587
rect 5993 1533 6007 1547
rect 5973 1513 5987 1527
rect 5993 1493 6007 1507
rect 5933 1453 5947 1467
rect 5953 1434 5967 1448
rect 6013 1453 6027 1467
rect 5993 1433 6007 1447
rect 5733 1373 5747 1387
rect 5753 1333 5767 1347
rect 5673 1253 5687 1267
rect 5573 1133 5587 1147
rect 5553 1113 5567 1127
rect 5433 1013 5447 1027
rect 5533 1013 5547 1027
rect 5393 993 5407 1007
rect 5373 953 5387 967
rect 5433 973 5447 987
rect 5493 933 5507 947
rect 5413 872 5427 886
rect 5453 872 5467 886
rect 5493 873 5507 887
rect 5473 833 5487 847
rect 5373 813 5387 827
rect 5413 813 5427 827
rect 5393 773 5407 787
rect 5373 733 5387 747
rect 5353 713 5367 727
rect 5233 694 5247 708
rect 5293 694 5307 708
rect 5333 694 5347 708
rect 5013 652 5027 666
rect 5053 652 5067 666
rect 5093 652 5107 666
rect 4973 613 4987 627
rect 5133 632 5147 646
rect 5113 613 5127 627
rect 4933 573 4947 587
rect 4913 394 4927 408
rect 5093 573 5107 587
rect 5313 652 5327 666
rect 5193 573 5207 587
rect 5253 573 5267 587
rect 5333 633 5347 647
rect 5313 553 5327 567
rect 5133 433 5147 447
rect 4993 394 5007 408
rect 5053 394 5067 408
rect 5093 394 5107 408
rect 5273 413 5287 427
rect 5233 394 5247 408
rect 4813 352 4827 366
rect 4893 352 4907 366
rect 4953 352 4967 366
rect 5013 352 5027 366
rect 4853 313 4867 327
rect 5353 573 5367 587
rect 5413 713 5427 727
rect 5473 713 5487 727
rect 5553 993 5567 1007
rect 5533 913 5547 927
rect 5593 973 5607 987
rect 5693 1153 5707 1167
rect 5653 1033 5667 1047
rect 5613 953 5627 967
rect 5653 953 5667 967
rect 5613 853 5627 867
rect 5573 813 5587 827
rect 5553 773 5567 787
rect 5533 753 5547 767
rect 5513 694 5527 708
rect 5633 813 5647 827
rect 5613 733 5627 747
rect 5593 694 5607 708
rect 5673 933 5687 947
rect 5653 773 5667 787
rect 5733 1153 5747 1167
rect 5713 1113 5727 1127
rect 5853 1333 5867 1347
rect 5833 1313 5847 1327
rect 5773 1273 5787 1287
rect 5813 1273 5827 1287
rect 5833 1253 5847 1267
rect 5813 1172 5827 1186
rect 5853 1172 5867 1186
rect 5913 1373 5927 1387
rect 5953 1373 5967 1387
rect 5933 1273 5947 1287
rect 5973 1353 5987 1367
rect 5973 1313 5987 1327
rect 5953 1253 5967 1267
rect 5993 1293 6007 1307
rect 5913 1213 5927 1227
rect 5993 1214 6007 1228
rect 6073 1653 6087 1667
rect 6073 1573 6087 1587
rect 6053 1493 6067 1507
rect 6293 2713 6307 2727
rect 6273 2693 6287 2707
rect 6273 2513 6287 2527
rect 6293 2413 6307 2427
rect 6273 2273 6287 2287
rect 6253 2254 6267 2268
rect 6313 2253 6327 2267
rect 6253 2193 6267 2207
rect 6313 2213 6327 2227
rect 6233 2073 6247 2087
rect 6273 2053 6287 2067
rect 6253 1973 6267 1987
rect 6233 1954 6247 1968
rect 6293 1953 6307 1967
rect 6213 1912 6227 1926
rect 6253 1912 6267 1926
rect 6193 1853 6207 1867
rect 6173 1813 6187 1827
rect 6133 1793 6147 1807
rect 6173 1734 6187 1748
rect 6293 1893 6307 1907
rect 6233 1813 6247 1827
rect 6213 1733 6227 1747
rect 6113 1673 6127 1687
rect 6113 1533 6127 1547
rect 6093 1453 6107 1467
rect 6193 1692 6207 1706
rect 6213 1693 6227 1707
rect 6173 1673 6187 1687
rect 6153 1452 6167 1466
rect 6053 1392 6067 1406
rect 6093 1392 6107 1406
rect 6153 1392 6167 1406
rect 6053 1353 6067 1367
rect 6133 1352 6147 1366
rect 6073 1313 6087 1327
rect 6113 1313 6127 1327
rect 6113 1273 6127 1287
rect 6153 1333 6167 1347
rect 6193 1653 6207 1667
rect 6193 1433 6207 1447
rect 6253 1773 6267 1787
rect 6313 1773 6327 1787
rect 6293 1753 6307 1767
rect 6313 1733 6327 1747
rect 6233 1633 6247 1647
rect 6233 1573 6247 1587
rect 6273 1692 6287 1706
rect 6313 1693 6327 1707
rect 6293 1653 6307 1667
rect 6293 1533 6307 1547
rect 6253 1473 6267 1487
rect 6293 1473 6307 1487
rect 6293 1433 6307 1447
rect 6193 1393 6207 1407
rect 6193 1353 6207 1367
rect 6253 1353 6267 1367
rect 6233 1333 6247 1347
rect 5913 1173 5927 1187
rect 5773 1113 5787 1127
rect 5753 1073 5767 1087
rect 5693 913 5707 927
rect 5773 933 5787 947
rect 5693 873 5707 887
rect 5453 652 5467 666
rect 5533 652 5547 666
rect 5573 652 5587 666
rect 5473 633 5487 647
rect 5553 633 5567 647
rect 5413 413 5427 427
rect 5373 394 5387 408
rect 5753 853 5767 867
rect 5833 1053 5847 1067
rect 5893 1033 5907 1047
rect 5853 953 5867 967
rect 5853 913 5867 927
rect 5933 1153 5947 1167
rect 5913 953 5927 967
rect 6073 1214 6087 1228
rect 6213 1273 6227 1287
rect 6172 1253 6186 1267
rect 6193 1253 6207 1267
rect 6153 1213 6167 1227
rect 6033 1153 6047 1167
rect 5973 1113 5987 1127
rect 5993 1013 6007 1027
rect 5933 914 5947 928
rect 5973 914 5987 928
rect 5713 833 5727 847
rect 5793 694 5807 708
rect 5733 673 5747 687
rect 5813 652 5827 666
rect 5693 633 5707 647
rect 5773 633 5787 647
rect 5953 873 5967 887
rect 5873 813 5887 827
rect 5913 813 5927 827
rect 5853 753 5867 767
rect 5953 793 5967 807
rect 6073 1153 6087 1167
rect 6053 993 6067 1007
rect 6033 914 6047 928
rect 6093 1113 6107 1127
rect 6153 1173 6167 1187
rect 6133 953 6147 967
rect 6013 872 6027 886
rect 6053 872 6067 886
rect 6093 872 6107 886
rect 5993 813 6007 827
rect 5893 733 5907 747
rect 5933 713 5947 727
rect 5613 513 5627 527
rect 5513 493 5527 507
rect 5693 473 5707 487
rect 5553 394 5567 408
rect 5633 394 5647 408
rect 5753 453 5767 467
rect 5713 413 5727 427
rect 5733 394 5747 408
rect 5113 313 5127 327
rect 5052 293 5066 307
rect 5073 293 5087 307
rect 4813 253 4827 267
rect 4633 213 4647 227
rect 4713 213 4727 227
rect 4793 213 4807 227
rect 4753 174 4767 188
rect 4533 132 4547 146
rect 4573 132 4587 146
rect 4773 113 4787 127
rect 4913 233 4927 247
rect 5033 233 5047 247
rect 4833 173 4847 187
rect 4873 174 4887 188
rect 5173 233 5187 247
rect 5113 173 5127 187
rect 5253 352 5267 366
rect 5333 352 5347 366
rect 5373 333 5387 347
rect 5213 193 5227 207
rect 4573 93 4587 107
rect 4613 93 4627 107
rect 4733 93 4747 107
rect 4813 93 4827 107
rect 4453 73 4467 87
rect 4513 73 4527 87
rect 4093 53 4107 67
rect 4893 132 4907 146
rect 4933 132 4947 146
rect 5013 132 5027 146
rect 5053 113 5067 127
rect 5153 132 5167 146
rect 5273 174 5287 188
rect 5333 174 5347 188
rect 5413 293 5427 307
rect 5193 113 5207 127
rect 5113 73 5127 87
rect 5313 132 5327 146
rect 5353 113 5367 127
rect 5313 73 5327 87
rect 5473 353 5487 367
rect 5533 352 5547 366
rect 5533 293 5547 307
rect 5433 253 5447 267
rect 5493 174 5507 188
rect 5793 413 5807 427
rect 5773 373 5787 387
rect 5673 352 5687 366
rect 5713 352 5727 366
rect 5753 352 5767 366
rect 5873 693 5887 707
rect 5913 693 5927 707
rect 5893 652 5907 666
rect 5933 613 5947 627
rect 5933 493 5947 507
rect 5813 393 5827 407
rect 5853 393 5867 407
rect 5913 393 5927 407
rect 5813 353 5827 367
rect 5653 313 5667 327
rect 5793 313 5807 327
rect 5633 293 5647 307
rect 5573 253 5587 267
rect 5673 293 5687 307
rect 5673 253 5687 267
rect 5873 313 5887 327
rect 5833 233 5847 247
rect 6173 1133 6187 1147
rect 6153 853 6167 867
rect 6013 453 6027 467
rect 5993 394 6007 408
rect 6293 1393 6307 1407
rect 6273 1273 6287 1287
rect 6293 1253 6307 1267
rect 6233 1214 6247 1228
rect 6313 1213 6327 1227
rect 6233 1153 6247 1167
rect 6253 1133 6267 1147
rect 6313 1153 6327 1167
rect 6293 1073 6307 1087
rect 6253 1013 6267 1027
rect 6213 914 6227 928
rect 6313 993 6327 1007
rect 6293 913 6307 927
rect 6173 833 6187 847
rect 6133 773 6147 787
rect 6073 753 6087 767
rect 6173 613 6187 627
rect 6113 573 6127 587
rect 6213 853 6227 867
rect 6193 493 6207 507
rect 6053 413 6067 427
rect 6133 413 6147 427
rect 6173 394 6187 408
rect 5973 293 5987 307
rect 6073 353 6087 367
rect 6113 352 6127 366
rect 6033 333 6047 347
rect 6013 273 6027 287
rect 5953 193 5967 207
rect 5593 153 5607 167
rect 5453 133 5467 147
rect 5473 113 5487 127
rect 6133 313 6147 327
rect 6093 273 6107 287
rect 6153 273 6167 287
rect 6273 872 6287 886
rect 6313 873 6327 887
rect 6293 853 6307 867
rect 6233 833 6247 847
rect 6253 813 6267 827
rect 6233 413 6247 427
rect 6213 213 6227 227
rect 6273 713 6287 727
rect 6253 313 6267 327
rect 6173 174 6187 188
rect 6233 174 6247 188
rect 5773 132 5787 146
rect 5633 113 5647 127
rect 5713 113 5727 127
rect 5513 92 5527 106
rect 5593 93 5607 107
rect 5413 53 5427 67
rect 5813 53 5827 67
rect 6033 132 6047 146
rect 6073 132 6087 146
rect 6113 132 6127 146
rect 5973 93 5987 107
rect 6213 132 6227 146
rect 6173 53 6187 67
rect 6293 93 6307 107
rect 3913 33 3927 47
rect 4833 33 4847 47
rect 5273 33 5287 47
rect 5933 33 5947 47
rect 6273 33 6287 47
rect 2913 13 2927 27
rect 3393 13 3407 27
rect 3433 13 3447 27
rect 3613 13 3627 27
<< metal3 >>
rect 1707 6256 1793 6264
rect 3347 6256 3673 6264
rect 5047 6256 5073 6264
rect 1647 6216 1833 6224
rect 1487 6196 1713 6204
rect 2367 6196 2953 6204
rect 5707 6196 5733 6204
rect 5747 6196 6033 6204
rect 127 6176 713 6184
rect 1927 6176 4393 6184
rect 5020 6184 5033 6187
rect 5016 6173 5033 6184
rect 387 6156 653 6164
rect 827 6156 1233 6164
rect 1247 6156 1673 6164
rect 687 6136 753 6144
rect 1367 6136 1433 6144
rect 2727 6137 2753 6145
rect 3327 6136 3373 6144
rect 3387 6136 3873 6144
rect 367 6117 413 6125
rect 467 6117 513 6125
rect 576 6116 713 6124
rect 356 6104 364 6114
rect 556 6104 564 6114
rect 356 6096 564 6104
rect 576 6086 584 6116
rect 927 6117 953 6125
rect 1007 6116 1053 6124
rect 1067 6117 1093 6125
rect 1407 6116 1513 6124
rect 1567 6117 1613 6125
rect 1836 6116 1873 6124
rect 667 6096 813 6104
rect 916 6104 924 6114
rect 1136 6104 1144 6114
rect 916 6096 1144 6104
rect 947 6075 973 6083
rect 1276 6084 1284 6114
rect 1127 6076 1284 6084
rect 1307 6075 1373 6083
rect 1427 6076 1473 6084
rect 1836 6084 1844 6116
rect 1987 6117 2073 6125
rect 2287 6120 2344 6124
rect 2287 6116 2347 6120
rect 2333 6107 2347 6116
rect 1747 6076 1844 6084
rect 1867 6075 1913 6083
rect 2167 6076 2253 6084
rect 2267 6076 2313 6084
rect 2556 6084 2564 6094
rect 2907 6096 2933 6104
rect 3007 6097 3153 6105
rect 3316 6107 3324 6134
rect 3887 6136 3973 6144
rect 5016 6144 5024 6173
rect 5047 6156 5293 6164
rect 6007 6156 6153 6164
rect 5016 6136 5053 6144
rect 5787 6136 5933 6144
rect 5947 6136 6093 6144
rect 6107 6136 6253 6144
rect 4507 6116 4633 6124
rect 5367 6117 5393 6125
rect 5487 6117 5553 6125
rect 5576 6116 5593 6124
rect 3307 6096 3324 6107
rect 3336 6096 3533 6104
rect 3307 6093 3320 6096
rect 2556 6076 2653 6084
rect 3336 6084 3344 6096
rect 3847 6097 4133 6105
rect 4667 6095 4793 6103
rect 3287 6076 3344 6084
rect 3727 6076 4293 6084
rect 4407 6076 4473 6084
rect 5053 6084 5067 6093
rect 5576 6087 5584 6116
rect 6047 6116 6073 6124
rect 5053 6080 5133 6084
rect 5056 6076 5133 6080
rect 5407 6076 5453 6084
rect 5627 6076 5713 6084
rect 5836 6084 5844 6113
rect 5727 6076 5853 6084
rect 5907 6075 5933 6083
rect 6187 6076 6273 6084
rect 6356 6084 6364 6124
rect 6287 6076 6364 6084
rect 607 6056 913 6064
rect 1267 6056 1613 6064
rect 3407 6056 3673 6064
rect 3787 6056 3893 6064
rect 4387 6056 4713 6064
rect 287 6036 373 6044
rect 747 6036 873 6044
rect 947 6036 1053 6044
rect 5347 6036 5673 6044
rect 5716 6036 6012 6044
rect 367 6016 452 6024
rect 487 6016 593 6024
rect 1027 6016 1353 6024
rect 1367 6016 1533 6024
rect 1627 6016 1993 6024
rect 2456 6020 2713 6024
rect 2453 6016 2713 6020
rect 2453 6007 2467 6016
rect 2727 6016 2853 6024
rect 3427 6016 3773 6024
rect 5716 6024 5724 6036
rect 6047 6036 6133 6044
rect 4807 6016 5724 6024
rect 5867 6016 5973 6024
rect 647 5996 673 6004
rect 687 5996 713 6004
rect 947 5996 1333 6004
rect 1387 5996 1593 6004
rect 2767 5996 3033 6004
rect 3047 5996 3293 6004
rect 4007 5996 4373 6004
rect 4687 5996 4833 6004
rect 5367 5996 5472 6004
rect 5507 5996 5593 6004
rect 5647 5996 5753 6004
rect 867 5976 893 5984
rect 2607 5976 2833 5984
rect 2847 5976 2913 5984
rect 3227 5976 3273 5984
rect 4127 5976 4853 5984
rect 627 5956 993 5964
rect 1327 5956 1453 5964
rect 1507 5956 1713 5964
rect 1767 5956 1973 5964
rect 2027 5956 2073 5964
rect 2087 5956 2193 5964
rect 3347 5956 3453 5964
rect 4907 5956 4973 5964
rect 4987 5956 5573 5964
rect 107 5936 433 5944
rect 587 5936 1113 5944
rect 1487 5936 1533 5944
rect 1547 5936 1733 5944
rect 2067 5936 2253 5944
rect 2736 5936 2993 5944
rect 836 5916 1033 5924
rect 187 5897 253 5905
rect 836 5907 844 5916
rect 2736 5924 2744 5936
rect 3107 5936 3313 5944
rect 3887 5936 3933 5944
rect 4587 5936 4733 5944
rect 5087 5936 5173 5944
rect 5187 5936 5253 5944
rect 5527 5936 5813 5944
rect 5827 5936 5953 5944
rect 2547 5916 2744 5924
rect 3587 5916 3713 5924
rect 3727 5916 4053 5924
rect 5647 5916 5913 5924
rect 6027 5916 6093 5924
rect 787 5896 833 5904
rect 136 5867 144 5894
rect 376 5867 384 5894
rect 676 5867 684 5894
rect 136 5856 153 5867
rect 140 5853 153 5856
rect 247 5855 313 5863
rect 367 5856 384 5867
rect 367 5853 380 5856
rect 407 5856 533 5864
rect 547 5856 573 5864
rect 676 5856 693 5867
rect 680 5853 693 5856
rect 887 5856 993 5864
rect 1007 5855 1033 5863
rect 1056 5847 1064 5894
rect 1076 5866 1084 5913
rect 1187 5896 1253 5904
rect 1267 5896 1373 5904
rect 1747 5896 1853 5904
rect 2087 5897 2113 5905
rect 2307 5896 2404 5904
rect 1127 5855 1193 5863
rect 1267 5855 1293 5863
rect 1436 5864 1444 5894
rect 1347 5856 1444 5864
rect 1547 5855 1573 5863
rect 2007 5856 2073 5864
rect 2156 5864 2164 5894
rect 2396 5866 2404 5896
rect 2427 5897 2513 5905
rect 2767 5897 2813 5905
rect 2867 5896 3133 5904
rect 3147 5897 3173 5905
rect 3327 5897 3373 5905
rect 3507 5896 3573 5904
rect 3627 5897 3653 5905
rect 3887 5896 3913 5904
rect 4167 5897 4653 5905
rect 2156 5856 2233 5864
rect 2287 5855 2353 5863
rect 2447 5856 2533 5864
rect 3247 5855 3293 5863
rect 3416 5864 3424 5893
rect 3416 5856 3433 5864
rect 3487 5856 3653 5864
rect 3927 5855 3973 5863
rect 4067 5855 4133 5863
rect 4196 5864 4204 5874
rect 4447 5876 4573 5884
rect 4147 5856 4204 5864
rect 847 5836 913 5844
rect 1387 5836 1453 5844
rect 2487 5836 2573 5844
rect 2667 5836 2733 5844
rect 2907 5836 3113 5844
rect 3367 5836 4533 5844
rect 4616 5844 4624 5873
rect 4767 5855 4793 5863
rect 4587 5836 4624 5844
rect 4876 5847 4884 5913
rect 4967 5896 5033 5904
rect 5227 5896 5364 5904
rect 5356 5884 5364 5896
rect 5387 5897 5433 5905
rect 5456 5896 5533 5904
rect 5356 5880 5424 5884
rect 5356 5876 5427 5880
rect 5413 5867 5427 5876
rect 4987 5855 5153 5863
rect 5267 5856 5313 5864
rect 5456 5866 5464 5896
rect 5587 5896 5613 5904
rect 5707 5897 5753 5905
rect 5916 5884 5924 5894
rect 6167 5896 6193 5904
rect 5916 5876 5944 5884
rect 5647 5856 5853 5864
rect 5867 5856 5893 5864
rect 5936 5864 5944 5876
rect 5936 5856 6093 5864
rect 6247 5856 6364 5864
rect 4876 5836 4893 5847
rect 4880 5833 4893 5836
rect 287 5816 433 5824
rect 507 5816 733 5824
rect 1047 5816 1153 5824
rect 1487 5816 1713 5824
rect 1727 5816 1933 5824
rect 1947 5816 2253 5824
rect 2347 5816 2693 5824
rect 3147 5816 3313 5824
rect 3667 5816 4013 5824
rect 4027 5816 4093 5824
rect 4536 5824 4544 5833
rect 4536 5816 5233 5824
rect 5247 5816 5613 5824
rect 5807 5816 5933 5824
rect 167 5796 353 5804
rect 436 5804 444 5813
rect 436 5796 793 5804
rect 2747 5796 3073 5804
rect 3607 5796 3853 5804
rect 4567 5796 4633 5804
rect 4727 5796 4873 5804
rect 5027 5796 5313 5804
rect 5427 5796 5693 5804
rect 307 5776 493 5784
rect 1067 5776 1473 5784
rect 2247 5776 2493 5784
rect 2507 5776 3133 5784
rect 3147 5776 5053 5784
rect 5067 5776 5393 5784
rect 1627 5756 1753 5764
rect 1767 5756 1793 5764
rect 1807 5756 2213 5764
rect 2267 5756 2733 5764
rect 2907 5756 3093 5764
rect 4647 5756 5373 5764
rect 5387 5756 5573 5764
rect 667 5736 1033 5744
rect 2887 5736 3193 5744
rect 3667 5736 4253 5744
rect 4307 5736 4493 5744
rect 5067 5736 5113 5744
rect 407 5716 453 5724
rect 467 5716 613 5724
rect 2467 5716 2853 5724
rect 3367 5716 3413 5724
rect 3556 5716 4584 5724
rect 2227 5696 2953 5704
rect 3556 5704 3564 5716
rect 3107 5696 3564 5704
rect 3707 5696 4093 5704
rect 4576 5704 4584 5716
rect 4607 5716 4853 5724
rect 5247 5716 5493 5724
rect 5507 5716 5833 5724
rect 4576 5696 4793 5704
rect 5027 5696 5153 5704
rect 5167 5696 5904 5704
rect 5896 5687 5904 5696
rect 367 5676 493 5684
rect 507 5676 693 5684
rect 1347 5676 2933 5684
rect 4267 5676 4633 5684
rect 4867 5676 4893 5684
rect 5087 5676 5233 5684
rect 5467 5676 5673 5684
rect 5907 5676 6153 5684
rect 2647 5656 2713 5664
rect 3947 5656 4193 5664
rect 4247 5656 4673 5664
rect 4687 5656 4833 5664
rect 5267 5656 5553 5664
rect 5567 5656 5753 5664
rect 5767 5656 6033 5664
rect 447 5636 593 5644
rect 716 5636 1313 5644
rect 127 5597 193 5605
rect 276 5564 284 5594
rect 527 5597 553 5605
rect 607 5597 653 5605
rect 316 5567 324 5593
rect 480 5584 493 5587
rect 476 5573 493 5584
rect 147 5556 284 5564
rect 476 5564 484 5573
rect 716 5566 724 5636
rect 1447 5636 1813 5644
rect 1887 5636 1973 5644
rect 2147 5636 2233 5644
rect 2987 5636 3253 5644
rect 3867 5636 4633 5644
rect 4936 5636 5193 5644
rect 2667 5616 2893 5624
rect 4936 5624 4944 5636
rect 4807 5616 4944 5624
rect 5567 5616 5613 5624
rect 5987 5616 6033 5624
rect 787 5597 813 5605
rect 1007 5596 1053 5604
rect 736 5584 744 5594
rect 856 5584 864 5594
rect 1287 5596 1393 5604
rect 1567 5596 1633 5604
rect 1767 5597 1813 5605
rect 1887 5596 1924 5604
rect 1916 5584 1924 5596
rect 1967 5596 2133 5604
rect 736 5576 764 5584
rect 856 5576 1204 5584
rect 1916 5576 2024 5584
rect 427 5556 484 5564
rect 756 5564 764 5576
rect 1196 5567 1204 5576
rect 756 5556 833 5564
rect 2016 5566 2024 5576
rect 1207 5556 1373 5564
rect 1427 5555 1633 5563
rect 167 5536 213 5544
rect 307 5536 353 5544
rect 367 5536 573 5544
rect 1907 5536 1973 5544
rect 2176 5544 2184 5594
rect 2307 5596 2364 5604
rect 2193 5584 2207 5593
rect 2356 5584 2364 5596
rect 2387 5597 2413 5605
rect 2507 5596 2544 5604
rect 2536 5584 2544 5596
rect 2587 5596 2884 5604
rect 2193 5580 2224 5584
rect 2196 5576 2224 5580
rect 2356 5576 2524 5584
rect 2536 5576 2584 5584
rect 2216 5564 2224 5576
rect 2216 5556 2312 5564
rect 2347 5556 2373 5564
rect 2516 5564 2524 5576
rect 2516 5556 2553 5564
rect 2576 5564 2584 5576
rect 2876 5584 2884 5596
rect 3047 5597 3193 5605
rect 3407 5597 3433 5605
rect 3547 5596 3572 5604
rect 2647 5576 2864 5584
rect 2876 5576 2904 5584
rect 2856 5566 2864 5576
rect 2896 5566 2904 5576
rect 2916 5567 2924 5594
rect 3607 5596 3653 5604
rect 3807 5596 3893 5604
rect 4087 5596 4133 5604
rect 4267 5596 4353 5604
rect 4576 5587 4584 5613
rect 4667 5597 4753 5605
rect 4947 5597 5113 5605
rect 5827 5596 5933 5604
rect 5947 5597 6013 5605
rect 6207 5596 6364 5604
rect 3987 5576 4233 5584
rect 4627 5576 4913 5584
rect 5587 5576 6093 5584
rect 2576 5556 2733 5564
rect 2916 5556 2933 5567
rect 2920 5553 2933 5556
rect 2987 5555 3013 5563
rect 3107 5555 3153 5563
rect 3207 5556 3513 5564
rect 3627 5556 3773 5564
rect 4747 5556 4993 5564
rect 5187 5556 5253 5564
rect 5687 5555 5733 5563
rect 5787 5555 5812 5563
rect 5847 5555 6053 5563
rect 2176 5536 2253 5544
rect 2487 5536 2513 5544
rect 3187 5536 3273 5544
rect 3927 5536 4033 5544
rect 4047 5536 4153 5544
rect 4167 5536 4613 5544
rect 5027 5536 5053 5544
rect 107 5516 193 5524
rect 467 5516 533 5524
rect 807 5516 873 5524
rect 887 5516 973 5524
rect 1127 5516 1333 5524
rect 1707 5516 1773 5524
rect 1867 5516 1953 5524
rect 2067 5516 2273 5524
rect 2667 5516 2733 5524
rect 3067 5516 3393 5524
rect 3447 5516 3993 5524
rect 4867 5516 5073 5524
rect 5147 5516 5873 5524
rect 267 5496 313 5504
rect 2387 5496 2593 5504
rect 2607 5496 2633 5504
rect 3047 5496 3253 5504
rect 3787 5496 3813 5504
rect 4087 5496 4384 5504
rect 4376 5487 4384 5496
rect 4927 5496 5213 5504
rect 567 5476 653 5484
rect 2167 5476 2273 5484
rect 2367 5476 2973 5484
rect 3027 5476 3073 5484
rect 3287 5476 3533 5484
rect 3587 5476 4193 5484
rect 4376 5476 4393 5487
rect 4380 5473 4393 5476
rect 4507 5476 4533 5484
rect 4547 5476 4753 5484
rect 5327 5476 5913 5484
rect 487 5456 753 5464
rect 2247 5456 2493 5464
rect 2547 5456 3053 5464
rect 3107 5456 3173 5464
rect 3267 5456 3573 5464
rect 4847 5456 4973 5464
rect 4987 5456 5173 5464
rect 5187 5456 5273 5464
rect 5287 5456 5304 5464
rect 127 5436 153 5444
rect 1187 5436 1573 5444
rect 1827 5436 2233 5444
rect 2727 5436 3713 5444
rect 4407 5436 5133 5444
rect 5296 5444 5304 5456
rect 5296 5436 5913 5444
rect 327 5416 373 5424
rect 647 5416 773 5424
rect 787 5416 853 5424
rect 1067 5416 1113 5424
rect 2167 5416 2653 5424
rect 2987 5416 3353 5424
rect 3447 5416 3653 5424
rect 4107 5416 4333 5424
rect 4427 5416 4493 5424
rect 4507 5416 4733 5424
rect 5987 5416 6173 5424
rect 287 5396 593 5404
rect 607 5396 913 5404
rect 927 5396 1193 5404
rect 1207 5396 1233 5404
rect 2247 5396 2633 5404
rect 3087 5396 3224 5404
rect 27 5377 153 5385
rect 167 5376 273 5384
rect 407 5377 513 5385
rect 727 5377 753 5385
rect 987 5377 1073 5385
rect 1287 5376 1324 5384
rect 1316 5364 1324 5376
rect 1347 5377 1373 5385
rect 1427 5376 1533 5384
rect 1647 5377 1673 5385
rect 1867 5376 2093 5384
rect 2187 5377 2213 5385
rect 2267 5376 2373 5384
rect 2387 5377 2413 5385
rect 2636 5376 2693 5384
rect 1316 5356 1384 5364
rect 207 5335 253 5343
rect 387 5335 413 5343
rect 827 5335 853 5343
rect 1027 5336 1093 5344
rect 1147 5335 1173 5343
rect 1307 5336 1333 5344
rect 1376 5344 1384 5356
rect 1436 5356 1524 5364
rect 1436 5346 1444 5356
rect 1376 5336 1433 5344
rect 1516 5344 1524 5356
rect 1516 5336 1593 5344
rect 1707 5336 1793 5344
rect 2127 5336 2173 5344
rect 2287 5335 2313 5343
rect 2636 5344 2644 5376
rect 2787 5376 2873 5384
rect 2567 5336 2644 5344
rect 196 5324 204 5332
rect 2936 5327 2944 5393
rect 2987 5357 3073 5365
rect 3216 5366 3224 5396
rect 3387 5396 3893 5404
rect 4907 5396 5053 5404
rect 5067 5396 5113 5404
rect 3467 5376 3853 5384
rect 3907 5376 3953 5384
rect 4067 5377 4093 5385
rect 4307 5376 4373 5384
rect 4747 5377 4813 5385
rect 3407 5356 3973 5364
rect 3353 5344 3367 5353
rect 3353 5340 3413 5344
rect 3356 5336 3413 5340
rect 3527 5336 3593 5344
rect 3607 5335 3673 5343
rect 3727 5335 3753 5343
rect 3807 5336 3832 5344
rect 3867 5336 3933 5344
rect 4367 5335 4392 5343
rect 4456 5344 4464 5374
rect 4827 5377 4873 5385
rect 6007 5377 6093 5385
rect 4427 5336 4464 5344
rect 4527 5336 4593 5344
rect 5553 5344 5567 5353
rect 5747 5355 5873 5363
rect 5516 5336 5584 5344
rect 107 5316 204 5324
rect 327 5316 353 5324
rect 667 5316 713 5324
rect 727 5316 753 5324
rect 767 5316 1053 5324
rect 2547 5316 2713 5324
rect 3227 5316 3313 5324
rect 3387 5315 3453 5323
rect 4187 5316 4313 5324
rect 4327 5316 4533 5324
rect 4547 5316 4653 5324
rect 4707 5316 4753 5324
rect 5027 5316 5053 5324
rect 5516 5326 5524 5336
rect 5576 5326 5584 5336
rect 6247 5336 6364 5344
rect 787 5296 893 5304
rect 1547 5296 2153 5304
rect 2467 5296 2873 5304
rect 2887 5296 3492 5304
rect 3527 5296 3573 5304
rect 3667 5296 4073 5304
rect 4267 5296 4473 5304
rect 247 5276 293 5284
rect 307 5276 393 5284
rect 567 5276 613 5284
rect 1067 5276 1253 5284
rect 1267 5276 1393 5284
rect 1767 5276 2384 5284
rect 647 5256 733 5264
rect 1687 5256 2353 5264
rect 2376 5264 2384 5276
rect 3067 5276 3373 5284
rect 3496 5284 3504 5293
rect 3496 5276 3873 5284
rect 3887 5276 4653 5284
rect 4667 5276 4913 5284
rect 5467 5276 5493 5284
rect 5967 5276 6113 5284
rect 2376 5256 2793 5264
rect 2927 5256 2953 5264
rect 2967 5256 3473 5264
rect 3547 5256 3613 5264
rect 3987 5256 4412 5264
rect 4447 5256 5113 5264
rect 6147 5256 6173 5264
rect 1707 5236 2004 5244
rect 1996 5224 2004 5236
rect 2527 5236 2813 5244
rect 2947 5236 3613 5244
rect 3887 5236 4224 5244
rect 1996 5216 2944 5224
rect 927 5196 1693 5204
rect 1847 5196 1873 5204
rect 1887 5196 1953 5204
rect 2236 5196 2753 5204
rect 907 5176 1753 5184
rect 2236 5184 2244 5196
rect 2936 5204 2944 5216
rect 3027 5216 3653 5224
rect 4216 5224 4224 5236
rect 4216 5216 4613 5224
rect 4636 5216 4953 5224
rect 2936 5196 3073 5204
rect 3087 5196 3233 5204
rect 3447 5196 3553 5204
rect 4636 5204 4644 5216
rect 5367 5216 5393 5224
rect 3907 5196 4644 5204
rect 4807 5196 4933 5204
rect 4947 5196 5433 5204
rect 5476 5196 6113 5204
rect 2027 5176 2244 5184
rect 2407 5176 2593 5184
rect 2867 5176 3873 5184
rect 4027 5176 4293 5184
rect 4307 5176 4413 5184
rect 4427 5176 4853 5184
rect 5476 5184 5484 5196
rect 4967 5176 5484 5184
rect 5527 5176 5653 5184
rect 647 5156 833 5164
rect 1567 5156 1853 5164
rect 2696 5156 2873 5164
rect 2696 5147 2704 5156
rect 3247 5156 3473 5164
rect 3487 5156 3533 5164
rect 3587 5156 3893 5164
rect 4007 5156 4573 5164
rect 4587 5156 4833 5164
rect 5087 5156 5333 5164
rect 5447 5156 5493 5164
rect 5507 5156 5733 5164
rect 347 5136 893 5144
rect 1307 5136 1353 5144
rect 2307 5136 2373 5144
rect 2387 5136 2693 5144
rect 2827 5136 3213 5144
rect 4347 5136 4693 5144
rect 5196 5136 5313 5144
rect 547 5116 593 5124
rect 707 5116 773 5124
rect 967 5116 1033 5124
rect 1647 5116 1713 5124
rect 1727 5116 1933 5124
rect 2487 5116 2684 5124
rect 456 5096 793 5104
rect 456 5088 464 5096
rect 1287 5096 1433 5104
rect 2676 5104 2684 5116
rect 3427 5116 3553 5124
rect 3567 5116 3593 5124
rect 3987 5116 4033 5124
rect 4127 5124 4140 5127
rect 4127 5113 4144 5124
rect 5196 5124 5204 5136
rect 5427 5136 5913 5144
rect 4787 5116 5204 5124
rect 5247 5116 5293 5124
rect 5387 5116 5793 5124
rect 5947 5116 6173 5124
rect 2676 5096 2773 5104
rect 3067 5096 3113 5104
rect 3227 5096 4053 5104
rect 47 5077 93 5085
rect 347 5077 373 5085
rect 427 5077 453 5085
rect 567 5076 653 5084
rect 136 5047 144 5074
rect 67 5035 113 5043
rect 136 5036 153 5047
rect 140 5033 153 5036
rect 376 5024 384 5074
rect 516 5044 524 5074
rect 407 5036 524 5044
rect 556 5047 564 5074
rect 807 5076 993 5084
rect 1207 5077 1273 5085
rect 1327 5077 1373 5085
rect 1487 5077 1513 5085
rect 1527 5076 1573 5084
rect 1627 5076 1693 5084
rect 1707 5077 1733 5085
rect 1987 5077 2032 5085
rect 556 5036 573 5047
rect 560 5033 573 5036
rect 736 5044 744 5073
rect 727 5036 744 5044
rect 776 5040 813 5044
rect 773 5036 813 5040
rect 773 5027 787 5036
rect 867 5036 933 5044
rect 1116 5044 1124 5074
rect 987 5036 1124 5044
rect 1156 5047 1164 5074
rect 2147 5077 2173 5085
rect 2487 5076 2553 5084
rect 2053 5064 2067 5073
rect 2016 5060 2067 5064
rect 2256 5064 2264 5074
rect 2607 5076 2653 5084
rect 2776 5076 2833 5084
rect 2016 5056 2064 5060
rect 2256 5056 2444 5064
rect 1156 5036 1173 5047
rect 1160 5033 1173 5036
rect 1227 5035 1253 5043
rect 1387 5036 1413 5044
rect 1607 5036 1713 5044
rect 1867 5036 1913 5044
rect 376 5016 513 5024
rect 567 5016 593 5024
rect 1047 5016 1093 5024
rect 1107 5016 1133 5024
rect 1836 5024 1844 5032
rect 2016 5027 2024 5056
rect 2047 5036 2073 5044
rect 2187 5036 2233 5044
rect 2347 5035 2393 5043
rect 2436 5044 2444 5056
rect 2436 5036 2493 5044
rect 2776 5044 2784 5076
rect 2926 5073 2927 5080
rect 2947 5077 2973 5085
rect 3367 5076 3484 5084
rect 2913 5064 2927 5073
rect 2913 5060 3093 5064
rect 2915 5056 3093 5060
rect 3116 5056 3213 5064
rect 2727 5036 2784 5044
rect 2807 5036 2953 5044
rect 1636 5016 1844 5024
rect 1636 5007 1644 5016
rect 2007 5016 2024 5027
rect 2007 5013 2020 5016
rect 2547 5016 2633 5024
rect 3116 5024 3124 5056
rect 3476 5064 3484 5076
rect 3536 5067 3544 5096
rect 3896 5080 3993 5084
rect 3893 5076 3993 5080
rect 3476 5056 3524 5064
rect 3516 5044 3524 5056
rect 3893 5067 3907 5076
rect 3516 5036 3593 5044
rect 2867 5016 3124 5024
rect 3427 5016 3453 5024
rect 3756 5024 3764 5054
rect 4116 5044 4124 5074
rect 4136 5046 4144 5113
rect 4167 5096 4273 5104
rect 4367 5096 4453 5104
rect 4567 5096 4593 5104
rect 5400 5104 5413 5107
rect 5396 5093 5413 5104
rect 4276 5076 4293 5084
rect 4276 5064 4284 5076
rect 4547 5076 4833 5084
rect 4196 5060 4284 5064
rect 4193 5056 4284 5060
rect 4836 5064 4844 5074
rect 4887 5076 4993 5084
rect 5007 5076 5213 5084
rect 5267 5077 5293 5085
rect 5396 5084 5404 5093
rect 5307 5076 5404 5084
rect 5447 5077 5473 5085
rect 5607 5077 5633 5085
rect 6067 5077 6233 5085
rect 4836 5056 5124 5064
rect 4193 5047 4207 5056
rect 4067 5036 4124 5044
rect 4287 5036 4353 5044
rect 4916 5046 4924 5056
rect 4967 5035 4993 5043
rect 5047 5035 5093 5043
rect 5116 5044 5124 5056
rect 5516 5047 5524 5073
rect 5116 5036 5193 5044
rect 5327 5035 5413 5043
rect 3587 5016 3764 5024
rect 4027 5016 4093 5024
rect 4427 5016 4773 5024
rect 4996 5024 5004 5032
rect 4996 5016 5253 5024
rect 5447 5016 5473 5024
rect 5556 5024 5564 5074
rect 5696 5047 5704 5074
rect 5687 5036 5704 5047
rect 5687 5033 5700 5036
rect 5836 5027 5844 5074
rect 6147 5036 6193 5044
rect 5556 5016 5593 5024
rect 5747 5016 5824 5024
rect 47 4996 113 5004
rect 367 4996 604 5004
rect 387 4976 573 4984
rect 596 4984 604 4996
rect 1467 4996 1633 5004
rect 1807 4996 1873 5004
rect 1987 4996 2153 5004
rect 3416 5004 3424 5013
rect 2967 4996 3424 5004
rect 4147 4996 4233 5004
rect 4447 4996 4473 5004
rect 4667 4996 4813 5004
rect 4947 4996 5293 5004
rect 5387 4996 5513 5004
rect 5647 4996 5713 5004
rect 5816 5004 5824 5016
rect 5927 5016 5973 5024
rect 5816 4996 5893 5004
rect 6047 4996 6113 5004
rect 6187 4996 6233 5004
rect 596 4976 1233 4984
rect 1307 4976 1513 4984
rect 2327 4976 2713 4984
rect 2787 4976 2873 4984
rect 3087 4976 3433 4984
rect 3607 4976 3853 4984
rect 3987 4976 5753 4984
rect 216 4956 253 4964
rect 216 4944 224 4956
rect 507 4956 613 4964
rect 807 4956 1073 4964
rect 1207 4956 1273 4964
rect 1647 4956 1833 4964
rect 1907 4956 2113 4964
rect 2167 4956 2973 4964
rect 3227 4956 3353 4964
rect 3487 4956 3833 4964
rect 4007 4956 4073 4964
rect 4167 4956 4413 4964
rect 4627 4956 5573 4964
rect 5667 4956 5733 4964
rect 5787 4956 6253 4964
rect 47 4936 224 4944
rect 747 4936 873 4944
rect 1407 4936 1533 4944
rect 2147 4936 2453 4944
rect 2996 4936 3113 4944
rect 1787 4916 1953 4924
rect 2067 4916 2113 4924
rect 2267 4916 2293 4924
rect 2367 4916 2413 4924
rect 2427 4916 2493 4924
rect 2607 4916 2693 4924
rect 2996 4924 3004 4936
rect 3367 4936 3593 4944
rect 3727 4936 4113 4944
rect 4207 4936 4233 4944
rect 4247 4936 4333 4944
rect 4727 4936 5153 4944
rect 5487 4936 5533 4944
rect 2907 4916 3004 4924
rect 3127 4916 3693 4924
rect 4393 4924 4407 4933
rect 4216 4920 4407 4924
rect 4216 4916 4404 4920
rect 4216 4907 4224 4916
rect 4927 4916 5073 4924
rect 5247 4916 5373 4924
rect 5387 4916 5573 4924
rect 5587 4916 5673 4924
rect 5967 4916 6133 4924
rect 247 4896 433 4904
rect 447 4896 793 4904
rect 847 4896 893 4904
rect 1167 4896 1373 4904
rect 1507 4896 1593 4904
rect 1887 4896 2013 4904
rect 2207 4896 2273 4904
rect 2547 4896 2853 4904
rect 3547 4896 3673 4904
rect 3956 4896 4213 4904
rect 3956 4887 3964 4896
rect 4767 4896 4893 4904
rect 5427 4896 5513 4904
rect 5767 4896 5873 4904
rect 307 4876 424 4884
rect 167 4857 213 4865
rect 227 4856 393 4864
rect 416 4864 424 4876
rect 1427 4876 1473 4884
rect 1867 4876 1893 4884
rect 1907 4876 2133 4884
rect 2216 4876 2353 4884
rect 416 4856 464 4864
rect 456 4844 464 4856
rect 487 4857 513 4865
rect 607 4856 713 4864
rect 767 4856 793 4864
rect 847 4857 873 4865
rect 947 4857 1193 4865
rect 456 4836 504 4844
rect 227 4816 253 4824
rect 496 4824 504 4836
rect 496 4816 533 4824
rect 687 4816 733 4824
rect 747 4816 853 4824
rect 927 4815 953 4823
rect 1316 4824 1324 4854
rect 1547 4857 1633 4865
rect 1967 4856 2093 4864
rect 1356 4827 1364 4853
rect 1873 4844 1887 4853
rect 2216 4844 2224 4876
rect 2507 4876 2813 4884
rect 2827 4876 2933 4884
rect 2947 4876 3113 4884
rect 3500 4884 3513 4887
rect 3496 4873 3513 4884
rect 3707 4876 3953 4884
rect 4127 4876 4564 4884
rect 2287 4864 2300 4867
rect 2287 4853 2304 4864
rect 1847 4840 1887 4844
rect 2016 4840 2224 4844
rect 1847 4836 1884 4840
rect 2013 4836 2224 4840
rect 2013 4827 2027 4836
rect 1187 4816 1324 4824
rect 1527 4815 1573 4823
rect 2216 4826 2224 4836
rect 2296 4826 2304 4853
rect 2487 4856 2552 4864
rect 2413 4844 2427 4853
rect 2573 4844 2587 4853
rect 2413 4840 2464 4844
rect 2416 4836 2464 4840
rect 2456 4826 2464 4836
rect 2496 4840 2587 4844
rect 2656 4856 2773 4864
rect 2496 4836 2584 4840
rect 2496 4826 2504 4836
rect 2656 4826 2664 4856
rect 2927 4856 3213 4864
rect 3496 4864 3504 4873
rect 3396 4856 3504 4864
rect 3516 4856 3552 4864
rect 2147 4816 2173 4824
rect 3007 4815 3053 4823
rect 3267 4816 3333 4824
rect 3396 4824 3404 4856
rect 3516 4826 3524 4856
rect 3587 4856 3613 4864
rect 3667 4856 3733 4864
rect 3787 4857 3853 4865
rect 3987 4857 4053 4865
rect 4556 4864 4564 4876
rect 4987 4876 5033 4884
rect 5507 4884 5520 4887
rect 5507 4873 5524 4884
rect 5687 4876 5773 4884
rect 4556 4856 4813 4864
rect 4836 4856 4853 4864
rect 3387 4816 3404 4824
rect 3447 4815 3473 4823
rect 3607 4815 3633 4823
rect 3687 4816 3753 4824
rect 3767 4816 3813 4824
rect 4136 4824 4144 4834
rect 4407 4836 4473 4844
rect 4836 4844 4844 4856
rect 5067 4856 5113 4864
rect 5187 4857 5253 4865
rect 5347 4856 5413 4864
rect 4696 4836 4844 4844
rect 4136 4816 4373 4824
rect 4696 4826 4704 4836
rect 5476 4827 5484 4873
rect 4767 4815 4793 4823
rect 4887 4816 4993 4824
rect 5247 4816 5264 4824
rect 67 4796 133 4804
rect 947 4796 993 4804
rect 2567 4796 2612 4804
rect 2647 4796 2792 4804
rect 2827 4796 2873 4804
rect 3107 4796 3233 4804
rect 4596 4796 4653 4804
rect 107 4776 233 4784
rect 447 4776 473 4784
rect 487 4776 693 4784
rect 707 4776 773 4784
rect 787 4776 893 4784
rect 996 4784 1004 4793
rect 996 4776 1333 4784
rect 1587 4776 1973 4784
rect 2207 4776 2253 4784
rect 2680 4784 2692 4787
rect 2676 4773 2692 4784
rect 4596 4784 4604 4796
rect 5147 4796 5213 4804
rect 5256 4804 5264 4816
rect 5516 4826 5524 4873
rect 5560 4864 5573 4867
rect 5556 4853 5573 4864
rect 5627 4856 5713 4864
rect 5796 4856 5953 4864
rect 5556 4826 5564 4853
rect 5796 4844 5804 4856
rect 5976 4856 5993 4864
rect 5976 4844 5984 4856
rect 6207 4857 6293 4865
rect 5736 4840 5804 4844
rect 5733 4836 5804 4840
rect 5816 4836 5984 4844
rect 5733 4827 5747 4836
rect 5816 4824 5824 4836
rect 5756 4816 5824 4824
rect 5256 4796 5353 4804
rect 5756 4804 5764 4816
rect 6027 4816 6053 4824
rect 5707 4796 5764 4804
rect 5947 4796 6013 4804
rect 2727 4776 4604 4784
rect 5407 4776 5653 4784
rect 5767 4776 6033 4784
rect 6076 4784 6084 4853
rect 6127 4816 6233 4824
rect 6287 4815 6313 4823
rect 6076 4776 6133 4784
rect 27 4756 413 4764
rect 527 4756 573 4764
rect 1107 4756 1153 4764
rect 1267 4756 1512 4764
rect 1547 4756 2093 4764
rect 2207 4756 2333 4764
rect 2676 4764 2684 4773
rect 2627 4756 2684 4764
rect 2747 4756 3533 4764
rect 3627 4756 3733 4764
rect 3927 4756 4553 4764
rect 4647 4756 4933 4764
rect 4947 4756 5053 4764
rect 5487 4756 5813 4764
rect 487 4736 753 4744
rect 1227 4736 1553 4744
rect 1687 4736 1733 4744
rect 1927 4736 2113 4744
rect 2467 4736 2533 4744
rect 2887 4736 3312 4744
rect 3347 4736 3413 4744
rect 3587 4736 3793 4744
rect 4247 4736 4473 4744
rect 4607 4736 5453 4744
rect 5507 4736 5593 4744
rect 67 4716 353 4724
rect 587 4716 653 4724
rect 907 4716 1193 4724
rect 1347 4716 2673 4724
rect 2807 4716 2833 4724
rect 2967 4716 3053 4724
rect 3207 4716 3973 4724
rect 5187 4716 5233 4724
rect 747 4696 833 4704
rect 1247 4696 1573 4704
rect 2707 4696 2833 4704
rect 2847 4696 2953 4704
rect 2967 4696 3253 4704
rect 3667 4696 3873 4704
rect 4107 4696 4233 4704
rect 4247 4696 4533 4704
rect 5347 4696 5473 4704
rect 5667 4696 5853 4704
rect 6067 4696 6193 4704
rect 507 4676 693 4684
rect 807 4676 973 4684
rect 1187 4676 1853 4684
rect 1867 4676 1933 4684
rect 1947 4676 2033 4684
rect 2107 4676 2673 4684
rect 2867 4676 2913 4684
rect 2987 4676 3493 4684
rect 3547 4676 3873 4684
rect 4767 4676 4833 4684
rect 5967 4676 6173 4684
rect 27 4656 313 4664
rect 327 4656 1013 4664
rect 1027 4656 1053 4664
rect 1207 4656 1253 4664
rect 1327 4656 1753 4664
rect 2956 4656 3993 4664
rect 627 4636 873 4644
rect 927 4636 953 4644
rect 967 4636 993 4644
rect 1007 4636 1253 4644
rect 2407 4636 2493 4644
rect 2956 4644 2964 4656
rect 5147 4656 5213 4664
rect 5227 4656 5333 4664
rect 2507 4636 2964 4644
rect 3527 4636 3913 4644
rect 4067 4636 4173 4644
rect 4387 4636 4653 4644
rect 87 4616 533 4624
rect 767 4616 1053 4624
rect 1067 4616 1213 4624
rect 1327 4616 1533 4624
rect 1547 4616 1613 4624
rect 2567 4616 2733 4624
rect 2807 4616 2833 4624
rect 5187 4616 5293 4624
rect 5867 4616 6053 4624
rect 107 4596 153 4604
rect 227 4596 293 4604
rect 307 4596 473 4604
rect 867 4596 1193 4604
rect 1207 4596 1273 4604
rect 1396 4596 1453 4604
rect 647 4576 793 4584
rect 987 4576 1033 4584
rect 1396 4584 1404 4596
rect 1647 4596 1773 4604
rect 1967 4596 2053 4604
rect 2687 4596 2853 4604
rect 2927 4596 3513 4604
rect 3567 4596 3813 4604
rect 3827 4596 3893 4604
rect 4967 4596 5133 4604
rect 5567 4596 5633 4604
rect 1376 4576 1404 4584
rect 1376 4568 1384 4576
rect 2047 4576 2224 4584
rect -24 4556 73 4564
rect 556 4527 564 4554
rect 840 4564 853 4567
rect 836 4553 853 4564
rect 907 4556 933 4564
rect 1107 4557 1133 4565
rect 1427 4557 1453 4565
rect 1627 4557 1673 4565
rect 127 4516 153 4524
rect 167 4516 193 4524
rect 247 4516 333 4524
rect 347 4516 433 4524
rect 556 4516 573 4527
rect 560 4513 573 4516
rect 696 4524 704 4553
rect 836 4526 844 4553
rect 1056 4527 1064 4553
rect 667 4516 704 4524
rect 1336 4524 1344 4554
rect 1516 4544 1524 4554
rect 1767 4556 1833 4564
rect 2216 4564 2224 4576
rect 2896 4576 3033 4584
rect 2216 4556 2393 4564
rect 1516 4536 1564 4544
rect 1127 4516 1344 4524
rect 1487 4516 1533 4524
rect 47 4496 73 4504
rect 1147 4496 1193 4504
rect 1556 4504 1564 4536
rect 1887 4536 2193 4544
rect 1807 4515 1853 4523
rect 2047 4515 2073 4523
rect 2127 4516 2673 4524
rect 2736 4524 2744 4554
rect 2896 4564 2904 4576
rect 4107 4576 4173 4584
rect 4547 4576 4593 4584
rect 5087 4576 5173 4584
rect 5927 4576 6013 4584
rect 2787 4556 2904 4564
rect 2916 4560 3053 4564
rect 2913 4556 3053 4560
rect 2913 4547 2927 4556
rect 3347 4556 3433 4564
rect 3607 4556 3693 4564
rect 3947 4557 3972 4565
rect 4007 4556 4373 4564
rect 5316 4556 5413 4564
rect 3356 4536 3413 4544
rect 2736 4516 2833 4524
rect 3356 4524 3364 4536
rect 3936 4536 4553 4544
rect 2947 4516 3364 4524
rect 3407 4516 3773 4524
rect 3887 4515 3913 4523
rect 1556 4496 1633 4504
rect 1687 4496 1733 4504
rect 1827 4496 1873 4504
rect 3247 4496 3413 4504
rect 3427 4496 3593 4504
rect 3936 4504 3944 4536
rect 5007 4535 5033 4543
rect 3987 4516 4033 4524
rect 5096 4524 5104 4553
rect 5316 4526 5324 4556
rect 5707 4556 5724 4564
rect 5096 4516 5113 4524
rect 5167 4515 5193 4523
rect 5447 4516 5453 4524
rect 5467 4516 5573 4524
rect 5596 4524 5604 4554
rect 5716 4544 5724 4556
rect 5787 4557 5813 4565
rect 5987 4556 6093 4564
rect 6187 4556 6213 4564
rect 6227 4557 6253 4565
rect 5716 4536 5933 4544
rect 5596 4516 5713 4524
rect 3807 4496 3944 4504
rect 4207 4496 4473 4504
rect 4487 4496 4933 4504
rect 5247 4496 5273 4504
rect 5667 4496 5693 4504
rect 5976 4504 5984 4554
rect 6296 4544 6304 4554
rect 6256 4536 6304 4544
rect 6007 4516 6053 4524
rect 6256 4524 6264 4536
rect 6167 4516 6264 4524
rect 6316 4524 6324 4553
rect 6287 4516 6324 4524
rect 5887 4496 5984 4504
rect 387 4476 613 4484
rect 887 4476 1073 4484
rect 1467 4476 1653 4484
rect 1727 4476 2093 4484
rect 2527 4476 2593 4484
rect 2727 4476 2773 4484
rect 3156 4476 3393 4484
rect 407 4456 633 4464
rect 656 4456 964 4464
rect 567 4436 593 4444
rect 656 4444 664 4456
rect 956 4447 964 4456
rect 1187 4456 1393 4464
rect 1547 4456 1593 4464
rect 1887 4456 1993 4464
rect 2147 4460 2484 4464
rect 2147 4456 2487 4460
rect 2473 4447 2487 4456
rect 2647 4456 2833 4464
rect 3156 4464 3164 4476
rect 4007 4476 4072 4484
rect 4107 4476 4473 4484
rect 4607 4476 4653 4484
rect 5387 4476 5413 4484
rect 5787 4476 5853 4484
rect 5927 4476 6033 4484
rect 6047 4476 6113 4484
rect 6227 4476 6273 4484
rect 2887 4456 3164 4464
rect 3247 4456 3353 4464
rect 607 4436 664 4444
rect 967 4436 1093 4444
rect 1367 4436 1793 4444
rect 1987 4436 2153 4444
rect 2267 4436 2293 4444
rect 2536 4436 3093 4444
rect 147 4416 284 4424
rect 276 4407 284 4416
rect 347 4416 493 4424
rect 547 4416 733 4424
rect 1207 4416 1713 4424
rect 2227 4416 2433 4424
rect 287 4396 593 4404
rect 1007 4396 1104 4404
rect 1096 4387 1104 4396
rect 1147 4396 1733 4404
rect 2536 4404 2544 4436
rect 3787 4436 4093 4444
rect 4147 4436 4273 4444
rect 4567 4436 4713 4444
rect 4807 4436 4893 4444
rect 5207 4436 5313 4444
rect 5367 4436 5473 4444
rect 5627 4436 5933 4444
rect 1747 4396 2544 4404
rect 2807 4416 2853 4424
rect 3407 4416 3633 4424
rect 3767 4416 4013 4424
rect 4187 4416 4353 4424
rect 4527 4416 5013 4424
rect 5087 4416 6173 4424
rect 2613 4404 2627 4413
rect 2613 4400 2733 4404
rect 2616 4396 2733 4400
rect 3167 4396 3333 4404
rect 3467 4396 3573 4404
rect 427 4376 453 4384
rect 587 4376 813 4384
rect 1096 4376 1113 4387
rect 1100 4373 1113 4376
rect 1227 4376 1253 4384
rect 1767 4376 1793 4384
rect 1927 4376 1993 4384
rect 2947 4376 2993 4384
rect 3387 4376 3533 4384
rect 4167 4376 4233 4384
rect 4447 4376 4493 4384
rect 4647 4376 4733 4384
rect 5167 4376 5673 4384
rect 5727 4376 5793 4384
rect 5807 4376 5833 4384
rect 496 4356 853 4364
rect -24 4336 13 4344
rect 27 4336 93 4344
rect 496 4306 504 4356
rect 947 4356 993 4364
rect 1256 4356 1473 4364
rect 1087 4336 1233 4344
rect 596 4307 604 4333
rect 1256 4327 1264 4356
rect 2027 4356 2093 4364
rect 2107 4356 2133 4364
rect 2927 4356 3013 4364
rect 3087 4356 3193 4364
rect 3287 4356 3333 4364
rect 3627 4356 4093 4364
rect 4307 4356 4513 4364
rect 5227 4356 5273 4364
rect 696 4316 913 4324
rect 647 4295 673 4303
rect 696 4284 704 4316
rect 1240 4326 1264 4327
rect 1247 4316 1264 4326
rect 1367 4336 1593 4344
rect 2960 4344 2973 4347
rect 1273 4324 1287 4333
rect 1273 4320 1364 4324
rect 1276 4316 1364 4320
rect 1247 4313 1260 4316
rect 787 4295 833 4303
rect 887 4295 953 4303
rect 1167 4296 1333 4304
rect 1356 4304 1364 4316
rect 1356 4296 1433 4304
rect 1547 4295 1573 4303
rect 307 4276 704 4284
rect 1267 4276 1293 4284
rect 1636 4284 1644 4334
rect 1916 4324 1924 4334
rect 2036 4324 2044 4334
rect 2156 4324 2164 4334
rect 2956 4333 2973 4344
rect 3227 4336 3373 4344
rect 4116 4336 4213 4344
rect 1916 4316 2044 4324
rect 2076 4320 2164 4324
rect 2196 4320 2393 4324
rect 2073 4316 2164 4320
rect 2193 4316 2393 4320
rect 1667 4296 1693 4304
rect 1916 4304 1924 4316
rect 2073 4307 2087 4316
rect 1916 4296 1953 4304
rect 2027 4295 2052 4303
rect 2193 4307 2207 4316
rect 2767 4316 2783 4324
rect 2476 4287 2484 4313
rect 2775 4287 2783 4316
rect 2956 4306 2964 4333
rect 3107 4316 3324 4324
rect 3176 4306 3184 4316
rect 3316 4306 3324 4316
rect 3416 4307 3424 4333
rect 3496 4307 3504 4334
rect 3496 4296 3513 4307
rect 3500 4293 3513 4296
rect 1467 4276 1753 4284
rect 1867 4276 1893 4284
rect 2807 4275 2933 4283
rect 2947 4275 3033 4283
rect 3207 4276 3253 4284
rect 3536 4284 3544 4314
rect 3807 4316 3913 4324
rect 3615 4287 3623 4313
rect 4116 4306 4124 4336
rect 4547 4336 4573 4344
rect 4587 4336 4633 4344
rect 4687 4336 4784 4344
rect 4776 4306 4784 4336
rect 5436 4336 5753 4344
rect 4027 4295 4073 4303
rect 4527 4296 4613 4304
rect 5267 4296 5353 4304
rect 5436 4306 5444 4336
rect 5776 4336 5973 4344
rect 5776 4306 5784 4336
rect 5987 4336 6073 4344
rect 6216 4304 6224 4334
rect 6107 4296 6224 4304
rect 3467 4276 3544 4284
rect 3647 4276 3933 4284
rect 3947 4275 4153 4283
rect 4227 4276 4393 4284
rect 5727 4276 5793 4284
rect 207 4256 432 4264
rect 467 4256 853 4264
rect 1007 4256 1472 4264
rect 1507 4256 1613 4264
rect 1627 4256 1713 4264
rect 1927 4256 2133 4264
rect 2147 4256 2233 4264
rect 3287 4256 3433 4264
rect 4087 4256 4193 4264
rect 4467 4256 4573 4264
rect 4587 4256 4813 4264
rect 5427 4256 5533 4264
rect 6147 4256 6233 4264
rect 487 4236 1033 4244
rect 1107 4236 1304 4244
rect 147 4216 393 4224
rect 547 4216 713 4224
rect 787 4216 933 4224
rect 947 4216 1113 4224
rect 1296 4224 1304 4236
rect 1447 4236 1773 4244
rect 1947 4236 2073 4244
rect 2207 4236 2393 4244
rect 2927 4236 3053 4244
rect 3587 4236 3773 4244
rect 3793 4244 3807 4253
rect 3793 4240 3973 4244
rect 3796 4236 3973 4240
rect 4067 4236 4273 4244
rect 4287 4236 4333 4244
rect 5007 4236 5073 4244
rect 5507 4236 5553 4244
rect 5727 4236 5813 4244
rect 5827 4236 5853 4244
rect 1296 4216 1873 4224
rect 2827 4216 3244 4224
rect 347 4196 493 4204
rect 1467 4196 2264 4204
rect 147 4176 313 4184
rect 327 4176 373 4184
rect 547 4176 613 4184
rect 847 4176 1333 4184
rect 1347 4176 1373 4184
rect 1487 4176 1813 4184
rect 1887 4176 2193 4184
rect 2256 4184 2264 4196
rect 2387 4196 2433 4204
rect 2447 4196 3033 4204
rect 3236 4204 3244 4216
rect 3307 4216 3913 4224
rect 4047 4216 4073 4224
rect 4167 4216 4293 4224
rect 3236 4196 3953 4204
rect 3967 4196 4273 4204
rect 4647 4196 4873 4204
rect 5827 4196 5913 4204
rect 5927 4196 6053 4204
rect 2256 4176 2913 4184
rect 4247 4176 4353 4184
rect 4787 4176 5213 4184
rect 827 4156 913 4164
rect 1067 4156 1253 4164
rect 1380 4164 1393 4167
rect 1376 4153 1393 4164
rect 2067 4156 2093 4164
rect 2687 4156 2733 4164
rect 2807 4156 3353 4164
rect 3367 4156 3473 4164
rect 3487 4156 4373 4164
rect 4473 4164 4487 4173
rect 4447 4160 4487 4164
rect 4447 4156 4484 4160
rect 4727 4156 4873 4164
rect 5067 4156 5204 4164
rect 507 4136 1233 4144
rect 1376 4144 1384 4153
rect 1247 4136 1384 4144
rect 1427 4136 1553 4144
rect 1847 4136 1873 4144
rect 2787 4136 2853 4144
rect 2927 4136 2993 4144
rect 3047 4136 3153 4144
rect 3627 4136 3653 4144
rect 5196 4144 5204 4156
rect 5196 4136 5393 4144
rect 5407 4136 5913 4144
rect 227 4116 412 4124
rect 447 4116 713 4124
rect 727 4116 813 4124
rect 996 4116 1393 4124
rect 996 4104 1004 4116
rect 1987 4116 2093 4124
rect 2267 4116 2493 4124
rect 2907 4116 3013 4124
rect 3767 4116 3993 4124
rect 916 4096 1004 4104
rect 407 4076 473 4084
rect 487 4076 633 4084
rect 67 4037 93 4045
rect 156 4004 164 4033
rect 127 3996 164 4004
rect 176 4004 184 4073
rect 567 4056 773 4064
rect 456 4036 533 4044
rect 256 4024 264 4033
rect 256 4016 313 4024
rect 456 4007 464 4036
rect 553 4044 567 4053
rect 553 4040 593 4044
rect 556 4036 593 4040
rect 807 4036 893 4044
rect 176 3996 233 4004
rect 676 3987 684 4034
rect 916 4006 924 4096
rect 2167 4096 2233 4104
rect 2247 4096 2313 4104
rect 2847 4096 4033 4104
rect 5107 4096 5453 4104
rect 5467 4096 5633 4104
rect 987 4076 1013 4084
rect 1487 4076 1513 4084
rect 1747 4076 2173 4084
rect 2187 4076 2353 4084
rect 2407 4076 2993 4084
rect 3427 4076 3513 4084
rect 3887 4076 3973 4084
rect 3987 4076 4213 4084
rect 4316 4076 4513 4084
rect 1147 4056 1193 4064
rect 1387 4056 1573 4064
rect 1587 4056 1613 4064
rect 2127 4056 2452 4064
rect 2487 4056 2593 4064
rect 3020 4064 3033 4067
rect 956 4036 1013 4044
rect 956 4006 964 4036
rect 1127 4037 1153 4045
rect 1287 4037 1373 4045
rect 1447 4037 1473 4045
rect 1076 4024 1084 4034
rect 1076 4020 1144 4024
rect 1076 4016 1147 4020
rect 1133 4007 1147 4016
rect 1067 3996 1112 4004
rect 1187 3996 1273 4004
rect 1367 3996 1433 4004
rect 1547 3995 1573 4003
rect 1676 3987 1684 4053
rect 1707 4037 1733 4045
rect 1776 4036 1793 4044
rect 1776 4007 1784 4036
rect 1947 4036 1984 4044
rect 1976 4024 1984 4036
rect 2327 4036 2413 4044
rect 2467 4036 2553 4044
rect 2276 4024 2284 4034
rect 2707 4036 2873 4044
rect 2893 4044 2907 4053
rect 3016 4053 3033 4064
rect 3367 4057 3393 4065
rect 3827 4057 3933 4065
rect 4007 4056 4113 4064
rect 4316 4064 4324 4076
rect 5067 4076 5173 4084
rect 4127 4056 4324 4064
rect 4687 4056 4773 4064
rect 2887 4040 2907 4044
rect 2887 4036 2904 4040
rect 1976 4016 2084 4024
rect 1887 3996 1953 4004
rect 2076 4004 2084 4016
rect 2176 4016 2284 4024
rect 2933 4024 2947 4033
rect 2933 4020 2973 4024
rect 2936 4016 2973 4020
rect 2176 4006 2184 4016
rect 3016 4026 3024 4053
rect 3496 4027 3504 4053
rect 4196 4036 4273 4044
rect 2076 3996 2104 4004
rect 567 3976 613 3984
rect 767 3976 853 3984
rect 867 3976 1313 3984
rect 1676 3976 1693 3987
rect 1680 3973 1693 3976
rect 1767 3976 1833 3984
rect 1927 3976 1993 3984
rect 2096 3984 2104 3996
rect 2627 3996 2673 4004
rect 2727 3996 2813 4004
rect 3196 4004 3204 4014
rect 3227 4016 3433 4024
rect 3787 4016 3893 4024
rect 4013 4024 4027 4033
rect 3956 4020 4027 4024
rect 3956 4016 4024 4020
rect 3047 3996 3204 4004
rect 3487 3996 3513 4004
rect 3807 3996 3873 4004
rect 3956 4004 3964 4016
rect 3927 3996 3964 4004
rect 4156 4004 4164 4033
rect 4196 4007 4204 4036
rect 4347 4037 4393 4045
rect 4507 4036 4553 4044
rect 4727 4036 4833 4044
rect 4947 4036 5133 4044
rect 5507 4037 5533 4045
rect 5887 4037 5973 4045
rect 6027 4037 6093 4045
rect 4596 4024 4604 4034
rect 4596 4016 4664 4024
rect 3987 3996 4164 4004
rect 4267 3996 4333 4004
rect 4587 3996 4633 4004
rect 4656 4004 4664 4016
rect 4656 3996 4693 4004
rect 4827 3996 4993 4004
rect 5107 3996 5153 4004
rect 2096 3976 2153 3984
rect 2227 3976 2313 3984
rect 2327 3976 2373 3984
rect 2527 3976 2593 3984
rect 4067 3976 4113 3984
rect 4247 3976 4473 3984
rect 5296 3984 5304 4034
rect 5596 4007 5604 4034
rect 5800 4024 5813 4027
rect 5367 3996 5413 4004
rect 5587 3996 5604 4007
rect 5796 4013 5813 4024
rect 5587 3993 5600 3996
rect 5796 4004 5804 4013
rect 5667 3996 5804 4004
rect 5947 3995 6073 4003
rect 5247 3976 5304 3984
rect 5507 3976 5533 3984
rect 5547 3976 5613 3984
rect 5787 3976 6013 3984
rect 287 3956 313 3964
rect 707 3956 773 3964
rect 787 3956 833 3964
rect 1067 3956 1093 3964
rect 1227 3956 1293 3964
rect 1347 3956 1393 3964
rect 1467 3956 1633 3964
rect 2307 3956 2653 3964
rect 2776 3956 2853 3964
rect 87 3936 153 3944
rect 167 3936 264 3944
rect 256 3924 264 3936
rect 307 3936 413 3944
rect 1687 3936 1733 3944
rect 1907 3936 2113 3944
rect 2167 3936 2333 3944
rect 2776 3944 2784 3956
rect 3947 3956 4013 3964
rect 4187 3956 4353 3964
rect 4427 3956 4493 3964
rect 4507 3956 4653 3964
rect 4847 3956 4913 3964
rect 5047 3956 5313 3964
rect 5327 3956 5433 3964
rect 5773 3964 5787 3973
rect 5667 3960 5787 3964
rect 5667 3956 5784 3960
rect 2347 3936 2784 3944
rect 2907 3936 3033 3944
rect 3856 3936 3913 3944
rect 256 3916 373 3924
rect 527 3916 713 3924
rect 736 3916 1013 3924
rect 447 3896 592 3904
rect 736 3904 744 3916
rect 1227 3916 1413 3924
rect 2107 3916 2333 3924
rect 2807 3916 2853 3924
rect 3067 3916 3113 3924
rect 3187 3916 3293 3924
rect 3507 3916 3633 3924
rect 3856 3924 3864 3936
rect 4016 3944 4024 3953
rect 4016 3936 4213 3944
rect 4727 3936 4813 3944
rect 5727 3936 5773 3944
rect 3747 3916 3864 3924
rect 4007 3916 4093 3924
rect 4887 3916 5673 3924
rect 5767 3916 5953 3924
rect 627 3896 744 3904
rect 1047 3896 1573 3904
rect 1747 3896 1853 3904
rect 2447 3896 2673 3904
rect 2967 3904 2980 3907
rect 2967 3893 2984 3904
rect 587 3876 653 3884
rect 667 3876 773 3884
rect 787 3876 1013 3884
rect 1427 3876 1513 3884
rect 1607 3876 1973 3884
rect 2976 3884 2984 3893
rect 4096 3904 4104 3913
rect 4096 3896 4293 3904
rect 4307 3896 4413 3904
rect 5707 3896 5893 3904
rect 2976 3876 3033 3884
rect 3047 3876 3093 3884
rect 3413 3884 3427 3893
rect 3413 3880 3773 3884
rect 3416 3876 3773 3880
rect 4147 3876 4193 3884
rect 4467 3876 4633 3884
rect 5487 3876 5633 3884
rect 5747 3876 5853 3884
rect 5987 3876 6113 3884
rect 27 3856 173 3864
rect 407 3856 553 3864
rect 567 3856 593 3864
rect 727 3856 993 3864
rect 1167 3856 1552 3864
rect 1587 3856 1833 3864
rect 2047 3856 2073 3864
rect 2247 3856 2273 3864
rect 2727 3856 2813 3864
rect 2827 3856 2893 3864
rect 3607 3856 3733 3864
rect 6107 3856 6133 3864
rect 6227 3856 6293 3864
rect 367 3836 513 3844
rect 527 3836 553 3844
rect 1027 3836 1213 3844
rect 1287 3836 1893 3844
rect 2627 3836 2773 3844
rect 2947 3836 3153 3844
rect 3787 3836 4173 3844
rect 4527 3836 4573 3844
rect 5907 3836 5933 3844
rect 6047 3836 6153 3844
rect 67 3817 113 3825
rect 227 3816 263 3824
rect 255 3787 263 3816
rect 487 3817 633 3825
rect 847 3817 932 3825
rect 967 3816 1084 3824
rect 47 3775 93 3783
rect 167 3776 193 3784
rect 287 3776 373 3784
rect 435 3784 443 3813
rect 756 3787 764 3813
rect 427 3776 443 3784
rect 587 3775 653 3783
rect 867 3776 993 3784
rect 1007 3775 1033 3783
rect 1076 3784 1084 3816
rect 1107 3816 1144 3824
rect 1076 3776 1113 3784
rect 1136 3784 1144 3816
rect 1327 3816 1373 3824
rect 1507 3816 1813 3824
rect 2007 3817 2033 3825
rect 3207 3816 3453 3824
rect 3587 3816 3673 3824
rect 3696 3816 3813 3824
rect 2076 3787 2084 3813
rect 2107 3797 2233 3805
rect 2487 3796 2613 3804
rect 1136 3776 1224 3784
rect 247 3756 293 3764
rect 507 3756 733 3764
rect 747 3756 833 3764
rect 1216 3764 1224 3776
rect 1287 3775 1312 3783
rect 1347 3776 1393 3784
rect 1487 3775 1533 3783
rect 1687 3776 1713 3784
rect 1847 3775 1893 3783
rect 2167 3776 2273 3784
rect 2687 3775 2753 3783
rect 2836 3784 2844 3813
rect 2836 3776 2873 3784
rect 3113 3784 3127 3793
rect 3167 3795 3293 3803
rect 3067 3780 3127 3784
rect 3456 3780 3573 3784
rect 3067 3776 3124 3780
rect 3453 3776 3573 3780
rect 3453 3767 3467 3776
rect 3696 3786 3704 3816
rect 4267 3817 4293 3825
rect 3936 3804 3944 3814
rect 4216 3804 4224 3814
rect 4907 3816 4973 3824
rect 4987 3816 5073 3824
rect 5187 3816 5293 3824
rect 5527 3817 5713 3825
rect 3887 3796 3944 3804
rect 4136 3796 4224 3804
rect 3767 3775 3833 3783
rect 4136 3784 4144 3796
rect 3987 3776 4144 3784
rect 4167 3776 4193 3784
rect 4327 3776 4433 3784
rect 4487 3775 4513 3783
rect 4536 3784 4544 3813
rect 5176 3804 5184 3814
rect 5967 3817 5993 3825
rect 6107 3824 6120 3827
rect 6107 3813 6124 3824
rect 6167 3817 6232 3825
rect 5107 3796 5184 3804
rect 4536 3776 4773 3784
rect 4787 3776 4873 3784
rect 4987 3775 5013 3783
rect 5167 3776 5213 3784
rect 5607 3776 5693 3784
rect 5776 3784 5784 3813
rect 5776 3776 5813 3784
rect 5887 3776 6013 3784
rect 6116 3784 6124 3813
rect 6253 3804 6267 3813
rect 6253 3800 6304 3804
rect 6256 3796 6304 3800
rect 6296 3787 6304 3796
rect 6116 3776 6133 3784
rect 6247 3776 6273 3784
rect 6296 3776 6313 3787
rect 6300 3773 6313 3776
rect 1216 3756 1293 3764
rect 2127 3756 2153 3764
rect 2667 3756 2713 3764
rect 2807 3756 2853 3764
rect 3756 3764 3764 3772
rect 3667 3756 3764 3764
rect 5067 3756 5093 3764
rect 5107 3756 5133 3764
rect 5387 3756 5833 3764
rect 927 3736 1433 3744
rect 1507 3736 1993 3744
rect 2267 3736 3133 3744
rect 3187 3736 3553 3744
rect 3567 3736 3664 3744
rect 427 3716 544 3724
rect 536 3707 544 3716
rect 607 3716 773 3724
rect 947 3716 1073 3724
rect 1207 3716 1252 3724
rect 1287 3716 1473 3724
rect 1547 3716 1913 3724
rect 1987 3716 2113 3724
rect 2727 3716 2833 3724
rect 3027 3716 3113 3724
rect 3167 3716 3593 3724
rect 3656 3724 3664 3736
rect 3967 3736 3993 3744
rect 4107 3736 4373 3744
rect 5747 3736 5793 3744
rect 5947 3736 6053 3744
rect 3656 3716 3893 3724
rect 4727 3716 4793 3724
rect 5027 3716 5273 3724
rect 547 3696 913 3704
rect 1307 3696 1424 3704
rect 1416 3687 1424 3696
rect 1507 3696 1753 3704
rect 1767 3696 1933 3704
rect 2787 3696 2873 3704
rect 3007 3696 4004 3704
rect 3996 3687 4004 3696
rect 4047 3696 4993 3704
rect 5307 3696 5593 3704
rect 5667 3696 5753 3704
rect 5967 3696 6193 3704
rect 727 3676 833 3684
rect 887 3676 1133 3684
rect 1427 3676 1553 3684
rect 1927 3676 1953 3684
rect 2067 3676 2653 3684
rect 2727 3676 2913 3684
rect 3127 3676 3293 3684
rect 3507 3676 3653 3684
rect 3767 3676 3933 3684
rect 4007 3676 4252 3684
rect 4287 3676 4553 3684
rect 4647 3676 4913 3684
rect 1867 3656 1973 3664
rect 2707 3656 2953 3664
rect 3267 3656 3433 3664
rect 3727 3656 4113 3664
rect 4607 3656 4633 3664
rect 4707 3656 4873 3664
rect 5127 3656 5633 3664
rect 6187 3656 6213 3664
rect 47 3636 433 3644
rect 507 3636 693 3644
rect 807 3636 1393 3644
rect 1407 3636 1653 3644
rect 1887 3636 2573 3644
rect 2587 3636 2673 3644
rect 2887 3636 3153 3644
rect 3607 3636 5373 3644
rect 327 3616 673 3624
rect 956 3616 1193 3624
rect 347 3596 644 3604
rect 467 3576 533 3584
rect 636 3584 644 3596
rect 767 3596 833 3604
rect 956 3604 964 3616
rect 1367 3616 1573 3624
rect 1967 3616 2573 3624
rect 2767 3616 2793 3624
rect 2907 3616 3033 3624
rect 3367 3616 3493 3624
rect 4027 3616 4293 3624
rect 4847 3616 5233 3624
rect 5247 3616 5413 3624
rect 927 3596 964 3604
rect 1007 3596 1233 3604
rect 1247 3596 1313 3604
rect 1807 3596 1933 3604
rect 2847 3596 3013 3604
rect 3147 3596 3273 3604
rect 636 3576 713 3584
rect 1087 3576 1353 3584
rect 2227 3576 2333 3584
rect 2747 3576 2993 3584
rect 3227 3576 3593 3584
rect 3687 3576 3793 3584
rect 4147 3576 4433 3584
rect 5347 3576 5373 3584
rect -24 3556 13 3564
rect 627 3556 713 3564
rect 787 3556 973 3564
rect 1047 3556 1373 3564
rect 2767 3556 2873 3564
rect 2896 3556 3173 3564
rect 147 3536 433 3544
rect 447 3536 493 3544
rect 1147 3536 1193 3544
rect 1480 3544 1493 3547
rect 1476 3533 1493 3544
rect 1547 3536 1604 3544
rect -24 3516 53 3524
rect 67 3516 93 3524
rect 227 3516 253 3524
rect 356 3516 373 3524
rect 356 3487 364 3516
rect 867 3517 913 3525
rect 967 3516 984 3524
rect 636 3484 644 3514
rect 976 3486 984 3516
rect 1380 3524 1393 3527
rect 1376 3513 1393 3524
rect 1116 3487 1124 3513
rect 567 3476 644 3484
rect 847 3475 893 3483
rect 987 3475 1053 3483
rect 287 3456 393 3464
rect 707 3456 853 3464
rect 1156 3464 1164 3513
rect 1227 3476 1273 3484
rect 1376 3486 1384 3513
rect 1476 3486 1484 3533
rect 1596 3524 1604 3536
rect 1827 3536 2144 3544
rect 1596 3516 1613 3524
rect 1767 3516 1884 3524
rect 1516 3487 1524 3513
rect 1576 3484 1584 3513
rect 1576 3476 1593 3484
rect 1716 3484 1724 3513
rect 1876 3486 1884 3516
rect 1907 3516 2013 3524
rect 1687 3476 1724 3484
rect 2056 3484 2064 3514
rect 2136 3504 2144 3536
rect 2667 3536 2704 3544
rect 2167 3516 2213 3524
rect 2256 3507 2264 3533
rect 2313 3524 2327 3533
rect 2296 3520 2327 3524
rect 2696 3524 2704 3536
rect 2727 3536 2772 3544
rect 2896 3544 2904 3556
rect 3607 3556 3833 3564
rect 3847 3556 3973 3564
rect 5947 3556 6233 3564
rect 2807 3536 2904 3544
rect 3147 3536 3213 3544
rect 3596 3544 3604 3552
rect 3287 3536 3604 3544
rect 4787 3536 4853 3544
rect 4967 3536 5053 3544
rect 5547 3536 5573 3544
rect 2296 3516 2324 3520
rect 2696 3516 2753 3524
rect 2136 3496 2232 3504
rect 2296 3504 2304 3516
rect 2767 3516 2824 3524
rect 2856 3520 2893 3524
rect 2276 3496 2304 3504
rect 2316 3500 2473 3504
rect 2313 3496 2473 3500
rect 1896 3480 2064 3484
rect 1893 3476 2064 3480
rect 1893 3467 1907 3476
rect 2107 3476 2193 3484
rect 1156 3456 1193 3464
rect 1767 3456 1793 3464
rect 2276 3467 2284 3496
rect 2313 3487 2327 3496
rect 2627 3496 2673 3504
rect 2816 3487 2824 3516
rect 2853 3516 2893 3520
rect 2853 3507 2867 3516
rect 3187 3495 3353 3503
rect 3676 3503 3684 3533
rect 3887 3517 3973 3525
rect 4147 3517 4233 3525
rect 4327 3517 4353 3525
rect 4547 3517 4633 3525
rect 4887 3517 4913 3525
rect 5127 3517 5153 3525
rect 5387 3517 5473 3525
rect 5807 3517 5933 3525
rect 3627 3495 3693 3503
rect 4056 3504 4064 3514
rect 3747 3496 4064 3504
rect 2587 3476 2733 3484
rect 2907 3476 3233 3484
rect 3827 3476 4184 3484
rect 4176 3467 4184 3476
rect 4227 3476 4273 3484
rect 2276 3456 2293 3467
rect 2280 3453 2293 3456
rect 3307 3456 3613 3464
rect 3887 3456 3933 3464
rect 4176 3456 4193 3467
rect 4180 3453 4193 3456
rect 4396 3464 4404 3514
rect 4816 3504 4824 3514
rect 4816 3496 4864 3504
rect 4567 3475 4613 3483
rect 4807 3476 4833 3484
rect 4856 3484 4864 3496
rect 5027 3500 5104 3504
rect 5027 3496 5107 3500
rect 5093 3487 5107 3496
rect 4856 3476 4893 3484
rect 5273 3484 5287 3493
rect 5273 3480 5353 3484
rect 5276 3476 5353 3480
rect 4367 3456 4404 3464
rect 4707 3456 4753 3464
rect 4767 3456 4872 3464
rect 4896 3464 4904 3473
rect 5676 3484 5684 3514
rect 6276 3487 6284 3514
rect 5627 3476 5684 3484
rect 5707 3476 5733 3484
rect 5787 3475 5853 3483
rect 6107 3476 6173 3484
rect 6276 3476 6293 3487
rect 6280 3473 6293 3476
rect 4896 3456 5013 3464
rect 5087 3456 5113 3464
rect 5407 3456 5533 3464
rect 167 3436 213 3444
rect 427 3436 513 3444
rect 887 3436 913 3444
rect 1087 3436 1233 3444
rect 1347 3436 1413 3444
rect 1727 3436 1853 3444
rect 2707 3436 2773 3444
rect 3227 3436 3633 3444
rect 3647 3436 3733 3444
rect 3847 3436 3953 3444
rect 3967 3436 4153 3444
rect 4947 3436 4973 3444
rect 5567 3436 5713 3444
rect 5767 3444 5780 3447
rect 5767 3433 5784 3444
rect 5827 3436 6273 3444
rect 416 3424 424 3433
rect 327 3416 424 3424
rect 687 3416 773 3424
rect 947 3416 993 3424
rect 1067 3416 1253 3424
rect 1687 3416 1913 3424
rect 1987 3416 2573 3424
rect 2767 3416 3193 3424
rect 3367 3416 3713 3424
rect 3896 3416 4173 3424
rect 947 3396 1013 3404
rect 1287 3396 1413 3404
rect 1716 3396 1753 3404
rect 67 3376 193 3384
rect 467 3376 673 3384
rect 987 3376 1173 3384
rect 1716 3384 1724 3396
rect 2007 3396 2253 3404
rect 2507 3396 2673 3404
rect 2847 3396 3133 3404
rect 3327 3396 3753 3404
rect 3896 3404 3904 3416
rect 4187 3416 4233 3424
rect 4387 3416 4533 3424
rect 4587 3416 4713 3424
rect 5287 3416 5353 3424
rect 5627 3416 5733 3424
rect 5776 3424 5784 3433
rect 5776 3416 5973 3424
rect 5987 3416 6133 3424
rect 3767 3396 3904 3404
rect 3947 3396 4053 3404
rect 4447 3396 4513 3404
rect 4767 3396 4853 3404
rect 4867 3396 4953 3404
rect 5047 3396 5213 3404
rect 6027 3396 6093 3404
rect 1676 3376 1724 3384
rect 1676 3367 1684 3376
rect 1847 3376 2033 3384
rect 2567 3376 2613 3384
rect 2907 3376 2953 3384
rect 3007 3376 3213 3384
rect 3447 3376 3913 3384
rect 4207 3376 4693 3384
rect 5667 3376 5913 3384
rect 5987 3376 6313 3384
rect 267 3356 533 3364
rect 547 3356 633 3364
rect 747 3356 793 3364
rect 867 3356 1093 3364
rect 1107 3356 1133 3364
rect 1227 3356 1413 3364
rect 1647 3356 1673 3364
rect 1747 3356 1853 3364
rect 2047 3356 2113 3364
rect 2587 3356 2693 3364
rect 2747 3356 3233 3364
rect 3527 3356 3593 3364
rect 3967 3356 4013 3364
rect 4027 3356 4073 3364
rect 5487 3356 5633 3364
rect 27 3336 133 3344
rect 1287 3336 1353 3344
rect 1447 3336 1933 3344
rect 1987 3336 2073 3344
rect 3027 3336 3253 3344
rect 3707 3336 3793 3344
rect 4207 3336 4473 3344
rect 4947 3336 5053 3344
rect 5147 3336 5213 3344
rect 5927 3336 6053 3344
rect 227 3316 313 3324
rect 907 3316 1093 3324
rect 1107 3316 1213 3324
rect 1436 3316 1533 3324
rect 187 3296 213 3304
rect 407 3296 504 3304
rect 496 3267 504 3296
rect 27 3255 373 3263
rect 556 3247 564 3313
rect 587 3296 624 3304
rect 616 3264 624 3296
rect 647 3296 684 3304
rect 616 3256 653 3264
rect 676 3264 684 3296
rect 727 3296 853 3304
rect 916 3296 972 3304
rect 916 3267 924 3296
rect 1007 3296 1033 3304
rect 1147 3296 1173 3304
rect 1436 3304 1444 3316
rect 1547 3316 1753 3324
rect 1767 3316 1813 3324
rect 2427 3316 2593 3324
rect 3247 3316 3353 3324
rect 3587 3316 3773 3324
rect 4087 3316 4113 3324
rect 4407 3316 4433 3324
rect 4887 3316 4973 3324
rect 5327 3316 5493 3324
rect 5507 3316 5553 3324
rect 6227 3316 6253 3324
rect 1327 3296 1444 3304
rect 1467 3296 1573 3304
rect 1867 3296 1884 3304
rect 1036 3267 1044 3293
rect 1636 3284 1644 3294
rect 1476 3276 1644 3284
rect 676 3256 833 3264
rect 1087 3256 1192 3264
rect 1476 3266 1484 3276
rect 1227 3255 1253 3263
rect 1527 3256 1593 3264
rect 1636 3264 1644 3276
rect 1876 3284 1884 3296
rect 2087 3297 2113 3305
rect 1687 3276 1804 3284
rect 1876 3280 1944 3284
rect 1876 3276 1947 3280
rect 1636 3256 1733 3264
rect 247 3236 313 3244
rect 556 3236 573 3247
rect 560 3233 573 3236
rect 807 3236 1013 3244
rect 1636 3236 1713 3244
rect 327 3216 413 3224
rect 847 3216 913 3224
rect 1636 3224 1644 3236
rect 1796 3244 1804 3276
rect 1933 3267 1947 3276
rect 2213 3284 2227 3293
rect 2293 3304 2307 3313
rect 2293 3300 2364 3304
rect 2296 3296 2364 3300
rect 2273 3284 2287 3293
rect 1967 3280 2227 3284
rect 1967 3276 2224 3280
rect 2236 3276 2344 3284
rect 1827 3255 1873 3263
rect 1987 3255 2013 3263
rect 2236 3264 2244 3276
rect 2336 3266 2344 3276
rect 2356 3267 2364 3296
rect 2387 3296 2453 3304
rect 2587 3296 2633 3304
rect 2867 3297 2933 3305
rect 2947 3296 3033 3304
rect 3047 3296 3153 3304
rect 3387 3296 3493 3304
rect 4033 3304 4047 3313
rect 4007 3300 4047 3304
rect 4007 3296 4044 3300
rect 4187 3296 4493 3304
rect 3736 3267 3744 3293
rect 4176 3284 4184 3294
rect 4507 3296 4524 3304
rect 5027 3296 5093 3304
rect 3976 3276 4184 3284
rect 2167 3256 2244 3264
rect 2267 3255 2293 3263
rect 2356 3256 2373 3267
rect 2360 3253 2373 3256
rect 2527 3255 2573 3263
rect 2667 3255 2813 3263
rect 3267 3256 3453 3264
rect 3907 3256 3933 3264
rect 3976 3266 3984 3276
rect 4167 3256 4393 3264
rect 4407 3256 4553 3264
rect 4887 3256 4993 3264
rect 5036 3264 5044 3296
rect 5187 3296 5273 3304
rect 5387 3296 5433 3304
rect 5607 3296 5624 3304
rect 5616 3267 5624 3296
rect 5676 3267 5684 3294
rect 5867 3296 5893 3304
rect 5947 3296 6053 3304
rect 5036 3256 5113 3264
rect 5467 3255 5493 3263
rect 5667 3256 5684 3267
rect 5667 3253 5680 3256
rect 5736 3264 5744 3293
rect 5776 3267 5784 3293
rect 5707 3256 5744 3264
rect 1796 3236 1913 3244
rect 2487 3236 2633 3244
rect 2807 3236 3153 3244
rect 3167 3236 3413 3244
rect 3487 3236 3513 3244
rect 3527 3236 3553 3244
rect 5207 3236 5293 3244
rect 5807 3236 5933 3244
rect 5947 3236 6053 3244
rect 6096 3244 6104 3293
rect 6176 3264 6184 3293
rect 6176 3256 6253 3264
rect 6096 3236 6133 3244
rect 1187 3216 1644 3224
rect 1667 3216 1693 3224
rect 1927 3216 1953 3224
rect 2427 3216 2473 3224
rect 2596 3216 2713 3224
rect 127 3196 453 3204
rect 507 3196 793 3204
rect 1156 3196 1433 3204
rect 1156 3187 1164 3196
rect 2596 3204 2604 3216
rect 3087 3216 3113 3224
rect 3127 3216 3293 3224
rect 3307 3216 3373 3224
rect 3647 3216 3713 3224
rect 3727 3216 3813 3224
rect 3887 3216 4013 3224
rect 4027 3216 4153 3224
rect 4227 3216 4253 3224
rect 4467 3216 4833 3224
rect 5427 3216 5473 3224
rect 5936 3224 5944 3232
rect 5936 3216 6113 3224
rect 2287 3196 2604 3204
rect 2627 3196 2953 3204
rect 3507 3196 3593 3204
rect 3787 3196 4193 3204
rect 4487 3196 4613 3204
rect 5627 3196 6153 3204
rect 6167 3196 6293 3204
rect 487 3176 873 3184
rect 987 3176 1153 3184
rect 1567 3176 1873 3184
rect 2227 3176 2353 3184
rect 2367 3176 2833 3184
rect 3087 3176 3433 3184
rect 4087 3176 4253 3184
rect 4327 3176 4373 3184
rect 4387 3176 4593 3184
rect 5636 3176 5753 3184
rect 467 3156 613 3164
rect 927 3156 1173 3164
rect 1267 3156 2393 3164
rect 3107 3156 3424 3164
rect 447 3136 733 3144
rect 1387 3136 1513 3144
rect 1627 3136 1973 3144
rect 2447 3136 3133 3144
rect 3416 3144 3424 3156
rect 3467 3156 3733 3164
rect 3747 3156 3893 3164
rect 5167 3156 5273 3164
rect 5636 3164 5644 3176
rect 6047 3176 6113 3184
rect 5467 3156 5644 3164
rect 5967 3156 6193 3164
rect 3416 3136 3444 3144
rect 67 3116 713 3124
rect 876 3116 1193 3124
rect 876 3107 884 3116
rect 1327 3116 1353 3124
rect 1367 3116 1593 3124
rect 1607 3116 2193 3124
rect 3247 3116 3273 3124
rect 3327 3116 3353 3124
rect 3436 3124 3444 3136
rect 3807 3136 5073 3144
rect 5087 3136 6073 3144
rect 6127 3136 6253 3144
rect 3436 3116 3693 3124
rect 5367 3116 5813 3124
rect 6107 3116 6313 3124
rect 47 3096 133 3104
rect 787 3096 873 3104
rect 1047 3096 1492 3104
rect 1527 3096 1613 3104
rect 1687 3096 1813 3104
rect 1827 3096 1933 3104
rect 1987 3096 2433 3104
rect 2507 3096 2733 3104
rect 2787 3096 2993 3104
rect 3187 3096 3393 3104
rect 3447 3096 3512 3104
rect 3547 3096 3593 3104
rect 4067 3096 4333 3104
rect 5187 3096 5213 3104
rect 5227 3096 5293 3104
rect 527 3076 633 3084
rect 727 3076 944 3084
rect 47 3056 273 3064
rect 387 3056 513 3064
rect 707 3056 913 3064
rect 936 3064 944 3076
rect 2467 3076 2573 3084
rect 3427 3076 3673 3084
rect 3687 3076 3773 3084
rect 4136 3076 4313 3084
rect 4136 3067 4144 3076
rect 4327 3076 4353 3084
rect 4687 3076 4753 3084
rect 5087 3076 5113 3084
rect 5927 3076 6053 3084
rect 936 3056 1372 3064
rect 1407 3056 1673 3064
rect 1847 3056 2093 3064
rect 2547 3056 3093 3064
rect 3147 3056 3253 3064
rect 3447 3056 3573 3064
rect 3927 3056 4133 3064
rect 4207 3056 4393 3064
rect 4507 3056 5253 3064
rect 5267 3056 5313 3064
rect 5387 3056 5873 3064
rect 6000 3064 6013 3067
rect 5996 3053 6013 3064
rect 27 3036 493 3044
rect 1127 3036 1313 3044
rect 1476 3036 1513 3044
rect 107 3016 173 3024
rect 287 3016 333 3024
rect 556 3016 673 3024
rect 147 2996 184 3004
rect 176 2984 184 2996
rect 207 2997 233 3005
rect 407 2997 453 3005
rect 556 2984 564 3016
rect 807 3016 924 3024
rect 916 3008 924 3016
rect 1476 3024 1484 3036
rect 2407 3036 2552 3044
rect 2587 3036 2753 3044
rect 3407 3036 3793 3044
rect 3867 3036 3953 3044
rect 4007 3036 4173 3044
rect 4727 3036 4933 3044
rect 4987 3036 5113 3044
rect 5996 3044 6004 3053
rect 5707 3036 6004 3044
rect 1027 3016 1484 3024
rect 2827 3016 2913 3024
rect 3527 3016 3653 3024
rect 6127 3016 6164 3024
rect 587 2996 793 3004
rect 816 2996 833 3004
rect 176 2976 544 2984
rect 556 2980 584 2984
rect 556 2976 587 2980
rect -24 2956 13 2964
rect 27 2956 73 2964
rect 127 2956 193 2964
rect 327 2956 373 2964
rect 536 2966 544 2976
rect 573 2967 587 2976
rect 467 2956 493 2964
rect 816 2984 824 2996
rect 927 2997 973 3005
rect 1127 2996 1173 3004
rect 1216 2996 1353 3004
rect 753 2964 767 2973
rect 667 2960 767 2964
rect 776 2976 824 2984
rect 667 2956 764 2960
rect 776 2944 784 2976
rect 1216 2984 1224 2996
rect 1447 2997 1472 3005
rect 1507 2997 1533 3005
rect 1587 2997 1613 3005
rect 1653 2984 1667 2993
rect 1067 2976 1224 2984
rect 1456 2980 1667 2984
rect 1456 2976 1664 2980
rect 867 2956 993 2964
rect 1156 2964 1164 2976
rect 1147 2956 1164 2964
rect 1187 2955 1233 2963
rect 1327 2955 1373 2963
rect 1456 2947 1464 2976
rect 1676 2966 1684 3013
rect 1747 2997 1773 3005
rect 1487 2956 1513 2964
rect 1567 2955 1593 2963
rect 1816 2964 1824 2993
rect 2156 2984 2164 2994
rect 2627 2997 2653 3005
rect 1936 2976 2164 2984
rect 1727 2956 1824 2964
rect 1936 2964 1944 2976
rect 2016 2966 2024 2976
rect 1907 2956 1944 2964
rect 2107 2956 2173 2964
rect 2387 2956 2413 2964
rect 2536 2964 2544 2993
rect 2696 2967 2704 2994
rect 2867 2997 2893 3005
rect 2947 2996 2973 3004
rect 3387 2996 3493 3004
rect 2753 2984 2767 2993
rect 2753 2980 2804 2984
rect 2756 2976 2804 2980
rect 2427 2956 2444 2964
rect 2536 2956 2553 2964
rect 707 2936 784 2944
rect 947 2936 973 2944
rect 1447 2936 1464 2947
rect 1447 2933 1460 2936
rect 1787 2936 1853 2944
rect 1967 2936 2013 2944
rect 2027 2936 2133 2944
rect 2436 2944 2444 2956
rect 2696 2956 2713 2967
rect 2700 2953 2713 2956
rect 2796 2966 2804 2976
rect 3096 2976 3153 2984
rect 3096 2966 3104 2976
rect 3207 2976 3313 2984
rect 3496 2967 3504 2994
rect 3827 2996 3973 3004
rect 2927 2955 2953 2963
rect 3487 2956 3504 2967
rect 3487 2953 3500 2956
rect 3576 2964 3584 2993
rect 3527 2956 3673 2964
rect 3787 2955 3833 2963
rect 4016 2964 4024 2994
rect 4156 2966 4164 3013
rect 4187 2996 4344 3004
rect 4336 2984 4344 2996
rect 4367 2996 4453 3004
rect 4527 3004 4540 3007
rect 4527 2993 4544 3004
rect 4567 2996 4733 3004
rect 4747 2996 4793 3004
rect 5047 2997 5233 3005
rect 5396 2996 5453 3004
rect 4536 2984 4544 2993
rect 5396 2984 5404 2996
rect 5627 2997 5693 3005
rect 4196 2976 4324 2984
rect 4336 2976 4444 2984
rect 4536 2976 4584 2984
rect 4196 2966 4204 2976
rect 3887 2956 4024 2964
rect 4056 2956 4113 2964
rect 2436 2936 2533 2944
rect 2647 2936 2793 2944
rect 3147 2936 3173 2944
rect 4056 2944 4064 2956
rect 4256 2956 4293 2964
rect 4007 2936 4064 2944
rect 4256 2944 4264 2956
rect 4316 2947 4324 2976
rect 4436 2966 4444 2976
rect 4576 2966 4584 2976
rect 5376 2976 5404 2984
rect 4667 2955 4733 2963
rect 4827 2956 4893 2964
rect 4907 2956 4953 2964
rect 5376 2964 5384 2976
rect 5516 2964 5524 2994
rect 5307 2956 5384 2964
rect 5436 2960 5524 2964
rect 5433 2956 5524 2960
rect 5736 2967 5744 2994
rect 5736 2956 5753 2967
rect 5433 2947 5447 2956
rect 5740 2953 5753 2956
rect 4127 2936 4264 2944
rect 4407 2936 4564 2944
rect 27 2916 173 2924
rect 187 2916 704 2924
rect 696 2907 704 2916
rect 1207 2916 1413 2924
rect 1527 2916 1653 2924
rect 1727 2916 1913 2924
rect 2687 2916 3173 2924
rect 3187 2916 3473 2924
rect 3627 2916 3653 2924
rect 3847 2916 3873 2924
rect 3967 2916 4073 2924
rect 4556 2924 4564 2936
rect 5487 2936 5573 2944
rect 5647 2936 5713 2944
rect 5816 2944 5824 2993
rect 5907 2956 5933 2964
rect 5956 2964 5964 2993
rect 6053 2984 6067 2993
rect 6053 2980 6104 2984
rect 6056 2976 6104 2980
rect 5956 2956 6013 2964
rect 6096 2964 6104 2976
rect 6156 2966 6164 3016
rect 6096 2956 6113 2964
rect 5816 2936 5873 2944
rect 6176 2944 6184 2994
rect 6147 2936 6184 2944
rect 6236 2947 6244 2993
rect 6236 2936 6253 2947
rect 6240 2933 6253 2936
rect 4556 2916 4693 2924
rect 4707 2916 4852 2924
rect 4887 2916 4993 2924
rect 5207 2916 5253 2924
rect 6187 2916 6313 2924
rect 347 2896 393 2904
rect 707 2896 1173 2904
rect 1467 2896 1893 2904
rect 2087 2896 2233 2904
rect 2767 2896 3013 2904
rect 3067 2896 3133 2904
rect 3267 2896 3453 2904
rect 3767 2896 3813 2904
rect 4247 2896 4533 2904
rect 4967 2896 5033 2904
rect 5607 2896 5833 2904
rect 5907 2896 6273 2904
rect 267 2876 573 2884
rect 647 2876 813 2884
rect 1087 2876 1213 2884
rect 1307 2876 1533 2884
rect 1807 2876 1953 2884
rect 1967 2876 2333 2884
rect 2376 2876 2513 2884
rect 607 2856 853 2864
rect 2376 2864 2384 2876
rect 2967 2876 3193 2884
rect 3287 2876 3353 2884
rect 3407 2876 3593 2884
rect 3767 2876 4033 2884
rect 5287 2876 5533 2884
rect 5896 2884 5904 2893
rect 5787 2876 5904 2884
rect 1987 2856 2384 2864
rect 2927 2856 3073 2864
rect 3727 2856 4053 2864
rect 4547 2856 4613 2864
rect 4767 2856 5093 2864
rect 747 2836 1413 2844
rect 1547 2836 1933 2844
rect 1947 2836 2453 2844
rect 2527 2836 2553 2844
rect 2807 2836 3273 2844
rect 3327 2836 3373 2844
rect 3567 2836 3673 2844
rect 3887 2836 4213 2844
rect 4347 2836 4373 2844
rect 4587 2836 4673 2844
rect 5547 2836 5613 2844
rect 5727 2836 5813 2844
rect 6087 2836 6153 2844
rect 287 2816 893 2824
rect 1067 2816 1173 2824
rect 1956 2816 2013 2824
rect 967 2796 1033 2804
rect 1047 2796 1093 2804
rect 1956 2804 1964 2816
rect 2847 2816 3093 2824
rect 3147 2816 3213 2824
rect 3327 2816 3413 2824
rect 3507 2816 3693 2824
rect 4047 2816 4224 2824
rect 1847 2796 1964 2804
rect 2127 2796 2173 2804
rect 2367 2796 2473 2804
rect 2727 2796 3153 2804
rect -24 2776 13 2784
rect 127 2777 213 2785
rect 327 2776 433 2784
rect 476 2776 513 2784
rect 476 2764 484 2776
rect 587 2776 633 2784
rect 727 2777 773 2785
rect 827 2776 1013 2784
rect 1427 2777 1473 2785
rect 1487 2776 1593 2784
rect 416 2756 484 2764
rect 416 2746 424 2756
rect 167 2736 373 2744
rect 627 2735 693 2743
rect 1336 2744 1344 2774
rect 1607 2776 1684 2784
rect 1676 2764 1684 2776
rect 1787 2777 1813 2785
rect 2207 2777 2233 2785
rect 2347 2777 2373 2785
rect 2396 2776 2533 2784
rect 1973 2764 1987 2773
rect 2396 2764 2404 2776
rect 2847 2776 2933 2784
rect 2947 2777 2973 2785
rect 3027 2776 3073 2784
rect 3096 2784 3104 2796
rect 3567 2796 3633 2804
rect 3927 2796 4073 2804
rect 4216 2804 4224 2816
rect 4247 2816 4293 2824
rect 4667 2816 4733 2824
rect 5087 2816 5393 2824
rect 5747 2816 5793 2824
rect 4216 2796 4313 2804
rect 4256 2788 4264 2796
rect 5327 2796 5373 2804
rect 5847 2796 5973 2804
rect 3096 2776 3184 2784
rect 1676 2760 1987 2764
rect 2356 2760 2404 2764
rect 1676 2756 1984 2760
rect 1267 2736 1392 2744
rect 1427 2736 1453 2744
rect 1507 2736 1633 2744
rect 1707 2736 1753 2744
rect 1827 2736 1873 2744
rect 1976 2744 1984 2756
rect 2353 2756 2404 2760
rect 2353 2747 2367 2756
rect 3176 2747 3184 2776
rect 3247 2776 3344 2784
rect 1976 2736 1993 2744
rect 2047 2735 2073 2743
rect 2707 2736 2813 2744
rect 2947 2736 3053 2744
rect 3176 2736 3193 2747
rect 3180 2733 3193 2736
rect 3336 2746 3344 2776
rect 3367 2776 3493 2784
rect 3547 2777 3593 2785
rect 4027 2776 4093 2784
rect 4447 2776 4593 2784
rect 4787 2776 4813 2784
rect 3833 2764 3847 2773
rect 3756 2760 3847 2764
rect 3756 2756 3844 2760
rect 3247 2735 3293 2743
rect 3627 2735 3673 2743
rect 227 2716 253 2724
rect 987 2716 1033 2724
rect 1247 2716 1793 2724
rect 1927 2716 1953 2724
rect 2027 2716 2293 2724
rect 2307 2716 2433 2724
rect 2447 2716 2473 2724
rect 2627 2716 3053 2724
rect 3756 2724 3764 2756
rect 3907 2735 3973 2743
rect 4136 2744 4144 2774
rect 4436 2764 4444 2774
rect 4887 2776 4933 2784
rect 5007 2777 5053 2785
rect 5067 2776 5213 2784
rect 5767 2777 5813 2785
rect 6047 2777 6093 2785
rect 6140 2784 6153 2787
rect 4227 2756 4444 2764
rect 5496 2747 5504 2774
rect 6136 2773 6153 2784
rect 6267 2776 6313 2784
rect 6136 2764 6144 2773
rect 6116 2756 6144 2764
rect 4047 2736 4144 2744
rect 4507 2736 4653 2744
rect 5067 2736 5153 2744
rect 5287 2735 5353 2743
rect 5407 2736 5433 2744
rect 5487 2736 5504 2747
rect 5487 2733 5500 2736
rect 5687 2735 5753 2743
rect 5847 2736 5873 2744
rect 5887 2736 5933 2744
rect 5947 2736 6053 2744
rect 6116 2746 6124 2756
rect 3687 2716 3764 2724
rect 3787 2716 3873 2724
rect 4007 2716 4113 2724
rect 4827 2716 4893 2724
rect 5027 2716 5173 2724
rect 6187 2716 6293 2724
rect 507 2696 1073 2704
rect 1407 2696 1833 2704
rect 2147 2696 2233 2704
rect 2247 2696 2313 2704
rect 2327 2696 2393 2704
rect 2687 2696 2733 2704
rect 2867 2696 2893 2704
rect 2907 2696 2993 2704
rect 3007 2696 3113 2704
rect 3207 2696 3253 2704
rect 3267 2696 3453 2704
rect 3527 2696 3853 2704
rect 4047 2696 4113 2704
rect 4187 2696 4753 2704
rect 5647 2696 5733 2704
rect 5867 2696 6073 2704
rect 6227 2696 6273 2704
rect 867 2676 1193 2684
rect 2007 2676 2493 2684
rect 3167 2676 3533 2684
rect 3927 2676 4613 2684
rect 4967 2676 5113 2684
rect 5727 2676 6053 2684
rect 727 2656 773 2664
rect 1107 2656 1373 2664
rect 1807 2656 2533 2664
rect 3087 2656 3133 2664
rect 3447 2656 3733 2664
rect 4087 2656 4153 2664
rect 4247 2656 4253 2664
rect 4267 2656 4313 2664
rect 4647 2656 4933 2664
rect 4947 2656 5033 2664
rect 5627 2656 5773 2664
rect 1827 2636 2013 2644
rect 2067 2636 2333 2644
rect 2407 2636 2624 2644
rect 367 2616 653 2624
rect 767 2616 793 2624
rect 807 2616 1353 2624
rect 2127 2616 2253 2624
rect 2616 2624 2624 2636
rect 3156 2636 3813 2644
rect 3156 2624 3164 2636
rect 3827 2636 3933 2644
rect 4627 2636 5593 2644
rect 2616 2616 3164 2624
rect 3287 2616 3593 2624
rect 3667 2616 3893 2624
rect 3987 2616 4193 2624
rect 4287 2616 4453 2624
rect 47 2596 1333 2604
rect 1387 2596 1713 2604
rect 1727 2596 1933 2604
rect 2367 2596 2473 2604
rect 2547 2596 2873 2604
rect 3076 2596 3133 2604
rect 3076 2587 3084 2596
rect 3196 2596 3913 2604
rect 207 2576 413 2584
rect 427 2576 1253 2584
rect 1967 2576 2393 2584
rect 2587 2576 3073 2584
rect 3196 2584 3204 2596
rect 4247 2596 4853 2604
rect 4967 2596 5373 2604
rect 3156 2576 3204 2584
rect 1367 2556 1493 2564
rect 1507 2556 1873 2564
rect 3156 2564 3164 2576
rect 3227 2576 3653 2584
rect 3747 2576 3793 2584
rect 3807 2576 3873 2584
rect 4107 2576 4493 2584
rect 2507 2556 3164 2564
rect 3207 2556 3353 2564
rect 3367 2556 3673 2564
rect 1347 2536 1513 2544
rect 1667 2536 1733 2544
rect 1747 2536 2033 2544
rect 2447 2536 2793 2544
rect 2807 2536 3133 2544
rect 3187 2536 3633 2544
rect 3647 2536 3693 2544
rect 3907 2536 3933 2544
rect 3947 2536 3993 2544
rect 4827 2536 5133 2544
rect 5147 2536 5253 2544
rect 5487 2536 5693 2544
rect 5707 2536 5973 2544
rect 47 2516 313 2524
rect 327 2516 653 2524
rect 1327 2516 1533 2524
rect 3227 2516 3373 2524
rect 3887 2516 4073 2524
rect 5227 2516 5413 2524
rect 5427 2516 5553 2524
rect 6167 2516 6273 2524
rect 1627 2496 1953 2504
rect 2607 2496 2913 2504
rect 3107 2496 3393 2504
rect 4047 2496 4093 2504
rect 5327 2504 5340 2507
rect 5327 2493 5344 2504
rect 5867 2496 5933 2504
rect 6107 2496 6193 2504
rect 267 2477 353 2485
rect 607 2476 713 2484
rect 116 2456 193 2464
rect 116 2446 124 2456
rect 456 2447 464 2474
rect 1227 2476 1353 2484
rect 456 2436 473 2447
rect 460 2433 473 2436
rect 776 2446 784 2473
rect 747 2435 773 2443
rect 936 2444 944 2474
rect 1076 2464 1084 2474
rect 1016 2456 1084 2464
rect 847 2436 944 2444
rect 1016 2444 1024 2456
rect 967 2436 1024 2444
rect 1047 2436 1093 2444
rect 1396 2444 1404 2474
rect 1787 2476 1813 2484
rect 2007 2476 2433 2484
rect 2747 2476 2833 2484
rect 1907 2456 2173 2464
rect 2096 2446 2104 2456
rect 2893 2464 2907 2473
rect 2876 2460 2907 2464
rect 2876 2456 2904 2460
rect 1396 2436 1553 2444
rect 1567 2436 1693 2444
rect 1707 2435 1793 2443
rect 1967 2435 2013 2443
rect 2647 2435 2713 2443
rect 2876 2444 2884 2456
rect 2867 2436 2884 2444
rect 2907 2436 2933 2444
rect 3016 2444 3024 2474
rect 3147 2476 3313 2484
rect 3787 2476 3853 2484
rect 3947 2476 4004 2484
rect 3053 2464 3067 2473
rect 3053 2460 3953 2464
rect 3056 2456 3953 2460
rect 3996 2447 4004 2476
rect 3016 2436 3113 2444
rect 3287 2436 3333 2444
rect 3467 2436 3573 2444
rect 3707 2435 3753 2443
rect 4156 2444 4164 2493
rect 4367 2477 4393 2485
rect 4507 2476 4593 2484
rect 4767 2476 4913 2484
rect 5007 2476 5093 2484
rect 5207 2477 5293 2485
rect 4156 2440 4184 2444
rect 4156 2436 4187 2440
rect 447 2416 513 2424
rect 1527 2416 1553 2424
rect 2147 2416 2173 2424
rect 2267 2416 2373 2424
rect 2636 2424 2644 2432
rect 4173 2427 4187 2436
rect 4236 2444 4244 2473
rect 5096 2447 5104 2474
rect 5336 2464 5344 2493
rect 5387 2484 5400 2487
rect 5387 2473 5404 2484
rect 4207 2436 4244 2444
rect 4267 2435 4453 2443
rect 4807 2435 4853 2443
rect 4867 2436 4933 2444
rect 5087 2436 5104 2447
rect 5316 2456 5344 2464
rect 5316 2444 5324 2456
rect 5396 2446 5404 2473
rect 5296 2440 5324 2444
rect 5293 2436 5324 2440
rect 5087 2433 5100 2436
rect 5293 2427 5307 2436
rect 5456 2444 5464 2474
rect 5787 2477 6013 2485
rect 5616 2447 5624 2473
rect 5416 2440 5464 2444
rect 5413 2436 5464 2440
rect 2587 2416 2644 2424
rect 3007 2416 3093 2424
rect 3516 2416 3833 2424
rect 3516 2407 3524 2416
rect 3907 2416 4053 2424
rect 4067 2416 4113 2424
rect 5016 2416 5213 2424
rect 87 2396 393 2404
rect 707 2396 833 2404
rect 947 2396 1013 2404
rect 1447 2396 1593 2404
rect 1947 2396 2013 2404
rect 3167 2396 3213 2404
rect 3307 2396 3493 2404
rect 3507 2396 3524 2407
rect 3507 2393 3520 2396
rect 3987 2396 4033 2404
rect 4107 2396 4153 2404
rect 4167 2396 4273 2404
rect 4347 2396 4613 2404
rect 5016 2404 5024 2416
rect 5413 2427 5427 2436
rect 6216 2444 6224 2473
rect 6147 2436 6224 2444
rect 5647 2416 5833 2424
rect 5887 2416 6073 2424
rect 6087 2416 6172 2424
rect 6207 2416 6293 2424
rect 4667 2396 5024 2404
rect 5047 2396 5253 2404
rect 5467 2396 5533 2404
rect 5707 2396 5773 2404
rect 5867 2396 5913 2404
rect 1647 2376 1913 2384
rect 1927 2376 2124 2384
rect 287 2356 553 2364
rect 1387 2356 1773 2364
rect 2116 2364 2124 2376
rect 2467 2376 2613 2384
rect 2807 2376 2833 2384
rect 3647 2376 3913 2384
rect 4987 2376 5113 2384
rect 5587 2376 5653 2384
rect 6047 2376 6093 2384
rect 2116 2356 2433 2364
rect 3627 2356 3804 2364
rect 736 2336 1293 2344
rect 147 2316 533 2324
rect 736 2324 744 2336
rect 1427 2336 1513 2344
rect 1887 2336 1953 2344
rect 2007 2336 2093 2344
rect 2367 2336 2953 2344
rect 3107 2336 3193 2344
rect 3347 2336 3593 2344
rect 3687 2336 3713 2344
rect 3796 2344 3804 2356
rect 3827 2356 3873 2364
rect 3947 2356 4113 2364
rect 4467 2356 4553 2364
rect 5116 2364 5124 2373
rect 5116 2356 5273 2364
rect 5447 2356 5993 2364
rect 3796 2336 4193 2344
rect 5387 2336 5493 2344
rect 5607 2336 5933 2344
rect 707 2316 744 2324
rect 1007 2316 1193 2324
rect 1267 2316 1433 2324
rect 1447 2316 1633 2324
rect 1687 2316 1853 2324
rect 2447 2316 2553 2324
rect 2667 2316 2973 2324
rect 2987 2316 3013 2324
rect 3647 2316 3773 2324
rect 3867 2316 4093 2324
rect 4367 2316 4993 2324
rect 5007 2316 5073 2324
rect 5407 2316 5453 2324
rect 287 2296 313 2304
rect 387 2296 453 2304
rect 1547 2296 1613 2304
rect 1807 2296 1893 2304
rect 2367 2296 2413 2304
rect 3047 2296 3093 2304
rect 3227 2296 3273 2304
rect 3667 2296 3733 2304
rect 4427 2296 4533 2304
rect 4667 2296 4893 2304
rect 4907 2296 4973 2304
rect 5227 2296 5273 2304
rect 5287 2296 5493 2304
rect 5547 2296 5633 2304
rect 5927 2296 5953 2304
rect 527 2276 593 2284
rect 1127 2276 1153 2284
rect 1167 2276 1293 2284
rect 1487 2276 1713 2284
rect 1727 2276 1933 2284
rect 1947 2276 1993 2284
rect 2047 2276 2433 2284
rect 2487 2276 2533 2284
rect 2927 2276 2993 2284
rect 3147 2276 3173 2284
rect 3736 2284 3744 2293
rect 3736 2276 3813 2284
rect 3876 2276 3933 2284
rect 147 2257 173 2265
rect 287 2256 372 2264
rect 207 2215 253 2223
rect 396 2224 404 2254
rect 827 2257 853 2265
rect 1027 2257 1073 2265
rect 493 2244 507 2253
rect 1167 2257 1193 2265
rect 1247 2256 1384 2264
rect 493 2240 524 2244
rect 496 2236 524 2240
rect 307 2216 404 2224
rect 427 2216 473 2224
rect 516 2226 524 2236
rect 1376 2227 1384 2256
rect 607 2215 753 2223
rect 1007 2215 1053 2223
rect 1267 2215 1293 2223
rect 167 2196 253 2204
rect 867 2196 973 2204
rect 1296 2204 1304 2212
rect 1436 2207 1444 2273
rect 3876 2268 3884 2276
rect 4127 2276 4293 2284
rect 5347 2276 5433 2284
rect 5447 2276 5473 2284
rect 5527 2276 5633 2284
rect 1867 2256 2013 2264
rect 2127 2256 2313 2264
rect 2327 2256 2373 2264
rect 2427 2257 2793 2265
rect 1556 2227 1564 2253
rect 1756 2227 1764 2253
rect 2936 2227 2944 2254
rect 3107 2256 3253 2264
rect 3467 2256 3593 2264
rect 3616 2256 3653 2264
rect 3007 2236 3164 2244
rect 1627 2216 1732 2224
rect 1887 2215 1933 2223
rect 2047 2215 2093 2223
rect 2267 2215 2293 2223
rect 2827 2215 2913 2223
rect 2936 2216 2953 2227
rect 2940 2213 2953 2216
rect 3156 2224 3164 2236
rect 3416 2227 3424 2253
rect 3616 2244 3624 2256
rect 3787 2264 3800 2267
rect 3787 2253 3804 2264
rect 3907 2256 3933 2264
rect 3596 2236 3624 2244
rect 3156 2216 3233 2224
rect 3247 2216 3313 2224
rect 3596 2224 3604 2236
rect 3587 2216 3604 2224
rect 3796 2207 3804 2253
rect 3836 2207 3844 2253
rect 3867 2216 3933 2224
rect 1296 2196 1393 2204
rect 2007 2196 2053 2204
rect 3007 2196 3353 2204
rect 3487 2196 3553 2204
rect 3747 2196 3772 2204
rect 3976 2204 3984 2273
rect 6107 2276 6173 2284
rect 4147 2256 4164 2264
rect 4156 2227 4164 2256
rect 4376 2256 4393 2264
rect 4007 2216 4073 2224
rect 4376 2226 4384 2256
rect 4407 2256 4473 2264
rect 4547 2257 4613 2265
rect 4627 2256 4773 2264
rect 4827 2256 4953 2264
rect 5007 2256 5084 2264
rect 5076 2226 5084 2256
rect 5127 2257 5173 2265
rect 5240 2264 5253 2267
rect 5236 2253 5253 2264
rect 5507 2256 5644 2264
rect 5236 2226 5244 2253
rect 5636 2226 5644 2256
rect 5827 2256 5893 2264
rect 5907 2256 5953 2264
rect 6007 2257 6053 2265
rect 6256 2244 6264 2254
rect 6216 2236 6264 2244
rect 4247 2216 4333 2224
rect 4447 2215 4493 2223
rect 4567 2215 4633 2223
rect 4927 2216 5033 2224
rect 5287 2215 5313 2223
rect 5367 2215 5393 2223
rect 6216 2224 6224 2236
rect 6276 2224 6284 2273
rect 6316 2227 6324 2253
rect 6047 2216 6224 2224
rect 6256 2220 6284 2224
rect 6253 2216 6284 2220
rect 6253 2207 6267 2216
rect 3907 2196 3984 2204
rect 4647 2196 4793 2204
rect 5907 2196 5993 2204
rect 6127 2196 6153 2204
rect 647 2176 793 2184
rect 1387 2176 1573 2184
rect 1996 2184 2004 2193
rect 1847 2176 2004 2184
rect 2747 2176 2953 2184
rect 3007 2176 3113 2184
rect 3287 2176 3613 2184
rect 4027 2176 4173 2184
rect 4347 2176 4413 2184
rect 4967 2176 5093 2184
rect 5147 2176 5433 2184
rect 5447 2176 5473 2184
rect 927 2156 1033 2164
rect 1227 2156 1293 2164
rect 1307 2156 1513 2164
rect 1787 2156 1993 2164
rect 2707 2156 2873 2164
rect 2947 2156 2973 2164
rect 2987 2156 3313 2164
rect 3487 2156 3673 2164
rect 3727 2156 3773 2164
rect 3787 2156 3892 2164
rect 3927 2156 4113 2164
rect 1567 2136 1693 2144
rect 3087 2136 3293 2144
rect 3987 2136 4253 2144
rect 4607 2136 4753 2144
rect 307 2116 833 2124
rect 987 2116 1413 2124
rect 1867 2116 1973 2124
rect 2027 2116 2393 2124
rect 2407 2116 2873 2124
rect 3607 2116 3804 2124
rect 927 2096 1493 2104
rect 1887 2096 2173 2104
rect 2427 2096 2633 2104
rect 3027 2096 3473 2104
rect 3727 2096 3753 2104
rect 3796 2104 3804 2116
rect 3827 2116 3873 2124
rect 3887 2116 4273 2124
rect 5927 2116 5993 2124
rect 3796 2096 3972 2104
rect 4007 2096 4033 2104
rect 4267 2096 4453 2104
rect 4467 2096 4533 2104
rect 4627 2096 4693 2104
rect 1627 2076 1653 2084
rect 1667 2076 2793 2084
rect 2987 2076 3373 2084
rect 3387 2076 3513 2084
rect 3527 2076 3612 2084
rect 3647 2076 3833 2084
rect 3847 2076 4013 2084
rect 4207 2076 4973 2084
rect 4987 2076 5033 2084
rect 5387 2076 5733 2084
rect 6107 2076 6233 2084
rect 567 2056 893 2064
rect 907 2056 1373 2064
rect 1947 2056 2333 2064
rect 2607 2056 2753 2064
rect 2887 2056 2953 2064
rect 3307 2056 3693 2064
rect 3807 2056 4673 2064
rect 6087 2056 6273 2064
rect 367 2036 993 2044
rect 1007 2036 1533 2044
rect 2487 2036 2973 2044
rect 3027 2036 3193 2044
rect 3207 2036 3813 2044
rect 4307 2036 4613 2044
rect 5067 2036 5273 2044
rect 5807 2036 6153 2044
rect 527 2016 773 2024
rect 787 2016 873 2024
rect 1167 2016 1973 2024
rect 2207 2016 2413 2024
rect 3327 2016 3753 2024
rect 3767 2016 3893 2024
rect 4687 2016 4873 2024
rect 107 1996 193 2004
rect 707 1996 753 2004
rect 1456 1996 1953 2004
rect 1456 1984 1464 1996
rect 2567 1996 2693 2004
rect 2847 1996 2993 2004
rect 3267 1996 3413 2004
rect 3547 1996 3573 2004
rect 3587 1996 3713 2004
rect 4047 1996 4373 2004
rect 4547 1996 5073 2004
rect 6087 1996 6113 2004
rect 1387 1976 1464 1984
rect 2027 1976 2073 1984
rect 2167 1976 2233 1984
rect 3646 1973 3647 1980
rect 3667 1976 4013 1984
rect 4167 1976 4713 1984
rect 4727 1976 4753 1984
rect 4896 1976 5004 1984
rect 127 1956 164 1964
rect 156 1927 164 1956
rect 347 1957 373 1965
rect 427 1956 473 1964
rect 487 1957 533 1965
rect 647 1957 713 1965
rect 727 1956 793 1964
rect 980 1964 993 1967
rect 296 1924 304 1954
rect 976 1953 993 1964
rect 1107 1956 1213 1964
rect 1267 1956 1284 1964
rect 227 1916 304 1924
rect 407 1915 493 1923
rect 647 1915 813 1923
rect 827 1916 913 1924
rect 976 1924 984 1953
rect 1276 1927 1284 1956
rect 1507 1956 1573 1964
rect 1616 1956 1693 1964
rect 1616 1944 1624 1956
rect 1707 1956 1853 1964
rect 2056 1944 2064 1954
rect 2287 1957 2313 1965
rect 2427 1956 2464 1964
rect 1596 1936 1624 1944
rect 1876 1936 2064 1944
rect 967 1916 984 1924
rect 1047 1916 1193 1924
rect 1596 1926 1604 1936
rect 1876 1927 1884 1936
rect 1316 1916 1593 1924
rect 1316 1907 1324 1916
rect 1867 1916 1884 1927
rect 1867 1913 1880 1916
rect 1907 1915 2013 1923
rect 2136 1924 2144 1953
rect 2456 1944 2464 1956
rect 2607 1957 2653 1965
rect 2456 1936 2504 1944
rect 2087 1916 2144 1924
rect 2267 1916 2333 1924
rect 2447 1916 2473 1924
rect 2496 1924 2504 1936
rect 2676 1926 2684 1973
rect 2976 1956 3053 1964
rect 2976 1944 2984 1956
rect 3146 1953 3147 1960
rect 3167 1956 3193 1964
rect 3133 1944 3147 1953
rect 2956 1936 2984 1944
rect 3096 1940 3147 1944
rect 3096 1936 3143 1940
rect 2956 1926 2964 1936
rect 2496 1916 2533 1924
rect 3096 1924 3104 1936
rect 3007 1916 3104 1924
rect 3127 1915 3153 1923
rect 3296 1924 3304 1954
rect 3316 1944 3324 1973
rect 3633 1964 3647 1973
rect 3347 1956 3404 1964
rect 3316 1936 3364 1944
rect 3356 1926 3364 1936
rect 3396 1927 3404 1956
rect 3616 1960 3647 1964
rect 3616 1956 3643 1960
rect 3227 1916 3304 1924
rect 3616 1924 3624 1956
rect 3707 1956 3793 1964
rect 3967 1957 3993 1965
rect 4247 1957 4333 1965
rect 4896 1964 4904 1976
rect 4567 1956 4904 1964
rect 4996 1964 5004 1976
rect 6140 1984 6153 1987
rect 5047 1976 5104 1984
rect 5096 1968 5104 1976
rect 6136 1973 6153 1984
rect 6267 1976 6324 1984
rect 4996 1956 5013 1964
rect 5027 1956 5084 1964
rect 5076 1944 5084 1956
rect 5227 1957 5313 1965
rect 5447 1956 5733 1964
rect 6136 1967 6144 1973
rect 5907 1956 6033 1964
rect 5076 1936 5204 1944
rect 3507 1916 3633 1924
rect 3827 1916 4033 1924
rect 4236 1916 4533 1924
rect 147 1896 173 1904
rect 187 1896 373 1904
rect 527 1896 653 1904
rect 1027 1896 1113 1904
rect 1300 1906 1324 1907
rect 1307 1896 1324 1906
rect 1307 1893 1320 1896
rect 1467 1896 1633 1904
rect 2127 1896 2173 1904
rect 2187 1896 2413 1904
rect 2567 1896 2613 1904
rect 3267 1896 3313 1904
rect 3327 1896 3433 1904
rect 3687 1896 3753 1904
rect 4236 1904 4244 1916
rect 4767 1915 4833 1923
rect 5007 1916 5053 1924
rect 5196 1926 5204 1936
rect 5347 1916 5533 1924
rect 5547 1916 5633 1924
rect 5816 1924 5824 1953
rect 5956 1944 5964 1956
rect 6087 1964 6100 1967
rect 6087 1953 6104 1964
rect 6187 1957 6233 1965
rect 5956 1936 5984 1944
rect 5816 1916 5833 1924
rect 5976 1924 5984 1936
rect 5976 1916 6073 1924
rect 6096 1924 6104 1953
rect 6096 1916 6113 1924
rect 6167 1915 6213 1923
rect 6296 1924 6304 1953
rect 6267 1916 6304 1924
rect 6316 1907 6324 1976
rect 3987 1896 4244 1904
rect 4267 1896 4824 1904
rect 107 1876 193 1884
rect 207 1876 693 1884
rect 767 1876 853 1884
rect 947 1876 1353 1884
rect 1727 1876 1893 1884
rect 1987 1876 2453 1884
rect 2527 1876 2773 1884
rect 3947 1876 4173 1884
rect 4816 1884 4824 1896
rect 5847 1896 5973 1904
rect 6307 1896 6324 1907
rect 6307 1893 6320 1896
rect 4816 1876 5333 1884
rect 167 1856 233 1864
rect 287 1856 333 1864
rect 347 1856 553 1864
rect 607 1856 1073 1864
rect 1087 1856 1253 1864
rect 1487 1856 1533 1864
rect 1967 1856 2084 1864
rect 667 1836 753 1844
rect 1427 1836 1573 1844
rect 1587 1836 1613 1844
rect 1627 1836 1813 1844
rect 1867 1836 2053 1844
rect 2076 1844 2084 1856
rect 2447 1856 2493 1864
rect 2907 1856 2973 1864
rect 3087 1856 3133 1864
rect 3467 1856 3833 1864
rect 4176 1864 4184 1873
rect 4176 1856 4293 1864
rect 4307 1856 4393 1864
rect 5167 1856 5213 1864
rect 5227 1856 5413 1864
rect 5607 1856 5653 1864
rect 5807 1856 5873 1864
rect 5947 1856 6013 1864
rect 6127 1856 6193 1864
rect 2076 1836 2633 1844
rect 2767 1836 3213 1844
rect 3567 1836 3713 1844
rect 4807 1836 4853 1844
rect 5307 1836 5373 1844
rect 447 1816 973 1824
rect 987 1816 1193 1824
rect 1207 1816 1233 1824
rect 1807 1816 2213 1824
rect 2787 1816 3053 1824
rect 3307 1816 3393 1824
rect 3687 1816 3733 1824
rect 4127 1816 4313 1824
rect 6187 1816 6233 1824
rect 727 1796 793 1804
rect 1047 1796 1133 1804
rect 1287 1796 1373 1804
rect 1387 1796 1593 1804
rect 1827 1796 1873 1804
rect 2007 1796 2513 1804
rect 2887 1796 3033 1804
rect 3096 1796 3873 1804
rect 3096 1787 3104 1796
rect 4007 1796 4113 1804
rect 4807 1796 5013 1804
rect 5907 1796 6053 1804
rect 6067 1796 6133 1804
rect 347 1776 493 1784
rect 627 1776 1513 1784
rect 1907 1776 1973 1784
rect 2407 1776 2593 1784
rect 2647 1776 2913 1784
rect 2967 1776 3093 1784
rect 3247 1776 3573 1784
rect 4247 1776 4433 1784
rect 5247 1776 5293 1784
rect 6267 1776 6313 1784
rect 140 1764 153 1767
rect 136 1753 153 1764
rect 207 1756 264 1764
rect 67 1737 113 1745
rect 136 1706 144 1753
rect 207 1737 233 1745
rect 256 1706 264 1756
rect 387 1756 573 1764
rect 667 1756 693 1764
rect 927 1756 1232 1764
rect 3047 1756 3193 1764
rect 3316 1756 3533 1764
rect 287 1736 353 1744
rect 766 1734 767 1748
rect 787 1737 813 1745
rect 307 1695 333 1703
rect 416 1704 424 1734
rect 756 1724 764 1734
rect 827 1737 872 1745
rect 1207 1744 1220 1747
rect 1207 1733 1224 1744
rect 756 1716 804 1724
rect 387 1696 424 1704
rect 447 1696 493 1704
rect 507 1696 533 1704
rect 607 1696 653 1704
rect 667 1695 693 1703
rect 796 1704 804 1716
rect 896 1707 904 1733
rect 796 1696 833 1704
rect 1216 1706 1224 1733
rect 1256 1706 1264 1753
rect 1287 1736 1344 1744
rect 1007 1696 1093 1704
rect 1336 1704 1344 1736
rect 1447 1737 1513 1745
rect 1787 1737 1833 1745
rect 2207 1737 2252 1745
rect 2287 1737 2353 1745
rect 1593 1724 1607 1733
rect 1593 1720 1644 1724
rect 1596 1716 1644 1720
rect 1636 1706 1644 1716
rect 1307 1696 1393 1704
rect 1647 1696 1753 1704
rect 1916 1704 1924 1734
rect 2467 1736 2713 1744
rect 2807 1737 2873 1745
rect 2927 1736 3233 1744
rect 2427 1716 2853 1724
rect 3316 1707 3324 1756
rect 3707 1756 3753 1764
rect 3927 1756 4153 1764
rect 4467 1756 4533 1764
rect 4547 1756 4573 1764
rect 4627 1756 4713 1764
rect 5087 1756 5153 1764
rect 5167 1756 5213 1764
rect 5407 1756 5453 1764
rect 5467 1756 5493 1764
rect 5687 1756 5744 1764
rect 3367 1736 3384 1744
rect 1896 1696 1924 1704
rect 1896 1684 1904 1696
rect 1987 1696 2133 1704
rect 2247 1696 2433 1704
rect 2447 1696 2813 1704
rect 2987 1695 3253 1703
rect 3376 1687 3384 1736
rect 3475 1736 3493 1744
rect 3407 1696 3433 1704
rect 3475 1687 3483 1736
rect 3587 1737 3613 1745
rect 3827 1737 3913 1745
rect 3967 1736 4013 1744
rect 4067 1736 4133 1744
rect 4296 1740 4333 1744
rect 4293 1736 4333 1740
rect 4293 1727 4307 1736
rect 4387 1736 4433 1744
rect 4507 1736 4524 1744
rect 4516 1724 4524 1736
rect 4647 1736 4684 1744
rect 4676 1724 4684 1736
rect 4707 1737 4753 1745
rect 4476 1720 4624 1724
rect 4473 1716 4624 1720
rect 4676 1720 4844 1724
rect 4676 1716 4847 1720
rect 4473 1707 4487 1716
rect 3547 1696 3653 1704
rect 3747 1696 3813 1704
rect 4327 1695 4353 1703
rect 4616 1704 4624 1716
rect 4833 1707 4847 1716
rect 4616 1696 4653 1704
rect 4896 1706 4904 1753
rect 5127 1736 5244 1744
rect 1667 1676 1904 1684
rect 1927 1676 2013 1684
rect 2087 1676 2173 1684
rect 2227 1676 2333 1684
rect 2487 1676 2513 1684
rect 2527 1676 2673 1684
rect 2747 1676 2793 1684
rect 2867 1676 3053 1684
rect 3307 1676 3352 1684
rect 3507 1676 3553 1684
rect 3847 1676 3873 1684
rect 3887 1676 4073 1684
rect 4147 1676 4393 1684
rect 4407 1676 4453 1684
rect 4527 1676 4773 1684
rect 67 1656 393 1664
rect 447 1656 793 1664
rect 1007 1656 1033 1664
rect 1147 1656 1233 1664
rect 1247 1656 1293 1664
rect 1647 1656 1692 1664
rect 1727 1656 1813 1664
rect 1887 1656 1924 1664
rect 87 1636 373 1644
rect 1327 1636 1393 1644
rect 1807 1636 1893 1644
rect 1916 1644 1924 1656
rect 2547 1656 2653 1664
rect 2727 1656 2773 1664
rect 2787 1656 3013 1664
rect 3027 1656 3293 1664
rect 3687 1656 3773 1664
rect 4956 1664 4964 1734
rect 5236 1724 5244 1736
rect 5267 1736 5413 1744
rect 5236 1716 5264 1724
rect 5256 1704 5264 1716
rect 5376 1706 5384 1736
rect 5547 1736 5593 1744
rect 5736 1707 5744 1756
rect 6047 1756 6093 1764
rect 5847 1737 5913 1745
rect 5953 1724 5967 1733
rect 5936 1720 5967 1724
rect 5936 1716 5964 1720
rect 5256 1696 5333 1704
rect 5467 1695 5553 1703
rect 5027 1676 5093 1684
rect 5727 1676 5773 1684
rect 5936 1684 5944 1716
rect 5996 1704 6004 1734
rect 6176 1724 6184 1734
rect 6087 1716 6184 1724
rect 6216 1707 6224 1733
rect 6296 1724 6304 1753
rect 6327 1744 6340 1747
rect 6327 1733 6344 1744
rect 6296 1720 6324 1724
rect 6296 1716 6327 1720
rect 6313 1707 6327 1716
rect 5967 1696 6004 1704
rect 6207 1696 6213 1704
rect 6227 1696 6273 1704
rect 5887 1676 5944 1684
rect 6127 1676 6173 1684
rect 4847 1656 4964 1664
rect 5667 1656 5733 1664
rect 5867 1656 5913 1664
rect 5927 1656 5973 1664
rect 6087 1656 6193 1664
rect 6336 1664 6344 1733
rect 6307 1656 6344 1664
rect 1916 1636 2333 1644
rect 2507 1636 2593 1644
rect 3707 1636 4064 1644
rect 207 1616 273 1624
rect 447 1616 833 1624
rect 1167 1616 1333 1624
rect 1347 1616 1373 1624
rect 1567 1616 1713 1624
rect 1767 1616 1853 1624
rect 2007 1616 2073 1624
rect 2827 1616 3193 1624
rect 3207 1616 3313 1624
rect 3436 1616 3973 1624
rect 47 1596 224 1604
rect 216 1587 224 1596
rect 487 1596 1173 1604
rect 1227 1596 1453 1604
rect 1547 1596 1973 1604
rect 2027 1596 2233 1604
rect 2307 1596 2533 1604
rect 3436 1604 3444 1616
rect 4056 1624 4064 1636
rect 5607 1636 5813 1644
rect 5827 1636 5913 1644
rect 5927 1636 5953 1644
rect 6027 1636 6233 1644
rect 4056 1616 4513 1624
rect 5107 1616 5233 1624
rect 2956 1596 3444 1604
rect 216 1576 233 1587
rect 220 1573 233 1576
rect 247 1576 593 1584
rect 747 1576 933 1584
rect 947 1576 1913 1584
rect 1927 1576 2373 1584
rect 2956 1584 2964 1596
rect 3467 1596 4113 1604
rect 4187 1596 4973 1604
rect 5847 1596 5993 1604
rect 2387 1576 2964 1584
rect 2987 1576 3173 1584
rect 3427 1576 5053 1584
rect 5067 1576 5193 1584
rect 5507 1576 5673 1584
rect 6047 1576 6073 1584
rect 6087 1576 6233 1584
rect 1307 1556 1433 1564
rect 1447 1556 1513 1564
rect 1747 1556 1953 1564
rect 2007 1556 2153 1564
rect 2267 1556 2392 1564
rect 2427 1556 3153 1564
rect 4147 1556 4293 1564
rect 5847 1556 5893 1564
rect 207 1536 633 1544
rect 647 1536 673 1544
rect 1087 1536 1273 1544
rect 1327 1536 2053 1544
rect 2547 1536 2613 1544
rect 2707 1536 2884 1544
rect 1447 1516 1793 1524
rect 2116 1516 2213 1524
rect 2116 1507 2124 1516
rect 2267 1516 2433 1524
rect 2627 1516 2853 1524
rect 2876 1524 2884 1536
rect 2907 1536 2953 1544
rect 2967 1536 3173 1544
rect 3347 1536 3453 1544
rect 3907 1536 3973 1544
rect 3987 1536 4073 1544
rect 6007 1536 6113 1544
rect 6127 1536 6293 1544
rect 2876 1516 2973 1524
rect 3227 1516 3533 1524
rect 3547 1516 3573 1524
rect 5907 1516 5973 1524
rect 347 1496 513 1504
rect 1427 1496 1673 1504
rect 1727 1496 1773 1504
rect 1827 1496 1944 1504
rect 367 1476 413 1484
rect 607 1476 733 1484
rect 1127 1476 1653 1484
rect 1936 1484 1944 1496
rect 1967 1496 2113 1504
rect 2167 1496 2413 1504
rect 3387 1496 3753 1504
rect 3767 1496 4033 1504
rect 4047 1496 4273 1504
rect 4447 1496 4553 1504
rect 4567 1496 4733 1504
rect 5167 1496 5233 1504
rect 5247 1496 5293 1504
rect 6007 1496 6053 1504
rect 1936 1476 2033 1484
rect 2187 1476 2353 1484
rect 2407 1476 2673 1484
rect 2867 1476 2933 1484
rect 2947 1476 2993 1484
rect 3076 1476 3333 1484
rect 827 1456 1033 1464
rect 1547 1456 1573 1464
rect 1787 1456 1833 1464
rect 2107 1456 2153 1464
rect 2567 1456 2664 1464
rect 247 1436 373 1444
rect 447 1444 460 1447
rect 447 1433 464 1444
rect 527 1437 553 1445
rect 647 1436 773 1444
rect 847 1437 873 1445
rect 927 1436 973 1444
rect 107 1396 213 1404
rect 227 1396 273 1404
rect 456 1406 464 1433
rect 567 1396 613 1404
rect 947 1396 993 1404
rect 1307 1396 1453 1404
rect 1476 1387 1484 1434
rect 1607 1436 1704 1444
rect 1516 1404 1524 1433
rect 1696 1406 1704 1436
rect 2187 1436 2253 1444
rect 1516 1396 1573 1404
rect 687 1376 1133 1384
rect 1476 1376 1493 1387
rect 1480 1373 1493 1376
rect 1756 1384 1764 1433
rect 1796 1404 1804 1433
rect 1956 1424 1964 1434
rect 2600 1444 2613 1447
rect 2367 1436 2613 1444
rect 2596 1433 2613 1436
rect 1936 1420 1964 1424
rect 1933 1416 1964 1420
rect 1933 1407 1947 1416
rect 1796 1396 1833 1404
rect 1956 1400 2013 1404
rect 1953 1396 2013 1400
rect 1727 1376 1764 1384
rect 1953 1387 1967 1396
rect 2093 1404 2107 1413
rect 2027 1400 2107 1404
rect 2027 1396 2104 1400
rect 2136 1396 2153 1404
rect 2136 1384 2144 1396
rect 2287 1396 2313 1404
rect 2367 1396 2473 1404
rect 2596 1406 2604 1433
rect 2656 1424 2664 1456
rect 3076 1464 3084 1476
rect 3387 1476 3413 1484
rect 3427 1476 3613 1484
rect 3867 1476 3953 1484
rect 5347 1476 5613 1484
rect 5627 1476 5793 1484
rect 6267 1476 6293 1484
rect 2867 1456 3084 1464
rect 3107 1456 3132 1464
rect 3167 1456 3284 1464
rect 2907 1436 2964 1444
rect 2656 1416 2724 1424
rect 2716 1404 2724 1416
rect 2716 1396 2733 1404
rect 2807 1396 2833 1404
rect 2956 1404 2964 1436
rect 3047 1436 3113 1444
rect 3187 1436 3253 1444
rect 3276 1444 3284 1456
rect 4247 1456 4313 1464
rect 4627 1456 4693 1464
rect 4947 1456 5153 1464
rect 5947 1456 6013 1464
rect 6107 1456 6153 1464
rect 3276 1436 3373 1444
rect 3446 1433 3447 1440
rect 3467 1437 3573 1445
rect 3707 1436 3733 1444
rect 3807 1436 3844 1444
rect 3116 1407 3124 1433
rect 3433 1424 3447 1433
rect 3396 1420 3447 1424
rect 3396 1416 3443 1420
rect 2956 1396 3013 1404
rect 3396 1406 3404 1416
rect 3227 1395 3313 1403
rect 3507 1395 3673 1403
rect 3836 1404 3844 1436
rect 3947 1436 3993 1444
rect 4167 1437 4193 1445
rect 4347 1436 4393 1444
rect 4036 1404 4044 1434
rect 4156 1424 4164 1434
rect 4547 1437 4573 1445
rect 4587 1436 4653 1444
rect 4436 1424 4444 1434
rect 4867 1437 4913 1445
rect 4927 1436 5033 1444
rect 5207 1436 5333 1444
rect 5387 1437 5433 1445
rect 5667 1436 5753 1444
rect 5813 1444 5827 1453
rect 5813 1440 5884 1444
rect 5816 1436 5884 1440
rect 4156 1416 4444 1424
rect 3836 1400 4044 1404
rect 4176 1400 4213 1404
rect 3836 1396 4047 1400
rect 4033 1387 4047 1396
rect 2087 1376 2144 1384
rect 2207 1376 2253 1384
rect 2507 1376 2693 1384
rect 2887 1376 2993 1384
rect 4173 1396 4213 1400
rect 4173 1387 4187 1396
rect 4307 1395 4353 1403
rect 4467 1396 4533 1404
rect 4707 1395 4753 1403
rect 4987 1395 5053 1403
rect 5307 1395 5353 1403
rect 5567 1396 5593 1404
rect 5647 1396 5773 1404
rect 4976 1384 4984 1392
rect 5733 1387 5747 1396
rect 5827 1396 5853 1404
rect 4927 1376 4984 1384
rect 5467 1376 5544 1384
rect 1307 1356 1533 1364
rect 1787 1356 1833 1364
rect 2007 1356 2053 1364
rect 2287 1356 2333 1364
rect 2587 1356 2653 1364
rect 2747 1356 2793 1364
rect 2807 1356 3144 1364
rect 607 1336 833 1344
rect 847 1336 953 1344
rect 1127 1336 1333 1344
rect 1427 1336 1473 1344
rect 1907 1336 1973 1344
rect 2027 1336 2353 1344
rect 3136 1344 3144 1356
rect 3167 1356 3453 1364
rect 4036 1364 4044 1373
rect 3767 1356 4044 1364
rect 4107 1356 4153 1364
rect 4167 1356 4313 1364
rect 5107 1356 5433 1364
rect 5447 1356 5473 1364
rect 5536 1364 5544 1376
rect 5876 1384 5884 1436
rect 5956 1387 5964 1434
rect 5996 1404 6004 1433
rect 6196 1407 6204 1433
rect 6296 1407 6304 1433
rect 5996 1396 6053 1404
rect 6107 1395 6153 1403
rect 5876 1376 5913 1384
rect 5536 1356 5633 1364
rect 5987 1356 6053 1364
rect 6147 1356 6193 1364
rect 6207 1356 6253 1364
rect 3136 1336 3284 1344
rect 767 1316 813 1324
rect 927 1316 1173 1324
rect 1187 1316 1533 1324
rect 2007 1316 2213 1324
rect 2307 1316 2373 1324
rect 2427 1316 2493 1324
rect 3127 1316 3153 1324
rect 3276 1324 3284 1336
rect 3687 1336 3733 1344
rect 3787 1336 3913 1344
rect 4427 1336 4573 1344
rect 4587 1336 4673 1344
rect 4996 1336 5384 1344
rect 4996 1327 5004 1336
rect 3276 1316 3293 1324
rect 3307 1316 3493 1324
rect 3567 1316 4313 1324
rect 4407 1316 4993 1324
rect 5376 1324 5384 1336
rect 5407 1336 5753 1344
rect 5767 1336 5853 1344
rect 6167 1336 6233 1344
rect 5376 1316 5453 1324
rect 5847 1316 5973 1324
rect 6087 1316 6113 1324
rect 1567 1296 1793 1304
rect 1947 1296 2233 1304
rect 2427 1296 2553 1304
rect 2727 1296 2893 1304
rect 3087 1296 3173 1304
rect 3347 1296 3393 1304
rect 3487 1296 3533 1304
rect 3747 1296 4133 1304
rect 4767 1296 4793 1304
rect 5227 1296 5513 1304
rect 5687 1296 5993 1304
rect 707 1276 1013 1284
rect 1507 1276 2633 1284
rect 2647 1276 3713 1284
rect 3727 1276 4353 1284
rect 4647 1276 5033 1284
rect 5547 1276 5773 1284
rect 5827 1276 5933 1284
rect 6127 1280 6183 1284
rect 6127 1276 6187 1280
rect 6173 1267 6187 1276
rect 6227 1276 6273 1284
rect 467 1256 653 1264
rect 747 1256 793 1264
rect 1087 1256 1173 1264
rect 1867 1256 1913 1264
rect 2047 1256 2213 1264
rect 2347 1256 2393 1264
rect 2447 1256 2613 1264
rect 2947 1256 3053 1264
rect 3107 1256 3133 1264
rect 3327 1256 3373 1264
rect 3387 1256 3493 1264
rect 3907 1256 3953 1264
rect 4007 1256 4173 1264
rect 4627 1256 4793 1264
rect 4947 1256 5133 1264
rect 5247 1256 5473 1264
rect 5687 1256 5833 1264
rect 6186 1260 6187 1267
rect 6207 1256 6293 1264
rect 167 1236 213 1244
rect 296 1236 413 1244
rect 47 1217 113 1225
rect 187 1216 224 1224
rect 216 1184 224 1216
rect 296 1186 304 1236
rect 856 1236 893 1244
rect 327 1217 353 1225
rect 527 1217 553 1225
rect 216 1176 253 1184
rect 367 1176 573 1184
rect 616 1167 624 1233
rect 696 1184 704 1214
rect 856 1186 864 1236
rect 1067 1236 1093 1244
rect 1627 1236 1693 1244
rect 1936 1236 2013 1244
rect 887 1217 973 1225
rect 1187 1217 1253 1225
rect 647 1176 704 1184
rect 907 1175 953 1183
rect 667 1156 753 1164
rect 1007 1156 1053 1164
rect 1136 1164 1144 1213
rect 1336 1184 1344 1214
rect 1496 1186 1504 1233
rect 1547 1216 1604 1224
rect 1596 1186 1604 1216
rect 1716 1187 1724 1213
rect 1227 1176 1344 1184
rect 1736 1186 1744 1233
rect 1767 1216 1784 1224
rect 1776 1204 1784 1216
rect 1807 1216 1913 1224
rect 1776 1200 1824 1204
rect 1776 1196 1827 1200
rect 1813 1187 1827 1196
rect 1936 1186 1944 1236
rect 2247 1236 2773 1244
rect 3367 1236 3433 1244
rect 3587 1236 3613 1244
rect 3747 1236 3833 1244
rect 3927 1236 4193 1244
rect 4247 1236 4293 1244
rect 4487 1236 4513 1244
rect 4776 1236 4833 1244
rect 1993 1204 2007 1213
rect 1993 1200 2024 1204
rect 1996 1196 2024 1200
rect 2016 1186 2024 1196
rect 2036 1167 2044 1214
rect 2127 1216 2173 1224
rect 2307 1216 2364 1224
rect 2076 1183 2084 1213
rect 2067 1175 2133 1183
rect 2267 1176 2293 1184
rect 2356 1186 2364 1216
rect 2387 1216 2404 1224
rect 2396 1187 2404 1216
rect 2467 1216 2544 1224
rect 2427 1196 2524 1204
rect 2516 1186 2524 1196
rect 2447 1175 2473 1183
rect 2536 1184 2544 1216
rect 2627 1216 2753 1224
rect 2867 1216 2964 1224
rect 2796 1187 2804 1213
rect 2536 1176 2633 1184
rect 2956 1186 2964 1216
rect 3027 1216 3093 1224
rect 3196 1216 3213 1224
rect 3136 1187 3144 1213
rect 3196 1187 3204 1216
rect 3307 1216 3364 1224
rect 1136 1156 1153 1164
rect 1167 1156 1332 1164
rect 1367 1156 1553 1164
rect 1667 1156 1833 1164
rect 867 1136 933 1144
rect 1047 1136 1233 1144
rect 1327 1136 1933 1144
rect 1987 1136 2473 1144
rect 2696 1144 2704 1173
rect 3356 1186 3364 1216
rect 3687 1216 3713 1224
rect 3767 1224 3780 1227
rect 3767 1213 3784 1224
rect 3867 1217 3913 1225
rect 3956 1216 3993 1224
rect 3287 1175 3313 1183
rect 3416 1184 3424 1213
rect 3776 1186 3784 1213
rect 3956 1204 3964 1216
rect 4047 1224 4060 1227
rect 4047 1213 4064 1224
rect 4260 1224 4273 1227
rect 4187 1216 4224 1224
rect 3936 1196 3964 1204
rect 3936 1186 3944 1196
rect 4056 1186 4064 1213
rect 4216 1186 4224 1216
rect 4256 1213 4273 1224
rect 4467 1217 4533 1225
rect 4776 1224 4784 1236
rect 4847 1236 4993 1244
rect 5007 1236 5084 1244
rect 4547 1216 4784 1224
rect 4807 1216 4873 1224
rect 5076 1224 5084 1236
rect 5427 1236 5453 1244
rect 5527 1236 5564 1244
rect 5076 1216 5093 1224
rect 5327 1217 5353 1225
rect 4256 1186 4264 1213
rect 5196 1204 5204 1214
rect 5507 1224 5520 1227
rect 5507 1213 5524 1224
rect 5196 1196 5293 1204
rect 3407 1176 3424 1184
rect 3527 1176 3613 1184
rect 3827 1175 3873 1183
rect 3987 1175 4013 1183
rect 4387 1176 4453 1184
rect 4567 1176 4613 1184
rect 4887 1175 4913 1183
rect 4967 1175 4992 1183
rect 5027 1180 5104 1184
rect 5027 1176 5107 1180
rect 3876 1164 3884 1172
rect 5093 1167 5107 1176
rect 5127 1176 5213 1184
rect 5347 1176 5433 1184
rect 5516 1186 5524 1213
rect 5556 1186 5564 1236
rect 5627 1236 5864 1244
rect 5587 1216 5704 1224
rect 5696 1204 5704 1216
rect 5696 1196 5824 1204
rect 5816 1186 5824 1196
rect 5856 1186 5864 1236
rect 5916 1187 5924 1213
rect 5956 1167 5964 1253
rect 6007 1216 6073 1224
rect 6140 1224 6153 1227
rect 6136 1213 6153 1224
rect 6136 1187 6144 1213
rect 6136 1176 6153 1187
rect 6140 1173 6153 1176
rect 6236 1167 6244 1214
rect 6327 1224 6340 1227
rect 6327 1213 6344 1224
rect 6336 1167 6344 1213
rect 3876 1156 4093 1164
rect 5707 1156 5733 1164
rect 5947 1156 5964 1167
rect 5947 1153 5960 1156
rect 6047 1156 6073 1164
rect 6327 1156 6344 1167
rect 6327 1153 6340 1156
rect 2607 1136 2704 1144
rect 2787 1136 2973 1144
rect 3027 1136 3233 1144
rect 3467 1136 3533 1144
rect 3587 1136 4593 1144
rect 4607 1136 4633 1144
rect 4887 1136 5013 1144
rect 5067 1136 5293 1144
rect 5307 1136 5373 1144
rect 5467 1136 5573 1144
rect 6187 1136 6253 1144
rect 107 1116 353 1124
rect 367 1116 493 1124
rect 587 1116 713 1124
rect 1267 1116 1453 1124
rect 1507 1116 2013 1124
rect 2127 1116 2313 1124
rect 2847 1116 2873 1124
rect 3047 1116 3113 1124
rect 4327 1116 4553 1124
rect 5567 1116 5713 1124
rect 5787 1116 5973 1124
rect 5987 1116 6093 1124
rect 1487 1096 1833 1104
rect 2147 1096 2793 1104
rect 2867 1096 2993 1104
rect 3567 1096 5173 1104
rect 5187 1096 5253 1104
rect 5267 1096 5313 1104
rect 147 1076 373 1084
rect 387 1076 533 1084
rect 827 1076 953 1084
rect 1347 1076 1453 1084
rect 1567 1076 1693 1084
rect 1907 1076 2033 1084
rect 2047 1076 2153 1084
rect 2267 1076 2413 1084
rect 2827 1076 3213 1084
rect 3227 1076 3693 1084
rect 4507 1076 5013 1084
rect 5387 1076 5744 1084
rect 287 1056 393 1064
rect 1027 1056 1173 1064
rect 1187 1056 1733 1064
rect 1867 1056 2193 1064
rect 2207 1056 3072 1064
rect 3107 1056 4484 1064
rect 267 1036 433 1044
rect 1307 1036 1333 1044
rect 1707 1036 2153 1044
rect 2247 1036 2273 1044
rect 2327 1036 2893 1044
rect 2987 1036 3393 1044
rect 4476 1044 4484 1056
rect 4687 1056 4953 1064
rect 5107 1056 5413 1064
rect 5736 1064 5744 1076
rect 5767 1076 6293 1084
rect 5736 1056 5833 1064
rect 4476 1036 4573 1044
rect 4987 1036 5353 1044
rect 5367 1036 5653 1044
rect 5667 1036 5893 1044
rect 807 1016 1233 1024
rect 1847 1016 2733 1024
rect 2747 1016 3293 1024
rect 5147 1016 5333 1024
rect 5447 1016 5533 1024
rect 6007 1016 6253 1024
rect 627 996 653 1004
rect 1367 996 1493 1004
rect 1647 996 1793 1004
rect 2287 996 2392 1004
rect 2427 996 3093 1004
rect 3207 996 3593 1004
rect 3727 996 3933 1004
rect 4187 996 4293 1004
rect 4487 996 4693 1004
rect 4767 996 5253 1004
rect 5267 996 5393 1004
rect 5407 996 5553 1004
rect 6067 996 6313 1004
rect 247 976 513 984
rect 527 976 713 984
rect 847 976 1253 984
rect 1327 976 1393 984
rect 1407 976 1544 984
rect 1536 967 1544 976
rect 2927 976 4593 984
rect 4607 976 4713 984
rect 4867 976 5213 984
rect 5227 976 5433 984
rect 5447 976 5593 984
rect 767 956 793 964
rect 807 956 873 964
rect 1547 956 1633 964
rect 1867 956 2053 964
rect 2147 956 2453 964
rect 2787 956 2813 964
rect 3187 956 3353 964
rect 3747 956 3913 964
rect 3927 956 3973 964
rect 5247 956 5373 964
rect 5627 956 5653 964
rect 5867 956 5913 964
rect 5927 956 6133 964
rect 647 936 973 944
rect 1167 936 1353 944
rect 1427 936 1673 944
rect 1847 936 2093 944
rect 2867 936 3533 944
rect 3547 936 3653 944
rect 4167 936 4253 944
rect 5507 936 5673 944
rect 5687 936 5773 944
rect 67 917 93 925
rect 147 916 213 924
rect 227 917 253 925
rect 316 916 333 924
rect 127 876 273 884
rect 316 867 324 916
rect 347 916 473 924
rect 767 916 833 924
rect 1013 924 1027 933
rect 996 920 1027 924
rect 996 916 1024 920
rect 367 876 453 884
rect 747 876 853 884
rect 907 876 933 884
rect 996 886 1004 916
rect 1047 917 1113 925
rect 1456 904 1464 914
rect 1367 896 1513 904
rect 1067 876 1213 884
rect 1227 876 1273 884
rect 1556 884 1564 913
rect 1487 876 1564 884
rect 1596 867 1604 914
rect 1656 884 1664 913
rect 1716 904 1724 933
rect 2007 916 2093 924
rect 2107 916 2213 924
rect 2240 924 2253 927
rect 2236 913 2253 924
rect 2367 917 2433 925
rect 2507 916 2544 924
rect 2236 904 2244 913
rect 1716 896 1764 904
rect 2176 900 2244 904
rect 1627 876 1664 884
rect 1687 875 1733 883
rect 1756 884 1764 896
rect 2173 896 2244 900
rect 2536 904 2544 916
rect 2567 917 2613 925
rect 2907 916 3133 924
rect 3147 916 3173 924
rect 3187 916 3313 924
rect 3367 916 3493 924
rect 3707 916 3793 924
rect 3847 916 3884 924
rect 3876 904 3884 916
rect 3907 916 4004 924
rect 2536 896 2664 904
rect 3876 900 3964 904
rect 3876 896 3967 900
rect 2173 887 2187 896
rect 1756 876 1773 884
rect 2047 876 2133 884
rect 2656 886 2664 896
rect 3953 887 3967 896
rect 2807 875 2853 883
rect 3007 875 3193 883
rect 3207 876 3333 884
rect 3447 875 3473 883
rect 3487 876 3633 884
rect 3867 875 3913 883
rect 3996 886 4004 916
rect 4107 917 4133 925
rect 4147 916 4333 924
rect 4407 917 4453 925
rect 4647 916 4773 924
rect 4827 916 4913 924
rect 4927 916 4944 924
rect 4496 904 4504 914
rect 4427 896 4504 904
rect 4936 887 4944 916
rect 5067 916 5133 924
rect 5160 924 5173 927
rect 5156 913 5173 924
rect 4167 876 4253 884
rect 4267 875 4313 883
rect 1347 856 1413 864
rect 2307 856 2333 864
rect 2487 856 2613 864
rect 2887 856 2913 864
rect 3116 856 3793 864
rect 1096 836 1493 844
rect 1096 827 1104 836
rect 1827 836 2173 844
rect 3116 844 3124 856
rect 4373 864 4387 873
rect 4567 875 4653 883
rect 4667 876 4753 884
rect 5156 886 5164 913
rect 5236 887 5244 913
rect 5047 875 5093 883
rect 5296 884 5304 914
rect 5347 916 5404 924
rect 5296 876 5333 884
rect 5396 884 5404 916
rect 5547 916 5624 924
rect 5396 876 5413 884
rect 5467 876 5493 884
rect 5616 867 5624 916
rect 5987 917 6033 925
rect 6096 916 6213 924
rect 5696 887 5704 913
rect 4227 860 4387 864
rect 4227 856 4384 860
rect 5856 864 5864 913
rect 5936 887 5944 914
rect 5936 876 5953 887
rect 5940 873 5953 876
rect 6096 886 6104 916
rect 6307 916 6344 924
rect 6027 875 6053 883
rect 6287 876 6313 884
rect 5767 856 5864 864
rect 6167 856 6213 864
rect 6336 864 6344 916
rect 6307 856 6344 864
rect 2467 836 3124 844
rect 3147 836 3173 844
rect 3387 836 3664 844
rect 67 816 193 824
rect 207 816 413 824
rect 607 816 713 824
rect 727 816 1093 824
rect 1547 816 1773 824
rect 1907 816 2293 824
rect 2587 816 3072 824
rect 3107 816 3413 824
rect 3656 824 3664 836
rect 3687 836 4093 844
rect 4207 836 4393 844
rect 4467 836 4593 844
rect 4767 836 4853 844
rect 4907 836 4993 844
rect 5487 836 5713 844
rect 6187 836 6233 844
rect 3656 816 3893 824
rect 4527 816 5333 824
rect 5387 816 5413 824
rect 5427 816 5573 824
rect 5647 816 5873 824
rect 5887 816 5913 824
rect 6007 816 6253 824
rect 1047 796 1353 804
rect 1407 796 1573 804
rect 1647 796 1733 804
rect 2207 796 2273 804
rect 2327 796 2373 804
rect 2447 796 2753 804
rect 2856 796 3193 804
rect 707 776 1073 784
rect 1367 776 1593 784
rect 1607 776 1753 784
rect 1767 776 1893 784
rect 1947 776 2013 784
rect 2087 776 2113 784
rect 2856 784 2864 796
rect 3347 796 4253 804
rect 4727 796 4893 804
rect 4947 796 5073 804
rect 5336 804 5344 813
rect 5336 796 5953 804
rect 2427 776 2864 784
rect 4967 776 5093 784
rect 5327 776 5393 784
rect 5567 776 5653 784
rect 5956 784 5964 793
rect 5956 776 6133 784
rect 347 756 733 764
rect 947 756 1333 764
rect 1627 756 1693 764
rect 1787 756 1913 764
rect 1987 756 2133 764
rect 2147 756 2233 764
rect 2387 756 2873 764
rect 2927 756 3213 764
rect 3607 756 3973 764
rect 3987 756 4073 764
rect 4296 756 4413 764
rect 4296 747 4304 756
rect 4427 756 4453 764
rect 4527 756 4873 764
rect 5027 756 5533 764
rect 5867 756 6073 764
rect 267 736 453 744
rect 547 736 593 744
rect 1107 736 1153 744
rect 1207 736 1433 744
rect 1447 736 1932 744
rect 1967 736 2253 744
rect 2607 736 2913 744
rect 3287 736 3492 744
rect 3527 736 3773 744
rect 3967 736 4293 744
rect 4387 736 4653 744
rect 4667 736 4713 744
rect 5287 736 5373 744
rect 5627 736 5893 744
rect 347 716 373 724
rect 1467 716 1533 724
rect 1767 724 1780 727
rect 1767 713 1784 724
rect 2127 716 2413 724
rect 2967 716 3113 724
rect 3247 716 3713 724
rect 3727 716 3813 724
rect 3827 716 3853 724
rect 4276 716 4333 724
rect 147 696 173 704
rect 287 696 404 704
rect 47 656 73 664
rect 87 656 213 664
rect 327 655 373 663
rect 396 664 404 696
rect 447 697 473 705
rect 607 696 653 704
rect 787 697 833 705
rect 936 696 993 704
rect 396 656 613 664
rect 936 664 944 696
rect 1167 697 1233 705
rect 1416 696 1593 704
rect 827 656 944 664
rect 1027 655 1073 663
rect 1187 656 1273 664
rect 1316 647 1324 694
rect 1416 687 1424 696
rect 1647 696 1713 704
rect 1407 676 1424 687
rect 1407 673 1420 676
rect 1776 666 1784 713
rect 1816 666 1824 713
rect 1993 704 2007 713
rect 1947 700 2007 704
rect 1947 696 2004 700
rect 2096 684 2104 694
rect 2267 696 2333 704
rect 2587 697 2653 705
rect 2747 697 2793 705
rect 2816 696 2833 704
rect 1867 676 2104 684
rect 1427 656 1653 664
rect 1827 656 1913 664
rect 2007 655 2153 663
rect 2176 664 2184 693
rect 2816 684 2824 696
rect 2847 696 3013 704
rect 3127 696 3373 704
rect 3427 697 3473 705
rect 3487 696 3553 704
rect 3647 696 3673 704
rect 3907 696 3924 704
rect 2727 676 2824 684
rect 3696 676 3804 684
rect 2176 656 2213 664
rect 2307 655 2353 663
rect 2487 656 2673 664
rect 2687 656 2732 664
rect 3696 666 3704 676
rect 3796 666 3804 676
rect 3916 667 3924 696
rect 3947 697 4013 705
rect 4027 696 4124 704
rect 2767 656 2813 664
rect 2827 655 2873 663
rect 2987 655 3013 663
rect 3027 656 3093 664
rect 3407 656 3533 664
rect 3747 655 3772 663
rect 3807 655 3833 663
rect 4116 666 4124 696
rect 4147 696 4204 704
rect 4196 667 4204 696
rect 4196 656 4213 667
rect 4200 653 4213 656
rect 4276 666 4284 716
rect 4347 716 4744 724
rect 4316 696 4413 704
rect 4316 667 4324 696
rect 4476 696 4553 704
rect 4347 676 4424 684
rect 4416 664 4424 676
rect 4476 667 4484 696
rect 4607 696 4704 704
rect 4696 667 4704 696
rect 4416 656 4433 664
rect 4627 655 4653 663
rect 4736 666 4744 716
rect 4927 716 4973 724
rect 5316 716 5353 724
rect 5007 704 5020 707
rect 5007 693 5024 704
rect 5047 696 5113 704
rect 5136 696 5173 704
rect 5016 666 5024 693
rect 4827 655 4893 663
rect 5067 655 5093 663
rect 767 636 893 644
rect 4180 644 4193 647
rect 4047 636 4193 644
rect 4176 633 4193 636
rect 5136 646 5144 696
rect 5247 697 5293 705
rect 5316 666 5324 716
rect 5427 716 5473 724
rect 5947 716 6273 724
rect 5347 696 5364 704
rect 5356 647 5364 696
rect 5456 696 5513 704
rect 5456 666 5464 696
rect 5527 697 5593 705
rect 5607 696 5793 704
rect 5887 696 5913 704
rect 5676 676 5733 684
rect 5547 655 5573 663
rect 5676 664 5684 676
rect 5587 656 5684 664
rect 5827 656 5893 664
rect 267 616 473 624
rect 487 616 693 624
rect 1187 616 1233 624
rect 1247 616 1293 624
rect 1727 616 2033 624
rect 2167 616 2193 624
rect 2207 616 2232 624
rect 2267 616 2473 624
rect 3207 616 3293 624
rect 3307 616 3433 624
rect 3447 616 3673 624
rect 4087 616 4153 624
rect 4176 624 4184 633
rect 5347 636 5364 647
rect 5347 633 5360 636
rect 5487 636 5553 644
rect 5707 636 5773 644
rect 4176 616 4393 624
rect 4707 616 4773 624
rect 4827 616 4973 624
rect 4987 616 5113 624
rect 5947 616 6173 624
rect 607 596 773 604
rect 787 596 973 604
rect 1367 596 1473 604
rect 1647 596 1853 604
rect 2107 596 2513 604
rect 2527 596 2573 604
rect 2587 596 2773 604
rect 2827 596 3164 604
rect 467 576 1133 584
rect 1147 576 1313 584
rect 2247 576 2393 584
rect 3156 584 3164 596
rect 3547 596 3573 604
rect 3156 576 3173 584
rect 3187 576 3253 584
rect 3727 576 3913 584
rect 4067 576 4493 584
rect 4507 576 4573 584
rect 4687 576 4933 584
rect 5107 576 5193 584
rect 5267 576 5353 584
rect 5756 576 6113 584
rect 127 556 413 564
rect 427 556 513 564
rect 787 556 813 564
rect 887 556 1093 564
rect 1547 556 1873 564
rect 2127 556 2813 564
rect 2947 556 3133 564
rect 3147 556 3473 564
rect 5756 564 5764 576
rect 5327 556 5764 564
rect 627 536 984 544
rect 976 527 984 536
rect 2867 536 3033 544
rect 3647 536 3953 544
rect 987 516 1133 524
rect 2147 516 2833 524
rect 2907 516 3393 524
rect 3687 516 3773 524
rect 4087 516 4693 524
rect 4807 516 5613 524
rect 527 496 873 504
rect 1207 496 1413 504
rect 2567 496 2753 504
rect 2867 496 3493 504
rect 3567 496 3873 504
rect 4007 496 4033 504
rect 4116 496 5513 504
rect 287 476 333 484
rect 487 476 853 484
rect 947 476 1173 484
rect 1236 476 1784 484
rect 1236 464 1244 476
rect 1107 456 1244 464
rect 1776 464 1784 476
rect 1807 476 2724 484
rect 2716 467 2724 476
rect 4116 484 4124 496
rect 5947 496 6193 504
rect 3687 476 4124 484
rect 4147 476 4273 484
rect 4696 476 5693 484
rect 1776 456 2213 464
rect 2287 456 2313 464
rect 2327 456 2373 464
rect 2727 456 2953 464
rect 2967 456 3033 464
rect 4696 464 4704 476
rect 3947 456 4704 464
rect 5767 456 6013 464
rect 407 436 693 444
rect 707 436 832 444
rect 867 436 1033 444
rect 1087 436 1193 444
rect 1407 436 1453 444
rect 1467 436 1653 444
rect 2247 436 2453 444
rect 2467 436 2613 444
rect 3187 436 3573 444
rect 4347 436 4473 444
rect 4567 436 4713 444
rect 4727 436 5133 444
rect 1707 416 1953 424
rect 1967 416 2013 424
rect 2027 416 2113 424
rect 2127 416 2213 424
rect 2316 416 2384 424
rect 167 397 353 405
rect 416 396 513 404
rect 396 384 404 394
rect 296 380 404 384
rect 293 376 404 380
rect 293 367 307 376
rect 416 366 424 396
rect 647 397 733 405
rect 556 364 564 394
rect 507 356 564 364
rect 587 356 613 364
rect 727 356 773 364
rect 936 364 944 393
rect 1087 396 1173 404
rect 1187 396 1213 404
rect 1327 396 1353 404
rect 1276 367 1284 394
rect 867 356 944 364
rect 1007 355 1073 363
rect 1167 356 1193 364
rect 1267 356 1284 367
rect 1267 353 1280 356
rect 127 336 213 344
rect 227 336 313 344
rect 807 336 984 344
rect 267 316 333 324
rect 447 316 493 324
rect 507 316 953 324
rect 976 324 984 336
rect 1247 336 1293 344
rect 976 316 1193 324
rect 1316 324 1324 394
rect 1507 396 1533 404
rect 1547 397 1573 405
rect 1627 396 1653 404
rect 1747 397 1813 405
rect 1836 396 1853 404
rect 1413 384 1427 393
rect 1413 380 1444 384
rect 1416 376 1444 380
rect 1436 366 1444 376
rect 1836 367 1844 396
rect 1907 396 1933 404
rect 2187 397 2273 405
rect 2316 404 2324 416
rect 2296 396 2324 404
rect 1347 355 1373 363
rect 1647 356 1753 364
rect 2076 364 2084 393
rect 2136 367 2144 393
rect 2296 384 2304 396
rect 2376 404 2384 416
rect 3147 416 3713 424
rect 4187 416 4213 424
rect 4227 416 4313 424
rect 5287 416 5413 424
rect 5727 416 5793 424
rect 6067 416 6133 424
rect 6147 416 6233 424
rect 2376 396 2464 404
rect 2276 380 2304 384
rect 2273 376 2304 380
rect 2273 367 2287 376
rect 2027 356 2084 364
rect 2207 356 2252 364
rect 2356 364 2364 394
rect 2456 384 2464 396
rect 2507 397 2553 405
rect 2667 397 2693 405
rect 2836 396 2913 404
rect 2456 376 2484 384
rect 2356 356 2433 364
rect 2476 364 2484 376
rect 2796 384 2804 394
rect 2836 384 2844 396
rect 2927 397 2992 405
rect 3027 397 3073 405
rect 3207 397 3253 405
rect 3267 396 3393 404
rect 3447 396 3533 404
rect 3547 396 3693 404
rect 3767 397 3833 405
rect 3967 397 4133 405
rect 4447 397 4493 405
rect 4607 397 4673 405
rect 4767 396 4913 404
rect 4927 396 4993 404
rect 5067 397 5093 405
rect 5247 396 5373 404
rect 5647 397 5733 405
rect 2727 376 2804 384
rect 2816 376 2844 384
rect 2476 356 2513 364
rect 2567 356 2633 364
rect 2707 356 2773 364
rect 2816 364 2824 376
rect 2796 360 2824 364
rect 2793 356 2824 360
rect 1376 344 1384 352
rect 2793 347 2807 356
rect 2867 355 2933 363
rect 2947 356 3012 364
rect 3047 355 3093 363
rect 3116 347 3124 393
rect 3187 355 3233 363
rect 3287 360 3324 364
rect 3287 356 3327 360
rect 3313 347 3327 356
rect 3427 356 3473 364
rect 3527 356 3633 364
rect 3787 355 3813 363
rect 3867 356 3933 364
rect 4027 355 4073 363
rect 4227 355 4293 363
rect 4396 364 4404 394
rect 5556 384 5564 394
rect 5867 396 5913 404
rect 5456 376 5564 384
rect 5696 376 5773 384
rect 4396 356 4533 364
rect 4587 355 4633 363
rect 4647 356 4733 364
rect 4827 355 4893 363
rect 4967 355 5013 363
rect 5267 355 5333 363
rect 1376 336 1593 344
rect 2127 336 2293 344
rect 3507 336 3553 344
rect 5456 344 5464 376
rect 5487 356 5533 364
rect 5696 364 5704 376
rect 5816 367 5824 393
rect 5687 356 5704 364
rect 5727 355 5753 363
rect 5996 344 6004 394
rect 6087 356 6113 364
rect 5387 336 5464 344
rect 5656 336 6033 344
rect 5656 327 5664 336
rect 6176 344 6184 394
rect 6047 336 6184 344
rect 1207 316 1324 324
rect 1487 316 1653 324
rect 1827 316 1873 324
rect 1927 316 2093 324
rect 2407 316 2593 324
rect 2827 316 3653 324
rect 4167 316 4353 324
rect 4547 316 4692 324
rect 4727 316 4853 324
rect 5127 316 5653 324
rect 5807 316 5873 324
rect 6147 316 6253 324
rect 387 296 473 304
rect 687 296 813 304
rect 827 296 1113 304
rect 1907 296 2433 304
rect 2507 296 2793 304
rect 3107 296 3193 304
rect 3207 296 3684 304
rect 407 276 453 284
rect 1327 276 1453 284
rect 1887 276 2393 284
rect 2407 276 2813 284
rect 3247 276 3373 284
rect 3676 284 3684 296
rect 3807 296 3973 304
rect 4507 296 4672 304
rect 4696 304 4704 313
rect 4696 296 5052 304
rect 5087 296 5413 304
rect 5547 296 5633 304
rect 5687 296 5973 304
rect 3467 276 3624 284
rect 3676 276 3753 284
rect 167 256 513 264
rect 867 256 913 264
rect 927 256 1473 264
rect 1536 256 1713 264
rect 1536 247 1544 256
rect 1727 256 1833 264
rect 2027 256 2213 264
rect 2227 256 2373 264
rect 2487 256 2693 264
rect 2807 256 2833 264
rect 3616 264 3624 276
rect 4607 276 6013 284
rect 6027 276 6093 284
rect 6107 276 6153 284
rect 3207 256 3604 264
rect 3616 256 3733 264
rect 627 236 813 244
rect 1147 236 1393 244
rect 1536 244 1553 247
rect 1467 236 1553 244
rect 1540 233 1553 236
rect 1976 236 2713 244
rect 1976 227 1984 236
rect 2727 236 3113 244
rect 3247 236 3453 244
rect 3596 244 3604 256
rect 3847 256 3913 264
rect 4007 256 4053 264
rect 4127 256 4273 264
rect 4827 256 5433 264
rect 5587 256 5673 264
rect 3596 236 3752 244
rect 3787 236 4324 244
rect 4316 227 4324 236
rect 4927 236 5033 244
rect 5047 236 5173 244
rect 5187 236 5833 244
rect 1127 216 1253 224
rect 1587 216 1653 224
rect 1767 216 1833 224
rect 1927 216 1973 224
rect 2087 216 2153 224
rect 2387 216 2413 224
rect 2467 216 2513 224
rect 2647 216 2973 224
rect 3147 216 3513 224
rect 3947 216 4193 224
rect 4327 216 4413 224
rect 4647 216 4713 224
rect 4727 216 4793 224
rect 6116 216 6213 224
rect 767 196 1333 204
rect 1727 196 1953 204
rect 2016 196 2053 204
rect 127 177 193 185
rect 267 176 353 184
rect 447 176 564 184
rect 207 136 233 144
rect 287 136 333 144
rect 467 136 513 144
rect 556 146 564 176
rect 587 177 633 185
rect 836 176 853 184
rect 596 156 653 164
rect 596 146 604 156
rect 716 144 724 174
rect 736 156 793 164
rect 736 146 744 156
rect 836 147 844 176
rect 876 176 993 184
rect 687 136 724 144
rect 876 146 884 176
rect 1007 176 1113 184
rect 1227 177 1273 185
rect 1367 177 1413 185
rect 1467 176 1513 184
rect 1027 136 1093 144
rect 1147 136 1193 144
rect 1556 146 1564 193
rect 1627 176 1733 184
rect 1807 184 1820 187
rect 1807 173 1824 184
rect 2016 184 2024 196
rect 2587 196 3113 204
rect 3567 196 3693 204
rect 3707 196 4253 204
rect 4487 196 4513 204
rect 5176 196 5213 204
rect 1947 176 2024 184
rect 2036 176 2133 184
rect 1307 136 1393 144
rect 1667 136 1693 144
rect 1707 136 1773 144
rect 1816 146 1824 173
rect 1856 156 1913 164
rect 1856 146 1864 156
rect 2036 146 2044 176
rect 2187 176 2284 184
rect 2276 146 2284 176
rect 2480 184 2493 187
rect 2407 176 2444 184
rect 2436 146 2444 176
rect 2476 173 2493 184
rect 2627 177 2672 185
rect 2707 177 2753 185
rect 2947 177 2993 185
rect 3067 177 3132 185
rect 3167 177 3373 185
rect 3427 176 3464 184
rect 2476 146 2484 173
rect 3456 164 3464 176
rect 3487 176 3513 184
rect 3627 176 3653 184
rect 3767 177 3873 185
rect 3887 176 4033 184
rect 4047 176 4144 184
rect 4136 164 4144 176
rect 4167 176 4233 184
rect 4353 184 4367 193
rect 4287 176 4344 184
rect 4353 180 4453 184
rect 4356 176 4453 180
rect 3456 156 3544 164
rect 2127 135 2213 143
rect 3536 146 3544 156
rect 3576 156 3784 164
rect 4136 156 4184 164
rect 3576 146 3584 156
rect 3776 146 3784 156
rect 4176 146 4184 156
rect 4336 146 4344 176
rect 4767 176 4833 184
rect 4887 176 5113 184
rect 5176 164 5184 196
rect 6116 204 6124 216
rect 5967 196 6124 204
rect 5287 177 5333 185
rect 5347 176 5493 184
rect 6187 177 6233 185
rect 5016 156 5184 164
rect 5016 146 5024 156
rect 2687 136 2733 144
rect 2747 135 2873 143
rect 2967 135 3133 143
rect 3196 136 3213 144
rect 107 116 173 124
rect 1247 116 1473 124
rect 2527 116 3153 124
rect 3196 124 3204 136
rect 3267 135 3313 143
rect 3787 135 3813 143
rect 3867 136 4013 144
rect 4027 135 4073 143
rect 4267 135 4293 143
rect 4487 135 4533 143
rect 4587 136 4893 144
rect 4947 136 5013 144
rect 5176 144 5184 156
rect 5607 156 5784 164
rect 5167 136 5184 144
rect 5327 136 5453 144
rect 5776 146 5784 156
rect 6047 135 6073 143
rect 6127 136 6213 144
rect 3167 116 3204 124
rect 3367 116 3453 124
rect 3547 116 3673 124
rect 3687 116 4133 124
rect 4416 116 4773 124
rect 247 96 673 104
rect 827 96 1213 104
rect 1227 96 1433 104
rect 1607 96 2073 104
rect 2127 96 2233 104
rect 2287 96 2853 104
rect 2927 96 3053 104
rect 3147 96 3273 104
rect 3387 96 3473 104
rect 3727 96 3933 104
rect 4416 104 4424 116
rect 4787 116 5053 124
rect 5067 116 5193 124
rect 5367 116 5473 124
rect 5487 116 5633 124
rect 5647 116 5713 124
rect 4247 96 4424 104
rect 4447 96 4573 104
rect 4627 96 4733 104
rect 4747 96 4813 104
rect 5527 96 5593 104
rect 5987 96 6293 104
rect 367 76 913 84
rect 1487 76 1573 84
rect 1627 76 1993 84
rect 2367 76 2893 84
rect 4467 76 4513 84
rect 5127 76 5313 84
rect 707 56 833 64
rect 1267 56 1373 64
rect 1387 56 1453 64
rect 1507 56 1553 64
rect 1647 56 1973 64
rect 2027 56 2193 64
rect 2247 56 2313 64
rect 2407 56 2593 64
rect 2607 56 2773 64
rect 3007 56 3033 64
rect 3047 56 4093 64
rect 5427 56 5813 64
rect 5827 56 6173 64
rect 1107 36 1353 44
rect 1407 36 1753 44
rect 2647 36 2693 44
rect 2707 36 2893 44
rect 3067 36 3373 44
rect 3427 36 3913 44
rect 4847 36 5273 44
rect 5947 36 6273 44
rect 2927 16 3393 24
rect 3447 16 3613 24
use INVX1  _889_
timestamp 0
transform -1 0 4050 0 1 5470
box -6 -8 46 268
use NOR2X1  _890_
timestamp 0
transform 1 0 3570 0 -1 5990
box -6 -8 66 268
use NAND2X1  _891_
timestamp 0
transform -1 0 4770 0 1 5470
box -6 -8 66 268
use INVX1  _892_
timestamp 0
transform 1 0 4990 0 1 5470
box -6 -8 46 268
use INVX1  _893_
timestamp 0
transform -1 0 3730 0 -1 5990
box -6 -8 46 268
use INVX2  _894_
timestamp 0
transform -1 0 4850 0 1 4950
box -6 -8 46 268
use NOR2X1  _895_
timestamp 0
transform -1 0 3930 0 1 5470
box -6 -8 66 268
use NAND2X1  _896_
timestamp 0
transform 1 0 3750 0 1 5470
box -6 -8 66 268
use INVX1  _897_
timestamp 0
transform 1 0 5610 0 -1 5990
box -6 -8 46 268
use NOR2X1  _898_
timestamp 0
transform -1 0 4170 0 1 5470
box -6 -8 66 268
use AOI21X1  _899_
timestamp 0
transform 1 0 5110 0 1 5470
box -6 -8 86 268
use NOR2X1  _900_
timestamp 0
transform -1 0 6190 0 1 5990
box -6 -8 66 268
use OAI21X1  _901_
timestamp 0
transform 1 0 5970 0 1 5990
box -6 -8 86 268
use INVX1  _902_
timestamp 0
transform -1 0 5630 0 1 5990
box -6 -8 46 268
use INVX4  _903_
timestamp 0
transform 1 0 4690 0 -1 5470
box -6 -8 66 268
use OAI21X1  _904_
timestamp 0
transform -1 0 4170 0 -1 5990
box -6 -8 86 268
use INVX1  _905_
timestamp 0
transform -1 0 5350 0 -1 5990
box -6 -8 46 268
use NOR2X1  _906_
timestamp 0
transform 1 0 4910 0 1 4950
box -6 -8 66 268
use INVX1  _907_
timestamp 0
transform -1 0 3170 0 1 5470
box -6 -8 46 268
use INVX1  _908_
timestamp 0
transform -1 0 6290 0 1 5990
box -6 -8 46 268
use OAI21X1  _909_
timestamp 0
transform 1 0 5870 0 1 5470
box -6 -8 86 268
use OAI21X1  _910_
timestamp 0
transform -1 0 5090 0 -1 5990
box -6 -8 86 268
use AOI22X1  _911_
timestamp 0
transform 1 0 4830 0 -1 5990
box -6 -8 106 268
use NAND2X1  _912_
timestamp 0
transform 1 0 4710 0 -1 5990
box -6 -8 66 268
use OAI21X1  _913_
timestamp 0
transform 1 0 5710 0 1 5990
box -6 -8 86 268
use OAI21X1  _914_
timestamp 0
transform -1 0 5510 0 1 5990
box -6 -8 86 268
use NAND2X1  _915_
timestamp 0
transform 1 0 4310 0 -1 5470
box -6 -8 66 268
use NOR2X1  _916_
timestamp 0
transform 1 0 5850 0 1 5990
box -6 -8 66 268
use NOR2X1  _917_
timestamp 0
transform 1 0 6070 0 -1 5990
box -6 -8 66 268
use OAI22X1  _918_
timestamp 0
transform -1 0 5530 0 -1 5990
box -6 -8 106 268
use OR2X2  _919_
timestamp 0
transform -1 0 5370 0 1 5990
box -6 -8 86 268
use INVX1  _920_
timestamp 0
transform -1 0 6070 0 1 5470
box -6 -8 46 268
use AOI22X1  _921_
timestamp 0
transform -1 0 5990 0 -1 5990
box -6 -8 106 268
use NAND3X1  _922_
timestamp 0
transform 1 0 5150 0 -1 5990
box -6 -8 86 268
use AND2X2  _923_
timestamp 0
transform -1 0 5810 0 -1 5990
box -6 -8 86 268
use OAI21X1  _924_
timestamp 0
transform -1 0 5790 0 1 5470
box -6 -8 86 268
use INVX8  _925_
timestamp 0
transform -1 0 2970 0 -1 5990
box -6 -8 106 268
use INVX1  _926_
timestamp 0
transform 1 0 2030 0 -1 3910
box -6 -8 46 268
use NAND2X1  _927_
timestamp 0
transform -1 0 2470 0 1 3910
box -6 -8 66 268
use OAI21X1  _928_
timestamp 0
transform -1 0 2830 0 -1 3910
box -6 -8 86 268
use INVX1  _929_
timestamp 0
transform 1 0 1230 0 1 2870
box -6 -8 46 268
use NAND2X1  _930_
timestamp 0
transform -1 0 2210 0 -1 3390
box -6 -8 66 268
use OAI21X1  _931_
timestamp 0
transform -1 0 2370 0 -1 3390
box -6 -8 86 268
use INVX1  _932_
timestamp 0
transform 1 0 3910 0 1 4430
box -6 -8 46 268
use NAND2X1  _933_
timestamp 0
transform 1 0 4330 0 -1 4430
box -6 -8 66 268
use OAI21X1  _934_
timestamp 0
transform 1 0 4030 0 1 4430
box -6 -8 86 268
use INVX1  _935_
timestamp 0
transform 1 0 1070 0 1 4430
box -6 -8 46 268
use NAND2X1  _936_
timestamp 0
transform 1 0 2030 0 -1 4950
box -6 -8 66 268
use OAI21X1  _937_
timestamp 0
transform -1 0 2130 0 1 4430
box -6 -8 86 268
use INVX1  _938_
timestamp 0
transform -1 0 130 0 -1 3910
box -6 -8 46 268
use NAND2X1  _939_
timestamp 0
transform 1 0 3310 0 -1 4430
box -6 -8 66 268
use OAI21X1  _940_
timestamp 0
transform -1 0 3510 0 -1 4430
box -6 -8 86 268
use INVX1  _941_
timestamp 0
transform 1 0 1910 0 1 3910
box -6 -8 46 268
use NAND2X1  _942_
timestamp 0
transform -1 0 2210 0 1 3910
box -6 -8 66 268
use OAI21X1  _943_
timestamp 0
transform -1 0 2350 0 1 3910
box -6 -8 86 268
use INVX1  _944_
timestamp 0
transform -1 0 2950 0 -1 5470
box -6 -8 46 268
use NAND2X1  _945_
timestamp 0
transform -1 0 2750 0 1 4950
box -6 -8 66 268
use OAI21X1  _946_
timestamp 0
transform -1 0 2910 0 1 4950
box -6 -8 86 268
use INVX4  _947_
timestamp 0
transform 1 0 3910 0 -1 4950
box -6 -8 66 268
use NAND2X1  _948_
timestamp 0
transform 1 0 4250 0 1 4950
box -6 -8 66 268
use OAI21X1  _949_
timestamp 0
transform 1 0 4390 0 1 4950
box -6 -8 86 268
use INVX1  _950_
timestamp 0
transform -1 0 4010 0 -1 5990
box -6 -8 46 268
use INVX1  _951_
timestamp 0
transform 1 0 950 0 1 1830
box -6 -8 46 268
use INVX2  _952_
timestamp 0
transform -1 0 2590 0 1 2870
box -6 -8 46 268
use NOR2X1  _953_
timestamp 0
transform 1 0 1610 0 -1 1830
box -6 -8 66 268
use AND2X2  _954_
timestamp 0
transform -1 0 1970 0 -1 1830
box -6 -8 86 268
use NAND2X1  _955_
timestamp 0
transform -1 0 1810 0 -1 1830
box -6 -8 66 268
use NAND2X1  _956_
timestamp 0
transform -1 0 730 0 1 1830
box -6 -8 66 268
use NAND2X1  _957_
timestamp 0
transform 1 0 510 0 -1 2350
box -6 -8 66 268
use OR2X2  _958_
timestamp 0
transform -1 0 610 0 -1 1830
box -6 -8 86 268
use NAND2X1  _959_
timestamp 0
transform -1 0 250 0 1 1310
box -6 -8 66 268
use AND2X2  _960_
timestamp 0
transform 1 0 90 0 -1 2350
box -6 -8 86 268
use OAI21X1  _961_
timestamp 0
transform 1 0 230 0 -1 1830
box -6 -8 86 268
use NAND2X1  _962_
timestamp 0
transform -1 0 390 0 1 1310
box -6 -8 66 268
use INVX1  _963_
timestamp 0
transform -1 0 130 0 1 270
box -6 -8 46 268
use NAND2X1  _964_
timestamp 0
transform 1 0 590 0 1 1310
box -6 -8 66 268
use NAND2X1  _965_
timestamp 0
transform 1 0 1030 0 1 1310
box -6 -8 66 268
use OR2X2  _966_
timestamp 0
transform -1 0 630 0 1 790
box -6 -8 86 268
use INVX1  _967_
timestamp 0
transform -1 0 890 0 -1 1830
box -6 -8 46 268
use INVX1  _968_
timestamp 0
transform -1 0 2810 0 -1 1830
box -6 -8 46 268
use OAI21X1  _969_
timestamp 0
transform 1 0 450 0 1 1310
box -6 -8 86 268
use NAND3X1  _970_
timestamp 0
transform 1 0 90 0 -1 1310
box -6 -8 86 268
use NOR2X1  _971_
timestamp 0
transform 1 0 670 0 -1 790
box -6 -8 66 268
use AND2X2  _972_
timestamp 0
transform -1 0 590 0 -1 790
box -6 -8 86 268
use OAI21X1  _973_
timestamp 0
transform -1 0 450 0 -1 790
box -6 -8 86 268
use NAND3X1  _974_
timestamp 0
transform 1 0 390 0 -1 1310
box -6 -8 86 268
use INVX1  _975_
timestamp 0
transform 1 0 1370 0 -1 1830
box -6 -8 46 268
use NAND2X1  _976_
timestamp 0
transform -1 0 1210 0 -1 1310
box -6 -8 66 268
use INVX2  _977_
timestamp 0
transform -1 0 1750 0 1 1830
box -6 -8 46 268
use NAND2X1  _978_
timestamp 0
transform -1 0 1950 0 -1 1310
box -6 -8 66 268
use OAI21X1  _979_
timestamp 0
transform 1 0 1290 0 -1 1310
box -6 -8 86 268
use OAI21X1  _980_
timestamp 0
transform -1 0 1070 0 -1 1310
box -6 -8 86 268
use AOI21X1  _981_
timestamp 0
transform 1 0 250 0 -1 1310
box -6 -8 86 268
use OAI21X1  _982_
timestamp 0
transform 1 0 690 0 -1 1310
box -6 -8 86 268
use OAI21X1  _983_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 86 268
use AND2X2  _984_
timestamp 0
transform -1 0 1750 0 1 2350
box -6 -8 86 268
use NAND3X1  _985_
timestamp 0
transform 1 0 1570 0 1 1830
box -6 -8 86 268
use AOI22X1  _986_
timestamp 0
transform -1 0 1590 0 1 2350
box -6 -8 106 268
use INVX1  _987_
timestamp 0
transform -1 0 1610 0 1 270
box -6 -8 46 268
use NAND2X1  _988_
timestamp 0
transform 1 0 730 0 1 1310
box -6 -8 66 268
use INVX1  _989_
timestamp 0
transform 1 0 850 0 -1 270
box -6 -8 46 268
use NAND3X1  _990_
timestamp 0
transform -1 0 1030 0 -1 270
box -6 -8 86 268
use NAND2X1  _991_
timestamp 0
transform 1 0 1350 0 1 2350
box -6 -8 66 268
use NOR2X1  _992_
timestamp 0
transform -1 0 1510 0 -1 790
box -6 -8 66 268
use OAI21X1  _993_
timestamp 0
transform -1 0 770 0 -1 270
box -6 -8 86 268
use NAND3X1  _994_
timestamp 0
transform 1 0 90 0 -1 270
box -6 -8 86 268
use AOI21X1  _995_
timestamp 0
transform 1 0 210 0 -1 790
box -6 -8 86 268
use OAI21X1  _996_
timestamp 0
transform -1 0 1350 0 1 270
box -6 -8 86 268
use NAND3X1  _997_
timestamp 0
transform -1 0 1510 0 1 270
box -6 -8 86 268
use NAND3X1  _998_
timestamp 0
transform -1 0 1030 0 1 270
box -6 -8 86 268
use NAND2X1  _999_
timestamp 0
transform 1 0 1490 0 -1 1830
box -6 -8 66 268
use INVX1  _1000_
timestamp 0
transform 1 0 1570 0 1 1310
box -6 -8 46 268
use AND2X2  _1001_
timestamp 0
transform 1 0 2690 0 1 1310
box -6 -8 86 268
use NAND2X1  _1002_
timestamp 0
transform 1 0 1810 0 1 1310
box -6 -8 66 268
use INVX1  _1003_
timestamp 0
transform 1 0 3670 0 1 1310
box -6 -8 46 268
use OAI21X1  _1004_
timestamp 0
transform -1 0 1530 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1005_
timestamp 0
transform 1 0 1670 0 1 1310
box -6 -8 86 268
use OAI21X1  _1006_
timestamp 0
transform -1 0 1510 0 1 1310
box -6 -8 86 268
use INVX1  _1007_
timestamp 0
transform 1 0 3390 0 1 1310
box -6 -8 46 268
use OAI21X1  _1008_
timestamp 0
transform -1 0 2030 0 1 1310
box -6 -8 86 268
use NAND3X1  _1009_
timestamp 0
transform 1 0 1270 0 1 1310
box -6 -8 86 268
use AND2X2  _1010_
timestamp 0
transform -1 0 1050 0 1 790
box -6 -8 86 268
use NAND3X1  _1011_
timestamp 0
transform -1 0 470 0 -1 270
box -6 -8 86 268
use AOI21X1  _1012_
timestamp 0
transform -1 0 1190 0 1 270
box -6 -8 86 268
use AOI21X1  _1013_
timestamp 0
transform 1 0 230 0 -1 270
box -6 -8 86 268
use NAND2X1  _1014_
timestamp 0
transform -1 0 1190 0 1 790
box -6 -8 66 268
use OAI21X1  _1015_
timestamp 0
transform 1 0 810 0 1 270
box -6 -8 86 268
use NAND3X1  _1016_
timestamp 0
transform 1 0 1130 0 -1 790
box -6 -8 86 268
use AOI21X1  _1017_
timestamp 0
transform 1 0 1290 0 -1 790
box -6 -8 86 268
use OAI21X1  _1018_
timestamp 0
transform 1 0 2330 0 -1 790
box -6 -8 86 268
use AOI21X1  _1019_
timestamp 0
transform 1 0 550 0 -1 270
box -6 -8 86 268
use OAI21X1  _1020_
timestamp 0
transform 1 0 1590 0 -1 790
box -6 -8 86 268
use AND2X2  _1021_
timestamp 0
transform -1 0 3090 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1022_
timestamp 0
transform 1 0 2790 0 1 1830
box -6 -8 66 268
use INVX1  _1023_
timestamp 0
transform -1 0 3230 0 1 1830
box -6 -8 46 268
use INVX2  _1024_
timestamp 0
transform 1 0 3290 0 -1 3390
box -6 -8 46 268
use NAND2X1  _1025_
timestamp 0
transform -1 0 2990 0 1 1830
box -6 -8 66 268
use OAI21X1  _1026_
timestamp 0
transform -1 0 3130 0 1 1830
box -6 -8 86 268
use NAND2X1  _1027_
timestamp 0
transform 1 0 2850 0 1 1310
box -6 -8 66 268
use INVX1  _1028_
timestamp 0
transform 1 0 2910 0 1 790
box -6 -8 46 268
use NAND3X1  _1029_
timestamp 0
transform 1 0 3170 0 1 790
box -6 -8 86 268
use NOR2X1  _1030_
timestamp 0
transform 1 0 3050 0 -1 1830
box -6 -8 66 268
use AOI22X1  _1031_
timestamp 0
transform -1 0 3390 0 1 1830
box -6 -8 106 268
use OAI21X1  _1032_
timestamp 0
transform 1 0 3470 0 1 790
box -6 -8 86 268
use AOI21X1  _1033_
timestamp 0
transform -1 0 3750 0 -1 790
box -6 -8 86 268
use AOI21X1  _1034_
timestamp 0
transform 1 0 1090 0 -1 270
box -6 -8 86 268
use OAI21X1  _1035_
timestamp 0
transform -1 0 3110 0 1 790
box -6 -8 86 268
use NAND3X1  _1036_
timestamp 0
transform -1 0 2830 0 1 790
box -6 -8 86 268
use AOI21X1  _1037_
timestamp 0
transform -1 0 2050 0 -1 270
box -6 -8 86 268
use NAND2X1  _1038_
timestamp 0
transform -1 0 2790 0 -1 1310
box -6 -8 66 268
use INVX1  _1039_
timestamp 0
transform 1 0 2610 0 -1 1310
box -6 -8 46 268
use AND2X2  _1040_
timestamp 0
transform 1 0 2110 0 1 1310
box -6 -8 86 268
use AND2X2  _1041_
timestamp 0
transform -1 0 2690 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1042_
timestamp 0
transform 1 0 2250 0 1 1310
box -6 -8 66 268
use INVX2  _1043_
timestamp 0
transform -1 0 1390 0 1 1830
box -6 -8 46 268
use NAND2X1  _1044_
timestamp 0
transform 1 0 2010 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1045_
timestamp 0
transform -1 0 2230 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1046_
timestamp 0
transform 1 0 2310 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1047_
timestamp 0
transform 1 0 2370 0 1 1310
box -6 -8 86 268
use OAI21X1  _1048_
timestamp 0
transform -1 0 2610 0 1 1310
box -6 -8 86 268
use NAND3X1  _1049_
timestamp 0
transform 1 0 2470 0 -1 1310
box -6 -8 86 268
use AND2X2  _1050_
timestamp 0
transform 1 0 2610 0 1 790
box -6 -8 86 268
use OAI21X1  _1051_
timestamp 0
transform -1 0 1890 0 -1 270
box -6 -8 86 268
use NAND3X1  _1052_
timestamp 0
transform 1 0 2110 0 -1 270
box -6 -8 86 268
use NAND3X1  _1053_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 86 268
use NAND2X1  _1054_
timestamp 0
transform 1 0 2490 0 1 790
box -6 -8 66 268
use NAND3X1  _1055_
timestamp 0
transform -1 0 2330 0 -1 270
box -6 -8 86 268
use NAND3X1  _1056_
timestamp 0
transform 1 0 1250 0 -1 270
box -6 -8 86 268
use OAI21X1  _1057_
timestamp 0
transform -1 0 430 0 1 270
box -6 -8 86 268
use NAND3X1  _1058_
timestamp 0
transform 1 0 2910 0 1 270
box -6 -8 86 268
use OAI21X1  _1059_
timestamp 0
transform -1 0 2830 0 1 270
box -6 -8 86 268
use NAND3X1  _1060_
timestamp 0
transform -1 0 2510 0 1 270
box -6 -8 86 268
use INVX4  _1061_
timestamp 0
transform -1 0 2770 0 1 3910
box -6 -8 66 268
use NOR2X1  _1062_
timestamp 0
transform -1 0 2250 0 1 790
box -6 -8 66 268
use OAI21X1  _1063_
timestamp 0
transform -1 0 1810 0 -1 1310
box -6 -8 86 268
use XNOR2X1  _1064_
timestamp 0
transform 1 0 1870 0 1 790
box -6 -8 126 268
use INVX1  _1065_
timestamp 0
transform -1 0 1730 0 -1 270
box -6 -8 46 268
use NAND3X1  _1066_
timestamp 0
transform 1 0 1850 0 1 270
box -6 -8 86 268
use AOI21X1  _1067_
timestamp 0
transform -1 0 2670 0 1 270
box -6 -8 86 268
use AOI21X1  _1068_
timestamp 0
transform 1 0 1390 0 -1 270
box -6 -8 86 268
use OAI21X1  _1069_
timestamp 0
transform 1 0 2150 0 1 270
box -6 -8 86 268
use NAND3X1  _1070_
timestamp 0
transform 1 0 2770 0 -1 790
box -6 -8 86 268
use NAND2X1  _1071_
timestamp 0
transform -1 0 2110 0 1 790
box -6 -8 66 268
use INVX1  _1072_
timestamp 0
transform -1 0 3730 0 1 270
box -6 -8 46 268
use OAI21X1  _1073_
timestamp 0
transform 1 0 2290 0 1 270
box -6 -8 86 268
use AOI21X1  _1074_
timestamp 0
transform 1 0 3070 0 1 270
box -6 -8 86 268
use OAI21X1  _1075_
timestamp 0
transform 1 0 3630 0 1 790
box -6 -8 86 268
use NAND3X1  _1076_
timestamp 0
transform -1 0 3530 0 1 1830
box -6 -8 86 268
use AOI22X1  _1077_
timestamp 0
transform 1 0 3610 0 1 1830
box -6 -8 106 268
use INVX1  _1078_
timestamp 0
transform -1 0 3830 0 1 1310
box -6 -8 46 268
use NAND2X1  _1079_
timestamp 0
transform 1 0 3330 0 -1 1830
box -6 -8 66 268
use INVX1  _1080_
timestamp 0
transform 1 0 3910 0 1 1310
box -6 -8 46 268
use NAND3X1  _1081_
timestamp 0
transform 1 0 4050 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1082_
timestamp 0
transform 1 0 3790 0 1 1830
box -6 -8 66 268
use NOR2X1  _1083_
timestamp 0
transform 1 0 3870 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1084_
timestamp 0
transform 1 0 4190 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1085_
timestamp 0
transform 1 0 4290 0 1 790
box -6 -8 86 268
use OAI21X1  _1086_
timestamp 0
transform 1 0 3910 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1087_
timestamp 0
transform 1 0 3770 0 -1 1310
box -6 -8 86 268
use AOI22X1  _1088_
timestamp 0
transform 1 0 3790 0 1 790
box -6 -8 106 268
use NAND2X1  _1089_
timestamp 0
transform -1 0 3410 0 -1 1310
box -6 -8 66 268
use INVX1  _1090_
timestamp 0
transform 1 0 3490 0 -1 1310
box -6 -8 46 268
use AND2X2  _1091_
timestamp 0
transform -1 0 2970 0 -1 1830
box -6 -8 86 268
use AND2X2  _1092_
timestamp 0
transform 1 0 2970 0 1 1310
box -6 -8 86 268
use NAND2X1  _1093_
timestamp 0
transform -1 0 3190 0 1 1310
box -6 -8 66 268
use AOI22X1  _1094_
timestamp 0
transform 1 0 3170 0 -1 1830
box -6 -8 106 268
use INVX1  _1095_
timestamp 0
transform 1 0 3610 0 -1 1830
box -6 -8 46 268
use NAND3X1  _1096_
timestamp 0
transform 1 0 3610 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1097_
timestamp 0
transform -1 0 3330 0 1 1310
box -6 -8 86 268
use OAI21X1  _1098_
timestamp 0
transform 1 0 3050 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1099_
timestamp 0
transform -1 0 3290 0 -1 1310
box -6 -8 86 268
use AND2X2  _1100_
timestamp 0
transform 1 0 3970 0 -1 790
box -6 -8 86 268
use OAI21X1  _1101_
timestamp 0
transform -1 0 4470 0 -1 790
box -6 -8 86 268
use AOI21X1  _1102_
timestamp 0
transform 1 0 3310 0 1 790
box -6 -8 86 268
use NAND3X1  _1103_
timestamp 0
transform 1 0 3970 0 1 790
box -6 -8 86 268
use NAND3X1  _1104_
timestamp 0
transform 1 0 4130 0 1 790
box -6 -8 86 268
use NAND2X1  _1105_
timestamp 0
transform 1 0 4110 0 -1 790
box -6 -8 66 268
use NAND3X1  _1106_
timestamp 0
transform -1 0 4630 0 -1 790
box -6 -8 86 268
use NAND3X1  _1107_
timestamp 0
transform -1 0 4330 0 1 270
box -6 -8 86 268
use OAI21X1  _1108_
timestamp 0
transform 1 0 2410 0 -1 270
box -6 -8 86 268
use NAND3X1  _1109_
timestamp 0
transform -1 0 4050 0 1 270
box -6 -8 86 268
use OAI21X1  _1110_
timestamp 0
transform -1 0 4310 0 -1 790
box -6 -8 86 268
use NAND3X1  _1111_
timestamp 0
transform 1 0 3350 0 -1 270
box -6 -8 86 268
use NAND2X1  _1112_
timestamp 0
transform -1 0 3790 0 -1 1830
box -6 -8 66 268
use INVX1  _1113_
timestamp 0
transform -1 0 5030 0 1 270
box -6 -8 46 268
use AOI22X1  _1114_
timestamp 0
transform -1 0 2970 0 -1 1310
box -6 -8 106 268
use INVX1  _1115_
timestamp 0
transform 1 0 4890 0 1 790
box -6 -8 46 268
use OAI21X1  _1116_
timestamp 0
transform 1 0 4750 0 1 790
box -6 -8 86 268
use NOR2X1  _1117_
timestamp 0
transform -1 0 4710 0 -1 1310
box -6 -8 66 268
use NAND2X1  _1118_
timestamp 0
transform -1 0 5070 0 -1 790
box -6 -8 66 268
use NAND3X1  _1119_
timestamp 0
transform -1 0 4930 0 1 270
box -6 -8 86 268
use NAND2X1  _1120_
timestamp 0
transform -1 0 5210 0 -1 790
box -6 -8 66 268
use OAI21X1  _1121_
timestamp 0
transform -1 0 4670 0 1 790
box -6 -8 86 268
use NAND3X1  _1122_
timestamp 0
transform -1 0 4610 0 1 270
box -6 -8 86 268
use NAND2X1  _1123_
timestamp 0
transform 1 0 4390 0 1 270
box -6 -8 66 268
use NAND3X1  _1124_
timestamp 0
transform -1 0 3590 0 -1 270
box -6 -8 86 268
use AOI21X1  _1125_
timestamp 0
transform -1 0 3270 0 -1 270
box -6 -8 86 268
use AOI21X1  _1126_
timestamp 0
transform -1 0 4190 0 1 270
box -6 -8 86 268
use NAND3X1  _1127_
timestamp 0
transform -1 0 4770 0 1 270
box -6 -8 86 268
use NAND3X1  _1128_
timestamp 0
transform -1 0 4950 0 -1 790
box -6 -8 86 268
use NAND2X1  _1129_
timestamp 0
transform -1 0 4490 0 -1 270
box -6 -8 66 268
use OAI21X1  _1130_
timestamp 0
transform -1 0 4050 0 -1 270
box -6 -8 86 268
use AOI21X1  _1131_
timestamp 0
transform 1 0 3030 0 -1 270
box -6 -8 86 268
use AOI21X1  _1132_
timestamp 0
transform 1 0 1550 0 -1 270
box -6 -8 86 268
use OAI21X1  _1133_
timestamp 0
transform -1 0 3890 0 -1 270
box -6 -8 86 268
use NAND3X1  _1134_
timestamp 0
transform -1 0 3730 0 -1 270
box -6 -8 86 268
use AOI21X1  _1135_
timestamp 0
transform -1 0 2650 0 -1 270
box -6 -8 86 268
use OAI21X1  _1136_
timestamp 0
transform 1 0 3370 0 1 270
box -6 -8 86 268
use NAND3X1  _1137_
timestamp 0
transform 1 0 2730 0 -1 270
box -6 -8 86 268
use NAND3X1  _1138_
timestamp 0
transform -1 0 2970 0 -1 270
box -6 -8 86 268
use NAND3X1  _1139_
timestamp 0
transform -1 0 3450 0 -1 790
box -6 -8 86 268
use AOI21X1  _1140_
timestamp 0
transform -1 0 3150 0 -1 790
box -6 -8 86 268
use INVX1  _1141_
timestamp 0
transform 1 0 2530 0 1 1830
box -6 -8 46 268
use INVX1  _1142_
timestamp 0
transform -1 0 2270 0 -1 790
box -6 -8 46 268
use NOR2X1  _1143_
timestamp 0
transform 1 0 90 0 1 1830
box -6 -8 66 268
use INVX1  _1144_
timestamp 0
transform -1 0 110 0 1 1310
box -6 -8 46 268
use OAI21X1  _1145_
timestamp 0
transform -1 0 770 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1146_
timestamp 0
transform 1 0 90 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1147_
timestamp 0
transform -1 0 150 0 -1 790
box -6 -8 86 268
use NAND3X1  _1148_
timestamp 0
transform -1 0 490 0 1 790
box -6 -8 86 268
use AOI21X1  _1149_
timestamp 0
transform 1 0 90 0 1 790
box -6 -8 86 268
use AND2X2  _1150_
timestamp 0
transform -1 0 1330 0 1 790
box -6 -8 86 268
use NAND3X1  _1151_
timestamp 0
transform 1 0 250 0 1 790
box -6 -8 86 268
use AOI21X1  _1152_
timestamp 0
transform -1 0 770 0 1 790
box -6 -8 86 268
use OAI21X1  _1153_
timestamp 0
transform 1 0 670 0 1 270
box -6 -8 86 268
use NAND3X1  _1154_
timestamp 0
transform 1 0 510 0 1 270
box -6 -8 86 268
use NAND3X1  _1155_
timestamp 0
transform 1 0 970 0 -1 790
box -6 -8 86 268
use NAND3X1  _1156_
timestamp 0
transform 1 0 1910 0 -1 790
box -6 -8 86 268
use OAI21X1  _1157_
timestamp 0
transform -1 0 2070 0 1 270
box -6 -8 86 268
use NAND3X1  _1158_
timestamp 0
transform 1 0 1690 0 1 270
box -6 -8 86 268
use AOI22X1  _1159_
timestamp 0
transform -1 0 2170 0 -1 790
box -6 -8 106 268
use NAND3X1  _1160_
timestamp 0
transform -1 0 3590 0 -1 790
box -6 -8 86 268
use OAI21X1  _1161_
timestamp 0
transform 1 0 3230 0 1 270
box -6 -8 86 268
use AOI21X1  _1162_
timestamp 0
transform -1 0 3310 0 -1 790
box -6 -8 86 268
use NAND3X1  _1163_
timestamp 0
transform 1 0 830 0 1 790
box -6 -8 86 268
use NAND3X1  _1164_
timestamp 0
transform 1 0 390 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1165_
timestamp 0
transform -1 0 2050 0 -1 2870
box -6 -8 66 268
use OR2X2  _1166_
timestamp 0
transform 1 0 90 0 1 2350
box -6 -8 86 268
use NAND2X1  _1167_
timestamp 0
transform 1 0 250 0 1 2350
box -6 -8 66 268
use AOI22X1  _1168_
timestamp 0
transform -1 0 890 0 1 1830
box -6 -8 106 268
use OAI21X1  _1169_
timestamp 0
transform -1 0 330 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1170_
timestamp 0
transform 1 0 230 0 1 1830
box -6 -8 86 268
use NAND3X1  _1171_
timestamp 0
transform 1 0 370 0 1 1830
box -6 -8 86 268
use AOI21X1  _1172_
timestamp 0
transform 1 0 530 0 1 1830
box -6 -8 86 268
use OAI21X1  _1173_
timestamp 0
transform -1 0 1290 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1174_
timestamp 0
transform 1 0 550 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1175_
timestamp 0
transform 1 0 850 0 -1 1310
box -6 -8 86 268
use INVX1  _1176_
timestamp 0
transform -1 0 1190 0 1 1310
box -6 -8 46 268
use AOI22X1  _1177_
timestamp 0
transform -1 0 910 0 -1 790
box -6 -8 106 268
use OAI21X1  _1178_
timestamp 0
transform 1 0 1570 0 1 790
box -6 -8 86 268
use NAND3X1  _1179_
timestamp 0
transform 1 0 1710 0 1 790
box -6 -8 86 268
use AOI21X1  _1180_
timestamp 0
transform -1 0 2690 0 -1 790
box -6 -8 86 268
use NOR3X1  _1181_
timestamp 0
transform 1 0 1810 0 1 1830
box -6 -8 166 268
use INVX1  _1182_
timestamp 0
transform 1 0 1070 0 1 1830
box -6 -8 46 268
use NAND3X1  _1183_
timestamp 0
transform -1 0 1270 0 1 1830
box -6 -8 86 268
use INVX1  _1184_
timestamp 0
transform 1 0 390 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1185_
timestamp 0
transform 1 0 390 0 1 2350
box -6 -8 86 268
use OR2X2  _1186_
timestamp 0
transform 1 0 530 0 1 2350
box -6 -8 86 268
use NAND2X1  _1187_
timestamp 0
transform -1 0 1930 0 -1 2870
box -6 -8 66 268
use NOR2X1  _1188_
timestamp 0
transform 1 0 1330 0 -1 2870
box -6 -8 66 268
use INVX1  _1189_
timestamp 0
transform -1 0 670 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1190_
timestamp 0
transform -1 0 830 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1191_
timestamp 0
transform -1 0 770 0 1 2350
box -6 -8 86 268
use INVX1  _1192_
timestamp 0
transform 1 0 830 0 1 2350
box -6 -8 46 268
use INVX1  _1193_
timestamp 0
transform 1 0 970 0 -1 1830
box -6 -8 46 268
use OAI21X1  _1194_
timestamp 0
transform 1 0 1070 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1195_
timestamp 0
transform 1 0 1050 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1196_
timestamp 0
transform 1 0 870 0 1 1310
box -6 -8 86 268
use NOR3X1  _1197_
timestamp 0
transform 1 0 1330 0 -1 2350
box -6 -8 166 268
use OAI21X1  _1198_
timestamp 0
transform 1 0 1750 0 -1 790
box -6 -8 86 268
use NAND3X1  _1199_
timestamp 0
transform 1 0 1410 0 1 790
box -6 -8 86 268
use NAND3X1  _1200_
timestamp 0
transform 1 0 1590 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1201_
timestamp 0
transform 1 0 1830 0 -1 2350
box -6 -8 86 268
use INVX1  _1202_
timestamp 0
transform 1 0 2110 0 -1 2870
box -6 -8 46 268
use OAI21X1  _1203_
timestamp 0
transform -1 0 2130 0 1 1830
box -6 -8 86 268
use AOI21X1  _1204_
timestamp 0
transform 1 0 2290 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1205_
timestamp 0
transform -1 0 2950 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1206_
timestamp 0
transform 1 0 3530 0 1 270
box -6 -8 86 268
use NAND2X1  _1207_
timestamp 0
transform -1 0 5150 0 1 270
box -6 -8 66 268
use OAI21X1  _1208_
timestamp 0
transform -1 0 4210 0 -1 270
box -6 -8 86 268
use NAND2X1  _1209_
timestamp 0
transform -1 0 3530 0 -1 1830
box -6 -8 66 268
use INVX1  _1210_
timestamp 0
transform -1 0 5170 0 1 790
box -6 -8 46 268
use NOR2X1  _1211_
timestamp 0
transform 1 0 4350 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1212_
timestamp 0
transform 1 0 3510 0 1 1310
box -6 -8 86 268
use NAND2X1  _1213_
timestamp 0
transform -1 0 4970 0 -1 1310
box -6 -8 66 268
use OR2X2  _1214_
timestamp 0
transform -1 0 4570 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1215_
timestamp 0
transform -1 0 5070 0 1 790
box -6 -8 86 268
use AND2X2  _1216_
timestamp 0
transform 1 0 5050 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1217_
timestamp 0
transform -1 0 4850 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1218_
timestamp 0
transform 1 0 5190 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1219_
timestamp 0
transform 1 0 5450 0 -1 790
box -6 -8 66 268
use AOI21X1  _1220_
timestamp 0
transform 1 0 4450 0 1 790
box -6 -8 86 268
use NAND2X1  _1221_
timestamp 0
transform 1 0 3710 0 -1 2350
box -6 -8 66 268
use AND2X2  _1222_
timestamp 0
transform -1 0 2450 0 1 2350
box -6 -8 86 268
use OAI21X1  _1223_
timestamp 0
transform -1 0 3510 0 -1 2350
box -6 -8 86 268
use AND2X2  _1224_
timestamp 0
transform 1 0 2530 0 1 2350
box -6 -8 86 268
use OAI21X1  _1225_
timestamp 0
transform 1 0 3170 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1226_
timestamp 0
transform 1 0 3570 0 -1 2350
box -6 -8 86 268
use INVX1  _1227_
timestamp 0
transform 1 0 3970 0 -1 2350
box -6 -8 46 268
use NAND2X1  _1228_
timestamp 0
transform -1 0 3370 0 -1 2350
box -6 -8 66 268
use AOI22X1  _1229_
timestamp 0
transform -1 0 3230 0 1 2350
box -6 -8 106 268
use INVX1  _1230_
timestamp 0
transform 1 0 3750 0 1 2350
box -6 -8 46 268
use NAND3X1  _1231_
timestamp 0
transform 1 0 4070 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1232_
timestamp 0
transform -1 0 4730 0 1 1830
box -6 -8 66 268
use AOI21X1  _1233_
timestamp 0
transform 1 0 4030 0 1 1310
box -6 -8 86 268
use NAND2X1  _1234_
timestamp 0
transform -1 0 3970 0 1 1830
box -6 -8 66 268
use XOR2X1  _1235_
timestamp 0
transform 1 0 4170 0 -1 1830
box -6 -8 126 268
use NAND2X1  _1236_
timestamp 0
transform -1 0 4490 0 1 1310
box -6 -8 66 268
use OAI21X1  _1237_
timestamp 0
transform 1 0 4010 0 -1 1830
box -6 -8 86 268
use XNOR2X1  _1238_
timestamp 0
transform 1 0 4050 0 1 1830
box -6 -8 126 268
use NAND2X1  _1239_
timestamp 0
transform -1 0 4410 0 -1 1830
box -6 -8 66 268
use NAND3X1  _1240_
timestamp 0
transform 1 0 4730 0 1 1310
box -6 -8 86 268
use AND2X2  _1241_
timestamp 0
transform -1 0 4890 0 1 1830
box -6 -8 86 268
use NAND2X1  _1242_
timestamp 0
transform 1 0 4610 0 -1 1830
box -6 -8 66 268
use NAND2X1  _1243_
timestamp 0
transform -1 0 4250 0 1 1310
box -6 -8 66 268
use NAND3X1  _1244_
timestamp 0
transform 1 0 4870 0 1 1310
box -6 -8 86 268
use NAND3X1  _1245_
timestamp 0
transform 1 0 5250 0 1 790
box -6 -8 86 268
use OAI21X1  _1246_
timestamp 0
transform 1 0 4710 0 -1 790
box -6 -8 86 268
use AOI22X1  _1247_
timestamp 0
transform 1 0 4890 0 -1 1830
box -6 -8 106 268
use AOI21X1  _1248_
timestamp 0
transform 1 0 4570 0 1 1310
box -6 -8 86 268
use OAI21X1  _1249_
timestamp 0
transform 1 0 5290 0 -1 790
box -6 -8 86 268
use NAND3X1  _1250_
timestamp 0
transform -1 0 5290 0 1 270
box -6 -8 86 268
use AND2X2  _1251_
timestamp 0
transform 1 0 5750 0 -1 790
box -6 -8 86 268
use NAND3X1  _1252_
timestamp 0
transform 1 0 5390 0 1 790
box -6 -8 86 268
use OAI21X1  _1253_
timestamp 0
transform 1 0 5870 0 1 790
box -6 -8 86 268
use NAND3X1  _1254_
timestamp 0
transform -1 0 5910 0 1 270
box -6 -8 86 268
use NAND3X1  _1255_
timestamp 0
transform 1 0 5010 0 -1 270
box -6 -8 86 268
use AOI21X1  _1256_
timestamp 0
transform 1 0 4290 0 -1 270
box -6 -8 86 268
use AOI22X1  _1257_
timestamp 0
transform 1 0 5570 0 -1 790
box -6 -8 106 268
use AOI21X1  _1258_
timestamp 0
transform 1 0 5370 0 1 270
box -6 -8 86 268
use OAI21X1  _1259_
timestamp 0
transform -1 0 4650 0 -1 270
box -6 -8 86 268
use AOI21X1  _1260_
timestamp 0
transform -1 0 6050 0 1 270
box -6 -8 86 268
use INVX1  _1261_
timestamp 0
transform -1 0 5670 0 -1 270
box -6 -8 46 268
use NAND3X1  _1262_
timestamp 0
transform -1 0 4950 0 -1 270
box -6 -8 86 268
use OAI21X1  _1263_
timestamp 0
transform 1 0 4710 0 -1 270
box -6 -8 86 268
use AOI21X1  _1264_
timestamp 0
transform 1 0 5310 0 -1 270
box -6 -8 86 268
use OAI21X1  _1265_
timestamp 0
transform -1 0 5590 0 1 270
box -6 -8 86 268
use OAI21X1  _1266_
timestamp 0
transform 1 0 3810 0 1 270
box -6 -8 86 268
use NAND3X1  _1267_
timestamp 0
transform 1 0 5470 0 -1 270
box -6 -8 86 268
use NAND3X1  _1268_
timestamp 0
transform -1 0 6190 0 1 270
box -6 -8 86 268
use NAND3X1  _1269_
timestamp 0
transform -1 0 5750 0 1 270
box -6 -8 86 268
use AND2X2  _1270_
timestamp 0
transform 1 0 5770 0 -1 2870
box -6 -8 86 268
use XOR2X1  _1271_
timestamp 0
transform 1 0 5150 0 1 3390
box -6 -8 126 268
use NOR2X1  _1272_
timestamp 0
transform -1 0 2690 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1273_
timestamp 0
transform -1 0 2630 0 1 4950
box -6 -8 66 268
use OAI21X1  _1274_
timestamp 0
transform -1 0 2830 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1275_
timestamp 0
transform 1 0 2550 0 1 3910
box -6 -8 86 268
use OAI21X1  _1276_
timestamp 0
transform 1 0 2430 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1277_
timestamp 0
transform 1 0 2590 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1278_
timestamp 0
transform -1 0 3810 0 -1 5470
box -6 -8 66 268
use OAI21X1  _1279_
timestamp 0
transform -1 0 3890 0 -1 5990
box -6 -8 86 268
use INVX1  _1280_
timestamp 0
transform 1 0 2250 0 1 5990
box -6 -8 46 268
use INVX1  _1281_
timestamp 0
transform 1 0 4010 0 1 4950
box -6 -8 46 268
use OAI21X1  _1282_
timestamp 0
transform 1 0 5190 0 1 4950
box -6 -8 86 268
use OAI21X1  _1283_
timestamp 0
transform -1 0 5770 0 1 4950
box -6 -8 86 268
use NAND3X1  _1284_
timestamp 0
transform -1 0 2990 0 -1 790
box -6 -8 86 268
use INVX1  _1285_
timestamp 0
transform 1 0 2050 0 -1 1830
box -6 -8 46 268
use NAND2X1  _1286_
timestamp 0
transform -1 0 2530 0 -1 790
box -6 -8 66 268
use NAND3X1  _1287_
timestamp 0
transform -1 0 2410 0 1 790
box -6 -8 86 268
use NAND3X1  _1288_
timestamp 0
transform -1 0 2390 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1289_
timestamp 0
transform -1 0 2230 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1290_
timestamp 0
transform 1 0 2210 0 1 1830
box -6 -8 86 268
use AOI21X1  _1291_
timestamp 0
transform 1 0 2370 0 1 1830
box -6 -8 86 268
use NAND2X1  _1292_
timestamp 0
transform -1 0 5690 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1293_
timestamp 0
transform 1 0 5670 0 1 2870
box -6 -8 86 268
use INVX1  _1294_
timestamp 0
transform -1 0 6250 0 -1 270
box -6 -8 46 268
use AOI21X1  _1295_
timestamp 0
transform 1 0 6070 0 -1 270
box -6 -8 86 268
use OAI21X1  _1296_
timestamp 0
transform 1 0 5350 0 -1 1310
box -6 -8 86 268
use INVX1  _1297_
timestamp 0
transform -1 0 6310 0 -1 1830
box -6 -8 46 268
use AOI21X1  _1298_
timestamp 0
transform 1 0 5550 0 1 790
box -6 -8 86 268
use OAI21X1  _1299_
timestamp 0
transform 1 0 5710 0 1 790
box -6 -8 86 268
use NAND2X1  _1300_
timestamp 0
transform 1 0 4230 0 1 1830
box -6 -8 66 268
use NOR2X1  _1301_
timestamp 0
transform 1 0 4530 0 1 1830
box -6 -8 66 268
use NAND2X1  _1302_
timestamp 0
transform 1 0 3430 0 1 2350
box -6 -8 66 268
use NAND2X1  _1303_
timestamp 0
transform -1 0 3370 0 1 2350
box -6 -8 66 268
use OAI22X1  _1304_
timestamp 0
transform 1 0 3570 0 1 2350
box -6 -8 106 268
use XNOR2X1  _1305_
timestamp 0
transform 1 0 5090 0 1 1830
box -6 -8 126 268
use XNOR2X1  _1306_
timestamp 0
transform 1 0 5430 0 1 1830
box -6 -8 126 268
use NOR2X1  _1307_
timestamp 0
transform -1 0 4370 0 1 1310
box -6 -8 66 268
use AOI21X1  _1308_
timestamp 0
transform 1 0 5030 0 1 1310
box -6 -8 86 268
use NAND2X1  _1309_
timestamp 0
transform 1 0 3230 0 1 2870
box -6 -8 66 268
use NAND2X1  _1310_
timestamp 0
transform -1 0 2710 0 1 2870
box -6 -8 66 268
use INVX1  _1311_
timestamp 0
transform 1 0 2670 0 -1 2870
box -6 -8 46 268
use AND2X2  _1312_
timestamp 0
transform -1 0 3150 0 1 2870
box -6 -8 86 268
use AND2X2  _1313_
timestamp 0
transform 1 0 2670 0 1 2350
box -6 -8 86 268
use NAND2X1  _1314_
timestamp 0
transform -1 0 2890 0 1 2350
box -6 -8 66 268
use AOI22X1  _1315_
timestamp 0
transform 1 0 2770 0 1 2870
box -6 -8 106 268
use INVX1  _1316_
timestamp 0
transform 1 0 2950 0 1 2870
box -6 -8 46 268
use AOI21X1  _1317_
timestamp 0
transform -1 0 2870 0 -1 2870
box -6 -8 86 268
use INVX2  _1318_
timestamp 0
transform 1 0 4050 0 1 3390
box -6 -8 46 268
use OAI21X1  _1319_
timestamp 0
transform -1 0 3730 0 1 2870
box -6 -8 86 268
use OAI21X1  _1320_
timestamp 0
transform -1 0 3050 0 1 2350
box -6 -8 86 268
use AOI21X1  _1321_
timestamp 0
transform -1 0 3430 0 1 2870
box -6 -8 86 268
use OAI22X1  _1322_
timestamp 0
transform -1 0 3370 0 -1 2870
box -6 -8 106 268
use NAND3X1  _1323_
timestamp 0
transform 1 0 3490 0 1 2870
box -6 -8 86 268
use NAND3X1  _1324_
timestamp 0
transform 1 0 2950 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1325_
timestamp 0
transform 1 0 3450 0 -1 2870
box -6 -8 66 268
use NAND3X1  _1326_
timestamp 0
transform 1 0 3570 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1327_
timestamp 0
transform -1 0 5250 0 1 1310
box -6 -8 66 268
use NOR2X1  _1328_
timestamp 0
transform -1 0 5530 0 1 1310
box -6 -8 66 268
use NOR2X1  _1329_
timestamp 0
transform -1 0 4550 0 -1 1830
box -6 -8 66 268
use OAI21X1  _1330_
timestamp 0
transform 1 0 4750 0 -1 1830
box -6 -8 86 268
use AOI21X1  _1331_
timestamp 0
transform 1 0 5190 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1332_
timestamp 0
transform 1 0 5490 0 -1 1830
box -6 -8 86 268
use XOR2X1  _1333_
timestamp 0
transform -1 0 5750 0 1 1830
box -6 -8 126 268
use NAND3X1  _1334_
timestamp 0
transform 1 0 5050 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1335_
timestamp 0
transform -1 0 5570 0 -1 1310
box -6 -8 66 268
use NAND3X1  _1336_
timestamp 0
transform 1 0 5750 0 1 1310
box -6 -8 86 268
use NAND3X1  _1337_
timestamp 0
transform 1 0 5970 0 -1 1830
box -6 -8 86 268
use NOR3X1  _1338_
timestamp 0
transform 1 0 6050 0 -1 790
box -6 -8 166 268
use AOI21X1  _1339_
timestamp 0
transform 1 0 5890 0 -1 790
box -6 -8 86 268
use AOI21X1  _1340_
timestamp 0
transform 1 0 5610 0 1 1310
box -6 -8 86 268
use NAND3X1  _1341_
timestamp 0
transform 1 0 5330 0 1 1310
box -6 -8 86 268
use OAI21X1  _1342_
timestamp 0
transform 1 0 5630 0 -1 1310
box -6 -8 86 268
use AOI21X1  _1343_
timestamp 0
transform -1 0 5870 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1344_
timestamp 0
transform -1 0 6010 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1345_
timestamp 0
transform 1 0 6210 0 1 1310
box -6 -8 86 268
use NAND3X1  _1346_
timestamp 0
transform 1 0 5910 0 1 1310
box -6 -8 86 268
use OAI21X1  _1347_
timestamp 0
transform 1 0 6070 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1348_
timestamp 0
transform -1 0 6310 0 -1 1310
box -6 -8 86 268
use NAND3X1  _1349_
timestamp 0
transform 1 0 6210 0 1 790
box -6 -8 86 268
use AOI21X1  _1350_
timestamp 0
transform 1 0 5150 0 -1 270
box -6 -8 86 268
use OAI21X1  _1351_
timestamp 0
transform 1 0 5750 0 -1 270
box -6 -8 86 268
use NAND3X1  _1352_
timestamp 0
transform -1 0 6130 0 1 1310
box -6 -8 86 268
use NAND3X1  _1353_
timestamp 0
transform -1 0 6210 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1354_
timestamp 0
transform -1 0 6030 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1355_
timestamp 0
transform 1 0 6090 0 -1 2350
box -6 -8 66 268
use AND2X2  _1356_
timestamp 0
transform 1 0 5490 0 1 3390
box -6 -8 86 268
use OAI21X1  _1357_
timestamp 0
transform -1 0 5410 0 1 3390
box -6 -8 86 268
use OAI21X1  _1358_
timestamp 0
transform 1 0 5530 0 1 4950
box -6 -8 86 268
use AND2X2  _1359_
timestamp 0
transform 1 0 1970 0 1 2870
box -6 -8 86 268
use NAND2X1  _1360_
timestamp 0
transform 1 0 2010 0 1 3910
box -6 -8 66 268
use OAI21X1  _1361_
timestamp 0
transform 1 0 2130 0 1 2870
box -6 -8 86 268
use OAI21X1  _1362_
timestamp 0
transform -1 0 2090 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1363_
timestamp 0
transform 1 0 2750 0 -1 5470
box -6 -8 86 268
use AOI22X1  _1364_
timestamp 0
transform 1 0 2690 0 -1 5990
box -6 -8 106 268
use OAI21X1  _1365_
timestamp 0
transform -1 0 3510 0 -1 5990
box -6 -8 86 268
use AOI21X1  _1366_
timestamp 0
transform -1 0 5910 0 1 1830
box -6 -8 86 268
use AOI22X1  _1367_
timestamp 0
transform 1 0 6030 0 1 790
box -6 -8 106 268
use NOR2X1  _1368_
timestamp 0
transform -1 0 6030 0 1 1830
box -6 -8 66 268
use NAND3X1  _1369_
timestamp 0
transform 1 0 6070 0 -1 2870
box -6 -8 86 268
use AOI21X1  _1370_
timestamp 0
transform 1 0 5790 0 -1 2350
box -6 -8 86 268
use INVX1  _1371_
timestamp 0
transform -1 0 6290 0 1 2870
box -6 -8 46 268
use NAND2X1  _1372_
timestamp 0
transform -1 0 5030 0 1 1830
box -6 -8 66 268
use OAI21X1  _1373_
timestamp 0
transform -1 0 5350 0 1 1830
box -6 -8 86 268
use INVX1  _1374_
timestamp 0
transform -1 0 5730 0 1 2350
box -6 -8 46 268
use AOI21X1  _1375_
timestamp 0
transform -1 0 5730 0 -1 1830
box -6 -8 86 268
use NAND2X1  _1376_
timestamp 0
transform 1 0 3850 0 -1 2870
box -6 -8 66 268
use INVX1  _1377_
timestamp 0
transform 1 0 4590 0 -1 2870
box -6 -8 46 268
use NOR2X1  _1378_
timestamp 0
transform 1 0 3830 0 -1 2350
box -6 -8 66 268
use OAI21X1  _1379_
timestamp 0
transform -1 0 3190 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1380_
timestamp 0
transform -1 0 4050 0 -1 2870
box -6 -8 66 268
use OR2X2  _1381_
timestamp 0
transform 1 0 4110 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1382_
timestamp 0
transform 1 0 4710 0 -1 2870
box -6 -8 86 268
use AND2X2  _1383_
timestamp 0
transform -1 0 3950 0 1 2350
box -6 -8 86 268
use NOR2X1  _1384_
timestamp 0
transform -1 0 4070 0 1 2350
box -6 -8 66 268
use OAI21X1  _1385_
timestamp 0
transform 1 0 4150 0 1 2350
box -6 -8 86 268
use NAND2X1  _1386_
timestamp 0
transform 1 0 4850 0 -1 2870
box -6 -8 66 268
use OR2X2  _1387_
timestamp 0
transform 1 0 4370 0 1 1830
box -6 -8 86 268
use NAND2X1  _1388_
timestamp 0
transform 1 0 3730 0 -1 2870
box -6 -8 66 268
use NAND2X1  _1389_
timestamp 0
transform 1 0 3970 0 1 2870
box -6 -8 66 268
use NAND2X1  _1390_
timestamp 0
transform -1 0 3470 0 -1 3390
box -6 -8 66 268
use AOI22X1  _1391_
timestamp 0
transform -1 0 3910 0 1 2870
box -6 -8 106 268
use INVX1  _1392_
timestamp 0
transform 1 0 4430 0 1 2870
box -6 -8 46 268
use OAI21X1  _1393_
timestamp 0
transform 1 0 4290 0 1 2870
box -6 -8 86 268
use XNOR2X1  _1394_
timestamp 0
transform -1 0 4370 0 -1 2870
box -6 -8 126 268
use AOI21X1  _1395_
timestamp 0
transform 1 0 4750 0 -1 2350
box -6 -8 86 268
use NAND3X1  _1396_
timestamp 0
transform 1 0 4590 0 -1 2350
box -6 -8 86 268
use INVX1  _1397_
timestamp 0
transform 1 0 4890 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1398_
timestamp 0
transform 1 0 5170 0 -1 2350
box -6 -8 86 268
use AND2X2  _1399_
timestamp 0
transform 1 0 4750 0 1 2350
box -6 -8 86 268
use NAND2X1  _1400_
timestamp 0
transform -1 0 4510 0 -1 2350
box -6 -8 66 268
use INVX1  _1401_
timestamp 0
transform -1 0 4270 0 -1 2350
box -6 -8 46 268
use NAND2X1  _1402_
timestamp 0
transform -1 0 4390 0 -1 2350
box -6 -8 66 268
use NAND3X1  _1403_
timestamp 0
transform 1 0 5090 0 1 2350
box -6 -8 86 268
use NAND3X1  _1404_
timestamp 0
transform 1 0 5630 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1405_
timestamp 0
transform -1 0 5410 0 -1 1830
box -6 -8 86 268
use AOI22X1  _1406_
timestamp 0
transform 1 0 4910 0 1 2350
box -6 -8 106 268
use OR2X2  _1407_
timestamp 0
transform 1 0 4430 0 1 2350
box -6 -8 86 268
use NAND2X1  _1408_
timestamp 0
transform 1 0 4310 0 1 2350
box -6 -8 66 268
use AOI21X1  _1409_
timestamp 0
transform 1 0 4590 0 1 2350
box -6 -8 86 268
use OAI21X1  _1410_
timestamp 0
transform 1 0 5390 0 1 2350
box -6 -8 86 268
use NAND3X1  _1411_
timestamp 0
transform 1 0 5970 0 1 2350
box -6 -8 86 268
use NAND3X1  _1412_
timestamp 0
transform 1 0 5470 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1413_
timestamp 0
transform 1 0 5530 0 1 2350
box -6 -8 86 268
use NAND3X1  _1414_
timestamp 0
transform 1 0 5810 0 1 2350
box -6 -8 86 268
use NAND2X1  _1415_
timestamp 0
transform -1 0 6290 0 1 1830
box -6 -8 66 268
use NAND3X1  _1416_
timestamp 0
transform 1 0 6230 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1417_
timestamp 0
transform 1 0 5810 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1418_
timestamp 0
transform -1 0 6170 0 1 1830
box -6 -8 86 268
use NAND3X1  _1419_
timestamp 0
transform -1 0 6210 0 1 2350
box -6 -8 86 268
use NAND2X1  _1420_
timestamp 0
transform -1 0 6290 0 -1 2870
box -6 -8 66 268
use AOI21X1  _1421_
timestamp 0
transform -1 0 6190 0 1 2870
box -6 -8 86 268
use NAND2X1  _1422_
timestamp 0
transform 1 0 5930 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1423_
timestamp 0
transform 1 0 5970 0 1 2870
box -6 -8 86 268
use INVX1  _1424_
timestamp 0
transform -1 0 6310 0 -1 3910
box -6 -8 46 268
use NOR2X1  _1425_
timestamp 0
transform -1 0 6050 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1426_
timestamp 0
transform -1 0 5910 0 -1 3910
box -6 -8 86 268
use NOR2X1  _1427_
timestamp 0
transform -1 0 2330 0 1 5470
box -6 -8 66 268
use NOR2X1  _1428_
timestamp 0
transform 1 0 2550 0 1 5470
box -6 -8 66 268
use AOI21X1  _1429_
timestamp 0
transform 1 0 750 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1430_
timestamp 0
transform 1 0 1170 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1431_
timestamp 0
transform 1 0 2450 0 1 4950
box -6 -8 66 268
use NOR2X1  _1432_
timestamp 0
transform 1 0 2690 0 1 5470
box -6 -8 66 268
use AOI22X1  _1433_
timestamp 0
transform 1 0 2830 0 1 5470
box -6 -8 106 268
use OAI21X1  _1434_
timestamp 0
transform 1 0 3170 0 -1 5990
box -6 -8 86 268
use INVX1  _1435_
timestamp 0
transform -1 0 6210 0 1 4950
box -6 -8 46 268
use INVX1  _1436_
timestamp 0
transform 1 0 4470 0 1 5990
box -6 -8 46 268
use OAI21X1  _1437_
timestamp 0
transform 1 0 5490 0 -1 4950
box -6 -8 86 268
use INVX1  _1438_
timestamp 0
transform -1 0 6150 0 1 3390
box -6 -8 46 268
use OAI21X1  _1439_
timestamp 0
transform 1 0 4430 0 -1 2870
box -6 -8 86 268
use INVX1  _1440_
timestamp 0
transform 1 0 5370 0 -1 2870
box -6 -8 46 268
use AOI21X1  _1441_
timestamp 0
transform 1 0 5250 0 1 2350
box -6 -8 86 268
use NAND2X1  _1442_
timestamp 0
transform 1 0 3790 0 1 3390
box -6 -8 66 268
use INVX1  _1443_
timestamp 0
transform 1 0 4690 0 -1 3390
box -6 -8 46 268
use NOR2X1  _1444_
timestamp 0
transform 1 0 4530 0 1 2870
box -6 -8 66 268
use OAI22X1  _1445_
timestamp 0
transform 1 0 4110 0 1 2870
box -6 -8 106 268
use NAND2X1  _1446_
timestamp 0
transform 1 0 4790 0 1 2870
box -6 -8 66 268
use NOR2X1  _1447_
timestamp 0
transform 1 0 4650 0 1 2870
box -6 -8 66 268
use INVX1  _1448_
timestamp 0
transform 1 0 5090 0 1 2870
box -6 -8 46 268
use NAND3X1  _1449_
timestamp 0
transform 1 0 4930 0 1 2870
box -6 -8 86 268
use INVX1  _1450_
timestamp 0
transform -1 0 5090 0 1 3390
box -6 -8 46 268
use OAI21X1  _1451_
timestamp 0
transform -1 0 4990 0 1 3390
box -6 -8 86 268
use NAND2X1  _1452_
timestamp 0
transform -1 0 3730 0 -1 3390
box -6 -8 66 268
use NAND2X1  _1453_
timestamp 0
transform 1 0 3930 0 1 3390
box -6 -8 66 268
use OR2X2  _1454_
timestamp 0
transform 1 0 3810 0 -1 3390
box -6 -8 86 268
use INVX1  _1455_
timestamp 0
transform 1 0 4290 0 -1 3910
box -6 -8 46 268
use OAI21X1  _1456_
timestamp 0
transform 1 0 4330 0 1 3390
box -6 -8 86 268
use AND2X2  _1457_
timestamp 0
transform 1 0 4390 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1458_
timestamp 0
transform -1 0 4890 0 -1 3390
box -6 -8 86 268
use INVX1  _1459_
timestamp 0
transform 1 0 4990 0 -1 2870
box -6 -8 46 268
use NAND3X1  _1460_
timestamp 0
transform 1 0 4950 0 -1 3390
box -6 -8 86 268
use NAND3X1  _1461_
timestamp 0
transform 1 0 5370 0 1 2870
box -6 -8 86 268
use OAI21X1  _1462_
timestamp 0
transform 1 0 5010 0 -1 2350
box -6 -8 86 268
use INVX1  _1463_
timestamp 0
transform 1 0 5090 0 -1 2870
box -6 -8 46 268
use OAI21X1  _1464_
timestamp 0
transform 1 0 5210 0 1 2870
box -6 -8 86 268
use NAND3X1  _1465_
timestamp 0
transform 1 0 5510 0 1 2870
box -6 -8 86 268
use NAND3X1  _1466_
timestamp 0
transform 1 0 5110 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1467_
timestamp 0
transform 1 0 5210 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1468_
timestamp 0
transform 1 0 5250 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1469_
timestamp 0
transform -1 0 5470 0 -1 3390
box -6 -8 66 268
use NAND3X1  _1470_
timestamp 0
transform 1 0 5830 0 1 2870
box -6 -8 86 268
use AOI21X1  _1471_
timestamp 0
transform 1 0 5310 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1472_
timestamp 0
transform 1 0 5490 0 -1 2870
box -6 -8 86 268
use NAND3X1  _1473_
timestamp 0
transform 1 0 5530 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1474_
timestamp 0
transform -1 0 6170 0 -1 3390
box -6 -8 66 268
use NOR3X1  _1475_
timestamp 0
transform -1 0 6170 0 1 3910
box -6 -8 166 268
use AOI21X1  _1476_
timestamp 0
transform -1 0 6190 0 -1 3910
box -6 -8 86 268
use INVX1  _1477_
timestamp 0
transform -1 0 5790 0 1 3910
box -6 -8 46 268
use OAI21X1  _1478_
timestamp 0
transform 1 0 5850 0 1 3910
box -6 -8 86 268
use OAI21X1  _1479_
timestamp 0
transform -1 0 5890 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1480_
timestamp 0
transform 1 0 910 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1481_
timestamp 0
transform 1 0 930 0 1 2350
box -6 -8 66 268
use NAND2X1  _1482_
timestamp 0
transform -1 0 1130 0 1 2350
box -6 -8 66 268
use NAND2X1  _1483_
timestamp 0
transform 1 0 2170 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1484_
timestamp 0
transform -1 0 2370 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1485_
timestamp 0
transform 1 0 4650 0 -1 4950
box -6 -8 86 268
use AOI22X1  _1486_
timestamp 0
transform -1 0 5930 0 1 4950
box -6 -8 106 268
use INVX1  _1487_
timestamp 0
transform -1 0 2610 0 -1 5990
box -6 -8 46 268
use OAI21X1  _1488_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 86 268
use INVX1  _1489_
timestamp 0
transform 1 0 4910 0 1 3910
box -6 -8 46 268
use INVX1  _1490_
timestamp 0
transform 1 0 3930 0 -1 3910
box -6 -8 46 268
use NAND2X1  _1491_
timestamp 0
transform -1 0 3610 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1492_
timestamp 0
transform 1 0 3950 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1493_
timestamp 0
transform -1 0 4190 0 -1 3390
box -6 -8 86 268
use OR2X2  _1494_
timestamp 0
transform 1 0 4250 0 -1 3390
box -6 -8 86 268
use INVX1  _1495_
timestamp 0
transform -1 0 4230 0 -1 3910
box -6 -8 46 268
use OAI21X1  _1496_
timestamp 0
transform 1 0 4170 0 1 3390
box -6 -8 86 268
use NAND2X1  _1497_
timestamp 0
transform 1 0 4550 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1498_
timestamp 0
transform 1 0 4410 0 -1 3910
box -6 -8 86 268
use INVX1  _1499_
timestamp 0
transform 1 0 4470 0 1 3390
box -6 -8 46 268
use NAND3X1  _1500_
timestamp 0
transform 1 0 4590 0 1 3390
box -6 -8 86 268
use NAND2X1  _1501_
timestamp 0
transform 1 0 4870 0 -1 3910
box -6 -8 66 268
use NOR2X1  _1502_
timestamp 0
transform -1 0 5190 0 -1 3910
box -6 -8 66 268
use NAND2X1  _1503_
timestamp 0
transform -1 0 5070 0 -1 3910
box -6 -8 66 268
use INVX1  _1504_
timestamp 0
transform 1 0 5030 0 1 3910
box -6 -8 46 268
use OAI21X1  _1505_
timestamp 0
transform -1 0 5210 0 1 3910
box -6 -8 86 268
use OR2X2  _1506_
timestamp 0
transform 1 0 5270 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1507_
timestamp 0
transform 1 0 5410 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1508_
timestamp 0
transform -1 0 5510 0 1 3910
box -6 -8 66 268
use NAND3X1  _1509_
timestamp 0
transform 1 0 5690 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1510_
timestamp 0
transform -1 0 5610 0 -1 3910
box -6 -8 66 268
use NAND3X1  _1511_
timestamp 0
transform 1 0 5590 0 1 3910
box -6 -8 86 268
use NAND2X1  _1512_
timestamp 0
transform -1 0 6030 0 1 4430
box -6 -8 66 268
use NOR2X1  _1513_
timestamp 0
transform 1 0 5670 0 -1 3390
box -6 -8 66 268
use NOR2X1  _1514_
timestamp 0
transform 1 0 5970 0 1 3390
box -6 -8 66 268
use NAND3X1  _1515_
timestamp 0
transform 1 0 5630 0 1 3390
box -6 -8 86 268
use NAND2X1  _1516_
timestamp 0
transform -1 0 6310 0 -1 3390
box -6 -8 66 268
use AOI22X1  _1517_
timestamp 0
transform 1 0 5790 0 1 3390
box -6 -8 106 268
use AOI21X1  _1518_
timestamp 0
transform 1 0 5810 0 1 4430
box -6 -8 86 268
use NAND2X1  _1519_
timestamp 0
transform 1 0 6230 0 1 3390
box -6 -8 66 268
use OAI21X1  _1520_
timestamp 0
transform 1 0 5910 0 -1 270
box -6 -8 86 268
use AOI21X1  _1521_
timestamp 0
transform 1 0 5790 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1522_
timestamp 0
transform -1 0 6030 0 -1 3390
box -6 -8 86 268
use AOI22X1  _1523_
timestamp 0
transform 1 0 6090 0 1 4430
box -6 -8 106 268
use OAI21X1  _1524_
timestamp 0
transform -1 0 6090 0 1 4950
box -6 -8 86 268
use OR2X2  _1525_
timestamp 0
transform 1 0 1970 0 1 5990
box -6 -8 86 268
use NAND3X1  _1526_
timestamp 0
transform 1 0 2230 0 -1 5990
box -6 -8 86 268
use INVX1  _1527_
timestamp 0
transform 1 0 1710 0 -1 2350
box -6 -8 46 268
use OAI21X1  _1528_
timestamp 0
transform 1 0 1190 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1529_
timestamp 0
transform 1 0 1570 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1530_
timestamp 0
transform 1 0 2130 0 1 5470
box -6 -8 66 268
use OAI21X1  _1531_
timestamp 0
transform -1 0 2390 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1532_
timestamp 0
transform 1 0 2410 0 1 5470
box -6 -8 86 268
use AOI22X1  _1533_
timestamp 0
transform -1 0 2490 0 -1 5990
box -6 -8 106 268
use INVX1  _1534_
timestamp 0
transform 1 0 5050 0 -1 5470
box -6 -8 46 268
use INVX1  _1535_
timestamp 0
transform 1 0 5370 0 -1 4950
box -6 -8 46 268
use NAND2X1  _1536_
timestamp 0
transform -1 0 6310 0 1 4430
box -6 -8 66 268
use INVX1  _1537_
timestamp 0
transform 1 0 6090 0 -1 5470
box -6 -8 46 268
use AOI21X1  _1538_
timestamp 0
transform 1 0 5290 0 1 3910
box -6 -8 86 268
use OAI21X1  _1539_
timestamp 0
transform 1 0 4530 0 -1 3390
box -6 -8 86 268
use NOR2X1  _1540_
timestamp 0
transform 1 0 4090 0 1 3910
box -6 -8 66 268
use NAND3X1  _1541_
timestamp 0
transform 1 0 4470 0 -1 4430
box -6 -8 86 268
use OAI22X1  _1542_
timestamp 0
transform -1 0 4310 0 1 3910
box -6 -8 106 268
use NAND2X1  _1543_
timestamp 0
transform 1 0 4390 0 1 3910
box -6 -8 66 268
use XNOR2X1  _1544_
timestamp 0
transform -1 0 4790 0 -1 3910
box -6 -8 126 268
use XOR2X1  _1545_
timestamp 0
transform 1 0 5090 0 -1 4430
box -6 -8 126 268
use XOR2X1  _1546_
timestamp 0
transform 1 0 5550 0 -1 4430
box -6 -8 126 268
use NOR2X1  _1547_
timestamp 0
transform -1 0 6150 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1548_
timestamp 0
transform -1 0 6310 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1549_
timestamp 0
transform 1 0 5950 0 -1 4950
box -6 -8 86 268
use NAND3X1  _1550_
timestamp 0
transform 1 0 5650 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1551_
timestamp 0
transform 1 0 1990 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1552_
timestamp 0
transform 1 0 2370 0 -1 2870
box -6 -8 86 268
use INVX1  _1553_
timestamp 0
transform 1 0 3510 0 1 5470
box -6 -8 46 268
use AOI21X1  _1554_
timestamp 0
transform -1 0 4230 0 -1 5470
box -6 -8 86 268
use AOI21X1  _1555_
timestamp 0
transform 1 0 4110 0 1 4950
box -6 -8 86 268
use AOI22X1  _1556_
timestamp 0
transform 1 0 5350 0 1 4950
box -6 -8 106 268
use INVX1  _1557_
timestamp 0
transform -1 0 4630 0 -1 5470
box -6 -8 46 268
use NAND3X1  _1558_
timestamp 0
transform 1 0 5910 0 -1 4430
box -6 -8 86 268
use INVX1  _1559_
timestamp 0
transform 1 0 6070 0 -1 4430
box -6 -8 46 268
use NAND3X1  _1560_
timestamp 0
transform -1 0 6250 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1561_
timestamp 0
transform -1 0 5750 0 1 4430
box -6 -8 66 268
use OAI21X1  _1562_
timestamp 0
transform 1 0 5530 0 1 4430
box -6 -8 86 268
use INVX1  _1563_
timestamp 0
transform -1 0 5450 0 1 4430
box -6 -8 46 268
use INVX1  _1564_
timestamp 0
transform 1 0 4810 0 1 3910
box -6 -8 46 268
use NAND2X1  _1565_
timestamp 0
transform 1 0 4670 0 1 3910
box -6 -8 66 268
use OAI21X1  _1566_
timestamp 0
transform 1 0 4530 0 1 3910
box -6 -8 86 268
use OAI21X1  _1567_
timestamp 0
transform 1 0 3930 0 1 3910
box -6 -8 86 268
use XOR2X1  _1568_
timestamp 0
transform 1 0 4890 0 -1 4430
box -6 -8 126 268
use NAND3X1  _1569_
timestamp 0
transform -1 0 5350 0 1 4430
box -6 -8 86 268
use AOI21X1  _1570_
timestamp 0
transform -1 0 5830 0 -1 4430
box -6 -8 86 268
use INVX1  _1571_
timestamp 0
transform 1 0 5270 0 -1 4430
box -6 -8 46 268
use OAI21X1  _1572_
timestamp 0
transform -1 0 5470 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1573_
timestamp 0
transform -1 0 5290 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1574_
timestamp 0
transform 1 0 2150 0 -1 2350
box -6 -8 66 268
use NOR2X1  _1575_
timestamp 0
transform 1 0 2090 0 1 2350
box -6 -8 66 268
use AOI21X1  _1576_
timestamp 0
transform -1 0 2290 0 1 2350
box -6 -8 86 268
use OAI21X1  _1577_
timestamp 0
transform 1 0 2230 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1578_
timestamp 0
transform -1 0 2030 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1579_
timestamp 0
transform 1 0 2110 0 -1 5990
box -6 -8 66 268
use AOI21X1  _1580_
timestamp 0
transform 1 0 2470 0 -1 5470
box -6 -8 86 268
use AOI22X1  _1581_
timestamp 0
transform -1 0 4530 0 -1 5470
box -6 -8 106 268
use INVX1  _1582_
timestamp 0
transform 1 0 4970 0 -1 4950
box -6 -8 46 268
use AOI21X1  _1583_
timestamp 0
transform -1 0 5190 0 1 4430
box -6 -8 86 268
use NAND3X1  _1584_
timestamp 0
transform 1 0 4610 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1585_
timestamp 0
transform -1 0 4830 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1586_
timestamp 0
transform 1 0 5070 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1587_
timestamp 0
transform 1 0 2650 0 1 1830
box -6 -8 66 268
use XNOR2X1  _1588_
timestamp 0
transform 1 0 2690 0 -1 2350
box -6 -8 126 268
use NAND2X1  _1589_
timestamp 0
transform -1 0 3030 0 1 4950
box -6 -8 66 268
use OAI21X1  _1590_
timestamp 0
transform -1 0 3130 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1591_
timestamp 0
transform 1 0 3470 0 -1 4950
box -6 -8 86 268
use AOI22X1  _1592_
timestamp 0
transform -1 0 4890 0 -1 4950
box -6 -8 106 268
use NAND2X1  _1593_
timestamp 0
transform -1 0 2810 0 1 3390
box -6 -8 66 268
use OAI21X1  _1594_
timestamp 0
transform 1 0 2890 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1595_
timestamp 0
transform 1 0 2610 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1596_
timestamp 0
transform 1 0 2450 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1597_
timestamp 0
transform -1 0 4250 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1598_
timestamp 0
transform 1 0 4050 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1599_
timestamp 0
transform -1 0 2870 0 1 4430
box -6 -8 66 268
use OAI21X1  _1600_
timestamp 0
transform 1 0 2670 0 1 4430
box -6 -8 86 268
use NAND2X1  _1601_
timestamp 0
transform 1 0 3790 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1602_
timestamp 0
transform 1 0 3630 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1603_
timestamp 0
transform 1 0 2910 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1604_
timestamp 0
transform 1 0 2850 0 1 3910
box -6 -8 86 268
use NAND2X1  _1605_
timestamp 0
transform 1 0 3630 0 -1 5470
box -6 -8 66 268
use OAI21X1  _1606_
timestamp 0
transform 1 0 3490 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1607_
timestamp 0
transform -1 0 3390 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1608_
timestamp 0
transform -1 0 3710 0 -1 4950
box -6 -8 86 268
use DFFSR  _1609_
timestamp 0
transform -1 0 2670 0 -1 3910
box -6 -8 466 268
use DFFSR  _1610_
timestamp 0
transform -1 0 2670 0 1 3390
box -6 -8 466 268
use DFFSR  _1611_
timestamp 0
transform -1 0 4570 0 1 4430
box -6 -8 466 268
use DFFSR  _1612_
timestamp 0
transform -1 0 2590 0 1 4430
box -6 -8 466 268
use DFFSR  _1613_
timestamp 0
transform -1 0 3970 0 -1 4430
box -6 -8 466 268
use DFFSR  _1614_
timestamp 0
transform -1 0 2830 0 -1 4430
box -6 -8 466 268
use DFFSR  _1615_
timestamp 0
transform 1 0 3030 0 1 4950
box -6 -8 466 268
use DFFSR  _1616_
timestamp 0
transform -1 0 4570 0 -1 4950
box -6 -8 466 268
use DFFSR  _1617_
timestamp 0
transform 1 0 3950 0 1 5990
box -6 -8 466 268
use DFFSR  _1618_
timestamp 0
transform -1 0 2750 0 1 5990
box -6 -8 466 268
use DFFSR  _1619_
timestamp 0
transform 1 0 3350 0 1 5990
box -6 -8 466 268
use DFFSR  _1620_
timestamp 0
transform 1 0 5550 0 -1 5470
box -6 -8 466 268
use DFFSR  _1621_
timestamp 0
transform -1 0 3350 0 1 5990
box -6 -8 466 268
use DFFSR  _1622_
timestamp 0
transform -1 0 5550 0 -1 5470
box -6 -8 466 268
use DFFSR  _1623_
timestamp 0
transform 1 0 4170 0 1 5470
box -6 -8 466 268
use DFFSR  _1624_
timestamp 0
transform 1 0 4570 0 1 4430
box -6 -8 466 268
use DFFSR  _1625_
timestamp 0
transform 1 0 3110 0 -1 3910
box -6 -8 466 268
use DFFSR  _1626_
timestamp 0
transform 1 0 2810 0 1 3390
box -6 -8 466 268
use DFFSR  _1627_
timestamp 0
transform -1 0 3850 0 1 3910
box -6 -8 466 268
use DFFSR  _1628_
timestamp 0
transform 1 0 2870 0 1 4430
box -6 -8 466 268
use DFFSR  _1629_
timestamp 0
transform 1 0 3270 0 1 3390
box -6 -8 466 268
use DFFSR  _1630_
timestamp 0
transform -1 0 3390 0 1 3910
box -6 -8 466 268
use DFFSR  _1631_
timestamp 0
transform -1 0 3410 0 -1 5470
box -6 -8 466 268
use DFFSR  _1632_
timestamp 0
transform -1 0 3950 0 1 4950
box -6 -8 466 268
use DFFSR  _1633_
timestamp 0
transform -1 0 4630 0 -1 5990
box -6 -8 466 268
use DFFSR  _1634_
timestamp 0
transform -1 0 5230 0 1 5990
box -6 -8 466 268
use DFFSR  _1635_
timestamp 0
transform -1 0 5650 0 1 5470
box -6 -8 466 268
use INVX1  _1636_
timestamp 0
transform -1 0 290 0 1 3390
box -6 -8 46 268
use INVX4  _1637_
timestamp 0
transform 1 0 70 0 1 4430
box -6 -8 66 268
use OAI21X1  _1638_
timestamp 0
transform -1 0 170 0 1 3390
box -6 -8 86 268
use NOR2X1  _1639_
timestamp 0
transform -1 0 150 0 -1 3390
box -6 -8 66 268
use INVX1  _1640_
timestamp 0
transform 1 0 770 0 1 3390
box -6 -8 46 268
use INVX2  _1641_
timestamp 0
transform 1 0 1110 0 1 2870
box -6 -8 46 268
use NAND2X1  _1642_
timestamp 0
transform 1 0 490 0 -1 3910
box -6 -8 66 268
use INVX2  _1643_
timestamp 0
transform -1 0 1030 0 -1 3390
box -6 -8 46 268
use NAND2X1  _1644_
timestamp 0
transform 1 0 970 0 1 2870
box -6 -8 66 268
use NAND2X1  _1645_
timestamp 0
transform -1 0 670 0 -1 2870
box -6 -8 66 268
use AOI22X1  _1646_
timestamp 0
transform 1 0 790 0 1 2870
box -6 -8 106 268
use INVX2  _1647_
timestamp 0
transform 1 0 210 0 1 4430
box -6 -8 46 268
use INVX1  _1648_
timestamp 0
transform -1 0 290 0 -1 2870
box -6 -8 46 268
use INVX1  _1649_
timestamp 0
transform -1 0 570 0 1 3910
box -6 -8 46 268
use OAI21X1  _1650_
timestamp 0
transform 1 0 70 0 1 2870
box -6 -8 86 268
use NAND2X1  _1651_
timestamp 0
transform -1 0 290 0 1 2870
box -6 -8 66 268
use NAND2X1  _1652_
timestamp 0
transform -1 0 430 0 -1 3390
box -6 -8 66 268
use OAI21X1  _1653_
timestamp 0
transform -1 0 710 0 1 2870
box -6 -8 86 268
use OAI21X1  _1654_
timestamp 0
transform -1 0 570 0 1 3390
box -6 -8 86 268
use AOI21X1  _1655_
timestamp 0
transform 1 0 630 0 1 3390
box -6 -8 86 268
use NOR2X1  _1656_
timestamp 0
transform 1 0 390 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1657_
timestamp 0
transform 1 0 890 0 1 3390
box -6 -8 86 268
use OAI21X1  _1658_
timestamp 0
transform 1 0 1170 0 1 3390
box -6 -8 86 268
use XOR2X1  _1659_
timestamp 0
transform 1 0 1530 0 -1 3910
box -6 -8 126 268
use NOR2X1  _1660_
timestamp 0
transform -1 0 1110 0 1 3390
box -6 -8 66 268
use OAI21X1  _1661_
timestamp 0
transform -1 0 1390 0 1 3390
box -6 -8 86 268
use NAND2X1  _1662_
timestamp 0
transform 1 0 1830 0 1 2870
box -6 -8 66 268
use NAND3X1  _1663_
timestamp 0
transform -1 0 1590 0 1 2870
box -6 -8 86 268
use AOI22X1  _1664_
timestamp 0
transform 1 0 1350 0 1 2870
box -6 -8 106 268
use INVX1  _1665_
timestamp 0
transform -1 0 1790 0 -1 2870
box -6 -8 46 268
use NOR2X1  _1666_
timestamp 0
transform 1 0 1610 0 -1 2870
box -6 -8 66 268
use OAI21X1  _1667_
timestamp 0
transform 1 0 1470 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1668_
timestamp 0
transform 1 0 1670 0 1 2870
box -6 -8 86 268
use OAI21X1  _1669_
timestamp 0
transform 1 0 1090 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1670_
timestamp 0
transform 1 0 1250 0 -1 3390
box -6 -8 86 268
use INVX1  _1671_
timestamp 0
transform -1 0 1770 0 -1 3390
box -6 -8 46 268
use OAI21X1  _1672_
timestamp 0
transform 1 0 1410 0 -1 3390
box -6 -8 86 268
use MUX2X1  _1673_
timestamp 0
transform -1 0 1670 0 -1 3390
box -6 -8 106 268
use NAND2X1  _1674_
timestamp 0
transform -1 0 1510 0 1 3390
box -6 -8 66 268
use INVX1  _1675_
timestamp 0
transform -1 0 410 0 1 3390
box -6 -8 46 268
use OAI21X1  _1676_
timestamp 0
transform 1 0 210 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1677_
timestamp 0
transform -1 0 910 0 -1 3390
box -6 -8 86 268
use MUX2X1  _1678_
timestamp 0
transform 1 0 90 0 -1 2870
box -6 -8 106 268
use NAND2X1  _1679_
timestamp 0
transform 1 0 490 0 -1 2870
box -6 -8 66 268
use NAND2X1  _1680_
timestamp 0
transform -1 0 430 0 -1 2870
box -6 -8 66 268
use AOI21X1  _1681_
timestamp 0
transform -1 0 570 0 1 2870
box -6 -8 86 268
use NAND2X1  _1682_
timestamp 0
transform -1 0 410 0 1 2870
box -6 -8 66 268
use NAND3X1  _1683_
timestamp 0
transform 1 0 510 0 -1 3390
box -6 -8 86 268
use AOI22X1  _1684_
timestamp 0
transform -1 0 750 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1685_
timestamp 0
transform 1 0 1590 0 1 3390
box -6 -8 86 268
use OAI21X1  _1686_
timestamp 0
transform 1 0 1850 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1687_
timestamp 0
transform 1 0 2010 0 1 3390
box -6 -8 66 268
use NAND2X1  _1688_
timestamp 0
transform 1 0 1890 0 -1 3910
box -6 -8 66 268
use INVX1  _1689_
timestamp 0
transform 1 0 2030 0 -1 4430
box -6 -8 46 268
use NOR2X1  _1690_
timestamp 0
transform -1 0 1790 0 1 3390
box -6 -8 66 268
use OAI21X1  _1691_
timestamp 0
transform 1 0 1870 0 1 3390
box -6 -8 86 268
use NAND2X1  _1692_
timestamp 0
transform 1 0 1030 0 1 3910
box -6 -8 66 268
use NAND3X1  _1693_
timestamp 0
transform -1 0 1450 0 -1 3910
box -6 -8 86 268
use AOI22X1  _1694_
timestamp 0
transform 1 0 1190 0 -1 3910
box -6 -8 106 268
use INVX1  _1695_
timestamp 0
transform 1 0 770 0 -1 3910
box -6 -8 46 268
use NOR2X1  _1696_
timestamp 0
transform -1 0 950 0 -1 3910
box -6 -8 66 268
use OAI21X1  _1697_
timestamp 0
transform -1 0 1110 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1698_
timestamp 0
transform -1 0 1230 0 1 3910
box -6 -8 86 268
use OAI21X1  _1699_
timestamp 0
transform 1 0 630 0 -1 3910
box -6 -8 86 268
use AOI21X1  _1700_
timestamp 0
transform 1 0 630 0 1 3910
box -6 -8 86 268
use OAI21X1  _1701_
timestamp 0
transform 1 0 1310 0 1 3910
box -6 -8 86 268
use OAI21X1  _1702_
timestamp 0
transform -1 0 1550 0 1 3910
box -6 -8 86 268
use XOR2X1  _1703_
timestamp 0
transform -1 0 2370 0 -1 4430
box -6 -8 126 268
use INVX1  _1704_
timestamp 0
transform 1 0 2230 0 1 4950
box -6 -8 46 268
use INVX1  _1705_
timestamp 0
transform 1 0 770 0 1 3910
box -6 -8 46 268
use OAI21X1  _1706_
timestamp 0
transform -1 0 970 0 1 3910
box -6 -8 86 268
use INVX1  _1707_
timestamp 0
transform -1 0 1830 0 1 3910
box -6 -8 46 268
use AOI22X1  _1708_
timestamp 0
transform 1 0 1610 0 1 3910
box -6 -8 106 268
use NAND2X1  _1709_
timestamp 0
transform -1 0 1570 0 1 4430
box -6 -8 66 268
use AND2X2  _1710_
timestamp 0
transform -1 0 1850 0 1 4430
box -6 -8 86 268
use NAND2X1  _1711_
timestamp 0
transform -1 0 1690 0 1 4430
box -6 -8 66 268
use AOI22X1  _1712_
timestamp 0
transform 1 0 1330 0 1 4430
box -6 -8 106 268
use OAI21X1  _1713_
timestamp 0
transform -1 0 1650 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1714_
timestamp 0
transform 1 0 1430 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1715_
timestamp 0
transform -1 0 1210 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1716_
timestamp 0
transform -1 0 1350 0 -1 4950
box -6 -8 86 268
use OAI21X1  _1717_
timestamp 0
transform 1 0 1250 0 1 4950
box -6 -8 86 268
use OAI21X1  _1718_
timestamp 0
transform 1 0 1410 0 1 4950
box -6 -8 86 268
use XOR2X1  _1719_
timestamp 0
transform 1 0 1710 0 -1 4950
box -6 -8 126 268
use XNOR2X1  _1720_
timestamp 0
transform 1 0 1730 0 1 4950
box -6 -8 126 268
use NAND2X1  _1721_
timestamp 0
transform 1 0 2130 0 -1 4430
box -6 -8 66 268
use NAND3X1  _1722_
timestamp 0
transform -1 0 1810 0 -1 3910
box -6 -8 86 268
use NAND3X1  _1723_
timestamp 0
transform -1 0 1950 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1724_
timestamp 0
transform -1 0 2130 0 -1 5470
box -6 -8 66 268
use OAI21X1  _1725_
timestamp 0
transform -1 0 1650 0 1 4950
box -6 -8 86 268
use INVX1  _1726_
timestamp 0
transform 1 0 1670 0 -1 5470
box -6 -8 46 268
use OAI21X1  _1727_
timestamp 0
transform -1 0 1870 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1728_
timestamp 0
transform -1 0 1250 0 1 4430
box -6 -8 66 268
use AND2X2  _1729_
timestamp 0
transform -1 0 1790 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1730_
timestamp 0
transform 1 0 1450 0 -1 4430
box -6 -8 66 268
use AOI22X1  _1731_
timestamp 0
transform 1 0 1110 0 -1 4430
box -6 -8 106 268
use OAI21X1  _1732_
timestamp 0
transform -1 0 1650 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1733_
timestamp 0
transform -1 0 1370 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1734_
timestamp 0
transform 1 0 930 0 1 4950
box -6 -8 86 268
use AOI21X1  _1735_
timestamp 0
transform -1 0 1170 0 1 4950
box -6 -8 86 268
use OAI21X1  _1736_
timestamp 0
transform 1 0 1230 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1737_
timestamp 0
transform 1 0 1370 0 -1 5470
box -6 -8 86 268
use INVX1  _1738_
timestamp 0
transform 1 0 1530 0 1 5470
box -6 -8 46 268
use XOR2X1  _1739_
timestamp 0
transform -1 0 1770 0 1 5470
box -6 -8 126 268
use INVX1  _1740_
timestamp 0
transform 1 0 1250 0 1 5470
box -6 -8 46 268
use AOI21X1  _1741_
timestamp 0
transform -1 0 1450 0 1 5470
box -6 -8 86 268
use NAND2X1  _1742_
timestamp 0
transform 1 0 370 0 -1 4430
box -6 -8 66 268
use AND2X2  _1743_
timestamp 0
transform -1 0 1010 0 1 4430
box -6 -8 86 268
use NAND2X1  _1744_
timestamp 0
transform 1 0 830 0 -1 4430
box -6 -8 66 268
use AOI22X1  _1745_
timestamp 0
transform -1 0 590 0 -1 4430
box -6 -8 106 268
use OAI21X1  _1746_
timestamp 0
transform -1 0 850 0 1 4430
box -6 -8 86 268
use OAI21X1  _1747_
timestamp 0
transform -1 0 750 0 -1 4430
box -6 -8 86 268
use OAI21X1  _1748_
timestamp 0
transform -1 0 870 0 1 4950
box -6 -8 86 268
use AOI21X1  _1749_
timestamp 0
transform 1 0 650 0 1 4950
box -6 -8 86 268
use OAI21X1  _1750_
timestamp 0
transform 1 0 590 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1751_
timestamp 0
transform 1 0 750 0 -1 5470
box -6 -8 86 268
use INVX1  _1752_
timestamp 0
transform 1 0 970 0 1 5470
box -6 -8 46 268
use XOR2X1  _1753_
timestamp 0
transform -1 0 1190 0 1 5470
box -6 -8 126 268
use INVX1  _1754_
timestamp 0
transform 1 0 3010 0 1 5470
box -6 -8 46 268
use OAI21X1  _1755_
timestamp 0
transform -1 0 890 0 1 5470
box -6 -8 86 268
use INVX1  _1756_
timestamp 0
transform -1 0 270 0 1 4950
box -6 -8 46 268
use AND2X2  _1757_
timestamp 0
transform -1 0 930 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1758_
timestamp 0
transform 1 0 630 0 1 4430
box -6 -8 66 268
use AOI22X1  _1759_
timestamp 0
transform -1 0 570 0 1 4430
box -6 -8 106 268
use OAI21X1  _1760_
timestamp 0
transform -1 0 770 0 -1 4950
box -6 -8 86 268
use OAI22X1  _1761_
timestamp 0
transform 1 0 510 0 -1 4950
box -6 -8 106 268
use OAI21X1  _1762_
timestamp 0
transform 1 0 350 0 1 4950
box -6 -8 86 268
use AOI21X1  _1763_
timestamp 0
transform -1 0 570 0 1 4950
box -6 -8 86 268
use OAI21X1  _1764_
timestamp 0
transform -1 0 630 0 1 5470
box -6 -8 86 268
use OAI21X1  _1765_
timestamp 0
transform -1 0 470 0 1 5470
box -6 -8 86 268
use NAND2X1  _1766_
timestamp 0
transform 1 0 690 0 1 5470
box -6 -8 66 268
use INVX1  _1767_
timestamp 0
transform 1 0 2210 0 -1 5470
box -6 -8 46 268
use AOI21X1  _1768_
timestamp 0
transform -1 0 2150 0 1 4950
box -6 -8 86 268
use AOI21X1  _1769_
timestamp 0
transform -1 0 1990 0 1 4950
box -6 -8 86 268
use OAI21X1  _1770_
timestamp 0
transform 1 0 1530 0 -1 5470
box -6 -8 86 268
use OR2X2  _1771_
timestamp 0
transform 1 0 890 0 -1 5470
box -6 -8 86 268
use AOI22X1  _1772_
timestamp 0
transform 1 0 1050 0 -1 5470
box -6 -8 106 268
use INVX1  _1773_
timestamp 0
transform 1 0 370 0 -1 5990
box -6 -8 46 268
use NAND2X1  _1774_
timestamp 0
transform -1 0 1210 0 -1 5990
box -6 -8 66 268
use NAND2X1  _1775_
timestamp 0
transform -1 0 1350 0 -1 5990
box -6 -8 66 268
use OAI21X1  _1776_
timestamp 0
transform -1 0 690 0 -1 5990
box -6 -8 86 268
use NAND2X1  _1777_
timestamp 0
transform -1 0 150 0 1 3910
box -6 -8 66 268
use AND2X2  _1778_
timestamp 0
transform -1 0 310 0 -1 4430
box -6 -8 86 268
use NAND2X1  _1779_
timestamp 0
transform 1 0 190 0 -1 3910
box -6 -8 66 268
use AOI22X1  _1780_
timestamp 0
transform -1 0 430 0 -1 3910
box -6 -8 106 268
use OAI21X1  _1781_
timestamp 0
transform 1 0 370 0 1 3910
box -6 -8 86 268
use OAI21X1  _1782_
timestamp 0
transform -1 0 290 0 1 3910
box -6 -8 86 268
use OAI21X1  _1783_
timestamp 0
transform -1 0 170 0 -1 4950
box -6 -8 86 268
use AOI21X1  _1784_
timestamp 0
transform -1 0 150 0 1 4950
box -6 -8 86 268
use OAI21X1  _1785_
timestamp 0
transform -1 0 170 0 -1 5470
box -6 -8 86 268
use OAI21X1  _1786_
timestamp 0
transform 1 0 90 0 1 5470
box -6 -8 86 268
use NAND2X1  _1787_
timestamp 0
transform -1 0 810 0 -1 5990
box -6 -8 66 268
use NAND2X1  _1788_
timestamp 0
transform -1 0 550 0 -1 5990
box -6 -8 66 268
use INVX1  _1789_
timestamp 0
transform 1 0 90 0 1 5990
box -6 -8 46 268
use NAND3X1  _1790_
timestamp 0
transform 1 0 550 0 1 5990
box -6 -8 86 268
use NAND2X1  _1791_
timestamp 0
transform 1 0 1030 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1792_
timestamp 0
transform 1 0 1890 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1793_
timestamp 0
transform 1 0 1950 0 -1 5470
box -6 -8 66 268
use NOR2X1  _1794_
timestamp 0
transform -1 0 1910 0 1 5470
box -6 -8 66 268
use NAND3X1  _1795_
timestamp 0
transform 1 0 1410 0 -1 5990
box -6 -8 86 268
use NOR2X1  _1796_
timestamp 0
transform 1 0 1850 0 -1 5990
box -6 -8 66 268
use AND2X2  _1797_
timestamp 0
transform 1 0 1970 0 1 5470
box -6 -8 86 268
use NAND3X1  _1798_
timestamp 0
transform 1 0 410 0 1 5990
box -6 -8 86 268
use NAND2X1  _1799_
timestamp 0
transform 1 0 710 0 1 5990
box -6 -8 66 268
use NAND2X1  _1800_
timestamp 0
transform -1 0 1150 0 1 5990
box -6 -8 66 268
use NAND2X1  _1801_
timestamp 0
transform -1 0 1630 0 -1 5990
box -6 -8 66 268
use NOR2X1  _1802_
timestamp 0
transform -1 0 390 0 1 4430
box -6 -8 66 268
use OAI21X1  _1803_
timestamp 0
transform -1 0 310 0 1 5470
box -6 -8 86 268
use NOR2X1  _1804_
timestamp 0
transform 1 0 90 0 -1 5990
box -6 -8 66 268
use AOI21X1  _1805_
timestamp 0
transform -1 0 290 0 -1 5990
box -6 -8 86 268
use XOR2X1  _1806_
timestamp 0
transform 1 0 210 0 1 5990
box -6 -8 126 268
use OAI21X1  _1807_
timestamp 0
transform -1 0 1310 0 1 5990
box -6 -8 86 268
use NAND3X1  _1808_
timestamp 0
transform -1 0 1770 0 -1 5990
box -6 -8 86 268
use AOI21X1  _1809_
timestamp 0
transform 1 0 250 0 -1 5470
box -6 -8 86 268
use XOR2X1  _1810_
timestamp 0
transform 1 0 410 0 -1 5470
box -6 -8 126 268
use NAND3X1  _1811_
timestamp 0
transform 1 0 870 0 -1 5990
box -6 -8 86 268
use INVX1  _1812_
timestamp 0
transform 1 0 850 0 1 5990
box -6 -8 46 268
use NAND3X1  _1813_
timestamp 0
transform 1 0 950 0 1 5990
box -6 -8 86 268
use NAND2X1  _1814_
timestamp 0
transform 1 0 1390 0 1 5990
box -6 -8 66 268
use NAND3X1  _1815_
timestamp 0
transform 1 0 1670 0 1 5990
box -6 -8 86 268
use NAND3X1  _1816_
timestamp 0
transform 1 0 1510 0 1 5990
box -6 -8 86 268
use NAND2X1  _1817_
timestamp 0
transform -1 0 1890 0 1 5990
box -6 -8 66 268
use BUFX2  _1818_
timestamp 0
transform 1 0 4710 0 1 5990
box -6 -8 66 268
use BUFX2  _1819_
timestamp 0
transform -1 0 2170 0 1 5990
box -6 -8 66 268
use BUFX2  _1820_
timestamp 0
transform 1 0 3890 0 1 5990
box -6 -8 66 268
use BUFX2  _1821_
timestamp 0
transform 1 0 6190 0 -1 5470
box -6 -8 66 268
use BUFX2  _1822_
timestamp 0
transform 1 0 2830 0 1 5990
box -6 -8 66 268
use BUFX2  _1823_
timestamp 0
transform -1 0 4910 0 1 5470
box -6 -8 66 268
use BUFX2  _1824_
timestamp 0
transform -1 0 4630 0 1 5990
box -6 -8 66 268
use BUFX2  _1825_
timestamp 0
transform -1 0 5110 0 1 4950
box -6 -8 66 268
use BUFX2  _1826_
timestamp 0
transform 1 0 6190 0 -1 5990
box -6 -8 66 268
use BUFX2  _1827_
timestamp 0
transform 1 0 6150 0 1 5470
box -6 -8 66 268
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 2470 0 -1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert1
timestamp 0
transform -1 0 1990 0 1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 2410 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 2530 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert4
timestamp 0
transform -1 0 970 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 1030 0 -1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 2210 0 1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 2430 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 3770 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 2910 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 3610 0 1 5470
box -6 -8 66 268
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 3210 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert17
timestamp 0
transform 1 0 4050 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 3090 0 -1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 3110 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 3310 0 -1 5990
box -6 -8 66 268
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 3890 0 -1 5470
box -6 -8 66 268
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 2950 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 3150 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 3030 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert25
timestamp 0
transform -1 0 3110 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert26
timestamp 0
transform -1 0 4070 0 -1 5470
box -6 -8 66 268
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 2210 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert28
timestamp 0
transform 1 0 2330 0 1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert29
timestamp 0
transform 1 0 4050 0 -1 3910
box -6 -8 66 268
use BUFX2  BUFX2_insert30
timestamp 0
transform 1 0 2750 0 -1 3390
box -6 -8 66 268
use BUFX2  BUFX2_insert31
timestamp 0
transform -1 0 1870 0 1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert32
timestamp 0
transform 1 0 1950 0 1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert33
timestamp 0
transform -1 0 3230 0 -1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert34
timestamp 0
transform 1 0 2550 0 -1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert35
timestamp 0
transform -1 0 2350 0 1 2870
box -6 -8 66 268
use BUFX2  BUFX2_insert36
timestamp 0
transform 1 0 1450 0 1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert37
timestamp 0
transform -1 0 1270 0 1 2350
box -6 -8 66 268
use BUFX2  BUFX2_insert38
timestamp 0
transform -1 0 310 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert39
timestamp 0
transform -1 0 1050 0 -1 4950
box -6 -8 66 268
use BUFX2  BUFX2_insert40
timestamp 0
transform -1 0 1030 0 -1 4430
box -6 -8 66 268
use BUFX2  BUFX2_insert41
timestamp 0
transform 1 0 90 0 -1 4430
box -6 -8 66 268
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 3850 0 1 4430
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform 1 0 4550 0 1 4950
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform 1 0 4810 0 -1 5470
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert11
timestamp 0
transform -1 0 3430 0 1 5470
box -6 -8 186 268
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform -1 0 3590 0 1 4430
box -6 -8 186 268
use FILL  FILL92550x58650
timestamp 0
transform 1 0 6170 0 1 3910
box -6 -8 26 268
use FILL  FILL92850x4050
timestamp 0
transform 1 0 6190 0 1 270
box -6 -8 26 268
use FILL  FILL92850x58650
timestamp 0
transform 1 0 6190 0 1 3910
box -6 -8 26 268
use FILL  FILL93150x4050
timestamp 0
transform 1 0 6210 0 1 270
box -6 -8 26 268
use FILL  FILL93150x7950
timestamp 0
transform -1 0 6230 0 -1 790
box -6 -8 26 268
use FILL  FILL93150x35250
timestamp 0
transform 1 0 6210 0 1 2350
box -6 -8 26 268
use FILL  FILL93150x58650
timestamp 0
transform 1 0 6210 0 1 3910
box -6 -8 26 268
use FILL  FILL93150x74250
timestamp 0
transform 1 0 6210 0 1 4950
box -6 -8 26 268
use FILL  FILL93150x82050
timestamp 0
transform 1 0 6210 0 1 5470
box -6 -8 26 268
use FILL  FILL93450x4050
timestamp 0
transform 1 0 6230 0 1 270
box -6 -8 26 268
use FILL  FILL93450x7950
timestamp 0
transform -1 0 6250 0 -1 790
box -6 -8 26 268
use FILL  FILL93450x35250
timestamp 0
transform 1 0 6230 0 1 2350
box -6 -8 26 268
use FILL  FILL93450x58650
timestamp 0
transform 1 0 6230 0 1 3910
box -6 -8 26 268
use FILL  FILL93450x74250
timestamp 0
transform 1 0 6230 0 1 4950
box -6 -8 26 268
use FILL  FILL93450x82050
timestamp 0
transform 1 0 6230 0 1 5470
box -6 -8 26 268
use FILL  FILL93750x150
timestamp 0
transform -1 0 6270 0 -1 270
box -6 -8 26 268
use FILL  FILL93750x4050
timestamp 0
transform 1 0 6250 0 1 270
box -6 -8 26 268
use FILL  FILL93750x7950
timestamp 0
transform -1 0 6270 0 -1 790
box -6 -8 26 268
use FILL  FILL93750x35250
timestamp 0
transform 1 0 6250 0 1 2350
box -6 -8 26 268
use FILL  FILL93750x58650
timestamp 0
transform 1 0 6250 0 1 3910
box -6 -8 26 268
use FILL  FILL93750x62550
timestamp 0
transform -1 0 6270 0 -1 4430
box -6 -8 26 268
use FILL  FILL93750x74250
timestamp 0
transform 1 0 6250 0 1 4950
box -6 -8 26 268
use FILL  FILL93750x78150
timestamp 0
transform -1 0 6270 0 -1 5470
box -6 -8 26 268
use FILL  FILL93750x82050
timestamp 0
transform 1 0 6250 0 1 5470
box -6 -8 26 268
use FILL  FILL93750x85950
timestamp 0
transform -1 0 6270 0 -1 5990
box -6 -8 26 268
use FILL  FILL94050x150
timestamp 0
transform -1 0 6290 0 -1 270
box -6 -8 26 268
use FILL  FILL94050x4050
timestamp 0
transform 1 0 6270 0 1 270
box -6 -8 26 268
use FILL  FILL94050x7950
timestamp 0
transform -1 0 6290 0 -1 790
box -6 -8 26 268
use FILL  FILL94050x35250
timestamp 0
transform 1 0 6270 0 1 2350
box -6 -8 26 268
use FILL  FILL94050x58650
timestamp 0
transform 1 0 6270 0 1 3910
box -6 -8 26 268
use FILL  FILL94050x62550
timestamp 0
transform -1 0 6290 0 -1 4430
box -6 -8 26 268
use FILL  FILL94050x74250
timestamp 0
transform 1 0 6270 0 1 4950
box -6 -8 26 268
use FILL  FILL94050x78150
timestamp 0
transform -1 0 6290 0 -1 5470
box -6 -8 26 268
use FILL  FILL94050x82050
timestamp 0
transform 1 0 6270 0 1 5470
box -6 -8 26 268
use FILL  FILL94050x85950
timestamp 0
transform -1 0 6290 0 -1 5990
box -6 -8 26 268
use FILL  FILL94350x150
timestamp 0
transform -1 0 6310 0 -1 270
box -6 -8 26 268
use FILL  FILL94350x4050
timestamp 0
transform 1 0 6290 0 1 270
box -6 -8 26 268
use FILL  FILL94350x7950
timestamp 0
transform -1 0 6310 0 -1 790
box -6 -8 26 268
use FILL  FILL94350x11850
timestamp 0
transform 1 0 6290 0 1 790
box -6 -8 26 268
use FILL  FILL94350x19650
timestamp 0
transform 1 0 6290 0 1 1310
box -6 -8 26 268
use FILL  FILL94350x27450
timestamp 0
transform 1 0 6290 0 1 1830
box -6 -8 26 268
use FILL  FILL94350x35250
timestamp 0
transform 1 0 6290 0 1 2350
box -6 -8 26 268
use FILL  FILL94350x39150
timestamp 0
transform -1 0 6310 0 -1 2870
box -6 -8 26 268
use FILL  FILL94350x43050
timestamp 0
transform 1 0 6290 0 1 2870
box -6 -8 26 268
use FILL  FILL94350x50850
timestamp 0
transform 1 0 6290 0 1 3390
box -6 -8 26 268
use FILL  FILL94350x58650
timestamp 0
transform 1 0 6290 0 1 3910
box -6 -8 26 268
use FILL  FILL94350x62550
timestamp 0
transform -1 0 6310 0 -1 4430
box -6 -8 26 268
use FILL  FILL94350x74250
timestamp 0
transform 1 0 6290 0 1 4950
box -6 -8 26 268
use FILL  FILL94350x78150
timestamp 0
transform -1 0 6310 0 -1 5470
box -6 -8 26 268
use FILL  FILL94350x82050
timestamp 0
transform 1 0 6290 0 1 5470
box -6 -8 26 268
use FILL  FILL94350x85950
timestamp 0
transform -1 0 6310 0 -1 5990
box -6 -8 26 268
use FILL  FILL94350x89850
timestamp 0
transform 1 0 6290 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__889_
timestamp 0
transform -1 0 3950 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__890_
timestamp 0
transform 1 0 3510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__891_
timestamp 0
transform -1 0 4650 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__892_
timestamp 0
transform 1 0 4910 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__893_
timestamp 0
transform -1 0 3650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__894_
timestamp 0
transform -1 0 4750 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__895_
timestamp 0
transform -1 0 3830 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__896_
timestamp 0
transform 1 0 3670 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__897_
timestamp 0
transform 1 0 5530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__898_
timestamp 0
transform -1 0 4070 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__899_
timestamp 0
transform 1 0 5030 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__900_
timestamp 0
transform -1 0 6070 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__901_
timestamp 0
transform 1 0 5910 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__902_
timestamp 0
transform -1 0 5530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__903_
timestamp 0
transform 1 0 4630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__904_
timestamp 0
transform -1 0 4030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__905_
timestamp 0
transform -1 0 5250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__906_
timestamp 0
transform 1 0 4850 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__907_
timestamp 0
transform -1 0 3070 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__908_
timestamp 0
transform -1 0 6210 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__909_
timestamp 0
transform 1 0 5790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__910_
timestamp 0
transform -1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__911_
timestamp 0
transform 1 0 4770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__912_
timestamp 0
transform 1 0 4630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__913_
timestamp 0
transform 1 0 5630 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__914_
timestamp 0
transform -1 0 5390 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__915_
timestamp 0
transform 1 0 4230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__916_
timestamp 0
transform 1 0 5790 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__917_
timestamp 0
transform 1 0 5990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__918_
timestamp 0
transform -1 0 5370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__919_
timestamp 0
transform -1 0 5250 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__920_
timestamp 0
transform -1 0 5970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__921_
timestamp 0
transform -1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform 1 0 5090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform -1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform -1 0 5670 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform -1 0 2810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform 1 0 1950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform -1 0 2370 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform -1 0 2690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform 1 0 1150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform -1 0 2110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform -1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform 1 0 3850 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform 1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform 1 0 3950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform 1 0 1010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform 1 0 1950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform -1 0 2010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__938_
timestamp 0
transform -1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__939_
timestamp 0
transform 1 0 3230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__940_
timestamp 0
transform -1 0 3390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__941_
timestamp 0
transform 1 0 1830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__942_
timestamp 0
transform -1 0 2090 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__943_
timestamp 0
transform -1 0 2230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__944_
timestamp 0
transform -1 0 2850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__945_
timestamp 0
transform -1 0 2650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__946_
timestamp 0
transform -1 0 2770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__947_
timestamp 0
transform 1 0 3830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__948_
timestamp 0
transform 1 0 4190 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__949_
timestamp 0
transform 1 0 4310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__950_
timestamp 0
transform -1 0 3910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__951_
timestamp 0
transform 1 0 890 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__952_
timestamp 0
transform -1 0 2490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__953_
timestamp 0
transform 1 0 1550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__954_
timestamp 0
transform -1 0 1830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__955_
timestamp 0
transform -1 0 1690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__956_
timestamp 0
transform -1 0 630 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform 1 0 430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform -1 0 490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform 1 0 10 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform 1 0 170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform -1 0 270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform -1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform 1 0 530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform 1 0 950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform -1 0 510 0 1 790
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform -1 0 790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform -1 0 2710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform 1 0 390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform 1 0 10 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform 1 0 590 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform -1 0 470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform -1 0 310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform 1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform 1 0 1290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform -1 0 1090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform -1 0 1670 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform -1 0 1830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform 1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform -1 0 950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform 1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform 1 0 630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform 1 0 130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform -1 0 1610 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform 1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform -1 0 1430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform -1 0 1530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform 1 0 650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform 1 0 770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform -1 0 910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform 1 0 1270 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform -1 0 1390 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform -1 0 650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform 1 0 10 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform 1 0 150 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform -1 0 1210 0 1 270
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform -1 0 1370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform -1 0 910 0 1 270
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform 1 0 1410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform 1 0 1510 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform 1 0 2610 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform 1 0 1750 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 3590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform -1 0 1390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform 1 0 1610 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 1370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 3330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform 1 0 1190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform -1 0 1050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform 1 0 750 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform 1 0 1050 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform 1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform 1 0 2270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform 1 0 470 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform 1 0 1510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform 1 0 2710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 3150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 3210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform -1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform -1 0 3010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 2770 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform 1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 3110 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform 1 0 2970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 3250 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 3390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform -1 0 3610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 1030 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform -1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform -1 0 2710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform -1 0 1910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform -1 0 2670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 2030 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform -1 0 2550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 2190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 1290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform 1 0 1950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform -1 0 2090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform 1 0 2230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform -1 0 2470 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform 1 0 2390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 2550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform -1 0 1750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform 1 0 2050 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform 1 0 3750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 2410 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform -1 0 2210 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform 1 0 1170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform -1 0 310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform 1 0 2830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 2690 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 2390 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 2650 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform -1 0 2130 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform -1 0 1690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 1790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 1650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 1770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform -1 0 2530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform 1 0 1330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 2070 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 2690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform -1 0 2010 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 3630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 2230 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform 1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform 1 0 3550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 3410 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 3530 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform -1 0 3730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 3270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform 1 0 3830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 3710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform 1 0 3790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform 1 0 4130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform 1 0 4210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform 1 0 3850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform 1 0 3690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform -1 0 3310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform 1 0 3410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform -1 0 2830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 2910 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform -1 0 3070 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 3110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 3530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform 1 0 3530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform -1 0 3210 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform 1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 3150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 3910 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 4330 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform 1 0 3250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform 1 0 3890 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform 1 0 4050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform 1 0 4050 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform -1 0 4490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform 1 0 2330 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 3910 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 4190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 3270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 3670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform -1 0 4950 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform -1 0 2810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 4830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 4670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform -1 0 4590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform -1 0 4970 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform -1 0 4790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform -1 0 5090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 4550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 4470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 4330 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform -1 0 3450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform -1 0 3130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform -1 0 4070 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 4630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform -1 0 4810 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform -1 0 4390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform -1 0 3910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform 1 0 1470 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform -1 0 3750 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform -1 0 3610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform -1 0 2510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform 1 0 3310 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform 1 0 2650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform -1 0 2830 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform -1 0 3330 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform -1 0 3010 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 2450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 2190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform 1 0 10 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform -1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform -1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 10 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform -1 0 350 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform 1 0 10 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform -1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform 1 0 170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform 1 0 590 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform 1 0 430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 910 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform 1 0 1830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 1950 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform 1 0 1610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 2010 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform -1 0 3470 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform 1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 3170 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform 1 0 770 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform 1 0 310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform -1 0 1950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform 1 0 10 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform 1 0 170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform -1 0 750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform -1 0 190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 310 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform -1 0 1170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform -1 0 1110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform -1 0 750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform 1 0 1490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform 1 0 1650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform -1 0 2550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 1750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform 1 0 990 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform -1 0 1130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform 1 0 310 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform 1 0 470 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 1810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform 1 0 1250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform -1 0 630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform 1 0 770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform 1 0 890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform 1 0 1010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform 1 0 970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform 1 0 790 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 1270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform 1 0 1670 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform 1 0 1330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform 1 0 1530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 1750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 2050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 1990 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform 1 0 2210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform -1 0 2830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 3450 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 5050 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 4070 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 3410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform -1 0 5090 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 4270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform 1 0 3430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform -1 0 4870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 4430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform -1 0 4950 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform 1 0 4970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform -1 0 4730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform 1 0 5130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform 1 0 5370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 4370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 3650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform -1 0 2310 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform -1 0 3390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 2450 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 3090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform 1 0 3510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 3890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform -1 0 3270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 3070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 3670 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 4010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 4610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform 1 0 3950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform -1 0 3870 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform 1 0 4090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform -1 0 4390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 3930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform 1 0 3970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 4310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 4650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform -1 0 4750 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 4550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform -1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 4810 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform 1 0 5170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 4630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform 1 0 4830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 4490 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform 1 0 5210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform -1 0 5170 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 5670 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform 1 0 5330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform 1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform -1 0 5770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform 1 0 4950 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform 1 0 4210 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 5510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform -1 0 4510 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform -1 0 5930 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform -1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform -1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform 1 0 4650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform 1 0 5230 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 5470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 3730 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 5390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform -1 0 6070 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 5610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform 1 0 5690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform -1 0 2570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform -1 0 2530 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform -1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform 1 0 2470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform 1 0 2370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 2510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform -1 0 3710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 3750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 2170 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform 1 0 3950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform 1 0 5110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform -1 0 5630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform -1 0 2870 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform 1 0 1970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 2430 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 2270 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform -1 0 2250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 2110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 2130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 2290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform -1 0 5590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 5590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 6170 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform 1 0 5990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 5270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform -1 0 6230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform 1 0 5470 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform 1 0 5630 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform 1 0 4170 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 4450 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform 1 0 3370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform -1 0 3250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform 1 0 3490 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform 1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 5350 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform -1 0 4270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 4950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform 1 0 3150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform -1 0 2610 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform 1 0 2590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform -1 0 3010 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 2610 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform -1 0 2770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 2710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 2870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform -1 0 2730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 3990 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform -1 0 3590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 2910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 3310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 3210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 3430 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform 1 0 2870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 3370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 3510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform -1 0 5130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform -1 0 5430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 4670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 5130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 5410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform -1 0 5570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform 1 0 4990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform -1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform 1 0 5690 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform 1 0 5890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 5970 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform 1 0 5830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform 1 0 5530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform 1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 5570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform -1 0 5730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 5890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 6130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform 1 0 5830 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 6010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 6170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 6130 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform 1 0 5090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 5670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 6010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform -1 0 6070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform -1 0 5890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 6030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform 1 0 5410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 5290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 5450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 1890 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 1950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform 1 0 2050 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform -1 0 1950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform 1 0 2690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform 1 0 2610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 3390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 5770 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 5930 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform 1 0 5990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform 1 0 5710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform -1 0 6210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 4910 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 5230 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform -1 0 5630 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 5590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 3790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform 1 0 4510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform 1 0 3770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 3050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform -1 0 3930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform 1 0 4050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform 1 0 4630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 3810 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform -1 0 3970 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform 1 0 4070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform 1 0 4790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 4290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 3650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform 1 0 3910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform -1 0 3350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform -1 0 3750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform 1 0 4370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform 1 0 4210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 4210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform 1 0 4670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform 1 0 4510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform 1 0 4830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 5090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 4670 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform -1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 4170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 4290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform 1 0 5010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform 1 0 5550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 5290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform 1 0 4830 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 4370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 4230 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform 1 0 4510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform 1 0 5330 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform 1 0 5890 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 5390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 5470 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform -1 0 6190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 6150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform 1 0 5730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 6050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform -1 0 6070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform -1 0 6170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 6070 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 5850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform 1 0 5910 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform -1 0 6210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform -1 0 5930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform -1 0 5790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform -1 0 2210 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform 1 0 2490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 1090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform 1 0 2390 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 2610 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform 1 0 2750 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 3110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform -1 0 6110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 4410 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 5410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 6050 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform 1 0 4370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform 1 0 5290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform 1 0 5170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform 1 0 3730 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 4610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 4470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform 1 0 4030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform 1 0 4710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform 1 0 4590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 5010 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform 1 0 4850 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 5010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform -1 0 4850 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1452_
timestamp 0
transform -1 0 3630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1453_
timestamp 0
transform 1 0 3850 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1454_
timestamp 0
transform 1 0 3730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1455_
timestamp 0
transform 1 0 4230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1456_
timestamp 0
transform 1 0 4250 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1457_
timestamp 0
transform 1 0 4330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1458_
timestamp 0
transform -1 0 4750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1459_
timestamp 0
transform 1 0 4910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 4890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 5290 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1462_
timestamp 0
transform 1 0 4930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1463_
timestamp 0
transform 1 0 5030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1464_
timestamp 0
transform 1 0 5130 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 5450 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1466_
timestamp 0
transform 1 0 5030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1467_
timestamp 0
transform 1 0 5130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1468_
timestamp 0
transform 1 0 5190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1469_
timestamp 0
transform -1 0 5350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1470_
timestamp 0
transform 1 0 5750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1471_
timestamp 0
transform 1 0 5250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1472_
timestamp 0
transform 1 0 5410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1473_
timestamp 0
transform 1 0 5470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1474_
timestamp 0
transform -1 0 6050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1475_
timestamp 0
transform -1 0 5950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1476_
timestamp 0
transform -1 0 6070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1477_
timestamp 0
transform -1 0 5690 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1478_
timestamp 0
transform 1 0 5790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1479_
timestamp 0
transform -1 0 5750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1480_
timestamp 0
transform 1 0 830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 870 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1482_
timestamp 0
transform -1 0 1010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1483_
timestamp 0
transform 1 0 2090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1485_
timestamp 0
transform 1 0 4570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1486_
timestamp 0
transform -1 0 5790 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1487_
timestamp 0
transform -1 0 2510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 4670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 4850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1490_
timestamp 0
transform 1 0 3850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 3490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1492_
timestamp 0
transform 1 0 3890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1493_
timestamp 0
transform -1 0 4050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1494_
timestamp 0
transform 1 0 4190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1495_
timestamp 0
transform -1 0 4130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1496_
timestamp 0
transform 1 0 4090 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1497_
timestamp 0
transform 1 0 4490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 4330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1499_
timestamp 0
transform 1 0 4410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1500_
timestamp 0
transform 1 0 4510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1501_
timestamp 0
transform 1 0 4790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1502_
timestamp 0
transform -1 0 5090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1503_
timestamp 0
transform -1 0 4950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1504_
timestamp 0
transform 1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1505_
timestamp 0
transform -1 0 5090 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1506_
timestamp 0
transform 1 0 5190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 5350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1508_
timestamp 0
transform -1 0 5390 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1509_
timestamp 0
transform 1 0 5610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1510_
timestamp 0
transform -1 0 5510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1511_
timestamp 0
transform 1 0 5510 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1512_
timestamp 0
transform -1 0 5910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1513_
timestamp 0
transform 1 0 5610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1514_
timestamp 0
transform 1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1515_
timestamp 0
transform 1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1516_
timestamp 0
transform -1 0 6190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1517_
timestamp 0
transform 1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1518_
timestamp 0
transform 1 0 5750 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1519_
timestamp 0
transform 1 0 6150 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1520_
timestamp 0
transform 1 0 5830 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1521_
timestamp 0
transform 1 0 5730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1522_
timestamp 0
transform -1 0 5890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 6030 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1524_
timestamp 0
transform -1 0 5950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1525_
timestamp 0
transform 1 0 1890 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1526_
timestamp 0
transform 1 0 2170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 1630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 1130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1529_
timestamp 0
transform 1 0 1490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 2050 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1531_
timestamp 0
transform -1 0 2270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1532_
timestamp 0
transform 1 0 2330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 2330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1534_
timestamp 0
transform 1 0 4990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1535_
timestamp 0
transform 1 0 5290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1536_
timestamp 0
transform -1 0 6210 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1537_
timestamp 0
transform 1 0 6010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1538_
timestamp 0
transform 1 0 5210 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1539_
timestamp 0
transform 1 0 4470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1540_
timestamp 0
transform 1 0 4010 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1541_
timestamp 0
transform 1 0 4390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1542_
timestamp 0
transform -1 0 4170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1543_
timestamp 0
transform 1 0 4310 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1544_
timestamp 0
transform -1 0 4630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1545_
timestamp 0
transform 1 0 5010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 5470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1547_
timestamp 0
transform -1 0 6050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1548_
timestamp 0
transform -1 0 6170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1549_
timestamp 0
transform 1 0 5890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1550_
timestamp 0
transform 1 0 5570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1551_
timestamp 0
transform 1 0 1910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1552_
timestamp 0
transform 1 0 2310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1553_
timestamp 0
transform 1 0 3430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1554_
timestamp 0
transform -1 0 4090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1555_
timestamp 0
transform 1 0 4050 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1556_
timestamp 0
transform 1 0 5270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1557_
timestamp 0
transform -1 0 4550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1558_
timestamp 0
transform 1 0 5830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1559_
timestamp 0
transform 1 0 5990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1560_
timestamp 0
transform -1 0 6130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1561_
timestamp 0
transform -1 0 5630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1562_
timestamp 0
transform 1 0 5450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 5370 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1564_
timestamp 0
transform 1 0 4730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 4610 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1566_
timestamp 0
transform 1 0 4450 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1567_
timestamp 0
transform 1 0 3850 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1568_
timestamp 0
transform 1 0 4830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 5210 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1570_
timestamp 0
transform -1 0 5690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1571_
timestamp 0
transform 1 0 5210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1572_
timestamp 0
transform -1 0 5330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1573_
timestamp 0
transform -1 0 5170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1574_
timestamp 0
transform 1 0 2070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1575_
timestamp 0
transform 1 0 2010 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1576_
timestamp 0
transform -1 0 2170 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1577_
timestamp 0
transform 1 0 2150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1578_
timestamp 0
transform -1 0 1930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1579_
timestamp 0
transform 1 0 2030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 2390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 4390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1582_
timestamp 0
transform 1 0 4890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 5050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1584_
timestamp 0
transform 1 0 4550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1585_
timestamp 0
transform -1 0 4710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1586_
timestamp 0
transform 1 0 5010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1587_
timestamp 0
transform 1 0 2570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1588_
timestamp 0
transform 1 0 2610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 2930 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1590_
timestamp 0
transform -1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1591_
timestamp 0
transform 1 0 3390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1592_
timestamp 0
transform -1 0 4750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1593_
timestamp 0
transform -1 0 2690 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1594_
timestamp 0
transform 1 0 2830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1595_
timestamp 0
transform 1 0 2530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1596_
timestamp 0
transform 1 0 2370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1597_
timestamp 0
transform -1 0 4150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1598_
timestamp 0
transform 1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1599_
timestamp 0
transform -1 0 2770 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1600_
timestamp 0
transform 1 0 2590 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1601_
timestamp 0
transform 1 0 3710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1602_
timestamp 0
transform 1 0 3570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1603_
timestamp 0
transform 1 0 2830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1604_
timestamp 0
transform 1 0 2770 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 3570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1606_
timestamp 0
transform 1 0 3410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1607_
timestamp 0
transform -1 0 3290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1608_
timestamp 0
transform -1 0 3570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1636_
timestamp 0
transform -1 0 190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1637_
timestamp 0
transform 1 0 10 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1638_
timestamp 0
transform -1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1639_
timestamp 0
transform -1 0 30 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 710 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1641_
timestamp 0
transform 1 0 1030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1642_
timestamp 0
transform 1 0 430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1643_
timestamp 0
transform -1 0 930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1644_
timestamp 0
transform 1 0 890 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1645_
timestamp 0
transform -1 0 570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1646_
timestamp 0
transform 1 0 710 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1647_
timestamp 0
transform 1 0 130 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1648_
timestamp 0
transform -1 0 210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1649_
timestamp 0
transform -1 0 470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1650_
timestamp 0
transform 1 0 10 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1651_
timestamp 0
transform -1 0 170 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1652_
timestamp 0
transform -1 0 310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1653_
timestamp 0
transform -1 0 590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1654_
timestamp 0
transform -1 0 430 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1655_
timestamp 0
transform 1 0 570 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1656_
timestamp 0
transform 1 0 310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1657_
timestamp 0
transform 1 0 810 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 1110 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1659_
timestamp 0
transform 1 0 1450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1660_
timestamp 0
transform -1 0 990 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1661_
timestamp 0
transform -1 0 1270 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1662_
timestamp 0
transform 1 0 1750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1663_
timestamp 0
transform -1 0 1470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1664_
timestamp 0
transform 1 0 1270 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1665_
timestamp 0
transform -1 0 1690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1666_
timestamp 0
transform 1 0 1550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1667_
timestamp 0
transform 1 0 1390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1668_
timestamp 0
transform 1 0 1590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1669_
timestamp 0
transform 1 0 1030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1670_
timestamp 0
transform 1 0 1170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1671_
timestamp 0
transform -1 0 1690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1672_
timestamp 0
transform 1 0 1330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1673_
timestamp 0
transform -1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1674_
timestamp 0
transform -1 0 1410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1675_
timestamp 0
transform -1 0 310 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1676_
timestamp 0
transform 1 0 150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1677_
timestamp 0
transform -1 0 770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1678_
timestamp 0
transform 1 0 10 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1679_
timestamp 0
transform 1 0 430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1680_
timestamp 0
transform -1 0 310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1681_
timestamp 0
transform -1 0 430 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1682_
timestamp 0
transform -1 0 310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1683_
timestamp 0
transform 1 0 430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1684_
timestamp 0
transform -1 0 610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1685_
timestamp 0
transform 1 0 1510 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1686_
timestamp 0
transform 1 0 1770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1687_
timestamp 0
transform 1 0 1950 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1688_
timestamp 0
transform 1 0 1810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1689_
timestamp 0
transform 1 0 1950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1690_
timestamp 0
transform -1 0 1690 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1691_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1692_
timestamp 0
transform 1 0 970 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1693_
timestamp 0
transform -1 0 1310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1694_
timestamp 0
transform 1 0 1110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1695_
timestamp 0
transform 1 0 710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1696_
timestamp 0
transform -1 0 830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1698_
timestamp 0
transform -1 0 1110 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1699_
timestamp 0
transform 1 0 550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1700_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1701_
timestamp 0
transform 1 0 1230 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1702_
timestamp 0
transform -1 0 1410 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1703_
timestamp 0
transform -1 0 2210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1704_
timestamp 0
transform 1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1705_
timestamp 0
transform 1 0 710 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1706_
timestamp 0
transform -1 0 830 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1707_
timestamp 0
transform -1 0 1730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1708_
timestamp 0
transform 1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1709_
timestamp 0
transform -1 0 1450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1710_
timestamp 0
transform -1 0 1710 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1711_
timestamp 0
transform -1 0 1590 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1712_
timestamp 0
transform 1 0 1250 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1714_
timestamp 0
transform 1 0 1350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1715_
timestamp 0
transform -1 0 1070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1716_
timestamp 0
transform -1 0 1230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1717_
timestamp 0
transform 1 0 1170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1718_
timestamp 0
transform 1 0 1330 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1719_
timestamp 0
transform 1 0 1650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1720_
timestamp 0
transform 1 0 1650 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1721_
timestamp 0
transform 1 0 2070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1722_
timestamp 0
transform -1 0 1670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1723_
timestamp 0
transform -1 0 1810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1724_
timestamp 0
transform -1 0 2030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1725_
timestamp 0
transform -1 0 1510 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1726_
timestamp 0
transform 1 0 1610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1727_
timestamp 0
transform -1 0 1730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1728_
timestamp 0
transform -1 0 1130 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1729_
timestamp 0
transform -1 0 1670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1730_
timestamp 0
transform 1 0 1370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1731_
timestamp 0
transform 1 0 1030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1732_
timestamp 0
transform -1 0 1530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1733_
timestamp 0
transform -1 0 1230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1734_
timestamp 0
transform 1 0 870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1735_
timestamp 0
transform -1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1736_
timestamp 0
transform 1 0 1150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1737_
timestamp 0
transform 1 0 1310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1738_
timestamp 0
transform 1 0 1450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1739_
timestamp 0
transform -1 0 1590 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1740_
timestamp 0
transform 1 0 1190 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1741_
timestamp 0
transform -1 0 1310 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1742_
timestamp 0
transform 1 0 310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1743_
timestamp 0
transform -1 0 870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1744_
timestamp 0
transform 1 0 750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1745_
timestamp 0
transform -1 0 450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1746_
timestamp 0
transform -1 0 710 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1747_
timestamp 0
transform -1 0 610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1748_
timestamp 0
transform -1 0 750 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1749_
timestamp 0
transform 1 0 570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1750_
timestamp 0
transform 1 0 530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1751_
timestamp 0
transform 1 0 670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1752_
timestamp 0
transform 1 0 890 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1753_
timestamp 0
transform -1 0 1030 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1754_
timestamp 0
transform 1 0 2930 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1755_
timestamp 0
transform -1 0 770 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1756_
timestamp 0
transform -1 0 170 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1757_
timestamp 0
transform -1 0 790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1758_
timestamp 0
transform 1 0 570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1759_
timestamp 0
transform -1 0 410 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1760_
timestamp 0
transform -1 0 630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1761_
timestamp 0
transform 1 0 450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1762_
timestamp 0
transform 1 0 270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1763_
timestamp 0
transform -1 0 450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1764_
timestamp 0
transform -1 0 490 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1765_
timestamp 0
transform -1 0 330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1766_
timestamp 0
transform 1 0 630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1767_
timestamp 0
transform 1 0 2130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1768_
timestamp 0
transform -1 0 2010 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1769_
timestamp 0
transform -1 0 1870 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1770_
timestamp 0
transform 1 0 1450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1771_
timestamp 0
transform 1 0 830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1772_
timestamp 0
transform 1 0 970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1773_
timestamp 0
transform 1 0 290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1774_
timestamp 0
transform -1 0 1110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1775_
timestamp 0
transform -1 0 1230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1776_
timestamp 0
transform -1 0 570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1777_
timestamp 0
transform -1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1778_
timestamp 0
transform -1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1779_
timestamp 0
transform 1 0 130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1780_
timestamp 0
transform -1 0 270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1781_
timestamp 0
transform 1 0 290 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1782_
timestamp 0
transform -1 0 170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1783_
timestamp 0
transform -1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1784_
timestamp 0
transform -1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1785_
timestamp 0
transform -1 0 30 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1786_
timestamp 0
transform 1 0 10 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1787_
timestamp 0
transform -1 0 710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1788_
timestamp 0
transform -1 0 430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1789_
timestamp 0
transform 1 0 10 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1790_
timestamp 0
transform 1 0 490 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1791_
timestamp 0
transform 1 0 950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1792_
timestamp 0
transform 1 0 1830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1793_
timestamp 0
transform 1 0 1870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1794_
timestamp 0
transform -1 0 1790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1795_
timestamp 0
transform 1 0 1350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1796_
timestamp 0
transform 1 0 1770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1797_
timestamp 0
transform 1 0 1910 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1798_
timestamp 0
transform 1 0 330 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1799_
timestamp 0
transform 1 0 630 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1800_
timestamp 0
transform -1 0 1050 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1801_
timestamp 0
transform -1 0 1510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1802_
timestamp 0
transform -1 0 270 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1803_
timestamp 0
transform -1 0 190 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1804_
timestamp 0
transform 1 0 10 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1805_
timestamp 0
transform -1 0 170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 130 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1807_
timestamp 0
transform -1 0 1170 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1808_
timestamp 0
transform -1 0 1650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1809_
timestamp 0
transform 1 0 170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1810_
timestamp 0
transform 1 0 330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1811_
timestamp 0
transform 1 0 810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1812_
timestamp 0
transform 1 0 770 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 890 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1814_
timestamp 0
transform 1 0 1310 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 1590 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1816_
timestamp 0
transform 1 0 1450 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1817_
timestamp 0
transform -1 0 1770 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1818_
timestamp 0
transform 1 0 4630 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1819_
timestamp 0
transform -1 0 2070 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1820_
timestamp 0
transform 1 0 3810 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1821_
timestamp 0
transform 1 0 6130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1822_
timestamp 0
transform 1 0 2750 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1823_
timestamp 0
transform -1 0 4790 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1824_
timestamp 0
transform -1 0 4530 0 1 5990
box -6 -8 26 268
use FILL  FILL_0__1825_
timestamp 0
transform -1 0 4990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1826_
timestamp 0
transform 1 0 6130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1827_
timestamp 0
transform 1 0 6070 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 2390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform -1 0 1870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 2350 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 2450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform -1 0 850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 2090 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 2370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 3710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 2830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 3550 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 3130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform 1 0 3970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 2990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 3250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 3810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 2830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform 1 0 3090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 2950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform -1 0 2990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform -1 0 3970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 2090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform 1 0 2270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert29
timestamp 0
transform 1 0 3970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert30
timestamp 0
transform 1 0 2670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform -1 0 1770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert32
timestamp 0
transform 1 0 1870 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert33
timestamp 0
transform -1 0 3110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert34
timestamp 0
transform 1 0 2490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert35
timestamp 0
transform -1 0 2230 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert36
timestamp 0
transform 1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert37
timestamp 0
transform -1 0 1150 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert38
timestamp 0
transform -1 0 190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert39
timestamp 0
transform -1 0 950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert40
timestamp 0
transform -1 0 910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert41
timestamp 0
transform 1 0 10 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert8
timestamp 0
transform -1 0 3610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert9
timestamp 0
transform 1 0 4470 0 1 4950
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert10
timestamp 0
transform 1 0 4750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert11
timestamp 0
transform -1 0 3190 0 1 5470
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert12
timestamp 0
transform -1 0 3350 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__889_
timestamp 0
transform -1 0 3970 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__890_
timestamp 0
transform 1 0 3530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__891_
timestamp 0
transform -1 0 4670 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__892_
timestamp 0
transform 1 0 4930 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__893_
timestamp 0
transform -1 0 3670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__894_
timestamp 0
transform -1 0 4770 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__895_
timestamp 0
transform -1 0 3850 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__896_
timestamp 0
transform 1 0 3690 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__897_
timestamp 0
transform 1 0 5550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__898_
timestamp 0
transform -1 0 4090 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__899_
timestamp 0
transform 1 0 5050 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__900_
timestamp 0
transform -1 0 6090 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__901_
timestamp 0
transform 1 0 5930 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__902_
timestamp 0
transform -1 0 5550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__903_
timestamp 0
transform 1 0 4650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__904_
timestamp 0
transform -1 0 4050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__905_
timestamp 0
transform -1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__906_
timestamp 0
transform 1 0 4870 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__907_
timestamp 0
transform -1 0 3090 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__908_
timestamp 0
transform -1 0 6230 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__909_
timestamp 0
transform 1 0 5810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__910_
timestamp 0
transform -1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__911_
timestamp 0
transform 1 0 4790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__912_
timestamp 0
transform 1 0 4650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__913_
timestamp 0
transform 1 0 5650 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__914_
timestamp 0
transform -1 0 5410 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__915_
timestamp 0
transform 1 0 4250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__916_
timestamp 0
transform 1 0 5810 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__917_
timestamp 0
transform 1 0 6010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__918_
timestamp 0
transform -1 0 5390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__919_
timestamp 0
transform -1 0 5270 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__920_
timestamp 0
transform -1 0 5990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__921_
timestamp 0
transform -1 0 5850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform 1 0 5110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform -1 0 5690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform -1 0 5690 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform -1 0 2830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform 1 0 1970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform -1 0 2390 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform -1 0 2710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform 1 0 1170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform -1 0 2130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform -1 0 2250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform 1 0 3870 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform 1 0 4270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform 1 0 3970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform 1 0 1030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform 1 0 1970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform -1 0 2030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__938_
timestamp 0
transform -1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__939_
timestamp 0
transform 1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__940_
timestamp 0
transform -1 0 3410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__941_
timestamp 0
transform 1 0 1850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__942_
timestamp 0
transform -1 0 2110 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__943_
timestamp 0
transform -1 0 2250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__944_
timestamp 0
transform -1 0 2870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__945_
timestamp 0
transform -1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__946_
timestamp 0
transform -1 0 2790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__947_
timestamp 0
transform 1 0 3850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__948_
timestamp 0
transform 1 0 4210 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__949_
timestamp 0
transform 1 0 4330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__950_
timestamp 0
transform -1 0 3930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__951_
timestamp 0
transform 1 0 910 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__952_
timestamp 0
transform -1 0 2510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__953_
timestamp 0
transform 1 0 1570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__954_
timestamp 0
transform -1 0 1850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__955_
timestamp 0
transform -1 0 1710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__956_
timestamp 0
transform -1 0 650 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform 1 0 450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform -1 0 510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform 1 0 30 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform 1 0 190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform -1 0 290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform -1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform 1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform 1 0 970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform -1 0 530 0 1 790
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform -1 0 810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform -1 0 2730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform 1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform 1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform 1 0 610 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform -1 0 490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform -1 0 330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform 1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform 1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform -1 0 1110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform -1 0 1690 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform -1 0 1850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform 1 0 1230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform 1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform 1 0 650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform 1 0 150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform -1 0 1630 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform 1 0 1530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform -1 0 1450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform -1 0 1550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform 1 0 670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform 1 0 790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform -1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform 1 0 1290 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform -1 0 1410 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform -1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform 1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform 1 0 170 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform -1 0 1230 0 1 270
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform -1 0 1390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform -1 0 930 0 1 270
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform 1 0 1430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform 1 0 1530 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform 1 0 2630 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform 1 0 1770 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform 1 0 3610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform -1 0 1410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform 1 0 1630 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 1390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform 1 0 3350 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform 1 0 1210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 950 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform -1 0 350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform -1 0 1070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform -1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform 1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform 1 0 1070 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform 1 0 1230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform 1 0 2290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform 1 0 490 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform 1 0 1530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 2990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform 1 0 2730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 3170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 3230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform -1 0 2890 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform -1 0 3030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 2790 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform 1 0 2850 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 3130 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform 1 0 2990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 3270 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 3410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform -1 0 3630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 1050 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform -1 0 2990 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform -1 0 2730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform -1 0 1930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform -1 0 2690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 2570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform -1 0 2570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 2210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 1310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform 1 0 1970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform -1 0 2110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform 1 0 2250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform -1 0 2490 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform 1 0 2410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 2570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform -1 0 1770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform 1 0 2070 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform 1 0 3770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform 1 0 2430 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform -1 0 2230 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform 1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform -1 0 330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform 1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 2710 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 2410 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 2670 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform -1 0 2150 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 1810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform -1 0 1670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform -1 0 2550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform 1 0 1350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform 1 0 2090 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 2710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform -1 0 2030 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 3650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 2250 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform 1 0 3010 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform 1 0 3570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 3430 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform 1 0 3550 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform -1 0 3750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 3290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform 1 0 3850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform 1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 3730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform 1 0 3810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform 1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform 1 0 4230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform 1 0 3870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform 1 0 3710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform 1 0 3730 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform -1 0 3330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform 1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform -1 0 2850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 2930 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform -1 0 3090 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 3130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 3550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform 1 0 3550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform -1 0 3230 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform 1 0 2990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 3170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 3930 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 4350 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform 1 0 3270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform 1 0 3910 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform 1 0 4070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform 1 0 4070 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform -1 0 4510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 4230 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform 1 0 2350 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 3930 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 4210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 3290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform -1 0 3690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform -1 0 4970 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform -1 0 2830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 4850 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 4690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform -1 0 4610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform -1 0 4990 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform -1 0 4810 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform -1 0 5110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 4570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 4490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 4350 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform -1 0 3470 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform -1 0 3150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform -1 0 4090 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 4650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform -1 0 4830 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform -1 0 4410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform -1 0 3930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform 1 0 1490 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform -1 0 3770 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform -1 0 3630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform -1 0 2530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform 1 0 3330 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform 1 0 2670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform -1 0 2850 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform -1 0 3350 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform -1 0 3030 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 2470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 2210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform 1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform -1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform -1 0 650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform -1 0 370 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform 1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform -1 0 1230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform 1 0 190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform 1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform 1 0 450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 930 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform 1 0 1850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 1970 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform 1 0 1630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 2030 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform -1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform 1 0 3170 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 3190 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform 1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform 1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform -1 0 1970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform 1 0 30 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform 1 0 190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform -1 0 770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform -1 0 210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 170 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 330 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform -1 0 1190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform -1 0 1130 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform -1 0 770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform 1 0 1510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform 1 0 1670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform -1 0 2570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 1770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform 1 0 1010 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform -1 0 1150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform 1 0 330 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform 1 0 490 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 1830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform 1 0 1270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform -1 0 650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform 1 0 790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform 1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform 1 0 1030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform 1 0 990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform 1 0 810 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 1290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform 1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform 1 0 1350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform 1 0 1550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 1770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 2070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 2010 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform 1 0 2230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform -1 0 2850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 3470 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 5070 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 4090 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 3430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform -1 0 5110 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 4290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform 1 0 3450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform -1 0 4890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 4450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform -1 0 4970 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform 1 0 4990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform -1 0 4750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform 1 0 5150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform 1 0 5390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 3670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform -1 0 2330 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform -1 0 3410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 2470 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 3110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform 1 0 3530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 3910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform -1 0 3290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 3090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 3690 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 4030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 4630 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform 1 0 3970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform -1 0 3890 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform 1 0 4110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform -1 0 4410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 3950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform 1 0 3990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 4330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform 1 0 4670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform -1 0 4770 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 4570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform -1 0 4150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 4830 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform 1 0 5190 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 4650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform 1 0 4850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 4510 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform 1 0 5230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform -1 0 5190 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 5690 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform 1 0 5350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform -1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform 1 0 4970 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform 1 0 4230 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 5530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 5310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform -1 0 4530 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform -1 0 5950 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform -1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform -1 0 4830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform 1 0 4670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform 1 0 5250 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 5490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 3750 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 5410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform -1 0 6090 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 5630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform 1 0 5710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 5110 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform -1 0 2590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform -1 0 2550 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform -1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform 1 0 2490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform 1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 2530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform -1 0 3730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform -1 0 3770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 2190 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform 1 0 3970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform 1 0 5130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform -1 0 5650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform -1 0 2890 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform 1 0 1990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 2450 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 2290 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform -1 0 2270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 2130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform 1 0 2150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 2310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform -1 0 5610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 5610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 6190 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform 1 0 6010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 5290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform -1 0 6250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform 1 0 5490 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform 1 0 5650 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform 1 0 4190 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 4470 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform 1 0 3390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform -1 0 3270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform 1 0 3510 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform 1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 5370 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform -1 0 4290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 4970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform 1 0 3170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform -1 0 2630 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform 1 0 2610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform -1 0 3030 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 2630 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform -1 0 2790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 2730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 2890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform -1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 4010 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform -1 0 3610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 2930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 3330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 3230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 3450 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform 1 0 2890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform 1 0 3390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 3530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform -1 0 5150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform -1 0 5450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 4690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 5150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 5430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform -1 0 5590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform 1 0 5010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform -1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform 1 0 5710 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform 1 0 5910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 5990 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform 1 0 5850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform 1 0 5550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform 1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 5590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform -1 0 5750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 5910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 6150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform 1 0 5850 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 6030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform -1 0 6190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 6150 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform 1 0 5110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 5690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 6030 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform -1 0 6090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform -1 0 5910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 6050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform 1 0 5430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 5310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 5470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 1910 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 1970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform 1 0 2070 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform -1 0 1970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform 1 0 2710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform 1 0 2630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 3410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform 1 0 5970 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 5950 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform 1 0 6010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform 1 0 5730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform -1 0 6230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 4930 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 5250 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform -1 0 5650 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 5610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 3810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform 1 0 4530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform 1 0 3790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 3070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform -1 0 3950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform 1 0 4070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform 1 0 4650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 3830 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform -1 0 3990 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform 1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform 1 0 4810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform 1 0 4310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 3670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform 1 0 3930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform -1 0 3370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform -1 0 3770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform 1 0 4390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform 1 0 4230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 4230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform 1 0 4690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform 1 0 4530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform 1 0 4850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 5110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 4690 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform -1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 4190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 4310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform 1 0 5030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform 1 0 5570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 5310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform 1 0 4850 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 4390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 4250 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform 1 0 4530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform 1 0 5350 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform 1 0 5910 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 5410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 5490 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 5750 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform -1 0 6210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 6170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform 1 0 5750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 6070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform -1 0 6090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform -1 0 6190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 6090 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 5870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform 1 0 5930 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform -1 0 6230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform -1 0 5950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform -1 0 5810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform -1 0 2230 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform 1 0 2510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform 1 0 1110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform 1 0 2410 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 2630 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform 1 0 2770 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 3130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform -1 0 6130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 4430 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 5430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 6070 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform 1 0 4390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform 1 0 5310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform 1 0 5190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform 1 0 3750 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 4630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 4490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform 1 0 4050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform 1 0 4730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform 1 0 4610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 5030 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform 1 0 4870 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 5030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform -1 0 4870 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1452_
timestamp 0
transform -1 0 3650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1453_
timestamp 0
transform 1 0 3870 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1454_
timestamp 0
transform 1 0 3750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1455_
timestamp 0
transform 1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1456_
timestamp 0
transform 1 0 4270 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1457_
timestamp 0
transform 1 0 4350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1458_
timestamp 0
transform -1 0 4770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1459_
timestamp 0
transform 1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 4910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1461_
timestamp 0
transform 1 0 5310 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1462_
timestamp 0
transform 1 0 4950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1463_
timestamp 0
transform 1 0 5050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1464_
timestamp 0
transform 1 0 5150 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 5470 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1466_
timestamp 0
transform 1 0 5050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1467_
timestamp 0
transform 1 0 5150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1468_
timestamp 0
transform 1 0 5210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1469_
timestamp 0
transform -1 0 5370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1470_
timestamp 0
transform 1 0 5770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1471_
timestamp 0
transform 1 0 5270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1472_
timestamp 0
transform 1 0 5430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1473_
timestamp 0
transform 1 0 5490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1474_
timestamp 0
transform -1 0 6070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1475_
timestamp 0
transform -1 0 5970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1476_
timestamp 0
transform -1 0 6090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1477_
timestamp 0
transform -1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1478_
timestamp 0
transform 1 0 5810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1479_
timestamp 0
transform -1 0 5770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1480_
timestamp 0
transform 1 0 850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 890 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1482_
timestamp 0
transform -1 0 1030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1483_
timestamp 0
transform 1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1485_
timestamp 0
transform 1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1486_
timestamp 0
transform -1 0 5810 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1487_
timestamp 0
transform -1 0 2530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1488_
timestamp 0
transform 1 0 4690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 4870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1490_
timestamp 0
transform 1 0 3870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 3510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1492_
timestamp 0
transform 1 0 3910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1493_
timestamp 0
transform -1 0 4070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1494_
timestamp 0
transform 1 0 4210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1495_
timestamp 0
transform -1 0 4150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1496_
timestamp 0
transform 1 0 4110 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1497_
timestamp 0
transform 1 0 4510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 4350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1499_
timestamp 0
transform 1 0 4430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1500_
timestamp 0
transform 1 0 4530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1501_
timestamp 0
transform 1 0 4810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1502_
timestamp 0
transform -1 0 5110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1503_
timestamp 0
transform -1 0 4970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1504_
timestamp 0
transform 1 0 4970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1505_
timestamp 0
transform -1 0 5110 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1506_
timestamp 0
transform 1 0 5210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1507_
timestamp 0
transform 1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1508_
timestamp 0
transform -1 0 5410 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1509_
timestamp 0
transform 1 0 5630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1510_
timestamp 0
transform -1 0 5530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1511_
timestamp 0
transform 1 0 5530 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1512_
timestamp 0
transform -1 0 5930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1513_
timestamp 0
transform 1 0 5630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1514_
timestamp 0
transform 1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1515_
timestamp 0
transform 1 0 5590 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1516_
timestamp 0
transform -1 0 6210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1517_
timestamp 0
transform 1 0 5730 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1518_
timestamp 0
transform 1 0 5770 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1519_
timestamp 0
transform 1 0 6170 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1520_
timestamp 0
transform 1 0 5850 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1521_
timestamp 0
transform 1 0 5750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1522_
timestamp 0
transform -1 0 5910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1523_
timestamp 0
transform 1 0 6050 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1524_
timestamp 0
transform -1 0 5970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1525_
timestamp 0
transform 1 0 1910 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1526_
timestamp 0
transform 1 0 2190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 1650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 1150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1529_
timestamp 0
transform 1 0 1510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 2070 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1531_
timestamp 0
transform -1 0 2290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1532_
timestamp 0
transform 1 0 2350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 2350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1534_
timestamp 0
transform 1 0 5010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1535_
timestamp 0
transform 1 0 5310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1536_
timestamp 0
transform -1 0 6230 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1537_
timestamp 0
transform 1 0 6030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1538_
timestamp 0
transform 1 0 5230 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1539_
timestamp 0
transform 1 0 4490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1540_
timestamp 0
transform 1 0 4030 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1541_
timestamp 0
transform 1 0 4410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1542_
timestamp 0
transform -1 0 4190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1543_
timestamp 0
transform 1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1544_
timestamp 0
transform -1 0 4650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1545_
timestamp 0
transform 1 0 5030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1546_
timestamp 0
transform 1 0 5490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1547_
timestamp 0
transform -1 0 6070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1548_
timestamp 0
transform -1 0 6190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1549_
timestamp 0
transform 1 0 5910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1550_
timestamp 0
transform 1 0 5590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1551_
timestamp 0
transform 1 0 1930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1552_
timestamp 0
transform 1 0 2330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1553_
timestamp 0
transform 1 0 3450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1554_
timestamp 0
transform -1 0 4110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1555_
timestamp 0
transform 1 0 4070 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1556_
timestamp 0
transform 1 0 5290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1557_
timestamp 0
transform -1 0 4570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1558_
timestamp 0
transform 1 0 5850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1559_
timestamp 0
transform 1 0 6010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1560_
timestamp 0
transform -1 0 6150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1561_
timestamp 0
transform -1 0 5650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1562_
timestamp 0
transform 1 0 5470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 5390 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1564_
timestamp 0
transform 1 0 4750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1566_
timestamp 0
transform 1 0 4470 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1567_
timestamp 0
transform 1 0 3870 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1568_
timestamp 0
transform 1 0 4850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1569_
timestamp 0
transform -1 0 5230 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1570_
timestamp 0
transform -1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1571_
timestamp 0
transform 1 0 5230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1572_
timestamp 0
transform -1 0 5350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1573_
timestamp 0
transform -1 0 5190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1574_
timestamp 0
transform 1 0 2090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1575_
timestamp 0
transform 1 0 2030 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1576_
timestamp 0
transform -1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1577_
timestamp 0
transform 1 0 2170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1578_
timestamp 0
transform -1 0 1950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1579_
timestamp 0
transform 1 0 2050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 2410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1581_
timestamp 0
transform -1 0 4410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1582_
timestamp 0
transform 1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 5070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1584_
timestamp 0
transform 1 0 4570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1585_
timestamp 0
transform -1 0 4730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1586_
timestamp 0
transform 1 0 5030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1587_
timestamp 0
transform 1 0 2590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1588_
timestamp 0
transform 1 0 2630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1589_
timestamp 0
transform -1 0 2950 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1590_
timestamp 0
transform -1 0 3010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1591_
timestamp 0
transform 1 0 3410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1592_
timestamp 0
transform -1 0 4770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1593_
timestamp 0
transform -1 0 2710 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1594_
timestamp 0
transform 1 0 2850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1595_
timestamp 0
transform 1 0 2550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1596_
timestamp 0
transform 1 0 2390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1597_
timestamp 0
transform -1 0 4170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1598_
timestamp 0
transform 1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1599_
timestamp 0
transform -1 0 2790 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1600_
timestamp 0
transform 1 0 2610 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1601_
timestamp 0
transform 1 0 3730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1602_
timestamp 0
transform 1 0 3590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1603_
timestamp 0
transform 1 0 2850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1604_
timestamp 0
transform 1 0 2790 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 3590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1606_
timestamp 0
transform 1 0 3430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1607_
timestamp 0
transform -1 0 3310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1608_
timestamp 0
transform -1 0 3590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1636_
timestamp 0
transform -1 0 210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1637_
timestamp 0
transform 1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1638_
timestamp 0
transform -1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1639_
timestamp 0
transform -1 0 50 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 730 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1641_
timestamp 0
transform 1 0 1050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1642_
timestamp 0
transform 1 0 450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1643_
timestamp 0
transform -1 0 950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1644_
timestamp 0
transform 1 0 910 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1645_
timestamp 0
transform -1 0 590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1646_
timestamp 0
transform 1 0 730 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1647_
timestamp 0
transform 1 0 150 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1648_
timestamp 0
transform -1 0 230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1649_
timestamp 0
transform -1 0 490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1650_
timestamp 0
transform 1 0 30 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1651_
timestamp 0
transform -1 0 190 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1652_
timestamp 0
transform -1 0 330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1653_
timestamp 0
transform -1 0 610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1654_
timestamp 0
transform -1 0 450 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1655_
timestamp 0
transform 1 0 590 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1656_
timestamp 0
transform 1 0 330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1657_
timestamp 0
transform 1 0 830 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1658_
timestamp 0
transform 1 0 1130 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1659_
timestamp 0
transform 1 0 1470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1660_
timestamp 0
transform -1 0 1010 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1661_
timestamp 0
transform -1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1662_
timestamp 0
transform 1 0 1770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1663_
timestamp 0
transform -1 0 1490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1664_
timestamp 0
transform 1 0 1290 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1665_
timestamp 0
transform -1 0 1710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1666_
timestamp 0
transform 1 0 1570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1667_
timestamp 0
transform 1 0 1410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1668_
timestamp 0
transform 1 0 1610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1669_
timestamp 0
transform 1 0 1050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1670_
timestamp 0
transform 1 0 1190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1671_
timestamp 0
transform -1 0 1710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1672_
timestamp 0
transform 1 0 1350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1673_
timestamp 0
transform -1 0 1530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1674_
timestamp 0
transform -1 0 1430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1675_
timestamp 0
transform -1 0 330 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1676_
timestamp 0
transform 1 0 170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1677_
timestamp 0
transform -1 0 790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1678_
timestamp 0
transform 1 0 30 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1679_
timestamp 0
transform 1 0 450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1680_
timestamp 0
transform -1 0 330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1681_
timestamp 0
transform -1 0 450 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1682_
timestamp 0
transform -1 0 330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1683_
timestamp 0
transform 1 0 450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1684_
timestamp 0
transform -1 0 630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1685_
timestamp 0
transform 1 0 1530 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1686_
timestamp 0
transform 1 0 1790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1687_
timestamp 0
transform 1 0 1970 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1688_
timestamp 0
transform 1 0 1830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1689_
timestamp 0
transform 1 0 1970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1690_
timestamp 0
transform -1 0 1710 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1691_
timestamp 0
transform 1 0 1810 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1692_
timestamp 0
transform 1 0 990 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1693_
timestamp 0
transform -1 0 1330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1694_
timestamp 0
transform 1 0 1130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1695_
timestamp 0
transform 1 0 730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1696_
timestamp 0
transform -1 0 850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1697_
timestamp 0
transform -1 0 990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1698_
timestamp 0
transform -1 0 1130 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1699_
timestamp 0
transform 1 0 570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1700_
timestamp 0
transform 1 0 590 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1701_
timestamp 0
transform 1 0 1250 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1702_
timestamp 0
transform -1 0 1430 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1703_
timestamp 0
transform -1 0 2230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1704_
timestamp 0
transform 1 0 2170 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1705_
timestamp 0
transform 1 0 730 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1706_
timestamp 0
transform -1 0 850 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1707_
timestamp 0
transform -1 0 1750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1708_
timestamp 0
transform 1 0 1570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1709_
timestamp 0
transform -1 0 1470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1710_
timestamp 0
transform -1 0 1730 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1711_
timestamp 0
transform -1 0 1610 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1712_
timestamp 0
transform 1 0 1270 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 1550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1714_
timestamp 0
transform 1 0 1370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1715_
timestamp 0
transform -1 0 1090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1716_
timestamp 0
transform -1 0 1250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1717_
timestamp 0
transform 1 0 1190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1718_
timestamp 0
transform 1 0 1350 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1719_
timestamp 0
transform 1 0 1670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1720_
timestamp 0
transform 1 0 1670 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1721_
timestamp 0
transform 1 0 2090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1722_
timestamp 0
transform -1 0 1690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1723_
timestamp 0
transform -1 0 1830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1724_
timestamp 0
transform -1 0 2050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1725_
timestamp 0
transform -1 0 1530 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1726_
timestamp 0
transform 1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1727_
timestamp 0
transform -1 0 1750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1728_
timestamp 0
transform -1 0 1150 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1729_
timestamp 0
transform -1 0 1690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1730_
timestamp 0
transform 1 0 1390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1731_
timestamp 0
transform 1 0 1050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1732_
timestamp 0
transform -1 0 1550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1733_
timestamp 0
transform -1 0 1250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1734_
timestamp 0
transform 1 0 890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1735_
timestamp 0
transform -1 0 1050 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1736_
timestamp 0
transform 1 0 1170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1737_
timestamp 0
transform 1 0 1330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1738_
timestamp 0
transform 1 0 1470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1739_
timestamp 0
transform -1 0 1610 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1740_
timestamp 0
transform 1 0 1210 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1741_
timestamp 0
transform -1 0 1330 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1742_
timestamp 0
transform 1 0 330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1743_
timestamp 0
transform -1 0 890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1744_
timestamp 0
transform 1 0 770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1745_
timestamp 0
transform -1 0 470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1746_
timestamp 0
transform -1 0 730 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1747_
timestamp 0
transform -1 0 630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1748_
timestamp 0
transform -1 0 770 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1749_
timestamp 0
transform 1 0 590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1750_
timestamp 0
transform 1 0 550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1751_
timestamp 0
transform 1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1752_
timestamp 0
transform 1 0 910 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1753_
timestamp 0
transform -1 0 1050 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1754_
timestamp 0
transform 1 0 2950 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1755_
timestamp 0
transform -1 0 790 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1756_
timestamp 0
transform -1 0 190 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1757_
timestamp 0
transform -1 0 810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1758_
timestamp 0
transform 1 0 590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1759_
timestamp 0
transform -1 0 430 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1760_
timestamp 0
transform -1 0 650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1761_
timestamp 0
transform 1 0 470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1762_
timestamp 0
transform 1 0 290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1763_
timestamp 0
transform -1 0 470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1764_
timestamp 0
transform -1 0 510 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1765_
timestamp 0
transform -1 0 350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1766_
timestamp 0
transform 1 0 650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1767_
timestamp 0
transform 1 0 2150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1768_
timestamp 0
transform -1 0 2030 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1769_
timestamp 0
transform -1 0 1890 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1770_
timestamp 0
transform 1 0 1470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1771_
timestamp 0
transform 1 0 850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1772_
timestamp 0
transform 1 0 990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1773_
timestamp 0
transform 1 0 310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1774_
timestamp 0
transform -1 0 1130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1775_
timestamp 0
transform -1 0 1250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1776_
timestamp 0
transform -1 0 590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1777_
timestamp 0
transform -1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1778_
timestamp 0
transform -1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1779_
timestamp 0
transform 1 0 150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1780_
timestamp 0
transform -1 0 290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1781_
timestamp 0
transform 1 0 310 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1782_
timestamp 0
transform -1 0 190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1783_
timestamp 0
transform -1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1784_
timestamp 0
transform -1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1785_
timestamp 0
transform -1 0 50 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1786_
timestamp 0
transform 1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1787_
timestamp 0
transform -1 0 730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1788_
timestamp 0
transform -1 0 450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1789_
timestamp 0
transform 1 0 30 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1790_
timestamp 0
transform 1 0 510 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1791_
timestamp 0
transform 1 0 970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1792_
timestamp 0
transform 1 0 1850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1793_
timestamp 0
transform 1 0 1890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1794_
timestamp 0
transform -1 0 1810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1795_
timestamp 0
transform 1 0 1370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1796_
timestamp 0
transform 1 0 1790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1797_
timestamp 0
transform 1 0 1930 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1798_
timestamp 0
transform 1 0 350 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1799_
timestamp 0
transform 1 0 650 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1800_
timestamp 0
transform -1 0 1070 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1801_
timestamp 0
transform -1 0 1530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1802_
timestamp 0
transform -1 0 290 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1803_
timestamp 0
transform -1 0 210 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1804_
timestamp 0
transform 1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1805_
timestamp 0
transform -1 0 190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1806_
timestamp 0
transform 1 0 150 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1807_
timestamp 0
transform -1 0 1190 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1808_
timestamp 0
transform -1 0 1670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1809_
timestamp 0
transform 1 0 190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1810_
timestamp 0
transform 1 0 350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1811_
timestamp 0
transform 1 0 830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1812_
timestamp 0
transform 1 0 790 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1813_
timestamp 0
transform 1 0 910 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1814_
timestamp 0
transform 1 0 1330 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 1610 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1816_
timestamp 0
transform 1 0 1470 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1817_
timestamp 0
transform -1 0 1790 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1818_
timestamp 0
transform 1 0 4650 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1819_
timestamp 0
transform -1 0 2090 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1820_
timestamp 0
transform 1 0 3830 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1821_
timestamp 0
transform 1 0 6150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1822_
timestamp 0
transform 1 0 2770 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1823_
timestamp 0
transform -1 0 4810 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1824_
timestamp 0
transform -1 0 4550 0 1 5990
box -6 -8 26 268
use FILL  FILL_1__1825_
timestamp 0
transform -1 0 5010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1826_
timestamp 0
transform 1 0 6150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1827_
timestamp 0
transform 1 0 6090 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform 1 0 2410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform -1 0 1890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 2370 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 2470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform -1 0 870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 2110 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 2390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 3730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 2850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 3570 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 3150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform 1 0 3990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 3010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform -1 0 3010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 3270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 3830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 2850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform 1 0 3110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 2970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform -1 0 3010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform -1 0 3990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 2110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform 1 0 2290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert29
timestamp 0
transform 1 0 3990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert30
timestamp 0
transform 1 0 2690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert31
timestamp 0
transform -1 0 1790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert32
timestamp 0
transform 1 0 1890 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert33
timestamp 0
transform -1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert34
timestamp 0
transform 1 0 2510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert35
timestamp 0
transform -1 0 2250 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert36
timestamp 0
transform 1 0 1410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert37
timestamp 0
transform -1 0 1170 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert38
timestamp 0
transform -1 0 210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert39
timestamp 0
transform -1 0 970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert40
timestamp 0
transform -1 0 930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert41
timestamp 0
transform 1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert8
timestamp 0
transform -1 0 3630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert9
timestamp 0
transform 1 0 4490 0 1 4950
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert10
timestamp 0
transform 1 0 4770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert11
timestamp 0
transform -1 0 3210 0 1 5470
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert12
timestamp 0
transform -1 0 3370 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__889_
timestamp 0
transform -1 0 3990 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__890_
timestamp 0
transform 1 0 3550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__891_
timestamp 0
transform -1 0 4690 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__892_
timestamp 0
transform 1 0 4950 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__893_
timestamp 0
transform -1 0 3690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__894_
timestamp 0
transform -1 0 4790 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__895_
timestamp 0
transform -1 0 3870 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__896_
timestamp 0
transform 1 0 3710 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__897_
timestamp 0
transform 1 0 5570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__898_
timestamp 0
transform -1 0 4110 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__899_
timestamp 0
transform 1 0 5070 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__900_
timestamp 0
transform -1 0 6110 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__901_
timestamp 0
transform 1 0 5950 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__902_
timestamp 0
transform -1 0 5570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__903_
timestamp 0
transform 1 0 4670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__904_
timestamp 0
transform -1 0 4070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__905_
timestamp 0
transform -1 0 5290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__906_
timestamp 0
transform 1 0 4890 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__907_
timestamp 0
transform -1 0 3110 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__908_
timestamp 0
transform -1 0 6250 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__909_
timestamp 0
transform 1 0 5830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__910_
timestamp 0
transform -1 0 4990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__911_
timestamp 0
transform 1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__912_
timestamp 0
transform 1 0 4670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__913_
timestamp 0
transform 1 0 5670 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__914_
timestamp 0
transform -1 0 5430 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__915_
timestamp 0
transform 1 0 4270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__916_
timestamp 0
transform 1 0 5830 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__917_
timestamp 0
transform 1 0 6030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__918_
timestamp 0
transform -1 0 5410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__919_
timestamp 0
transform -1 0 5290 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__920_
timestamp 0
transform -1 0 6010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__921_
timestamp 0
transform -1 0 5870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform 1 0 5130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform -1 0 5710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform -1 0 5710 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform -1 0 2850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform 1 0 1990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform -1 0 2410 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform -1 0 2730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform 1 0 1190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform -1 0 2150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform -1 0 2270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform 1 0 3890 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform 1 0 4290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform 1 0 3990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform 1 0 1050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform 1 0 1990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__938_
timestamp 0
transform -1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__939_
timestamp 0
transform 1 0 3270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__940_
timestamp 0
transform -1 0 3430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__941_
timestamp 0
transform 1 0 1870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__942_
timestamp 0
transform -1 0 2130 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__943_
timestamp 0
transform -1 0 2270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__944_
timestamp 0
transform -1 0 2890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__945_
timestamp 0
transform -1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__946_
timestamp 0
transform -1 0 2810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__947_
timestamp 0
transform 1 0 3870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__948_
timestamp 0
transform 1 0 4230 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__949_
timestamp 0
transform 1 0 4350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__950_
timestamp 0
transform -1 0 3950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__951_
timestamp 0
transform 1 0 930 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__952_
timestamp 0
transform -1 0 2530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__953_
timestamp 0
transform 1 0 1590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__954_
timestamp 0
transform -1 0 1870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__955_
timestamp 0
transform -1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__956_
timestamp 0
transform -1 0 670 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform 1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform -1 0 530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform 1 0 50 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform 1 0 210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform -1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform -1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform 1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform 1 0 990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform -1 0 550 0 1 790
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform -1 0 830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform -1 0 2750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform 1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform 1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform 1 0 630 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform -1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform -1 0 350 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform 1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform 1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform -1 0 1130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform -1 0 1710 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform -1 0 1870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform 1 0 1250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform -1 0 990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform 1 0 210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform 1 0 670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform 1 0 170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform -1 0 1650 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform 1 0 1550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform -1 0 1470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform -1 0 1570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform 1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform 1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform -1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform 1 0 1310 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform -1 0 1430 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform -1 0 690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform 1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform 1 0 190 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform -1 0 1250 0 1 270
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform -1 0 1410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform -1 0 950 0 1 270
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform 1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform 1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform 1 0 2650 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform 1 0 1790 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform 1 0 3630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform -1 0 1430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform 1 0 1650 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform -1 0 1410 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform 1 0 3370 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform -1 0 1930 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform 1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform -1 0 970 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform -1 0 370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform -1 0 1090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform -1 0 1110 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform 1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform 1 0 1090 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform 1 0 1250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform 1 0 2310 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform 1 0 510 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform 1 0 1550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform -1 0 3010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform 1 0 2750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform -1 0 3190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 3250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform -1 0 2910 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform -1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 2810 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform 1 0 2870 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform 1 0 3150 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform 1 0 3010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform -1 0 3290 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform 1 0 3430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform -1 0 3650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform 1 0 1070 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform -1 0 3010 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform -1 0 2750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform -1 0 1950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform -1 0 2710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform 1 0 2590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform 1 0 2070 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform -1 0 2590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform 1 0 2230 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 1330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform 1 0 1990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform -1 0 2130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform 1 0 2270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform 1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform -1 0 2510 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform 1 0 2430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform 1 0 2590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform -1 0 1790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform 1 0 2090 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform 1 0 2450 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform -1 0 2250 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform 1 0 1210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform -1 0 350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform 1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform -1 0 2730 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform -1 0 2430 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform -1 0 2690 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform -1 0 2170 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform -1 0 1730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform 1 0 1830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform -1 0 1690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform 1 0 1810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform -1 0 2570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform 1 0 1370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform 1 0 2110 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform 1 0 2730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform -1 0 2050 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform -1 0 3670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform 1 0 2270 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform 1 0 3030 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform 1 0 3590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform -1 0 3450 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform 1 0 3570 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform -1 0 3770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform 1 0 3310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform 1 0 3870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform 1 0 4030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 3750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform 1 0 3830 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform 1 0 4170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform 1 0 4250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform 1 0 3890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform 1 0 3730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform 1 0 3750 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform -1 0 3350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform 1 0 3450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform -1 0 2870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform 1 0 2950 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform -1 0 3110 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform 1 0 3150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 3570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform 1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform -1 0 3250 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform 1 0 3010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform -1 0 3190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform 1 0 3950 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 4370 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform 1 0 3290 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform 1 0 3930 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform 1 0 4090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform 1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform -1 0 4530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 4250 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform 1 0 2370 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform -1 0 3950 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform -1 0 4230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform 1 0 3310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform -1 0 3710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform -1 0 4990 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform -1 0 2850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform 1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform 1 0 4710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform -1 0 4630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform -1 0 5010 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform -1 0 4830 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform -1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 4590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform -1 0 4510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform 1 0 4370 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform -1 0 3490 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform -1 0 3170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform -1 0 4110 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform -1 0 4670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform -1 0 4850 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform -1 0 4430 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform -1 0 3950 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform 1 0 3010 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform 1 0 1510 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform -1 0 3790 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform -1 0 2550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform 1 0 3350 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform 1 0 2690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform -1 0 2870 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform -1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform -1 0 3050 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 2490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform -1 0 2230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform 1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform -1 0 70 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform -1 0 670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform -1 0 70 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform -1 0 390 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform 1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform -1 0 1250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform 1 0 210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform -1 0 690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform 1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform 1 0 470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform 1 0 950 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform 1 0 1870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform -1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform 1 0 1650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform -1 0 2050 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform -1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform 1 0 3190 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform -1 0 3210 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform 1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform 1 0 350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform -1 0 1990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform 1 0 50 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform 1 0 210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform -1 0 790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform -1 0 230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform 1 0 190 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform 1 0 350 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform 1 0 490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform -1 0 1210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform 1 0 810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform -1 0 1150 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform -1 0 790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform 1 0 1530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform 1 0 1690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform -1 0 2590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform 1 0 1790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform 1 0 1030 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform -1 0 1170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform 1 0 370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform 1 0 350 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform 1 0 510 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 1850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform 1 0 1290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform -1 0 630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform -1 0 730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform -1 0 670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform 1 0 810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform 1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform 1 0 1050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform 1 0 1010 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform 1 0 830 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform 1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform 1 0 1710 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform 1 0 1370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform 1 0 1570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform 1 0 1790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 2090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform -1 0 2030 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform -1 0 2870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform 1 0 3490 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform -1 0 5090 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform -1 0 4110 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform -1 0 3450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform -1 0 5130 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform 1 0 4310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform 1 0 3470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform -1 0 4910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform -1 0 4470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform -1 0 4990 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform 1 0 5010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform -1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform 1 0 5170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform 1 0 5410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform 1 0 4410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform 1 0 3690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform -1 0 2350 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform -1 0 3430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform 1 0 2490 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform 1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform 1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform 1 0 3930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform -1 0 3310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform -1 0 3110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 3710 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform 1 0 4050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform -1 0 4650 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform 1 0 3990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform -1 0 3910 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform 1 0 4130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform -1 0 4430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform 1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 4350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform 1 0 4690 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform -1 0 4790 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform 1 0 4590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform -1 0 4170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 4850 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform 1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 4670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform 1 0 4870 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 4530 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform 1 0 5250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform -1 0 5210 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform 1 0 5710 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform 1 0 5370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform 1 0 5830 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform -1 0 5810 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform 1 0 4990 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform 1 0 4250 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform 1 0 5550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 5330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform -1 0 4550 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform -1 0 5970 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform -1 0 5610 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform -1 0 4850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform 1 0 4690 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform 1 0 5270 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform -1 0 5510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform 1 0 3770 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform 1 0 5430 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform -1 0 6110 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform -1 0 5650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform 1 0 5730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 5130 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform -1 0 2610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform -1 0 2570 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform -1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform 1 0 2510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform 1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 2550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform -1 0 3750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform -1 0 3790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform 1 0 2210 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform 1 0 3990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform 1 0 5150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform -1 0 5670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform -1 0 2910 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform 1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform -1 0 2470 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform -1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform -1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform -1 0 2150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform 1 0 2170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform 1 0 2330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform -1 0 5630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform 1 0 5630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform -1 0 6210 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform 1 0 6030 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform 1 0 5310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform -1 0 6270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform 1 0 5510 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform 1 0 5670 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform 1 0 4210 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform 1 0 4490 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform 1 0 3410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform -1 0 3290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform 1 0 3530 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform 1 0 5070 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform 1 0 5390 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform -1 0 4310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform 1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform 1 0 3190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform -1 0 2650 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform 1 0 2630 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform -1 0 3050 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform 1 0 2650 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform -1 0 2810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform 1 0 2750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 2910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform -1 0 2770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 4030 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform -1 0 3630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform -1 0 2950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform -1 0 3350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform -1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 3470 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform 1 0 2910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform 1 0 3410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 3550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform -1 0 5170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform -1 0 5470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 4710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform 1 0 5170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform 1 0 5450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform -1 0 5610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform 1 0 5030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform -1 0 5490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform 1 0 5730 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform 1 0 5930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 6010 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform 1 0 5870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform 1 0 5570 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform 1 0 5290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 5610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform -1 0 5770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform 1 0 6170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform 1 0 5870 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform 1 0 6050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform -1 0 6210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform 1 0 6170 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform 1 0 5130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform 1 0 5710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform -1 0 6050 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform -1 0 6110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform -1 0 5930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform 1 0 6070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform 1 0 5450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 5330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform 1 0 5490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform 1 0 1930 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform 1 0 1990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform 1 0 2090 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform -1 0 1990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform 1 0 2730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform 1 0 2650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform -1 0 3430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform -1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform 1 0 5990 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform -1 0 5970 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform 1 0 6030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform -1 0 6250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform -1 0 4950 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform -1 0 5270 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform -1 0 5670 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform -1 0 5630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform 1 0 3830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform 1 0 4550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform 1 0 3810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform -1 0 3090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform -1 0 3970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform 1 0 4090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform 1 0 4670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 3850 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform -1 0 4010 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform 1 0 4110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform 1 0 4830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform 1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 3690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform 1 0 3950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform -1 0 3390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform -1 0 3790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform 1 0 4410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform 1 0 4250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform -1 0 4250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform 1 0 4710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform 1 0 4550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform 1 0 4870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform 1 0 5130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform 1 0 4710 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform -1 0 4450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform -1 0 4210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 4330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform 1 0 5050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform 1 0 5590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform -1 0 5330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform 1 0 4870 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform 1 0 4410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 4270 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform 1 0 4550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform 1 0 5370 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform 1 0 5930 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform 1 0 5510 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform 1 0 5770 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform -1 0 6230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform 1 0 6190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform 1 0 5770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform -1 0 6090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform -1 0 6110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform -1 0 6210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform -1 0 6110 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 5890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform 1 0 5950 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform -1 0 6250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform -1 0 5970 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform -1 0 5830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform -1 0 2250 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform 1 0 2530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform 1 0 710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform 1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform 1 0 2430 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform 1 0 2650 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform 1 0 2790 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform 1 0 3150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform -1 0 6150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform 1 0 4450 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform 1 0 5450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform -1 0 6090 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform 1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform 1 0 5330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform 1 0 5210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform 1 0 3770 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform 1 0 4650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform 1 0 4510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform 1 0 4070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform 1 0 4750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform 1 0 4630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 5050 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform 1 0 4890 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform -1 0 5050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform -1 0 4890 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1452_
timestamp 0
transform -1 0 3670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1453_
timestamp 0
transform 1 0 3890 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1454_
timestamp 0
transform 1 0 3770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1455_
timestamp 0
transform 1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1456_
timestamp 0
transform 1 0 4290 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1457_
timestamp 0
transform 1 0 4370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1458_
timestamp 0
transform -1 0 4790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1459_
timestamp 0
transform 1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1460_
timestamp 0
transform 1 0 4930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1461_
timestamp 0
transform 1 0 5330 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1462_
timestamp 0
transform 1 0 4970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1463_
timestamp 0
transform 1 0 5070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1464_
timestamp 0
transform 1 0 5170 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1465_
timestamp 0
transform 1 0 5490 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1466_
timestamp 0
transform 1 0 5070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1467_
timestamp 0
transform 1 0 5170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1468_
timestamp 0
transform 1 0 5230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1469_
timestamp 0
transform -1 0 5390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1470_
timestamp 0
transform 1 0 5790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1471_
timestamp 0
transform 1 0 5290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1472_
timestamp 0
transform 1 0 5450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1473_
timestamp 0
transform 1 0 5510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1474_
timestamp 0
transform -1 0 6090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1475_
timestamp 0
transform -1 0 5990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1476_
timestamp 0
transform -1 0 6110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1477_
timestamp 0
transform -1 0 5730 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1478_
timestamp 0
transform 1 0 5830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1479_
timestamp 0
transform -1 0 5790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1480_
timestamp 0
transform 1 0 870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1481_
timestamp 0
transform 1 0 910 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1482_
timestamp 0
transform -1 0 1050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1483_
timestamp 0
transform 1 0 2130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1484_
timestamp 0
transform -1 0 2290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1485_
timestamp 0
transform 1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1486_
timestamp 0
transform -1 0 5830 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1487_
timestamp 0
transform -1 0 2550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1488_
timestamp 0
transform 1 0 4710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1489_
timestamp 0
transform 1 0 4890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1490_
timestamp 0
transform 1 0 3890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1491_
timestamp 0
transform -1 0 3530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1492_
timestamp 0
transform 1 0 3930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1493_
timestamp 0
transform -1 0 4090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1494_
timestamp 0
transform 1 0 4230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1495_
timestamp 0
transform -1 0 4170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1496_
timestamp 0
transform 1 0 4130 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1497_
timestamp 0
transform 1 0 4530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1498_
timestamp 0
transform 1 0 4370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1499_
timestamp 0
transform 1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1500_
timestamp 0
transform 1 0 4550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1501_
timestamp 0
transform 1 0 4830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1502_
timestamp 0
transform -1 0 5130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1503_
timestamp 0
transform -1 0 4990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1504_
timestamp 0
transform 1 0 4990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1505_
timestamp 0
transform -1 0 5130 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1506_
timestamp 0
transform 1 0 5230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1507_
timestamp 0
transform 1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1508_
timestamp 0
transform -1 0 5430 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1509_
timestamp 0
transform 1 0 5650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1510_
timestamp 0
transform -1 0 5550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1511_
timestamp 0
transform 1 0 5550 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1512_
timestamp 0
transform -1 0 5950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1513_
timestamp 0
transform 1 0 5650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1514_
timestamp 0
transform 1 0 5930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1515_
timestamp 0
transform 1 0 5610 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1516_
timestamp 0
transform -1 0 6230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1517_
timestamp 0
transform 1 0 5750 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1518_
timestamp 0
transform 1 0 5790 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1519_
timestamp 0
transform 1 0 6190 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1520_
timestamp 0
transform 1 0 5870 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1521_
timestamp 0
transform 1 0 5770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1522_
timestamp 0
transform -1 0 5930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1523_
timestamp 0
transform 1 0 6070 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1524_
timestamp 0
transform -1 0 5990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1525_
timestamp 0
transform 1 0 1930 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1526_
timestamp 0
transform 1 0 2210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1527_
timestamp 0
transform 1 0 1670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1528_
timestamp 0
transform 1 0 1170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1529_
timestamp 0
transform 1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 2090 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1531_
timestamp 0
transform -1 0 2310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1532_
timestamp 0
transform 1 0 2370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1533_
timestamp 0
transform -1 0 2370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1534_
timestamp 0
transform 1 0 5030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1535_
timestamp 0
transform 1 0 5330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1536_
timestamp 0
transform -1 0 6250 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1537_
timestamp 0
transform 1 0 6050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1538_
timestamp 0
transform 1 0 5250 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1539_
timestamp 0
transform 1 0 4510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1540_
timestamp 0
transform 1 0 4050 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1541_
timestamp 0
transform 1 0 4430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1542_
timestamp 0
transform -1 0 4210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1543_
timestamp 0
transform 1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1544_
timestamp 0
transform -1 0 4670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1545_
timestamp 0
transform 1 0 5050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1546_
timestamp 0
transform 1 0 5510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1547_
timestamp 0
transform -1 0 6090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1548_
timestamp 0
transform -1 0 6210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1549_
timestamp 0
transform 1 0 5930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1550_
timestamp 0
transform 1 0 5610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1551_
timestamp 0
transform 1 0 1950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1552_
timestamp 0
transform 1 0 2350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1553_
timestamp 0
transform 1 0 3470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1554_
timestamp 0
transform -1 0 4130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1555_
timestamp 0
transform 1 0 4090 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1556_
timestamp 0
transform 1 0 5310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1557_
timestamp 0
transform -1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1558_
timestamp 0
transform 1 0 5870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1559_
timestamp 0
transform 1 0 6030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1560_
timestamp 0
transform -1 0 6170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1561_
timestamp 0
transform -1 0 5670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1562_
timestamp 0
transform 1 0 5490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1563_
timestamp 0
transform -1 0 5410 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1564_
timestamp 0
transform 1 0 4770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1565_
timestamp 0
transform 1 0 4650 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1566_
timestamp 0
transform 1 0 4490 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1567_
timestamp 0
transform 1 0 3890 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1568_
timestamp 0
transform 1 0 4870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1569_
timestamp 0
transform -1 0 5250 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1570_
timestamp 0
transform -1 0 5730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1571_
timestamp 0
transform 1 0 5250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1572_
timestamp 0
transform -1 0 5370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1573_
timestamp 0
transform -1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1574_
timestamp 0
transform 1 0 2110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1575_
timestamp 0
transform 1 0 2050 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1576_
timestamp 0
transform -1 0 2210 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1577_
timestamp 0
transform 1 0 2190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1578_
timestamp 0
transform -1 0 1970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1579_
timestamp 0
transform 1 0 2070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1580_
timestamp 0
transform 1 0 2430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1581_
timestamp 0
transform -1 0 4430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1582_
timestamp 0
transform 1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1583_
timestamp 0
transform -1 0 5090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1584_
timestamp 0
transform 1 0 4590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1585_
timestamp 0
transform -1 0 4750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1586_
timestamp 0
transform 1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1587_
timestamp 0
transform 1 0 2610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1588_
timestamp 0
transform 1 0 2650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1589_
timestamp 0
transform -1 0 2970 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1590_
timestamp 0
transform -1 0 3030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1591_
timestamp 0
transform 1 0 3430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1592_
timestamp 0
transform -1 0 4790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1593_
timestamp 0
transform -1 0 2730 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1594_
timestamp 0
transform 1 0 2870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1595_
timestamp 0
transform 1 0 2570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1596_
timestamp 0
transform 1 0 2410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1597_
timestamp 0
transform -1 0 4190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1598_
timestamp 0
transform 1 0 4010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1599_
timestamp 0
transform -1 0 2810 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1600_
timestamp 0
transform 1 0 2630 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1601_
timestamp 0
transform 1 0 3750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1602_
timestamp 0
transform 1 0 3610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1603_
timestamp 0
transform 1 0 2870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1604_
timestamp 0
transform 1 0 2810 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1605_
timestamp 0
transform 1 0 3610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1606_
timestamp 0
transform 1 0 3450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1607_
timestamp 0
transform -1 0 3330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1608_
timestamp 0
transform -1 0 3610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1636_
timestamp 0
transform -1 0 230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1637_
timestamp 0
transform 1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1638_
timestamp 0
transform -1 0 70 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1639_
timestamp 0
transform -1 0 70 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1640_
timestamp 0
transform 1 0 750 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1641_
timestamp 0
transform 1 0 1070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1642_
timestamp 0
transform 1 0 470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1643_
timestamp 0
transform -1 0 970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1644_
timestamp 0
transform 1 0 930 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1645_
timestamp 0
transform -1 0 610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1646_
timestamp 0
transform 1 0 750 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1647_
timestamp 0
transform 1 0 170 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1648_
timestamp 0
transform -1 0 250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1649_
timestamp 0
transform -1 0 510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1650_
timestamp 0
transform 1 0 50 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1651_
timestamp 0
transform -1 0 210 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1652_
timestamp 0
transform -1 0 350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1653_
timestamp 0
transform -1 0 630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1654_
timestamp 0
transform -1 0 470 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1655_
timestamp 0
transform 1 0 610 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1656_
timestamp 0
transform 1 0 350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1657_
timestamp 0
transform 1 0 850 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1658_
timestamp 0
transform 1 0 1150 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1659_
timestamp 0
transform 1 0 1490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1660_
timestamp 0
transform -1 0 1030 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1661_
timestamp 0
transform -1 0 1310 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1662_
timestamp 0
transform 1 0 1790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1663_
timestamp 0
transform -1 0 1510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1664_
timestamp 0
transform 1 0 1310 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1665_
timestamp 0
transform -1 0 1730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1666_
timestamp 0
transform 1 0 1590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1667_
timestamp 0
transform 1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1668_
timestamp 0
transform 1 0 1630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1669_
timestamp 0
transform 1 0 1070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1670_
timestamp 0
transform 1 0 1210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1671_
timestamp 0
transform -1 0 1730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1672_
timestamp 0
transform 1 0 1370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1673_
timestamp 0
transform -1 0 1550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1674_
timestamp 0
transform -1 0 1450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1675_
timestamp 0
transform -1 0 350 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1676_
timestamp 0
transform 1 0 190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1677_
timestamp 0
transform -1 0 810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1678_
timestamp 0
transform 1 0 50 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1679_
timestamp 0
transform 1 0 470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1680_
timestamp 0
transform -1 0 350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1681_
timestamp 0
transform -1 0 470 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1682_
timestamp 0
transform -1 0 350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1683_
timestamp 0
transform 1 0 470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1684_
timestamp 0
transform -1 0 650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1685_
timestamp 0
transform 1 0 1550 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1686_
timestamp 0
transform 1 0 1810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1687_
timestamp 0
transform 1 0 1990 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1688_
timestamp 0
transform 1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1689_
timestamp 0
transform 1 0 1990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1690_
timestamp 0
transform -1 0 1730 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1691_
timestamp 0
transform 1 0 1830 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1692_
timestamp 0
transform 1 0 1010 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1693_
timestamp 0
transform -1 0 1350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1694_
timestamp 0
transform 1 0 1150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1695_
timestamp 0
transform 1 0 750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1696_
timestamp 0
transform -1 0 870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1697_
timestamp 0
transform -1 0 1010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1698_
timestamp 0
transform -1 0 1150 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1699_
timestamp 0
transform 1 0 590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1700_
timestamp 0
transform 1 0 610 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1701_
timestamp 0
transform 1 0 1270 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1702_
timestamp 0
transform -1 0 1450 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1703_
timestamp 0
transform -1 0 2250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1704_
timestamp 0
transform 1 0 2190 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1705_
timestamp 0
transform 1 0 750 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1706_
timestamp 0
transform -1 0 870 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1707_
timestamp 0
transform -1 0 1770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1708_
timestamp 0
transform 1 0 1590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1709_
timestamp 0
transform -1 0 1490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1710_
timestamp 0
transform -1 0 1750 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1711_
timestamp 0
transform -1 0 1630 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1712_
timestamp 0
transform 1 0 1290 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1713_
timestamp 0
transform -1 0 1570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1714_
timestamp 0
transform 1 0 1390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1715_
timestamp 0
transform -1 0 1110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1716_
timestamp 0
transform -1 0 1270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1717_
timestamp 0
transform 1 0 1210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1718_
timestamp 0
transform 1 0 1370 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1719_
timestamp 0
transform 1 0 1690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1720_
timestamp 0
transform 1 0 1690 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1721_
timestamp 0
transform 1 0 2110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1722_
timestamp 0
transform -1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1723_
timestamp 0
transform -1 0 1850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1724_
timestamp 0
transform -1 0 2070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1725_
timestamp 0
transform -1 0 1550 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1726_
timestamp 0
transform 1 0 1650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1727_
timestamp 0
transform -1 0 1770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1728_
timestamp 0
transform -1 0 1170 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1729_
timestamp 0
transform -1 0 1710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1730_
timestamp 0
transform 1 0 1410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1731_
timestamp 0
transform 1 0 1070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1732_
timestamp 0
transform -1 0 1570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1733_
timestamp 0
transform -1 0 1270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1734_
timestamp 0
transform 1 0 910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1735_
timestamp 0
transform -1 0 1070 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1736_
timestamp 0
transform 1 0 1190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1737_
timestamp 0
transform 1 0 1350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1738_
timestamp 0
transform 1 0 1490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1739_
timestamp 0
transform -1 0 1630 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1740_
timestamp 0
transform 1 0 1230 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1741_
timestamp 0
transform -1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1742_
timestamp 0
transform 1 0 350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1743_
timestamp 0
transform -1 0 910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1744_
timestamp 0
transform 1 0 790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1745_
timestamp 0
transform -1 0 490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1746_
timestamp 0
transform -1 0 750 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1747_
timestamp 0
transform -1 0 650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1748_
timestamp 0
transform -1 0 790 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1749_
timestamp 0
transform 1 0 610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1750_
timestamp 0
transform 1 0 570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1751_
timestamp 0
transform 1 0 710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1752_
timestamp 0
transform 1 0 930 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1753_
timestamp 0
transform -1 0 1070 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1754_
timestamp 0
transform 1 0 2970 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1755_
timestamp 0
transform -1 0 810 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1756_
timestamp 0
transform -1 0 210 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1757_
timestamp 0
transform -1 0 830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1758_
timestamp 0
transform 1 0 610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1759_
timestamp 0
transform -1 0 450 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1760_
timestamp 0
transform -1 0 670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1761_
timestamp 0
transform 1 0 490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1762_
timestamp 0
transform 1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1763_
timestamp 0
transform -1 0 490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1764_
timestamp 0
transform -1 0 530 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1765_
timestamp 0
transform -1 0 370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1766_
timestamp 0
transform 1 0 670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1767_
timestamp 0
transform 1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1768_
timestamp 0
transform -1 0 2050 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1769_
timestamp 0
transform -1 0 1910 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1770_
timestamp 0
transform 1 0 1490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1771_
timestamp 0
transform 1 0 870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1772_
timestamp 0
transform 1 0 1010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1773_
timestamp 0
transform 1 0 330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1774_
timestamp 0
transform -1 0 1150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1775_
timestamp 0
transform -1 0 1270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1776_
timestamp 0
transform -1 0 610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1777_
timestamp 0
transform -1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1778_
timestamp 0
transform -1 0 210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1779_
timestamp 0
transform 1 0 170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1780_
timestamp 0
transform -1 0 310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1781_
timestamp 0
transform 1 0 330 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1782_
timestamp 0
transform -1 0 210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1783_
timestamp 0
transform -1 0 70 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1784_
timestamp 0
transform -1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1785_
timestamp 0
transform -1 0 70 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1786_
timestamp 0
transform 1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1787_
timestamp 0
transform -1 0 750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1788_
timestamp 0
transform -1 0 470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1789_
timestamp 0
transform 1 0 50 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1790_
timestamp 0
transform 1 0 530 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1791_
timestamp 0
transform 1 0 990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1792_
timestamp 0
transform 1 0 1870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1793_
timestamp 0
transform 1 0 1910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1794_
timestamp 0
transform -1 0 1830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1795_
timestamp 0
transform 1 0 1390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1796_
timestamp 0
transform 1 0 1810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1797_
timestamp 0
transform 1 0 1950 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1798_
timestamp 0
transform 1 0 370 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1799_
timestamp 0
transform 1 0 670 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1800_
timestamp 0
transform -1 0 1090 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1801_
timestamp 0
transform -1 0 1550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1802_
timestamp 0
transform -1 0 310 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1803_
timestamp 0
transform -1 0 230 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1804_
timestamp 0
transform 1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1805_
timestamp 0
transform -1 0 210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1806_
timestamp 0
transform 1 0 170 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1807_
timestamp 0
transform -1 0 1210 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1808_
timestamp 0
transform -1 0 1690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1809_
timestamp 0
transform 1 0 210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1810_
timestamp 0
transform 1 0 370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1811_
timestamp 0
transform 1 0 850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1812_
timestamp 0
transform 1 0 810 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1813_
timestamp 0
transform 1 0 930 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1814_
timestamp 0
transform 1 0 1350 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1815_
timestamp 0
transform 1 0 1630 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1816_
timestamp 0
transform 1 0 1490 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1817_
timestamp 0
transform -1 0 1810 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1818_
timestamp 0
transform 1 0 4670 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1819_
timestamp 0
transform -1 0 2110 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1820_
timestamp 0
transform 1 0 3850 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1821_
timestamp 0
transform 1 0 6170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1822_
timestamp 0
transform 1 0 2790 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1823_
timestamp 0
transform -1 0 4830 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1824_
timestamp 0
transform -1 0 4570 0 1 5990
box -6 -8 26 268
use FILL  FILL_2__1825_
timestamp 0
transform -1 0 5030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1826_
timestamp 0
transform 1 0 6170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1827_
timestamp 0
transform 1 0 6110 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform 1 0 2430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform -1 0 1910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform 1 0 2390 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform 1 0 2490 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform -1 0 890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform 1 0 1010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform -1 0 2130 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform 1 0 2410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 3750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 3590 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform 1 0 4010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform -1 0 3030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform -1 0 3030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 3290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform 1 0 3850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 2870 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform 1 0 3130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform 1 0 2990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform -1 0 3030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert26
timestamp 0
transform -1 0 4010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert27
timestamp 0
transform -1 0 2130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert28
timestamp 0
transform 1 0 2310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert29
timestamp 0
transform 1 0 4010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert30
timestamp 0
transform 1 0 2710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert31
timestamp 0
transform -1 0 1810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert32
timestamp 0
transform 1 0 1910 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert33
timestamp 0
transform -1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert34
timestamp 0
transform 1 0 2530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert35
timestamp 0
transform -1 0 2270 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert36
timestamp 0
transform 1 0 1430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert37
timestamp 0
transform -1 0 1190 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert38
timestamp 0
transform -1 0 230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert39
timestamp 0
transform -1 0 990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert40
timestamp 0
transform -1 0 950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert41
timestamp 0
transform 1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert8
timestamp 0
transform -1 0 3650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert9
timestamp 0
transform 1 0 4510 0 1 4950
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert10
timestamp 0
transform 1 0 4790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert11
timestamp 0
transform -1 0 3230 0 1 5470
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert12
timestamp 0
transform -1 0 3390 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__889_
timestamp 0
transform -1 0 4010 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__891_
timestamp 0
transform -1 0 4710 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__892_
timestamp 0
transform 1 0 4970 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__894_
timestamp 0
transform -1 0 4810 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__896_
timestamp 0
transform 1 0 3730 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__897_
timestamp 0
transform 1 0 5590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__899_
timestamp 0
transform 1 0 5090 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__900_
timestamp 0
transform -1 0 6130 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__902_
timestamp 0
transform -1 0 5590 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__904_
timestamp 0
transform -1 0 4090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__905_
timestamp 0
transform -1 0 5310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__907_
timestamp 0
transform -1 0 3130 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__909_
timestamp 0
transform 1 0 5850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__910_
timestamp 0
transform -1 0 5010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__912_
timestamp 0
transform 1 0 4690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__913_
timestamp 0
transform 1 0 5690 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__915_
timestamp 0
transform 1 0 4290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__917_
timestamp 0
transform 1 0 6050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__918_
timestamp 0
transform -1 0 5430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__920_
timestamp 0
transform -1 0 6030 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__921_
timestamp 0
transform -1 0 5890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__923_
timestamp 0
transform -1 0 5730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__925_
timestamp 0
transform -1 0 2870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__926_
timestamp 0
transform 1 0 2010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__928_
timestamp 0
transform -1 0 2750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__929_
timestamp 0
transform 1 0 1210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform -1 0 2290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__933_
timestamp 0
transform 1 0 4310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__934_
timestamp 0
transform 1 0 4010 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__936_
timestamp 0
transform 1 0 2010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__938_
timestamp 0
transform -1 0 90 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__939_
timestamp 0
transform 1 0 3290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__941_
timestamp 0
transform 1 0 1890 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__942_
timestamp 0
transform -1 0 2150 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__944_
timestamp 0
transform -1 0 2910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__946_
timestamp 0
transform -1 0 2830 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__947_
timestamp 0
transform 1 0 3890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__949_
timestamp 0
transform 1 0 4370 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__950_
timestamp 0
transform -1 0 3970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__952_
timestamp 0
transform -1 0 2550 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__954_
timestamp 0
transform -1 0 1890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__955_
timestamp 0
transform -1 0 1750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__957_
timestamp 0
transform 1 0 490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__959_
timestamp 0
transform -1 0 190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__960_
timestamp 0
transform 1 0 70 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__962_
timestamp 0
transform -1 0 330 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__963_
timestamp 0
transform -1 0 90 0 1 270
box -6 -8 26 268
use FILL  FILL_3__965_
timestamp 0
transform 1 0 1010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__967_
timestamp 0
transform -1 0 850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__968_
timestamp 0
transform -1 0 2770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__970_
timestamp 0
transform 1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__971_
timestamp 0
transform 1 0 650 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__973_
timestamp 0
transform -1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__975_
timestamp 0
transform 1 0 1350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__976_
timestamp 0
transform -1 0 1150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__978_
timestamp 0
transform -1 0 1890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__979_
timestamp 0
transform 1 0 1270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__981_
timestamp 0
transform 1 0 230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__983_
timestamp 0
transform 1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_3__984_
timestamp 0
transform -1 0 1670 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__986_
timestamp 0
transform -1 0 1490 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__988_
timestamp 0
transform 1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__989_
timestamp 0
transform 1 0 830 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__991_
timestamp 0
transform 1 0 1330 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__992_
timestamp 0
transform -1 0 1450 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__994_
timestamp 0
transform 1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__996_
timestamp 0
transform -1 0 1270 0 1 270
box -6 -8 26 268
use FILL  FILL_3__997_
timestamp 0
transform -1 0 1430 0 1 270
box -6 -8 26 268
use FILL  FILL_3__999_
timestamp 0
transform 1 0 1470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1001_
timestamp 0
transform 1 0 2670 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1003_
timestamp 0
transform 1 0 3650 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1004_
timestamp 0
transform -1 0 1450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1006_
timestamp 0
transform -1 0 1430 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1008_
timestamp 0
transform -1 0 1950 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1009_
timestamp 0
transform 1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1011_
timestamp 0
transform -1 0 390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1012_
timestamp 0
transform -1 0 1110 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1014_
timestamp 0
transform -1 0 1130 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1016_
timestamp 0
transform 1 0 1110 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1017_
timestamp 0
transform 1 0 1270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1019_
timestamp 0
transform 1 0 530 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1020_
timestamp 0
transform 1 0 1570 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1022_
timestamp 0
transform 1 0 2770 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1024_
timestamp 0
transform 1 0 3270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1025_
timestamp 0
transform -1 0 2930 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1027_
timestamp 0
transform 1 0 2830 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1028_
timestamp 0
transform 1 0 2890 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1030_
timestamp 0
transform 1 0 3030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1032_
timestamp 0
transform 1 0 3450 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1033_
timestamp 0
transform -1 0 3670 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1035_
timestamp 0
transform -1 0 3030 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1037_
timestamp 0
transform -1 0 1970 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1038_
timestamp 0
transform -1 0 2730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1040_
timestamp 0
transform 1 0 2090 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1041_
timestamp 0
transform -1 0 2610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1043_
timestamp 0
transform -1 0 1350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1045_
timestamp 0
transform -1 0 2150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1046_
timestamp 0
transform 1 0 2290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1048_
timestamp 0
transform -1 0 2530 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1049_
timestamp 0
transform 1 0 2450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1051_
timestamp 0
transform -1 0 1810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1053_
timestamp 0
transform 1 0 3810 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1054_
timestamp 0
transform 1 0 2470 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1056_
timestamp 0
transform 1 0 1230 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1058_
timestamp 0
transform 1 0 2890 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1059_
timestamp 0
transform -1 0 2750 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1061_
timestamp 0
transform -1 0 2710 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1062_
timestamp 0
transform -1 0 2190 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1064_
timestamp 0
transform 1 0 1850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1066_
timestamp 0
transform 1 0 1830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1067_
timestamp 0
transform -1 0 2590 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1069_
timestamp 0
transform 1 0 2130 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1070_
timestamp 0
transform 1 0 2750 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1072_
timestamp 0
transform -1 0 3690 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1074_
timestamp 0
transform 1 0 3050 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1075_
timestamp 0
transform 1 0 3610 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1077_
timestamp 0
transform 1 0 3590 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1078_
timestamp 0
transform -1 0 3790 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1080_
timestamp 0
transform 1 0 3890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1082_
timestamp 0
transform 1 0 3770 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1083_
timestamp 0
transform 1 0 3850 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1085_
timestamp 0
transform 1 0 4270 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1087_
timestamp 0
transform 1 0 3750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1088_
timestamp 0
transform 1 0 3770 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1090_
timestamp 0
transform 1 0 3470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1091_
timestamp 0
transform -1 0 2890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1093_
timestamp 0
transform -1 0 3130 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1095_
timestamp 0
transform 1 0 3590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1096_
timestamp 0
transform 1 0 3590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1098_
timestamp 0
transform 1 0 3030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1099_
timestamp 0
transform -1 0 3210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1101_
timestamp 0
transform -1 0 4390 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1103_
timestamp 0
transform 1 0 3950 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1104_
timestamp 0
transform 1 0 4110 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1106_
timestamp 0
transform -1 0 4550 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1108_
timestamp 0
transform 1 0 2390 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1109_
timestamp 0
transform -1 0 3970 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1111_
timestamp 0
transform 1 0 3330 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1112_
timestamp 0
transform -1 0 3730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1114_
timestamp 0
transform -1 0 2870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1116_
timestamp 0
transform 1 0 4730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1117_
timestamp 0
transform -1 0 4650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1119_
timestamp 0
transform -1 0 4850 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1120_
timestamp 0
transform -1 0 5150 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1122_
timestamp 0
transform -1 0 4530 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1124_
timestamp 0
transform -1 0 3510 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1125_
timestamp 0
transform -1 0 3190 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1127_
timestamp 0
transform -1 0 4690 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1128_
timestamp 0
transform -1 0 4870 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1130_
timestamp 0
transform -1 0 3970 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1132_
timestamp 0
transform 1 0 1530 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1133_
timestamp 0
transform -1 0 3810 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1135_
timestamp 0
transform -1 0 2570 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1137_
timestamp 0
transform 1 0 2710 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1138_
timestamp 0
transform -1 0 2890 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1140_
timestamp 0
transform -1 0 3070 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1141_
timestamp 0
transform 1 0 2510 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1143_
timestamp 0
transform 1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1145_
timestamp 0
transform -1 0 690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1146_
timestamp 0
transform 1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1148_
timestamp 0
transform -1 0 410 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1149_
timestamp 0
transform 1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1151_
timestamp 0
transform 1 0 230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1153_
timestamp 0
transform 1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1154_
timestamp 0
transform 1 0 490 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1156_
timestamp 0
transform 1 0 1890 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1158_
timestamp 0
transform 1 0 1670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1159_
timestamp 0
transform -1 0 2070 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1161_
timestamp 0
transform 1 0 3210 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1162_
timestamp 0
transform -1 0 3230 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1164_
timestamp 0
transform 1 0 370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1166_
timestamp 0
transform 1 0 70 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1167_
timestamp 0
transform 1 0 230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1169_
timestamp 0
transform -1 0 250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1170_
timestamp 0
transform 1 0 210 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1172_
timestamp 0
transform 1 0 510 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1174_
timestamp 0
transform 1 0 530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1175_
timestamp 0
transform 1 0 830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1177_
timestamp 0
transform -1 0 810 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1178_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1180_
timestamp 0
transform -1 0 2610 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1182_
timestamp 0
transform 1 0 1050 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1183_
timestamp 0
transform -1 0 1190 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform 1 0 370 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1187_
timestamp 0
transform -1 0 1870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1188_
timestamp 0
transform 1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1190_
timestamp 0
transform -1 0 750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1191_
timestamp 0
transform -1 0 690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1193_
timestamp 0
transform 1 0 950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1195_
timestamp 0
transform 1 0 1030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1196_
timestamp 0
transform 1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1198_
timestamp 0
transform 1 0 1730 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1199_
timestamp 0
transform 1 0 1390 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1201_
timestamp 0
transform 1 0 1810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1203_
timestamp 0
transform -1 0 2050 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1204_
timestamp 0
transform 1 0 2270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1206_
timestamp 0
transform 1 0 3510 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1208_
timestamp 0
transform -1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1209_
timestamp 0
transform -1 0 3470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1211_
timestamp 0
transform 1 0 4330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1212_
timestamp 0
transform 1 0 3490 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1214_
timestamp 0
transform -1 0 4490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1216_
timestamp 0
transform 1 0 5030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1217_
timestamp 0
transform -1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1219_
timestamp 0
transform 1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1220_
timestamp 0
transform 1 0 4430 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1222_
timestamp 0
transform -1 0 2370 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1224_
timestamp 0
transform 1 0 2510 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1225_
timestamp 0
transform 1 0 3150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1227_
timestamp 0
transform 1 0 3950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1229_
timestamp 0
transform -1 0 3130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1230_
timestamp 0
transform 1 0 3730 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1232_
timestamp 0
transform -1 0 4670 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1233_
timestamp 0
transform 1 0 4010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1235_
timestamp 0
transform 1 0 4150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1237_
timestamp 0
transform 1 0 3990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1238_
timestamp 0
transform 1 0 4030 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1240_
timestamp 0
transform 1 0 4710 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1241_
timestamp 0
transform -1 0 4810 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1243_
timestamp 0
transform -1 0 4190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1245_
timestamp 0
transform 1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1246_
timestamp 0
transform 1 0 4690 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1248_
timestamp 0
transform 1 0 4550 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1249_
timestamp 0
transform 1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1251_
timestamp 0
transform 1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1253_
timestamp 0
transform 1 0 5850 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1254_
timestamp 0
transform -1 0 5830 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1256_
timestamp 0
transform 1 0 4270 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1258_
timestamp 0
transform 1 0 5350 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1259_
timestamp 0
transform -1 0 4570 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1261_
timestamp 0
transform -1 0 5630 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1262_
timestamp 0
transform -1 0 4870 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1264_
timestamp 0
transform 1 0 5290 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1266_
timestamp 0
transform 1 0 3790 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1267_
timestamp 0
transform 1 0 5450 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1269_
timestamp 0
transform -1 0 5670 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1270_
timestamp 0
transform 1 0 5750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1272_
timestamp 0
transform -1 0 2630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1274_
timestamp 0
transform -1 0 2750 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1275_
timestamp 0
transform 1 0 2530 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1277_
timestamp 0
transform 1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1279_
timestamp 0
transform -1 0 3810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1280_
timestamp 0
transform 1 0 2230 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1282_
timestamp 0
transform 1 0 5170 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1283_
timestamp 0
transform -1 0 5690 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1285_
timestamp 0
transform 1 0 2030 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1287_
timestamp 0
transform -1 0 2330 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1288_
timestamp 0
transform -1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1290_
timestamp 0
transform 1 0 2190 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1291_
timestamp 0
transform 1 0 2350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1293_
timestamp 0
transform 1 0 5650 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1295_
timestamp 0
transform 1 0 6050 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1296_
timestamp 0
transform 1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1298_
timestamp 0
transform 1 0 5530 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1299_
timestamp 0
transform 1 0 5690 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1301_
timestamp 0
transform 1 0 4510 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1303_
timestamp 0
transform -1 0 3310 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1304_
timestamp 0
transform 1 0 3550 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1306_
timestamp 0
transform 1 0 5410 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1308_
timestamp 0
transform 1 0 5010 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1309_
timestamp 0
transform 1 0 3210 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1311_
timestamp 0
transform 1 0 2650 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1312_
timestamp 0
transform -1 0 3070 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1314_
timestamp 0
transform -1 0 2830 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1316_
timestamp 0
transform 1 0 2930 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1317_
timestamp 0
transform -1 0 2790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1319_
timestamp 0
transform -1 0 3650 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1320_
timestamp 0
transform -1 0 2970 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1322_
timestamp 0
transform -1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1324_
timestamp 0
transform 1 0 2930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1325_
timestamp 0
transform 1 0 3430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1327_
timestamp 0
transform -1 0 5190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1329_
timestamp 0
transform -1 0 4490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1330_
timestamp 0
transform 1 0 4730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1332_
timestamp 0
transform 1 0 5470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1333_
timestamp 0
transform -1 0 5630 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1335_
timestamp 0
transform -1 0 5510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1337_
timestamp 0
transform 1 0 5950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1338_
timestamp 0
transform 1 0 6030 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1340_
timestamp 0
transform 1 0 5590 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1341_
timestamp 0
transform 1 0 5310 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1343_
timestamp 0
transform -1 0 5790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1345_
timestamp 0
transform 1 0 6190 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1346_
timestamp 0
transform 1 0 5890 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1348_
timestamp 0
transform -1 0 6230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1349_
timestamp 0
transform 1 0 6190 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1351_
timestamp 0
transform 1 0 5730 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1353_
timestamp 0
transform -1 0 6130 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1354_
timestamp 0
transform -1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1356_
timestamp 0
transform 1 0 5470 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1358_
timestamp 0
transform 1 0 5510 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1359_
timestamp 0
transform 1 0 1950 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1361_
timestamp 0
transform 1 0 2110 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1362_
timestamp 0
transform -1 0 2010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1364_
timestamp 0
transform 1 0 2670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1366_
timestamp 0
transform -1 0 5830 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1367_
timestamp 0
transform 1 0 6010 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1369_
timestamp 0
transform 1 0 6050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1370_
timestamp 0
transform 1 0 5770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1372_
timestamp 0
transform -1 0 4970 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1374_
timestamp 0
transform -1 0 5690 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1375_
timestamp 0
transform -1 0 5650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1377_
timestamp 0
transform 1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1379_
timestamp 0
transform -1 0 3110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1380_
timestamp 0
transform -1 0 3990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1382_
timestamp 0
transform 1 0 4690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1383_
timestamp 0
transform -1 0 3870 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1385_
timestamp 0
transform 1 0 4130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1387_
timestamp 0
transform 1 0 4350 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1388_
timestamp 0
transform 1 0 3710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1390_
timestamp 0
transform -1 0 3410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1391_
timestamp 0
transform -1 0 3810 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1393_
timestamp 0
transform 1 0 4270 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1395_
timestamp 0
transform 1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1396_
timestamp 0
transform 1 0 4570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1398_
timestamp 0
transform 1 0 5150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1399_
timestamp 0
transform 1 0 4730 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1401_
timestamp 0
transform -1 0 4230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1403_
timestamp 0
transform 1 0 5070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1404_
timestamp 0
transform 1 0 5610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1406_
timestamp 0
transform 1 0 4890 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1408_
timestamp 0
transform 1 0 4290 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1409_
timestamp 0
transform 1 0 4570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1411_
timestamp 0
transform 1 0 5950 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1412_
timestamp 0
transform 1 0 5450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1414_
timestamp 0
transform 1 0 5790 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1416_
timestamp 0
transform 1 0 6210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1417_
timestamp 0
transform 1 0 5790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1419_
timestamp 0
transform -1 0 6130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform -1 0 6230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1422_
timestamp 0
transform 1 0 5910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1424_
timestamp 0
transform -1 0 6270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1425_
timestamp 0
transform -1 0 5990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1427_
timestamp 0
transform -1 0 2270 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1429_
timestamp 0
transform 1 0 730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1430_
timestamp 0
transform 1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1432_
timestamp 0
transform 1 0 2670 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1433_
timestamp 0
transform 1 0 2810 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1435_
timestamp 0
transform -1 0 6170 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1437_
timestamp 0
transform 1 0 5470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1438_
timestamp 0
transform -1 0 6110 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1440_
timestamp 0
transform 1 0 5350 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1441_
timestamp 0
transform 1 0 5230 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1443_
timestamp 0
transform 1 0 4670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1445_
timestamp 0
transform 1 0 4090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1446_
timestamp 0
transform 1 0 4770 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1448_
timestamp 0
transform 1 0 5070 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1449_
timestamp 0
transform 1 0 4910 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1451_
timestamp 0
transform -1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1453_
timestamp 0
transform 1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1454_
timestamp 0
transform 1 0 3790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1456_
timestamp 0
transform 1 0 4310 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1458_
timestamp 0
transform -1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1459_
timestamp 0
transform 1 0 4970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1461_
timestamp 0
transform 1 0 5350 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1462_
timestamp 0
transform 1 0 4990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1464_
timestamp 0
transform 1 0 5190 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1466_
timestamp 0
transform 1 0 5090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1467_
timestamp 0
transform 1 0 5190 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1469_
timestamp 0
transform -1 0 5410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1470_
timestamp 0
transform 1 0 5810 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1472_
timestamp 0
transform 1 0 5470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1474_
timestamp 0
transform -1 0 6110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1475_
timestamp 0
transform -1 0 6010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1477_
timestamp 0
transform -1 0 5750 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1479_
timestamp 0
transform -1 0 5810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1480_
timestamp 0
transform 1 0 890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1482_
timestamp 0
transform -1 0 1070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1483_
timestamp 0
transform 1 0 2150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1485_
timestamp 0
transform 1 0 4630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1487_
timestamp 0
transform -1 0 2570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1488_
timestamp 0
transform 1 0 4730 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1490_
timestamp 0
transform 1 0 3910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1491_
timestamp 0
transform -1 0 3550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1493_
timestamp 0
transform -1 0 4110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1495_
timestamp 0
transform -1 0 4190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1496_
timestamp 0
transform 1 0 4150 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1498_
timestamp 0
transform 1 0 4390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1500_
timestamp 0
transform 1 0 4570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1501_
timestamp 0
transform 1 0 4850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1503_
timestamp 0
transform -1 0 5010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1504_
timestamp 0
transform 1 0 5010 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1506_
timestamp 0
transform 1 0 5250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1508_
timestamp 0
transform -1 0 5450 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1509_
timestamp 0
transform 1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1511_
timestamp 0
transform 1 0 5570 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1512_
timestamp 0
transform -1 0 5970 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1514_
timestamp 0
transform 1 0 5950 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1516_
timestamp 0
transform -1 0 6250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1517_
timestamp 0
transform 1 0 5770 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1519_
timestamp 0
transform 1 0 6210 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1520_
timestamp 0
transform 1 0 5890 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__1522_
timestamp 0
transform -1 0 5950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1524_
timestamp 0
transform -1 0 6010 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1525_
timestamp 0
transform 1 0 1950 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1527_
timestamp 0
transform 1 0 1690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1529_
timestamp 0
transform 1 0 1550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1530_
timestamp 0
transform 1 0 2110 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1532_
timestamp 0
transform 1 0 2390 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1533_
timestamp 0
transform -1 0 2390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1535_
timestamp 0
transform 1 0 5350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1537_
timestamp 0
transform 1 0 6070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1538_
timestamp 0
transform 1 0 5270 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1540_
timestamp 0
transform 1 0 4070 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1541_
timestamp 0
transform 1 0 4450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1543_
timestamp 0
transform 1 0 4370 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1545_
timestamp 0
transform 1 0 5070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1546_
timestamp 0
transform 1 0 5530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1548_
timestamp 0
transform -1 0 6230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1550_
timestamp 0
transform 1 0 5630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1551_
timestamp 0
transform 1 0 1970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1553_
timestamp 0
transform 1 0 3490 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1554_
timestamp 0
transform -1 0 4150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1556_
timestamp 0
transform 1 0 5330 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1558_
timestamp 0
transform 1 0 5890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1559_
timestamp 0
transform 1 0 6050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1561_
timestamp 0
transform -1 0 5690 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1562_
timestamp 0
transform 1 0 5510 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1564_
timestamp 0
transform 1 0 4790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1566_
timestamp 0
transform 1 0 4510 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1567_
timestamp 0
transform 1 0 3910 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1569_
timestamp 0
transform -1 0 5270 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1570_
timestamp 0
transform -1 0 5750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1572_
timestamp 0
transform -1 0 5390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1574_
timestamp 0
transform 1 0 2130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1575_
timestamp 0
transform 1 0 2070 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1577_
timestamp 0
transform 1 0 2210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1579_
timestamp 0
transform 1 0 2090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1580_
timestamp 0
transform 1 0 2450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1582_
timestamp 0
transform 1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1583_
timestamp 0
transform -1 0 5110 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1585_
timestamp 0
transform -1 0 4770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1587_
timestamp 0
transform 1 0 2630 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1588_
timestamp 0
transform 1 0 2670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1590_
timestamp 0
transform -1 0 3050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1591_
timestamp 0
transform 1 0 3450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1593_
timestamp 0
transform -1 0 2750 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1595_
timestamp 0
transform 1 0 2590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1596_
timestamp 0
transform 1 0 2430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1598_
timestamp 0
transform 1 0 4030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1600_
timestamp 0
transform 1 0 2650 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1601_
timestamp 0
transform 1 0 3770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1603_
timestamp 0
transform 1 0 2890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1604_
timestamp 0
transform 1 0 2830 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1606_
timestamp 0
transform 1 0 3470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1608_
timestamp 0
transform -1 0 3630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1636_
timestamp 0
transform -1 0 250 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1638_
timestamp 0
transform -1 0 90 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1639_
timestamp 0
transform -1 0 90 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1641_
timestamp 0
transform 1 0 1090 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1643_
timestamp 0
transform -1 0 990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1644_
timestamp 0
transform 1 0 950 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1646_
timestamp 0
transform 1 0 770 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1647_
timestamp 0
transform 1 0 190 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1649_
timestamp 0
transform -1 0 530 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1651_
timestamp 0
transform -1 0 230 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1652_
timestamp 0
transform -1 0 370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1654_
timestamp 0
transform -1 0 490 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1656_
timestamp 0
transform 1 0 370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1657_
timestamp 0
transform 1 0 870 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1659_
timestamp 0
transform 1 0 1510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1660_
timestamp 0
transform -1 0 1050 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1662_
timestamp 0
transform 1 0 1810 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1664_
timestamp 0
transform 1 0 1330 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1665_
timestamp 0
transform -1 0 1750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1667_
timestamp 0
transform 1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1668_
timestamp 0
transform 1 0 1650 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1670_
timestamp 0
transform 1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1672_
timestamp 0
transform 1 0 1390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1673_
timestamp 0
transform -1 0 1570 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1675_
timestamp 0
transform -1 0 370 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1677_
timestamp 0
transform -1 0 830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1678_
timestamp 0
transform 1 0 70 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1680_
timestamp 0
transform -1 0 370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1681_
timestamp 0
transform -1 0 490 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__1683_
timestamp 0
transform 1 0 490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1685_
timestamp 0
transform 1 0 1570 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1686_
timestamp 0
transform 1 0 1830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1688_
timestamp 0
transform 1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1689_
timestamp 0
transform 1 0 2010 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1691_
timestamp 0
transform 1 0 1850 0 1 3390
box -6 -8 26 268
use FILL  FILL_3__1693_
timestamp 0
transform -1 0 1370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1694_
timestamp 0
transform 1 0 1170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1696_
timestamp 0
transform -1 0 890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1697_
timestamp 0
transform -1 0 1030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1699_
timestamp 0
transform 1 0 610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1701_
timestamp 0
transform 1 0 1290 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1702_
timestamp 0
transform -1 0 1470 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1704_
timestamp 0
transform 1 0 2210 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1706_
timestamp 0
transform -1 0 890 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1707_
timestamp 0
transform -1 0 1790 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1709_
timestamp 0
transform -1 0 1510 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1710_
timestamp 0
transform -1 0 1770 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1712_
timestamp 0
transform 1 0 1310 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1714_
timestamp 0
transform 1 0 1410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1715_
timestamp 0
transform -1 0 1130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1717_
timestamp 0
transform 1 0 1230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1718_
timestamp 0
transform 1 0 1390 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1720_
timestamp 0
transform 1 0 1710 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1722_
timestamp 0
transform -1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1723_
timestamp 0
transform -1 0 1870 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1725_
timestamp 0
transform -1 0 1570 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1727_
timestamp 0
transform -1 0 1790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1728_
timestamp 0
transform -1 0 1190 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1730_
timestamp 0
transform 1 0 1430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1731_
timestamp 0
transform 1 0 1090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1733_
timestamp 0
transform -1 0 1290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1735_
timestamp 0
transform -1 0 1090 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1736_
timestamp 0
transform 1 0 1210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1738_
timestamp 0
transform 1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1739_
timestamp 0
transform -1 0 1650 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1741_
timestamp 0
transform -1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1743_
timestamp 0
transform -1 0 930 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1744_
timestamp 0
transform 1 0 810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1746_
timestamp 0
transform -1 0 770 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1747_
timestamp 0
transform -1 0 670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1749_
timestamp 0
transform 1 0 630 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1751_
timestamp 0
transform 1 0 730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1752_
timestamp 0
transform 1 0 950 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1754_
timestamp 0
transform 1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1756_
timestamp 0
transform -1 0 230 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1757_
timestamp 0
transform -1 0 850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1759_
timestamp 0
transform -1 0 470 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1760_
timestamp 0
transform -1 0 690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1762_
timestamp 0
transform 1 0 330 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1764_
timestamp 0
transform -1 0 550 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1765_
timestamp 0
transform -1 0 390 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1767_
timestamp 0
transform 1 0 2190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1768_
timestamp 0
transform -1 0 2070 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1770_
timestamp 0
transform 1 0 1510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1772_
timestamp 0
transform 1 0 1030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1773_
timestamp 0
transform 1 0 350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1775_
timestamp 0
transform -1 0 1290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1777_
timestamp 0
transform -1 0 90 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1778_
timestamp 0
transform -1 0 230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1780_
timestamp 0
transform -1 0 330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1781_
timestamp 0
transform 1 0 350 0 1 3910
box -6 -8 26 268
use FILL  FILL_3__1783_
timestamp 0
transform -1 0 90 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1785_
timestamp 0
transform -1 0 90 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1786_
timestamp 0
transform 1 0 70 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1788_
timestamp 0
transform -1 0 490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1789_
timestamp 0
transform 1 0 70 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1791_
timestamp 0
transform 1 0 1010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1793_
timestamp 0
transform 1 0 1930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1794_
timestamp 0
transform -1 0 1850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1796_
timestamp 0
transform 1 0 1830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1798_
timestamp 0
transform 1 0 390 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1799_
timestamp 0
transform 1 0 690 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1801_
timestamp 0
transform -1 0 1570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1802_
timestamp 0
transform -1 0 330 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1804_
timestamp 0
transform 1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1806_
timestamp 0
transform 1 0 190 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1807_
timestamp 0
transform -1 0 1230 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1809_
timestamp 0
transform 1 0 230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1810_
timestamp 0
transform 1 0 390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__1812_
timestamp 0
transform 1 0 830 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1814_
timestamp 0
transform 1 0 1370 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1815_
timestamp 0
transform 1 0 1650 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1817_
timestamp 0
transform -1 0 1830 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1818_
timestamp 0
transform 1 0 4690 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1820_
timestamp 0
transform 1 0 3870 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1822_
timestamp 0
transform 1 0 2810 0 1 5990
box -6 -8 26 268
use FILL  FILL_3__1823_
timestamp 0
transform -1 0 4850 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1825_
timestamp 0
transform -1 0 5050 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1827_
timestamp 0
transform 1 0 6130 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert0
timestamp 0
transform 1 0 2450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert1
timestamp 0
transform -1 0 1930 0 1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform 1 0 2510 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert4
timestamp 0
transform -1 0 910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert6
timestamp 0
transform -1 0 2150 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform 1 0 2890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform 1 0 4030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform -1 0 3050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert21
timestamp 0
transform 1 0 3870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert22
timestamp 0
transform -1 0 2890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert24
timestamp 0
transform 1 0 3010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert25
timestamp 0
transform -1 0 3050 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert27
timestamp 0
transform -1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert29
timestamp 0
transform 1 0 4030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert30
timestamp 0
transform 1 0 2730 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert32
timestamp 0
transform 1 0 1930 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert33
timestamp 0
transform -1 0 3170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert35
timestamp 0
transform -1 0 2290 0 1 2870
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert37
timestamp 0
transform -1 0 1210 0 1 2350
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert38
timestamp 0
transform -1 0 250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert40
timestamp 0
transform -1 0 970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert41
timestamp 0
transform 1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert8
timestamp 0
transform -1 0 3670 0 1 4430
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert9
timestamp 0
transform 1 0 4530 0 1 4950
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert11
timestamp 0
transform -1 0 3250 0 1 5470
box -6 -8 26 268
use FILL  FILL_3_CLKBUF1_insert12
timestamp 0
transform -1 0 3410 0 1 4430
box -6 -8 26 268
<< labels >>
flabel metal1 s 6323 2 6383 2 0 FreeSans 48 0 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 0 FreeSans 48 0 0 0 vdd
port 1 nsew
flabel metal2 s 1957 6297 1963 6303 0 FreeSans 48 0 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 1697 6297 1703 6303 0 FreeSans 48 0 0 0 ABCmd_i[6]
port 3 nsew
flabel metal3 s -24 3556 -16 3564 0 FreeSans 64 0 0 0 ABCmd_i[5]
port 4 nsew
flabel metal3 s -24 3516 -16 3524 0 FreeSans 64 0 0 0 ABCmd_i[4]
port 5 nsew
flabel metal3 s -24 4556 -16 4564 0 FreeSans 64 0 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s -24 4336 -16 4344 0 FreeSans 64 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal3 s -24 2776 -16 2784 0 FreeSans 64 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s -24 2956 -16 2964 0 FreeSans 64 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal2 s 5077 6297 5083 6303 0 FreeSans 48 0 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 4597 6297 4603 6303 0 FreeSans 48 0 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 4877 6297 4883 6303 0 FreeSans 48 0 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 2857 6297 2863 6303 0 FreeSans 48 0 0 0 ACC_o[4]
port 13 nsew
flabel metal3 s 6356 5336 6364 5344 0 FreeSans 64 0 0 0 ACC_o[3]
port 14 nsew
flabel metal2 s 3917 6297 3923 6303 0 FreeSans 48 0 0 0 ACC_o[2]
port 15 nsew
flabel metal2 s 2137 6297 2143 6303 0 FreeSans 48 0 0 0 ACC_o[1]
port 16 nsew
flabel metal2 s 4737 6297 4743 6303 0 FreeSans 48 0 0 0 ACC_o[0]
port 17 nsew
flabel metal3 s 6356 5856 6364 5864 0 FreeSans 64 0 0 0 Done_LED
port 18 nsew
flabel metal3 s 6356 5596 6364 5604 0 FreeSans 64 0 0 0 Done_o
port 19 nsew
flabel metal2 s 5857 6297 5863 6303 0 FreeSans 48 0 0 0 LoadA_i
port 20 nsew
flabel metal2 s 5697 6297 5703 6303 0 FreeSans 48 0 0 0 LoadB_i
port 21 nsew
flabel metal3 s 6356 6116 6364 6124 0 FreeSans 64 0 0 0 LoadCmd_i
port 22 nsew
flabel metal2 s 3337 6297 3343 6303 0 FreeSans 48 0 0 0 clk
port 23 nsew
flabel metal2 s 2917 6297 2923 6303 0 FreeSans 48 0 0 0 reset
port 24 nsew
<< properties >>
string FIXED_BBOX -40 0 6360 6300
<< end >>
